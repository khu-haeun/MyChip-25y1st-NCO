magic
tech scmos
magscale 1 3
timestamp 1569533753
<< checkpaint >>
rect -60 -60 80 80
<< metal2 >>
rect 0 14 20 20
rect 0 6 6 14
rect 14 6 20 14
rect 0 0 20 6
<< m3contact >>
rect 6 6 14 14
<< metal3 >>
rect 0 14 20 20
rect 0 6 6 14
rect 14 6 20 14
rect 0 0 20 6
<< end >>
