magic
tech scmos
magscale 1 30
timestamp 1740920094
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 58800 142500 135100 145100
rect 48400 131200 50400 138500
rect 48400 129400 56200 131200
rect 133300 130900 135100 142500
<< m2contact >>
rect 50200 142500 58800 145100
rect 46200 132500 48400 138500
<< metal2 >>
rect 50200 145100 58800 145900
rect 44100 132500 46200 138500
rect 62400 133600 62900 145900
rect 75900 134600 76400 145900
rect 89400 136400 89900 145900
rect 102900 135400 103400 145900
rect 127200 142000 127700 145900
rect 140700 142000 141200 145900
rect 126600 141500 127700 142000
rect 130100 141600 141200 142000
rect 102900 135000 122300 135400
rect 75900 134100 121600 134600
rect 62400 133100 87900 133600
rect 87400 132000 87900 133100
rect 121200 131900 121600 134100
rect 121900 131900 122300 135000
rect 122600 131900 123000 135900
rect 126600 131700 127100 141500
rect 130100 131900 130500 141600
rect 138600 140800 145900 141200
rect 44100 116200 44800 116900
rect 44100 102700 46200 103400
rect 48100 89800 48500 122000
rect 44100 89400 48500 89800
rect 48900 76300 49300 125500
rect 44100 75900 49300 76300
rect 49700 62800 50100 126300
rect 44100 62400 50100 62800
rect 50500 49200 50900 127100
rect 138600 83600 139000 140800
rect 139400 127300 145900 127700
rect 139400 90800 139800 127300
rect 140200 113700 145900 114100
rect 142500 100300 145900 100700
rect 143300 86800 145900 87200
rect 144100 73300 145900 73700
rect 144900 59800 145900 60200
rect 58750 52750 59150 58900
rect 59450 53850 59750 58900
rect 60000 58700 60800 58900
rect 60300 54900 60800 58700
rect 63900 55900 64400 58900
rect 101400 56900 101900 58900
rect 113700 57900 114200 58900
rect 113700 57400 127700 57900
rect 101400 56400 114200 56900
rect 63900 55400 100700 55900
rect 60300 54400 87200 54900
rect 59450 53300 73700 53850
rect 58750 52200 60200 52750
rect 44100 48800 50900 49200
rect 59700 44100 60200 52200
rect 73200 44100 73700 53300
rect 86700 44100 87200 54400
rect 100200 44100 100700 55400
rect 113700 44100 114200 56400
rect 127200 44100 127700 57400
rect 129800 46000 130300 58900
rect 129800 45500 141200 46000
rect 140700 44100 141200 45500
<< m3contact >>
rect 89400 135900 90900 136400
rect 121500 135900 123000 136400
rect 50500 127100 50900 127500
rect 49700 126300 50100 126700
rect 48900 125500 49300 125900
rect 48100 122000 48500 122400
rect 44800 114800 45500 116900
rect 46200 101300 46900 103400
rect 140200 114100 140600 115200
rect 142100 100300 142500 101500
rect 139400 89600 139800 90800
rect 142900 86800 143300 88000
rect 138600 82400 139000 83600
rect 143700 73300 144100 74500
rect 144500 59800 144900 61000
<< metal3 >>
rect 90900 135900 121500 136400
rect 133700 131000 144900 131400
rect 133700 130300 144100 130700
rect 133700 129600 143300 130000
rect 133700 128900 142500 129300
rect 50900 127100 56400 127500
rect 50100 126300 56400 126700
rect 49300 125500 56400 125900
rect 48500 122000 56400 122400
rect 133700 114800 140200 115200
rect 44800 93800 45500 114800
rect 46200 95200 46900 101300
rect 142100 101500 142500 128900
rect 46200 94500 56500 95200
rect 55800 94100 56500 94500
rect 44800 93100 56500 93800
rect 133700 89600 139400 90000
rect 142900 88000 143300 129600
rect 133700 82400 138600 82800
rect 143700 74500 144100 130300
rect 144500 61000 144900 131000
<< end >>
