magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -127 -120 1127 5132
<< nwell >>
rect -7 4201 1007 4571
rect -7 2241 1007 3839
<< psubstratepdiff >>
rect 20 4680 980 5012
rect 20 0 980 1560
<< nsubstratendiff >>
rect 20 4220 980 4552
rect 20 2260 980 3820
<< metal1 >>
rect 24 4680 976 5012
rect 24 4220 976 4552
rect 24 2260 976 3820
rect 24 0 976 1560
<< metal2 >>
rect 24 4680 976 5012
rect 24 4220 976 4552
rect 24 2260 976 3820
rect 24 0 976 1560
<< metal3 >>
rect 0 4680 1000 5012
rect 0 4220 1000 4552
rect 0 2260 1000 3820
rect 0 0 1000 1560
use CONT$5  CONT$5_0
array 0 13 64 0 23 64
timestamp 1569543463
transform 1 0 104 0 1 22
box -6 -6 6 6
use CONT$5  CONT$5_1
array 0 14 64 0 23 64
timestamp 1569543463
transform 1 0 48 0 1 2300
box -6 -6 6 6
use CONT$5  CONT$5_2
array 0 14 64 0 3 64
timestamp 1569543463
transform 1 0 48 0 1 4264
box -6 -6 6 6
use CONT$5  CONT$5_3
array 0 14 64 0 3 64
timestamp 1569543463
transform 1 0 48 0 1 4740
box -6 -6 6 6
use VIA1$6  VIA1$6_0
array 0 13 64 0 22 64
timestamp 1569543463
transform 1 0 80 0 1 2332
box -8 -8 8 8
use VIA1$6  VIA1$6_1
array 0 13 64 0 22 64
timestamp 1569543463
transform 1 0 72 0 1 54
box -8 -8 8 8
use VIA1$6  VIA1$6_2
array 0 13 64 0 2 64
timestamp 1569543463
transform 1 0 80 0 1 4296
box -8 -8 8 8
use VIA1$6  VIA1$6_3
array 0 13 64 0 2 64
timestamp 1569543463
transform 1 0 80 0 1 4772
box -8 -8 8 8
use VIA2$6  VIA2$6_0
array 0 13 64 0 23 64
timestamp 1569543463
transform 1 0 104 0 1 22
box -8 -8 8 8
use VIA2$6  VIA2$6_1
array 0 14 64 0 23 64
timestamp 1569543463
transform 1 0 48 0 1 2300
box -8 -8 8 8
use VIA2$6  VIA2$6_2
array 0 14 64 0 3 64
timestamp 1569543463
transform 1 0 48 0 1 4264
box -8 -8 8 8
use VIA2$6  VIA2$6_3
array 0 14 64 0 3 64
timestamp 1569543463
transform 1 0 48 0 1 4740
box -8 -8 8 8
<< end >>
