magic
tech scmos
magscale 1 6
timestamp 1569536352
<< checkpaint >>
rect 8700 8700 29300 29300
<< metal1 >>
rect 11760 29019 27020 29020
rect 10041 29008 27020 29019
rect 10041 28992 10060 29008
rect 10076 28992 10092 29008
rect 10108 28992 10124 29008
rect 10140 28992 10156 29008
rect 10172 28992 10188 29008
rect 10204 28992 10220 29008
rect 10236 28992 10252 29008
rect 10268 28992 10284 29008
rect 10300 28992 10316 29008
rect 10332 28992 10348 29008
rect 10364 28992 10380 29008
rect 10396 28992 10412 29008
rect 10428 28992 10444 29008
rect 10460 28992 10476 29008
rect 10492 28992 10508 29008
rect 10524 28992 10540 29008
rect 10556 28992 10572 29008
rect 10588 28992 10604 29008
rect 10620 28992 10636 29008
rect 10652 28992 10668 29008
rect 10684 28992 10700 29008
rect 10716 28992 10732 29008
rect 10748 28992 10764 29008
rect 10780 28992 10796 29008
rect 10812 28992 10828 29008
rect 10844 28992 10860 29008
rect 10876 28992 10892 29008
rect 10908 28992 10924 29008
rect 10940 28992 10956 29008
rect 10972 28992 10988 29008
rect 11004 28992 11020 29008
rect 11036 28992 11052 29008
rect 11068 28992 11084 29008
rect 11100 28992 11116 29008
rect 11132 28992 11148 29008
rect 11164 28992 11180 29008
rect 11196 28992 11212 29008
rect 11228 28992 11244 29008
rect 11260 28992 11276 29008
rect 11292 28992 11308 29008
rect 11324 28992 11340 29008
rect 11356 28992 11372 29008
rect 11388 28992 11404 29008
rect 11420 28992 11436 29008
rect 11452 28992 11468 29008
rect 11484 28992 11500 29008
rect 11516 28992 11532 29008
rect 11548 28992 11564 29008
rect 11580 28992 11596 29008
rect 11612 28992 11628 29008
rect 11644 28992 11660 29008
rect 11676 28992 11692 29008
rect 11708 28992 11724 29008
rect 11740 28992 27020 29008
rect 10041 28976 27020 28992
rect 10041 28960 10060 28976
rect 10076 28960 10092 28976
rect 10108 28960 10124 28976
rect 10140 28960 10156 28976
rect 10172 28960 10188 28976
rect 10204 28960 10220 28976
rect 10236 28960 10252 28976
rect 10268 28960 10284 28976
rect 10300 28960 10316 28976
rect 10332 28960 10348 28976
rect 10364 28960 10380 28976
rect 10396 28960 10412 28976
rect 10428 28960 10444 28976
rect 10460 28960 10476 28976
rect 10492 28960 10508 28976
rect 10524 28960 10540 28976
rect 10556 28960 10572 28976
rect 10588 28960 10604 28976
rect 10620 28960 10636 28976
rect 10652 28960 10668 28976
rect 10684 28960 10700 28976
rect 10716 28960 10732 28976
rect 10748 28960 10764 28976
rect 10780 28960 10796 28976
rect 10812 28960 10828 28976
rect 10844 28960 10860 28976
rect 10876 28960 10892 28976
rect 10908 28960 10924 28976
rect 10940 28960 10956 28976
rect 10972 28960 10988 28976
rect 11004 28960 11020 28976
rect 11036 28960 11052 28976
rect 11068 28960 11084 28976
rect 11100 28960 11116 28976
rect 11132 28960 11148 28976
rect 11164 28960 11180 28976
rect 11196 28960 11212 28976
rect 11228 28960 11244 28976
rect 11260 28960 11276 28976
rect 11292 28960 11308 28976
rect 11324 28960 11340 28976
rect 11356 28960 11372 28976
rect 11388 28960 11404 28976
rect 11420 28960 11436 28976
rect 11452 28960 11468 28976
rect 11484 28960 11500 28976
rect 11516 28960 11532 28976
rect 11548 28960 11564 28976
rect 11580 28960 11596 28976
rect 11612 28960 11628 28976
rect 11644 28960 11660 28976
rect 11676 28960 11692 28976
rect 11708 28960 11724 28976
rect 11740 28960 27020 28976
rect 10041 28944 27020 28960
rect 10041 28928 10060 28944
rect 10076 28928 10092 28944
rect 10108 28928 10124 28944
rect 10140 28928 10156 28944
rect 10172 28928 10188 28944
rect 10204 28928 10220 28944
rect 10236 28928 10252 28944
rect 10268 28928 10284 28944
rect 10300 28928 10316 28944
rect 10332 28928 10348 28944
rect 10364 28928 10380 28944
rect 10396 28928 10412 28944
rect 10428 28928 10444 28944
rect 10460 28928 10476 28944
rect 10492 28928 10508 28944
rect 10524 28928 10540 28944
rect 10556 28928 10572 28944
rect 10588 28928 10604 28944
rect 10620 28928 10636 28944
rect 10652 28928 10668 28944
rect 10684 28928 10700 28944
rect 10716 28928 10732 28944
rect 10748 28928 10764 28944
rect 10780 28928 10796 28944
rect 10812 28928 10828 28944
rect 10844 28928 10860 28944
rect 10876 28928 10892 28944
rect 10908 28928 10924 28944
rect 10940 28928 10956 28944
rect 10972 28928 10988 28944
rect 11004 28928 11020 28944
rect 11036 28928 11052 28944
rect 11068 28928 11084 28944
rect 11100 28928 11116 28944
rect 11132 28928 11148 28944
rect 11164 28928 11180 28944
rect 11196 28928 11212 28944
rect 11228 28928 11244 28944
rect 11260 28928 11276 28944
rect 11292 28928 11308 28944
rect 11324 28928 11340 28944
rect 11356 28928 11372 28944
rect 11388 28928 11404 28944
rect 11420 28928 11436 28944
rect 11452 28928 11468 28944
rect 11484 28928 11500 28944
rect 11516 28928 11532 28944
rect 11548 28928 11564 28944
rect 11580 28928 11596 28944
rect 11612 28928 11628 28944
rect 11644 28928 11660 28944
rect 11676 28928 11692 28944
rect 11708 28928 11724 28944
rect 11740 28928 27020 28944
rect 10041 28912 27020 28928
rect 10041 28896 10060 28912
rect 10076 28896 10092 28912
rect 10108 28896 10124 28912
rect 10140 28896 10156 28912
rect 10172 28896 10188 28912
rect 10204 28896 10220 28912
rect 10236 28896 10252 28912
rect 10268 28896 10284 28912
rect 10300 28896 10316 28912
rect 10332 28896 10348 28912
rect 10364 28896 10380 28912
rect 10396 28896 10412 28912
rect 10428 28896 10444 28912
rect 10460 28896 10476 28912
rect 10492 28896 10508 28912
rect 10524 28896 10540 28912
rect 10556 28896 10572 28912
rect 10588 28896 10604 28912
rect 10620 28896 10636 28912
rect 10652 28896 10668 28912
rect 10684 28896 10700 28912
rect 10716 28896 10732 28912
rect 10748 28896 10764 28912
rect 10780 28896 10796 28912
rect 10812 28896 10828 28912
rect 10844 28896 10860 28912
rect 10876 28896 10892 28912
rect 10908 28896 10924 28912
rect 10940 28896 10956 28912
rect 10972 28896 10988 28912
rect 11004 28896 11020 28912
rect 11036 28896 11052 28912
rect 11068 28896 11084 28912
rect 11100 28896 11116 28912
rect 11132 28896 11148 28912
rect 11164 28896 11180 28912
rect 11196 28896 11212 28912
rect 11228 28896 11244 28912
rect 11260 28896 11276 28912
rect 11292 28896 11308 28912
rect 11324 28896 11340 28912
rect 11356 28896 11372 28912
rect 11388 28896 11404 28912
rect 11420 28896 11436 28912
rect 11452 28896 11468 28912
rect 11484 28896 11500 28912
rect 11516 28896 11532 28912
rect 11548 28896 11564 28912
rect 11580 28896 11596 28912
rect 11612 28896 11628 28912
rect 11644 28896 11660 28912
rect 11676 28896 11692 28912
rect 11708 28896 11724 28912
rect 11740 28896 27020 28912
rect 10041 28880 27020 28896
rect 10041 28864 10060 28880
rect 10076 28864 10092 28880
rect 10108 28864 10124 28880
rect 10140 28864 10156 28880
rect 10172 28864 10188 28880
rect 10204 28864 10220 28880
rect 10236 28864 10252 28880
rect 10268 28864 10284 28880
rect 10300 28864 10316 28880
rect 10332 28864 10348 28880
rect 10364 28864 10380 28880
rect 10396 28864 10412 28880
rect 10428 28864 10444 28880
rect 10460 28864 10476 28880
rect 10492 28864 10508 28880
rect 10524 28864 10540 28880
rect 10556 28864 10572 28880
rect 10588 28864 10604 28880
rect 10620 28864 10636 28880
rect 10652 28864 10668 28880
rect 10684 28864 10700 28880
rect 10716 28864 10732 28880
rect 10748 28864 10764 28880
rect 10780 28864 10796 28880
rect 10812 28864 10828 28880
rect 10844 28864 10860 28880
rect 10876 28864 10892 28880
rect 10908 28864 10924 28880
rect 10940 28864 10956 28880
rect 10972 28864 10988 28880
rect 11004 28864 11020 28880
rect 11036 28864 11052 28880
rect 11068 28864 11084 28880
rect 11100 28864 11116 28880
rect 11132 28864 11148 28880
rect 11164 28864 11180 28880
rect 11196 28864 11212 28880
rect 11228 28864 11244 28880
rect 11260 28864 11276 28880
rect 11292 28864 11308 28880
rect 11324 28864 11340 28880
rect 11356 28864 11372 28880
rect 11388 28864 11404 28880
rect 11420 28864 11436 28880
rect 11452 28864 11468 28880
rect 11484 28864 11500 28880
rect 11516 28864 11532 28880
rect 11548 28864 11564 28880
rect 11580 28864 11596 28880
rect 11612 28864 11628 28880
rect 11644 28864 11660 28880
rect 11676 28864 11692 28880
rect 11708 28864 11724 28880
rect 11740 28864 27020 28880
rect 10041 28848 27020 28864
rect 10041 28832 10060 28848
rect 10076 28832 10092 28848
rect 10108 28832 10124 28848
rect 10140 28832 10156 28848
rect 10172 28832 10188 28848
rect 10204 28832 10220 28848
rect 10236 28832 10252 28848
rect 10268 28832 10284 28848
rect 10300 28832 10316 28848
rect 10332 28832 10348 28848
rect 10364 28832 10380 28848
rect 10396 28832 10412 28848
rect 10428 28832 10444 28848
rect 10460 28832 10476 28848
rect 10492 28832 10508 28848
rect 10524 28832 10540 28848
rect 10556 28832 10572 28848
rect 10588 28832 10604 28848
rect 10620 28832 10636 28848
rect 10652 28832 10668 28848
rect 10684 28832 10700 28848
rect 10716 28832 10732 28848
rect 10748 28832 10764 28848
rect 10780 28832 10796 28848
rect 10812 28832 10828 28848
rect 10844 28832 10860 28848
rect 10876 28832 10892 28848
rect 10908 28832 10924 28848
rect 10940 28832 10956 28848
rect 10972 28832 10988 28848
rect 11004 28832 11020 28848
rect 11036 28832 11052 28848
rect 11068 28832 11084 28848
rect 11100 28832 11116 28848
rect 11132 28832 11148 28848
rect 11164 28832 11180 28848
rect 11196 28832 11212 28848
rect 11228 28832 11244 28848
rect 11260 28832 11276 28848
rect 11292 28832 11308 28848
rect 11324 28832 11340 28848
rect 11356 28832 11372 28848
rect 11388 28832 11404 28848
rect 11420 28832 11436 28848
rect 11452 28832 11468 28848
rect 11484 28832 11500 28848
rect 11516 28832 11532 28848
rect 11548 28832 11564 28848
rect 11580 28832 11596 28848
rect 11612 28832 11628 28848
rect 11644 28832 11660 28848
rect 11676 28832 11692 28848
rect 11708 28832 11724 28848
rect 11740 28832 27020 28848
rect 10041 28816 27020 28832
rect 10041 28800 10060 28816
rect 10076 28800 10092 28816
rect 10108 28800 10124 28816
rect 10140 28800 10156 28816
rect 10172 28800 10188 28816
rect 10204 28800 10220 28816
rect 10236 28800 10252 28816
rect 10268 28800 10284 28816
rect 10300 28800 10316 28816
rect 10332 28800 10348 28816
rect 10364 28800 10380 28816
rect 10396 28800 10412 28816
rect 10428 28800 10444 28816
rect 10460 28800 10476 28816
rect 10492 28800 10508 28816
rect 10524 28800 10540 28816
rect 10556 28800 10572 28816
rect 10588 28800 10604 28816
rect 10620 28800 10636 28816
rect 10652 28800 10668 28816
rect 10684 28800 10700 28816
rect 10716 28800 10732 28816
rect 10748 28800 10764 28816
rect 10780 28800 10796 28816
rect 10812 28800 10828 28816
rect 10844 28800 10860 28816
rect 10876 28800 10892 28816
rect 10908 28800 10924 28816
rect 10940 28800 10956 28816
rect 10972 28800 10988 28816
rect 11004 28800 11020 28816
rect 11036 28800 11052 28816
rect 11068 28800 11084 28816
rect 11100 28800 11116 28816
rect 11132 28800 11148 28816
rect 11164 28800 11180 28816
rect 11196 28800 11212 28816
rect 11228 28800 11244 28816
rect 11260 28800 11276 28816
rect 11292 28800 11308 28816
rect 11324 28800 11340 28816
rect 11356 28800 11372 28816
rect 11388 28800 11404 28816
rect 11420 28800 11436 28816
rect 11452 28800 11468 28816
rect 11484 28800 11500 28816
rect 11516 28800 11532 28816
rect 11548 28800 11564 28816
rect 11580 28800 11596 28816
rect 11612 28800 11628 28816
rect 11644 28800 11660 28816
rect 11676 28800 11692 28816
rect 11708 28800 11724 28816
rect 11740 28800 27020 28816
rect 10041 28784 27020 28800
rect 10041 28768 10060 28784
rect 10076 28768 10092 28784
rect 10108 28768 10124 28784
rect 10140 28768 10156 28784
rect 10172 28768 10188 28784
rect 10204 28768 10220 28784
rect 10236 28768 10252 28784
rect 10268 28768 10284 28784
rect 10300 28768 10316 28784
rect 10332 28768 10348 28784
rect 10364 28768 10380 28784
rect 10396 28768 10412 28784
rect 10428 28768 10444 28784
rect 10460 28768 10476 28784
rect 10492 28768 10508 28784
rect 10524 28768 10540 28784
rect 10556 28768 10572 28784
rect 10588 28768 10604 28784
rect 10620 28768 10636 28784
rect 10652 28768 10668 28784
rect 10684 28768 10700 28784
rect 10716 28768 10732 28784
rect 10748 28768 10764 28784
rect 10780 28768 10796 28784
rect 10812 28768 10828 28784
rect 10844 28768 10860 28784
rect 10876 28768 10892 28784
rect 10908 28768 10924 28784
rect 10940 28768 10956 28784
rect 10972 28768 10988 28784
rect 11004 28768 11020 28784
rect 11036 28768 11052 28784
rect 11068 28768 11084 28784
rect 11100 28768 11116 28784
rect 11132 28768 11148 28784
rect 11164 28768 11180 28784
rect 11196 28768 11212 28784
rect 11228 28768 11244 28784
rect 11260 28768 11276 28784
rect 11292 28768 11308 28784
rect 11324 28768 11340 28784
rect 11356 28768 11372 28784
rect 11388 28768 11404 28784
rect 11420 28768 11436 28784
rect 11452 28768 11468 28784
rect 11484 28768 11500 28784
rect 11516 28768 11532 28784
rect 11548 28768 11564 28784
rect 11580 28768 11596 28784
rect 11612 28768 11628 28784
rect 11644 28768 11660 28784
rect 11676 28768 11692 28784
rect 11708 28768 11724 28784
rect 11740 28768 27020 28784
rect 10041 28752 27020 28768
rect 10041 28736 10060 28752
rect 10076 28736 10092 28752
rect 10108 28736 10124 28752
rect 10140 28736 10156 28752
rect 10172 28736 10188 28752
rect 10204 28736 10220 28752
rect 10236 28736 10252 28752
rect 10268 28736 10284 28752
rect 10300 28736 10316 28752
rect 10332 28736 10348 28752
rect 10364 28736 10380 28752
rect 10396 28736 10412 28752
rect 10428 28736 10444 28752
rect 10460 28736 10476 28752
rect 10492 28736 10508 28752
rect 10524 28736 10540 28752
rect 10556 28736 10572 28752
rect 10588 28736 10604 28752
rect 10620 28736 10636 28752
rect 10652 28736 10668 28752
rect 10684 28736 10700 28752
rect 10716 28736 10732 28752
rect 10748 28736 10764 28752
rect 10780 28736 10796 28752
rect 10812 28736 10828 28752
rect 10844 28736 10860 28752
rect 10876 28736 10892 28752
rect 10908 28736 10924 28752
rect 10940 28736 10956 28752
rect 10972 28736 10988 28752
rect 11004 28736 11020 28752
rect 11036 28736 11052 28752
rect 11068 28736 11084 28752
rect 11100 28736 11116 28752
rect 11132 28736 11148 28752
rect 11164 28736 11180 28752
rect 11196 28736 11212 28752
rect 11228 28736 11244 28752
rect 11260 28736 11276 28752
rect 11292 28736 11308 28752
rect 11324 28736 11340 28752
rect 11356 28736 11372 28752
rect 11388 28736 11404 28752
rect 11420 28736 11436 28752
rect 11452 28736 11468 28752
rect 11484 28736 11500 28752
rect 11516 28736 11532 28752
rect 11548 28736 11564 28752
rect 11580 28736 11596 28752
rect 11612 28736 11628 28752
rect 11644 28736 11660 28752
rect 11676 28736 11692 28752
rect 11708 28736 11724 28752
rect 11740 28736 27020 28752
rect 10041 28720 27020 28736
rect 10041 28704 10060 28720
rect 10076 28704 10092 28720
rect 10108 28704 10124 28720
rect 10140 28704 10156 28720
rect 10172 28704 10188 28720
rect 10204 28704 10220 28720
rect 10236 28704 10252 28720
rect 10268 28704 10284 28720
rect 10300 28704 10316 28720
rect 10332 28704 10348 28720
rect 10364 28704 10380 28720
rect 10396 28704 10412 28720
rect 10428 28704 10444 28720
rect 10460 28704 10476 28720
rect 10492 28704 10508 28720
rect 10524 28704 10540 28720
rect 10556 28704 10572 28720
rect 10588 28704 10604 28720
rect 10620 28704 10636 28720
rect 10652 28704 10668 28720
rect 10684 28704 10700 28720
rect 10716 28704 10732 28720
rect 10748 28704 10764 28720
rect 10780 28704 10796 28720
rect 10812 28704 10828 28720
rect 10844 28704 10860 28720
rect 10876 28704 10892 28720
rect 10908 28704 10924 28720
rect 10940 28704 10956 28720
rect 10972 28704 10988 28720
rect 11004 28704 11020 28720
rect 11036 28704 11052 28720
rect 11068 28704 11084 28720
rect 11100 28704 11116 28720
rect 11132 28704 11148 28720
rect 11164 28704 11180 28720
rect 11196 28704 11212 28720
rect 11228 28704 11244 28720
rect 11260 28704 11276 28720
rect 11292 28704 11308 28720
rect 11324 28704 11340 28720
rect 11356 28704 11372 28720
rect 11388 28704 11404 28720
rect 11420 28704 11436 28720
rect 11452 28704 11468 28720
rect 11484 28704 11500 28720
rect 11516 28704 11532 28720
rect 11548 28704 11564 28720
rect 11580 28704 11596 28720
rect 11612 28704 11628 28720
rect 11644 28704 11660 28720
rect 11676 28704 11692 28720
rect 11708 28704 11724 28720
rect 11740 28704 27020 28720
rect 10041 28688 27020 28704
rect 10041 28672 10060 28688
rect 10076 28672 10092 28688
rect 10108 28672 10124 28688
rect 10140 28672 10156 28688
rect 10172 28672 10188 28688
rect 10204 28672 10220 28688
rect 10236 28672 10252 28688
rect 10268 28672 10284 28688
rect 10300 28672 10316 28688
rect 10332 28672 10348 28688
rect 10364 28672 10380 28688
rect 10396 28672 10412 28688
rect 10428 28672 10444 28688
rect 10460 28672 10476 28688
rect 10492 28672 10508 28688
rect 10524 28672 10540 28688
rect 10556 28672 10572 28688
rect 10588 28672 10604 28688
rect 10620 28672 10636 28688
rect 10652 28672 10668 28688
rect 10684 28672 10700 28688
rect 10716 28672 10732 28688
rect 10748 28672 10764 28688
rect 10780 28672 10796 28688
rect 10812 28672 10828 28688
rect 10844 28672 10860 28688
rect 10876 28672 10892 28688
rect 10908 28672 10924 28688
rect 10940 28672 10956 28688
rect 10972 28672 10988 28688
rect 11004 28672 11020 28688
rect 11036 28672 11052 28688
rect 11068 28672 11084 28688
rect 11100 28672 11116 28688
rect 11132 28672 11148 28688
rect 11164 28672 11180 28688
rect 11196 28672 11212 28688
rect 11228 28672 11244 28688
rect 11260 28672 11276 28688
rect 11292 28672 11308 28688
rect 11324 28672 11340 28688
rect 11356 28672 11372 28688
rect 11388 28672 11404 28688
rect 11420 28672 11436 28688
rect 11452 28672 11468 28688
rect 11484 28672 11500 28688
rect 11516 28672 11532 28688
rect 11548 28672 11564 28688
rect 11580 28672 11596 28688
rect 11612 28672 11628 28688
rect 11644 28672 11660 28688
rect 11676 28672 11692 28688
rect 11708 28672 11724 28688
rect 11740 28672 27020 28688
rect 10041 28656 27020 28672
rect 10041 28640 10060 28656
rect 10076 28640 10092 28656
rect 10108 28640 10124 28656
rect 10140 28640 10156 28656
rect 10172 28640 10188 28656
rect 10204 28640 10220 28656
rect 10236 28640 10252 28656
rect 10268 28640 10284 28656
rect 10300 28640 10316 28656
rect 10332 28640 10348 28656
rect 10364 28640 10380 28656
rect 10396 28640 10412 28656
rect 10428 28640 10444 28656
rect 10460 28640 10476 28656
rect 10492 28640 10508 28656
rect 10524 28640 10540 28656
rect 10556 28640 10572 28656
rect 10588 28640 10604 28656
rect 10620 28640 10636 28656
rect 10652 28640 10668 28656
rect 10684 28640 10700 28656
rect 10716 28640 10732 28656
rect 10748 28640 10764 28656
rect 10780 28640 10796 28656
rect 10812 28640 10828 28656
rect 10844 28640 10860 28656
rect 10876 28640 10892 28656
rect 10908 28640 10924 28656
rect 10940 28640 10956 28656
rect 10972 28640 10988 28656
rect 11004 28640 11020 28656
rect 11036 28640 11052 28656
rect 11068 28640 11084 28656
rect 11100 28640 11116 28656
rect 11132 28640 11148 28656
rect 11164 28640 11180 28656
rect 11196 28640 11212 28656
rect 11228 28640 11244 28656
rect 11260 28640 11276 28656
rect 11292 28640 11308 28656
rect 11324 28640 11340 28656
rect 11356 28640 11372 28656
rect 11388 28640 11404 28656
rect 11420 28640 11436 28656
rect 11452 28640 11468 28656
rect 11484 28640 11500 28656
rect 11516 28640 11532 28656
rect 11548 28640 11564 28656
rect 11580 28640 11596 28656
rect 11612 28640 11628 28656
rect 11644 28640 11660 28656
rect 11676 28640 11692 28656
rect 11708 28640 11724 28656
rect 11740 28640 27020 28656
rect 10041 28624 27020 28640
rect 10041 28608 10060 28624
rect 10076 28608 10092 28624
rect 10108 28608 10124 28624
rect 10140 28608 10156 28624
rect 10172 28608 10188 28624
rect 10204 28608 10220 28624
rect 10236 28608 10252 28624
rect 10268 28608 10284 28624
rect 10300 28608 10316 28624
rect 10332 28608 10348 28624
rect 10364 28608 10380 28624
rect 10396 28608 10412 28624
rect 10428 28608 10444 28624
rect 10460 28608 10476 28624
rect 10492 28608 10508 28624
rect 10524 28608 10540 28624
rect 10556 28608 10572 28624
rect 10588 28608 10604 28624
rect 10620 28608 10636 28624
rect 10652 28608 10668 28624
rect 10684 28608 10700 28624
rect 10716 28608 10732 28624
rect 10748 28608 10764 28624
rect 10780 28608 10796 28624
rect 10812 28608 10828 28624
rect 10844 28608 10860 28624
rect 10876 28608 10892 28624
rect 10908 28608 10924 28624
rect 10940 28608 10956 28624
rect 10972 28608 10988 28624
rect 11004 28608 11020 28624
rect 11036 28608 11052 28624
rect 11068 28608 11084 28624
rect 11100 28608 11116 28624
rect 11132 28608 11148 28624
rect 11164 28608 11180 28624
rect 11196 28608 11212 28624
rect 11228 28608 11244 28624
rect 11260 28608 11276 28624
rect 11292 28608 11308 28624
rect 11324 28608 11340 28624
rect 11356 28608 11372 28624
rect 11388 28608 11404 28624
rect 11420 28608 11436 28624
rect 11452 28608 11468 28624
rect 11484 28608 11500 28624
rect 11516 28608 11532 28624
rect 11548 28608 11564 28624
rect 11580 28608 11596 28624
rect 11612 28608 11628 28624
rect 11644 28608 11660 28624
rect 11676 28608 11692 28624
rect 11708 28608 11724 28624
rect 11740 28608 27020 28624
rect 10041 28592 27020 28608
rect 10041 28576 10060 28592
rect 10076 28576 10092 28592
rect 10108 28576 10124 28592
rect 10140 28576 10156 28592
rect 10172 28576 10188 28592
rect 10204 28576 10220 28592
rect 10236 28576 10252 28592
rect 10268 28576 10284 28592
rect 10300 28576 10316 28592
rect 10332 28576 10348 28592
rect 10364 28576 10380 28592
rect 10396 28576 10412 28592
rect 10428 28576 10444 28592
rect 10460 28576 10476 28592
rect 10492 28576 10508 28592
rect 10524 28576 10540 28592
rect 10556 28576 10572 28592
rect 10588 28576 10604 28592
rect 10620 28576 10636 28592
rect 10652 28576 10668 28592
rect 10684 28576 10700 28592
rect 10716 28576 10732 28592
rect 10748 28576 10764 28592
rect 10780 28576 10796 28592
rect 10812 28576 10828 28592
rect 10844 28576 10860 28592
rect 10876 28576 10892 28592
rect 10908 28576 10924 28592
rect 10940 28576 10956 28592
rect 10972 28576 10988 28592
rect 11004 28576 11020 28592
rect 11036 28576 11052 28592
rect 11068 28576 11084 28592
rect 11100 28576 11116 28592
rect 11132 28576 11148 28592
rect 11164 28576 11180 28592
rect 11196 28576 11212 28592
rect 11228 28576 11244 28592
rect 11260 28576 11276 28592
rect 11292 28576 11308 28592
rect 11324 28576 11340 28592
rect 11356 28576 11372 28592
rect 11388 28576 11404 28592
rect 11420 28576 11436 28592
rect 11452 28576 11468 28592
rect 11484 28576 11500 28592
rect 11516 28576 11532 28592
rect 11548 28576 11564 28592
rect 11580 28576 11596 28592
rect 11612 28576 11628 28592
rect 11644 28576 11660 28592
rect 11676 28576 11692 28592
rect 11708 28576 11724 28592
rect 11740 28576 27020 28592
rect 10041 28560 27020 28576
rect 10041 28544 10060 28560
rect 10076 28544 10092 28560
rect 10108 28544 10124 28560
rect 10140 28544 10156 28560
rect 10172 28544 10188 28560
rect 10204 28544 10220 28560
rect 10236 28544 10252 28560
rect 10268 28544 10284 28560
rect 10300 28544 10316 28560
rect 10332 28544 10348 28560
rect 10364 28544 10380 28560
rect 10396 28544 10412 28560
rect 10428 28544 10444 28560
rect 10460 28544 10476 28560
rect 10492 28544 10508 28560
rect 10524 28544 10540 28560
rect 10556 28544 10572 28560
rect 10588 28544 10604 28560
rect 10620 28544 10636 28560
rect 10652 28544 10668 28560
rect 10684 28544 10700 28560
rect 10716 28544 10732 28560
rect 10748 28544 10764 28560
rect 10780 28544 10796 28560
rect 10812 28544 10828 28560
rect 10844 28544 10860 28560
rect 10876 28544 10892 28560
rect 10908 28544 10924 28560
rect 10940 28544 10956 28560
rect 10972 28544 10988 28560
rect 11004 28544 11020 28560
rect 11036 28544 11052 28560
rect 11068 28544 11084 28560
rect 11100 28544 11116 28560
rect 11132 28544 11148 28560
rect 11164 28544 11180 28560
rect 11196 28544 11212 28560
rect 11228 28544 11244 28560
rect 11260 28544 11276 28560
rect 11292 28544 11308 28560
rect 11324 28544 11340 28560
rect 11356 28544 11372 28560
rect 11388 28544 11404 28560
rect 11420 28544 11436 28560
rect 11452 28544 11468 28560
rect 11484 28544 11500 28560
rect 11516 28544 11532 28560
rect 11548 28544 11564 28560
rect 11580 28544 11596 28560
rect 11612 28544 11628 28560
rect 11644 28544 11660 28560
rect 11676 28544 11692 28560
rect 11708 28544 11724 28560
rect 11740 28544 27020 28560
rect 10041 28528 27020 28544
rect 10041 28512 10060 28528
rect 10076 28512 10092 28528
rect 10108 28512 10124 28528
rect 10140 28512 10156 28528
rect 10172 28512 10188 28528
rect 10204 28512 10220 28528
rect 10236 28512 10252 28528
rect 10268 28512 10284 28528
rect 10300 28512 10316 28528
rect 10332 28512 10348 28528
rect 10364 28512 10380 28528
rect 10396 28512 10412 28528
rect 10428 28512 10444 28528
rect 10460 28512 10476 28528
rect 10492 28512 10508 28528
rect 10524 28512 10540 28528
rect 10556 28512 10572 28528
rect 10588 28512 10604 28528
rect 10620 28512 10636 28528
rect 10652 28512 10668 28528
rect 10684 28512 10700 28528
rect 10716 28512 10732 28528
rect 10748 28512 10764 28528
rect 10780 28512 10796 28528
rect 10812 28512 10828 28528
rect 10844 28512 10860 28528
rect 10876 28512 10892 28528
rect 10908 28512 10924 28528
rect 10940 28512 10956 28528
rect 10972 28512 10988 28528
rect 11004 28512 11020 28528
rect 11036 28512 11052 28528
rect 11068 28512 11084 28528
rect 11100 28512 11116 28528
rect 11132 28512 11148 28528
rect 11164 28512 11180 28528
rect 11196 28512 11212 28528
rect 11228 28512 11244 28528
rect 11260 28512 11276 28528
rect 11292 28512 11308 28528
rect 11324 28512 11340 28528
rect 11356 28512 11372 28528
rect 11388 28512 11404 28528
rect 11420 28512 11436 28528
rect 11452 28512 11468 28528
rect 11484 28512 11500 28528
rect 11516 28512 11532 28528
rect 11548 28512 11564 28528
rect 11580 28512 11596 28528
rect 11612 28512 11628 28528
rect 11644 28512 11660 28528
rect 11676 28512 11692 28528
rect 11708 28512 11724 28528
rect 11740 28512 27020 28528
rect 10041 28501 27020 28512
rect 11760 28500 27020 28501
rect 9680 27699 10080 27700
rect 9241 27684 10080 27699
rect 9241 27668 9260 27684
rect 9276 27668 9292 27684
rect 9308 27668 9324 27684
rect 9340 27668 9356 27684
rect 9372 27668 9388 27684
rect 9404 27668 9420 27684
rect 9436 27668 9452 27684
rect 9468 27668 9484 27684
rect 9500 27668 9516 27684
rect 9532 27668 9548 27684
rect 9564 27668 9580 27684
rect 9596 27668 9612 27684
rect 9628 27668 9644 27684
rect 9660 27668 10080 27684
rect 9241 27652 10080 27668
rect 9241 27636 9260 27652
rect 9276 27636 9292 27652
rect 9308 27636 9324 27652
rect 9340 27636 9356 27652
rect 9372 27636 9388 27652
rect 9404 27636 9420 27652
rect 9436 27636 9452 27652
rect 9468 27636 9484 27652
rect 9500 27636 9516 27652
rect 9532 27636 9548 27652
rect 9564 27636 9580 27652
rect 9596 27636 9612 27652
rect 9628 27636 9644 27652
rect 9660 27636 10080 27652
rect 9241 27620 10080 27636
rect 9241 27604 9260 27620
rect 9276 27604 9292 27620
rect 9308 27604 9324 27620
rect 9340 27604 9356 27620
rect 9372 27604 9388 27620
rect 9404 27604 9420 27620
rect 9436 27604 9452 27620
rect 9468 27604 9484 27620
rect 9500 27604 9516 27620
rect 9532 27604 9548 27620
rect 9564 27604 9580 27620
rect 9596 27604 9612 27620
rect 9628 27604 9644 27620
rect 9660 27604 10080 27620
rect 9241 27588 10080 27604
rect 9241 27572 9260 27588
rect 9276 27572 9292 27588
rect 9308 27572 9324 27588
rect 9340 27572 9356 27588
rect 9372 27572 9388 27588
rect 9404 27572 9420 27588
rect 9436 27572 9452 27588
rect 9468 27572 9484 27588
rect 9500 27572 9516 27588
rect 9532 27572 9548 27588
rect 9564 27572 9580 27588
rect 9596 27572 9612 27588
rect 9628 27572 9644 27588
rect 9660 27572 10080 27588
rect 9241 27556 10080 27572
rect 9241 27540 9260 27556
rect 9276 27540 9292 27556
rect 9308 27540 9324 27556
rect 9340 27540 9356 27556
rect 9372 27540 9388 27556
rect 9404 27540 9420 27556
rect 9436 27540 9452 27556
rect 9468 27540 9484 27556
rect 9500 27540 9516 27556
rect 9532 27540 9548 27556
rect 9564 27540 9580 27556
rect 9596 27540 9612 27556
rect 9628 27540 9644 27556
rect 9660 27540 10080 27556
rect 9241 27524 10080 27540
rect 9241 27508 9260 27524
rect 9276 27508 9292 27524
rect 9308 27508 9324 27524
rect 9340 27508 9356 27524
rect 9372 27508 9388 27524
rect 9404 27508 9420 27524
rect 9436 27508 9452 27524
rect 9468 27508 9484 27524
rect 9500 27508 9516 27524
rect 9532 27508 9548 27524
rect 9564 27508 9580 27524
rect 9596 27508 9612 27524
rect 9628 27508 9644 27524
rect 9660 27508 10080 27524
rect 9241 27492 10080 27508
rect 9241 27476 9260 27492
rect 9276 27476 9292 27492
rect 9308 27476 9324 27492
rect 9340 27476 9356 27492
rect 9372 27476 9388 27492
rect 9404 27476 9420 27492
rect 9436 27476 9452 27492
rect 9468 27476 9484 27492
rect 9500 27476 9516 27492
rect 9532 27476 9548 27492
rect 9564 27476 9580 27492
rect 9596 27476 9612 27492
rect 9628 27476 9644 27492
rect 9660 27476 10080 27492
rect 9241 27460 10080 27476
rect 9241 27444 9260 27460
rect 9276 27444 9292 27460
rect 9308 27444 9324 27460
rect 9340 27444 9356 27460
rect 9372 27444 9388 27460
rect 9404 27444 9420 27460
rect 9436 27444 9452 27460
rect 9468 27444 9484 27460
rect 9500 27444 9516 27460
rect 9532 27444 9548 27460
rect 9564 27444 9580 27460
rect 9596 27444 9612 27460
rect 9628 27444 9644 27460
rect 9660 27444 10080 27460
rect 9241 27428 10080 27444
rect 9241 27412 9260 27428
rect 9276 27412 9292 27428
rect 9308 27412 9324 27428
rect 9340 27412 9356 27428
rect 9372 27412 9388 27428
rect 9404 27412 9420 27428
rect 9436 27412 9452 27428
rect 9468 27412 9484 27428
rect 9500 27412 9516 27428
rect 9532 27412 9548 27428
rect 9564 27412 9580 27428
rect 9596 27412 9612 27428
rect 9628 27412 9644 27428
rect 9660 27412 10080 27428
rect 9241 27396 10080 27412
rect 9241 27380 9260 27396
rect 9276 27380 9292 27396
rect 9308 27380 9324 27396
rect 9340 27380 9356 27396
rect 9372 27380 9388 27396
rect 9404 27380 9420 27396
rect 9436 27380 9452 27396
rect 9468 27380 9484 27396
rect 9500 27380 9516 27396
rect 9532 27380 9548 27396
rect 9564 27380 9580 27396
rect 9596 27380 9612 27396
rect 9628 27380 9644 27396
rect 9660 27380 10080 27396
rect 9241 27364 10080 27380
rect 9241 27348 9260 27364
rect 9276 27348 9292 27364
rect 9308 27348 9324 27364
rect 9340 27348 9356 27364
rect 9372 27348 9388 27364
rect 9404 27348 9420 27364
rect 9436 27348 9452 27364
rect 9468 27348 9484 27364
rect 9500 27348 9516 27364
rect 9532 27348 9548 27364
rect 9564 27348 9580 27364
rect 9596 27348 9612 27364
rect 9628 27348 9644 27364
rect 9660 27348 10080 27364
rect 9241 27332 10080 27348
rect 9241 27316 9260 27332
rect 9276 27316 9292 27332
rect 9308 27316 9324 27332
rect 9340 27316 9356 27332
rect 9372 27316 9388 27332
rect 9404 27316 9420 27332
rect 9436 27316 9452 27332
rect 9468 27316 9484 27332
rect 9500 27316 9516 27332
rect 9532 27316 9548 27332
rect 9564 27316 9580 27332
rect 9596 27316 9612 27332
rect 9628 27316 9644 27332
rect 9660 27316 10080 27332
rect 9241 27300 10080 27316
rect 9241 27284 9260 27300
rect 9276 27284 9292 27300
rect 9308 27284 9324 27300
rect 9340 27284 9356 27300
rect 9372 27284 9388 27300
rect 9404 27284 9420 27300
rect 9436 27284 9452 27300
rect 9468 27284 9484 27300
rect 9500 27284 9516 27300
rect 9532 27284 9548 27300
rect 9564 27284 9580 27300
rect 9596 27284 9612 27300
rect 9628 27284 9644 27300
rect 9660 27284 10080 27300
rect 9241 27268 10080 27284
rect 9241 27252 9260 27268
rect 9276 27252 9292 27268
rect 9308 27252 9324 27268
rect 9340 27252 9356 27268
rect 9372 27252 9388 27268
rect 9404 27252 9420 27268
rect 9436 27252 9452 27268
rect 9468 27252 9484 27268
rect 9500 27252 9516 27268
rect 9532 27252 9548 27268
rect 9564 27252 9580 27268
rect 9596 27252 9612 27268
rect 9628 27252 9644 27268
rect 9660 27252 10080 27268
rect 9241 27236 10080 27252
rect 9241 27220 9260 27236
rect 9276 27220 9292 27236
rect 9308 27220 9324 27236
rect 9340 27220 9356 27236
rect 9372 27220 9388 27236
rect 9404 27220 9420 27236
rect 9436 27220 9452 27236
rect 9468 27220 9484 27236
rect 9500 27220 9516 27236
rect 9532 27220 9548 27236
rect 9564 27220 9580 27236
rect 9596 27220 9612 27236
rect 9628 27220 9644 27236
rect 9660 27220 10080 27236
rect 9241 27204 10080 27220
rect 9241 27188 9260 27204
rect 9276 27188 9292 27204
rect 9308 27188 9324 27204
rect 9340 27188 9356 27204
rect 9372 27188 9388 27204
rect 9404 27188 9420 27204
rect 9436 27188 9452 27204
rect 9468 27188 9484 27204
rect 9500 27188 9516 27204
rect 9532 27188 9548 27204
rect 9564 27188 9580 27204
rect 9596 27188 9612 27204
rect 9628 27188 9644 27204
rect 9660 27188 10080 27204
rect 9241 27172 10080 27188
rect 9241 27156 9260 27172
rect 9276 27156 9292 27172
rect 9308 27156 9324 27172
rect 9340 27156 9356 27172
rect 9372 27156 9388 27172
rect 9404 27156 9420 27172
rect 9436 27156 9452 27172
rect 9468 27156 9484 27172
rect 9500 27156 9516 27172
rect 9532 27156 9548 27172
rect 9564 27156 9580 27172
rect 9596 27156 9612 27172
rect 9628 27156 9644 27172
rect 9660 27156 10080 27172
rect 9241 27140 10080 27156
rect 9241 27124 9260 27140
rect 9276 27124 9292 27140
rect 9308 27124 9324 27140
rect 9340 27124 9356 27140
rect 9372 27124 9388 27140
rect 9404 27124 9420 27140
rect 9436 27124 9452 27140
rect 9468 27124 9484 27140
rect 9500 27124 9516 27140
rect 9532 27124 9548 27140
rect 9564 27124 9580 27140
rect 9596 27124 9612 27140
rect 9628 27124 9644 27140
rect 9660 27124 10080 27140
rect 9241 27108 10080 27124
rect 9241 27092 9260 27108
rect 9276 27092 9292 27108
rect 9308 27092 9324 27108
rect 9340 27092 9356 27108
rect 9372 27092 9388 27108
rect 9404 27092 9420 27108
rect 9436 27092 9452 27108
rect 9468 27092 9484 27108
rect 9500 27092 9516 27108
rect 9532 27092 9548 27108
rect 9564 27092 9580 27108
rect 9596 27092 9612 27108
rect 9628 27092 9644 27108
rect 9660 27092 10080 27108
rect 9241 27076 10080 27092
rect 9241 27060 9260 27076
rect 9276 27060 9292 27076
rect 9308 27060 9324 27076
rect 9340 27060 9356 27076
rect 9372 27060 9388 27076
rect 9404 27060 9420 27076
rect 9436 27060 9452 27076
rect 9468 27060 9484 27076
rect 9500 27060 9516 27076
rect 9532 27060 9548 27076
rect 9564 27060 9580 27076
rect 9596 27060 9612 27076
rect 9628 27060 9644 27076
rect 9660 27060 10080 27076
rect 9241 27044 10080 27060
rect 9241 27028 9260 27044
rect 9276 27028 9292 27044
rect 9308 27028 9324 27044
rect 9340 27028 9356 27044
rect 9372 27028 9388 27044
rect 9404 27028 9420 27044
rect 9436 27028 9452 27044
rect 9468 27028 9484 27044
rect 9500 27028 9516 27044
rect 9532 27028 9548 27044
rect 9564 27028 9580 27044
rect 9596 27028 9612 27044
rect 9628 27028 9644 27044
rect 9660 27028 10080 27044
rect 9241 27012 10080 27028
rect 9241 26996 9260 27012
rect 9276 26996 9292 27012
rect 9308 26996 9324 27012
rect 9340 26996 9356 27012
rect 9372 26996 9388 27012
rect 9404 26996 9420 27012
rect 9436 26996 9452 27012
rect 9468 26996 9484 27012
rect 9500 26996 9516 27012
rect 9532 26996 9548 27012
rect 9564 26996 9580 27012
rect 9596 26996 9612 27012
rect 9628 26996 9644 27012
rect 9660 26996 10080 27012
rect 9241 26980 10080 26996
rect 9241 26964 9260 26980
rect 9276 26964 9292 26980
rect 9308 26964 9324 26980
rect 9340 26964 9356 26980
rect 9372 26964 9388 26980
rect 9404 26964 9420 26980
rect 9436 26964 9452 26980
rect 9468 26964 9484 26980
rect 9500 26964 9516 26980
rect 9532 26964 9548 26980
rect 9564 26964 9580 26980
rect 9596 26964 9612 26980
rect 9628 26964 9644 26980
rect 9660 26964 10080 26980
rect 9241 26948 10080 26964
rect 9241 26932 9260 26948
rect 9276 26932 9292 26948
rect 9308 26932 9324 26948
rect 9340 26932 9356 26948
rect 9372 26932 9388 26948
rect 9404 26932 9420 26948
rect 9436 26932 9452 26948
rect 9468 26932 9484 26948
rect 9500 26932 9516 26948
rect 9532 26932 9548 26948
rect 9564 26932 9580 26948
rect 9596 26932 9612 26948
rect 9628 26932 9644 26948
rect 9660 26932 10080 26948
rect 9241 26916 10080 26932
rect 9241 26900 9260 26916
rect 9276 26900 9292 26916
rect 9308 26900 9324 26916
rect 9340 26900 9356 26916
rect 9372 26900 9388 26916
rect 9404 26900 9420 26916
rect 9436 26900 9452 26916
rect 9468 26900 9484 26916
rect 9500 26900 9516 26916
rect 9532 26900 9548 26916
rect 9564 26900 9580 26916
rect 9596 26900 9612 26916
rect 9628 26900 9644 26916
rect 9660 26900 10080 26916
rect 9241 26884 10080 26900
rect 9241 26868 9260 26884
rect 9276 26868 9292 26884
rect 9308 26868 9324 26884
rect 9340 26868 9356 26884
rect 9372 26868 9388 26884
rect 9404 26868 9420 26884
rect 9436 26868 9452 26884
rect 9468 26868 9484 26884
rect 9500 26868 9516 26884
rect 9532 26868 9548 26884
rect 9564 26868 9580 26884
rect 9596 26868 9612 26884
rect 9628 26868 9644 26884
rect 9660 26868 10080 26884
rect 9241 26852 10080 26868
rect 9241 26836 9260 26852
rect 9276 26836 9292 26852
rect 9308 26836 9324 26852
rect 9340 26836 9356 26852
rect 9372 26836 9388 26852
rect 9404 26836 9420 26852
rect 9436 26836 9452 26852
rect 9468 26836 9484 26852
rect 9500 26836 9516 26852
rect 9532 26836 9548 26852
rect 9564 26836 9580 26852
rect 9596 26836 9612 26852
rect 9628 26836 9644 26852
rect 9660 26836 10080 26852
rect 9241 26820 10080 26836
rect 9241 26804 9260 26820
rect 9276 26804 9292 26820
rect 9308 26804 9324 26820
rect 9340 26804 9356 26820
rect 9372 26804 9388 26820
rect 9404 26804 9420 26820
rect 9436 26804 9452 26820
rect 9468 26804 9484 26820
rect 9500 26804 9516 26820
rect 9532 26804 9548 26820
rect 9564 26804 9580 26820
rect 9596 26804 9612 26820
rect 9628 26804 9644 26820
rect 9660 26804 10080 26820
rect 9241 26788 10080 26804
rect 9241 26772 9260 26788
rect 9276 26772 9292 26788
rect 9308 26772 9324 26788
rect 9340 26772 9356 26788
rect 9372 26772 9388 26788
rect 9404 26772 9420 26788
rect 9436 26772 9452 26788
rect 9468 26772 9484 26788
rect 9500 26772 9516 26788
rect 9532 26772 9548 26788
rect 9564 26772 9580 26788
rect 9596 26772 9612 26788
rect 9628 26772 9644 26788
rect 9660 26772 10080 26788
rect 9241 26756 10080 26772
rect 9241 26740 9260 26756
rect 9276 26740 9292 26756
rect 9308 26740 9324 26756
rect 9340 26740 9356 26756
rect 9372 26740 9388 26756
rect 9404 26740 9420 26756
rect 9436 26740 9452 26756
rect 9468 26740 9484 26756
rect 9500 26740 9516 26756
rect 9532 26740 9548 26756
rect 9564 26740 9580 26756
rect 9596 26740 9612 26756
rect 9628 26740 9644 26756
rect 9660 26740 10080 26756
rect 9241 26724 10080 26740
rect 9241 26708 9260 26724
rect 9276 26708 9292 26724
rect 9308 26708 9324 26724
rect 9340 26708 9356 26724
rect 9372 26708 9388 26724
rect 9404 26708 9420 26724
rect 9436 26708 9452 26724
rect 9468 26708 9484 26724
rect 9500 26708 9516 26724
rect 9532 26708 9548 26724
rect 9564 26708 9580 26724
rect 9596 26708 9612 26724
rect 9628 26708 9644 26724
rect 9660 26708 10080 26724
rect 9241 26692 10080 26708
rect 9241 26676 9260 26692
rect 9276 26676 9292 26692
rect 9308 26676 9324 26692
rect 9340 26676 9356 26692
rect 9372 26676 9388 26692
rect 9404 26676 9420 26692
rect 9436 26676 9452 26692
rect 9468 26676 9484 26692
rect 9500 26676 9516 26692
rect 9532 26676 9548 26692
rect 9564 26676 9580 26692
rect 9596 26676 9612 26692
rect 9628 26676 9644 26692
rect 9660 26676 10080 26692
rect 9241 26660 10080 26676
rect 9241 26644 9260 26660
rect 9276 26644 9292 26660
rect 9308 26644 9324 26660
rect 9340 26644 9356 26660
rect 9372 26644 9388 26660
rect 9404 26644 9420 26660
rect 9436 26644 9452 26660
rect 9468 26644 9484 26660
rect 9500 26644 9516 26660
rect 9532 26644 9548 26660
rect 9564 26644 9580 26660
rect 9596 26644 9612 26660
rect 9628 26644 9644 26660
rect 9660 26644 10080 26660
rect 9241 26628 10080 26644
rect 9241 26612 9260 26628
rect 9276 26612 9292 26628
rect 9308 26612 9324 26628
rect 9340 26612 9356 26628
rect 9372 26612 9388 26628
rect 9404 26612 9420 26628
rect 9436 26612 9452 26628
rect 9468 26612 9484 26628
rect 9500 26612 9516 26628
rect 9532 26612 9548 26628
rect 9564 26612 9580 26628
rect 9596 26612 9612 26628
rect 9628 26612 9644 26628
rect 9660 26612 10080 26628
rect 9241 26596 10080 26612
rect 9241 26580 9260 26596
rect 9276 26580 9292 26596
rect 9308 26580 9324 26596
rect 9340 26580 9356 26596
rect 9372 26580 9388 26596
rect 9404 26580 9420 26596
rect 9436 26580 9452 26596
rect 9468 26580 9484 26596
rect 9500 26580 9516 26596
rect 9532 26580 9548 26596
rect 9564 26580 9580 26596
rect 9596 26580 9612 26596
rect 9628 26580 9644 26596
rect 9660 26580 10080 26596
rect 9241 26564 10080 26580
rect 9241 26548 9260 26564
rect 9276 26548 9292 26564
rect 9308 26548 9324 26564
rect 9340 26548 9356 26564
rect 9372 26548 9388 26564
rect 9404 26548 9420 26564
rect 9436 26548 9452 26564
rect 9468 26548 9484 26564
rect 9500 26548 9516 26564
rect 9532 26548 9548 26564
rect 9564 26548 9580 26564
rect 9596 26548 9612 26564
rect 9628 26548 9644 26564
rect 9660 26548 10080 26564
rect 9241 26532 10080 26548
rect 9241 26516 9260 26532
rect 9276 26516 9292 26532
rect 9308 26516 9324 26532
rect 9340 26516 9356 26532
rect 9372 26516 9388 26532
rect 9404 26516 9420 26532
rect 9436 26516 9452 26532
rect 9468 26516 9484 26532
rect 9500 26516 9516 26532
rect 9532 26516 9548 26532
rect 9564 26516 9580 26532
rect 9596 26516 9612 26532
rect 9628 26516 9644 26532
rect 9660 26516 10080 26532
rect 9241 26501 10080 26516
rect 9680 26240 10080 26501
rect 9680 25880 11240 26240
rect 26660 26180 27020 28500
<< m2contact >>
rect 10060 28992 10076 29008
rect 10092 28992 10108 29008
rect 10124 28992 10140 29008
rect 10156 28992 10172 29008
rect 10188 28992 10204 29008
rect 10220 28992 10236 29008
rect 10252 28992 10268 29008
rect 10284 28992 10300 29008
rect 10316 28992 10332 29008
rect 10348 28992 10364 29008
rect 10380 28992 10396 29008
rect 10412 28992 10428 29008
rect 10444 28992 10460 29008
rect 10476 28992 10492 29008
rect 10508 28992 10524 29008
rect 10540 28992 10556 29008
rect 10572 28992 10588 29008
rect 10604 28992 10620 29008
rect 10636 28992 10652 29008
rect 10668 28992 10684 29008
rect 10700 28992 10716 29008
rect 10732 28992 10748 29008
rect 10764 28992 10780 29008
rect 10796 28992 10812 29008
rect 10828 28992 10844 29008
rect 10860 28992 10876 29008
rect 10892 28992 10908 29008
rect 10924 28992 10940 29008
rect 10956 28992 10972 29008
rect 10988 28992 11004 29008
rect 11020 28992 11036 29008
rect 11052 28992 11068 29008
rect 11084 28992 11100 29008
rect 11116 28992 11132 29008
rect 11148 28992 11164 29008
rect 11180 28992 11196 29008
rect 11212 28992 11228 29008
rect 11244 28992 11260 29008
rect 11276 28992 11292 29008
rect 11308 28992 11324 29008
rect 11340 28992 11356 29008
rect 11372 28992 11388 29008
rect 11404 28992 11420 29008
rect 11436 28992 11452 29008
rect 11468 28992 11484 29008
rect 11500 28992 11516 29008
rect 11532 28992 11548 29008
rect 11564 28992 11580 29008
rect 11596 28992 11612 29008
rect 11628 28992 11644 29008
rect 11660 28992 11676 29008
rect 11692 28992 11708 29008
rect 11724 28992 11740 29008
rect 10060 28960 10076 28976
rect 10092 28960 10108 28976
rect 10124 28960 10140 28976
rect 10156 28960 10172 28976
rect 10188 28960 10204 28976
rect 10220 28960 10236 28976
rect 10252 28960 10268 28976
rect 10284 28960 10300 28976
rect 10316 28960 10332 28976
rect 10348 28960 10364 28976
rect 10380 28960 10396 28976
rect 10412 28960 10428 28976
rect 10444 28960 10460 28976
rect 10476 28960 10492 28976
rect 10508 28960 10524 28976
rect 10540 28960 10556 28976
rect 10572 28960 10588 28976
rect 10604 28960 10620 28976
rect 10636 28960 10652 28976
rect 10668 28960 10684 28976
rect 10700 28960 10716 28976
rect 10732 28960 10748 28976
rect 10764 28960 10780 28976
rect 10796 28960 10812 28976
rect 10828 28960 10844 28976
rect 10860 28960 10876 28976
rect 10892 28960 10908 28976
rect 10924 28960 10940 28976
rect 10956 28960 10972 28976
rect 10988 28960 11004 28976
rect 11020 28960 11036 28976
rect 11052 28960 11068 28976
rect 11084 28960 11100 28976
rect 11116 28960 11132 28976
rect 11148 28960 11164 28976
rect 11180 28960 11196 28976
rect 11212 28960 11228 28976
rect 11244 28960 11260 28976
rect 11276 28960 11292 28976
rect 11308 28960 11324 28976
rect 11340 28960 11356 28976
rect 11372 28960 11388 28976
rect 11404 28960 11420 28976
rect 11436 28960 11452 28976
rect 11468 28960 11484 28976
rect 11500 28960 11516 28976
rect 11532 28960 11548 28976
rect 11564 28960 11580 28976
rect 11596 28960 11612 28976
rect 11628 28960 11644 28976
rect 11660 28960 11676 28976
rect 11692 28960 11708 28976
rect 11724 28960 11740 28976
rect 10060 28928 10076 28944
rect 10092 28928 10108 28944
rect 10124 28928 10140 28944
rect 10156 28928 10172 28944
rect 10188 28928 10204 28944
rect 10220 28928 10236 28944
rect 10252 28928 10268 28944
rect 10284 28928 10300 28944
rect 10316 28928 10332 28944
rect 10348 28928 10364 28944
rect 10380 28928 10396 28944
rect 10412 28928 10428 28944
rect 10444 28928 10460 28944
rect 10476 28928 10492 28944
rect 10508 28928 10524 28944
rect 10540 28928 10556 28944
rect 10572 28928 10588 28944
rect 10604 28928 10620 28944
rect 10636 28928 10652 28944
rect 10668 28928 10684 28944
rect 10700 28928 10716 28944
rect 10732 28928 10748 28944
rect 10764 28928 10780 28944
rect 10796 28928 10812 28944
rect 10828 28928 10844 28944
rect 10860 28928 10876 28944
rect 10892 28928 10908 28944
rect 10924 28928 10940 28944
rect 10956 28928 10972 28944
rect 10988 28928 11004 28944
rect 11020 28928 11036 28944
rect 11052 28928 11068 28944
rect 11084 28928 11100 28944
rect 11116 28928 11132 28944
rect 11148 28928 11164 28944
rect 11180 28928 11196 28944
rect 11212 28928 11228 28944
rect 11244 28928 11260 28944
rect 11276 28928 11292 28944
rect 11308 28928 11324 28944
rect 11340 28928 11356 28944
rect 11372 28928 11388 28944
rect 11404 28928 11420 28944
rect 11436 28928 11452 28944
rect 11468 28928 11484 28944
rect 11500 28928 11516 28944
rect 11532 28928 11548 28944
rect 11564 28928 11580 28944
rect 11596 28928 11612 28944
rect 11628 28928 11644 28944
rect 11660 28928 11676 28944
rect 11692 28928 11708 28944
rect 11724 28928 11740 28944
rect 10060 28896 10076 28912
rect 10092 28896 10108 28912
rect 10124 28896 10140 28912
rect 10156 28896 10172 28912
rect 10188 28896 10204 28912
rect 10220 28896 10236 28912
rect 10252 28896 10268 28912
rect 10284 28896 10300 28912
rect 10316 28896 10332 28912
rect 10348 28896 10364 28912
rect 10380 28896 10396 28912
rect 10412 28896 10428 28912
rect 10444 28896 10460 28912
rect 10476 28896 10492 28912
rect 10508 28896 10524 28912
rect 10540 28896 10556 28912
rect 10572 28896 10588 28912
rect 10604 28896 10620 28912
rect 10636 28896 10652 28912
rect 10668 28896 10684 28912
rect 10700 28896 10716 28912
rect 10732 28896 10748 28912
rect 10764 28896 10780 28912
rect 10796 28896 10812 28912
rect 10828 28896 10844 28912
rect 10860 28896 10876 28912
rect 10892 28896 10908 28912
rect 10924 28896 10940 28912
rect 10956 28896 10972 28912
rect 10988 28896 11004 28912
rect 11020 28896 11036 28912
rect 11052 28896 11068 28912
rect 11084 28896 11100 28912
rect 11116 28896 11132 28912
rect 11148 28896 11164 28912
rect 11180 28896 11196 28912
rect 11212 28896 11228 28912
rect 11244 28896 11260 28912
rect 11276 28896 11292 28912
rect 11308 28896 11324 28912
rect 11340 28896 11356 28912
rect 11372 28896 11388 28912
rect 11404 28896 11420 28912
rect 11436 28896 11452 28912
rect 11468 28896 11484 28912
rect 11500 28896 11516 28912
rect 11532 28896 11548 28912
rect 11564 28896 11580 28912
rect 11596 28896 11612 28912
rect 11628 28896 11644 28912
rect 11660 28896 11676 28912
rect 11692 28896 11708 28912
rect 11724 28896 11740 28912
rect 10060 28864 10076 28880
rect 10092 28864 10108 28880
rect 10124 28864 10140 28880
rect 10156 28864 10172 28880
rect 10188 28864 10204 28880
rect 10220 28864 10236 28880
rect 10252 28864 10268 28880
rect 10284 28864 10300 28880
rect 10316 28864 10332 28880
rect 10348 28864 10364 28880
rect 10380 28864 10396 28880
rect 10412 28864 10428 28880
rect 10444 28864 10460 28880
rect 10476 28864 10492 28880
rect 10508 28864 10524 28880
rect 10540 28864 10556 28880
rect 10572 28864 10588 28880
rect 10604 28864 10620 28880
rect 10636 28864 10652 28880
rect 10668 28864 10684 28880
rect 10700 28864 10716 28880
rect 10732 28864 10748 28880
rect 10764 28864 10780 28880
rect 10796 28864 10812 28880
rect 10828 28864 10844 28880
rect 10860 28864 10876 28880
rect 10892 28864 10908 28880
rect 10924 28864 10940 28880
rect 10956 28864 10972 28880
rect 10988 28864 11004 28880
rect 11020 28864 11036 28880
rect 11052 28864 11068 28880
rect 11084 28864 11100 28880
rect 11116 28864 11132 28880
rect 11148 28864 11164 28880
rect 11180 28864 11196 28880
rect 11212 28864 11228 28880
rect 11244 28864 11260 28880
rect 11276 28864 11292 28880
rect 11308 28864 11324 28880
rect 11340 28864 11356 28880
rect 11372 28864 11388 28880
rect 11404 28864 11420 28880
rect 11436 28864 11452 28880
rect 11468 28864 11484 28880
rect 11500 28864 11516 28880
rect 11532 28864 11548 28880
rect 11564 28864 11580 28880
rect 11596 28864 11612 28880
rect 11628 28864 11644 28880
rect 11660 28864 11676 28880
rect 11692 28864 11708 28880
rect 11724 28864 11740 28880
rect 10060 28832 10076 28848
rect 10092 28832 10108 28848
rect 10124 28832 10140 28848
rect 10156 28832 10172 28848
rect 10188 28832 10204 28848
rect 10220 28832 10236 28848
rect 10252 28832 10268 28848
rect 10284 28832 10300 28848
rect 10316 28832 10332 28848
rect 10348 28832 10364 28848
rect 10380 28832 10396 28848
rect 10412 28832 10428 28848
rect 10444 28832 10460 28848
rect 10476 28832 10492 28848
rect 10508 28832 10524 28848
rect 10540 28832 10556 28848
rect 10572 28832 10588 28848
rect 10604 28832 10620 28848
rect 10636 28832 10652 28848
rect 10668 28832 10684 28848
rect 10700 28832 10716 28848
rect 10732 28832 10748 28848
rect 10764 28832 10780 28848
rect 10796 28832 10812 28848
rect 10828 28832 10844 28848
rect 10860 28832 10876 28848
rect 10892 28832 10908 28848
rect 10924 28832 10940 28848
rect 10956 28832 10972 28848
rect 10988 28832 11004 28848
rect 11020 28832 11036 28848
rect 11052 28832 11068 28848
rect 11084 28832 11100 28848
rect 11116 28832 11132 28848
rect 11148 28832 11164 28848
rect 11180 28832 11196 28848
rect 11212 28832 11228 28848
rect 11244 28832 11260 28848
rect 11276 28832 11292 28848
rect 11308 28832 11324 28848
rect 11340 28832 11356 28848
rect 11372 28832 11388 28848
rect 11404 28832 11420 28848
rect 11436 28832 11452 28848
rect 11468 28832 11484 28848
rect 11500 28832 11516 28848
rect 11532 28832 11548 28848
rect 11564 28832 11580 28848
rect 11596 28832 11612 28848
rect 11628 28832 11644 28848
rect 11660 28832 11676 28848
rect 11692 28832 11708 28848
rect 11724 28832 11740 28848
rect 10060 28800 10076 28816
rect 10092 28800 10108 28816
rect 10124 28800 10140 28816
rect 10156 28800 10172 28816
rect 10188 28800 10204 28816
rect 10220 28800 10236 28816
rect 10252 28800 10268 28816
rect 10284 28800 10300 28816
rect 10316 28800 10332 28816
rect 10348 28800 10364 28816
rect 10380 28800 10396 28816
rect 10412 28800 10428 28816
rect 10444 28800 10460 28816
rect 10476 28800 10492 28816
rect 10508 28800 10524 28816
rect 10540 28800 10556 28816
rect 10572 28800 10588 28816
rect 10604 28800 10620 28816
rect 10636 28800 10652 28816
rect 10668 28800 10684 28816
rect 10700 28800 10716 28816
rect 10732 28800 10748 28816
rect 10764 28800 10780 28816
rect 10796 28800 10812 28816
rect 10828 28800 10844 28816
rect 10860 28800 10876 28816
rect 10892 28800 10908 28816
rect 10924 28800 10940 28816
rect 10956 28800 10972 28816
rect 10988 28800 11004 28816
rect 11020 28800 11036 28816
rect 11052 28800 11068 28816
rect 11084 28800 11100 28816
rect 11116 28800 11132 28816
rect 11148 28800 11164 28816
rect 11180 28800 11196 28816
rect 11212 28800 11228 28816
rect 11244 28800 11260 28816
rect 11276 28800 11292 28816
rect 11308 28800 11324 28816
rect 11340 28800 11356 28816
rect 11372 28800 11388 28816
rect 11404 28800 11420 28816
rect 11436 28800 11452 28816
rect 11468 28800 11484 28816
rect 11500 28800 11516 28816
rect 11532 28800 11548 28816
rect 11564 28800 11580 28816
rect 11596 28800 11612 28816
rect 11628 28800 11644 28816
rect 11660 28800 11676 28816
rect 11692 28800 11708 28816
rect 11724 28800 11740 28816
rect 10060 28768 10076 28784
rect 10092 28768 10108 28784
rect 10124 28768 10140 28784
rect 10156 28768 10172 28784
rect 10188 28768 10204 28784
rect 10220 28768 10236 28784
rect 10252 28768 10268 28784
rect 10284 28768 10300 28784
rect 10316 28768 10332 28784
rect 10348 28768 10364 28784
rect 10380 28768 10396 28784
rect 10412 28768 10428 28784
rect 10444 28768 10460 28784
rect 10476 28768 10492 28784
rect 10508 28768 10524 28784
rect 10540 28768 10556 28784
rect 10572 28768 10588 28784
rect 10604 28768 10620 28784
rect 10636 28768 10652 28784
rect 10668 28768 10684 28784
rect 10700 28768 10716 28784
rect 10732 28768 10748 28784
rect 10764 28768 10780 28784
rect 10796 28768 10812 28784
rect 10828 28768 10844 28784
rect 10860 28768 10876 28784
rect 10892 28768 10908 28784
rect 10924 28768 10940 28784
rect 10956 28768 10972 28784
rect 10988 28768 11004 28784
rect 11020 28768 11036 28784
rect 11052 28768 11068 28784
rect 11084 28768 11100 28784
rect 11116 28768 11132 28784
rect 11148 28768 11164 28784
rect 11180 28768 11196 28784
rect 11212 28768 11228 28784
rect 11244 28768 11260 28784
rect 11276 28768 11292 28784
rect 11308 28768 11324 28784
rect 11340 28768 11356 28784
rect 11372 28768 11388 28784
rect 11404 28768 11420 28784
rect 11436 28768 11452 28784
rect 11468 28768 11484 28784
rect 11500 28768 11516 28784
rect 11532 28768 11548 28784
rect 11564 28768 11580 28784
rect 11596 28768 11612 28784
rect 11628 28768 11644 28784
rect 11660 28768 11676 28784
rect 11692 28768 11708 28784
rect 11724 28768 11740 28784
rect 10060 28736 10076 28752
rect 10092 28736 10108 28752
rect 10124 28736 10140 28752
rect 10156 28736 10172 28752
rect 10188 28736 10204 28752
rect 10220 28736 10236 28752
rect 10252 28736 10268 28752
rect 10284 28736 10300 28752
rect 10316 28736 10332 28752
rect 10348 28736 10364 28752
rect 10380 28736 10396 28752
rect 10412 28736 10428 28752
rect 10444 28736 10460 28752
rect 10476 28736 10492 28752
rect 10508 28736 10524 28752
rect 10540 28736 10556 28752
rect 10572 28736 10588 28752
rect 10604 28736 10620 28752
rect 10636 28736 10652 28752
rect 10668 28736 10684 28752
rect 10700 28736 10716 28752
rect 10732 28736 10748 28752
rect 10764 28736 10780 28752
rect 10796 28736 10812 28752
rect 10828 28736 10844 28752
rect 10860 28736 10876 28752
rect 10892 28736 10908 28752
rect 10924 28736 10940 28752
rect 10956 28736 10972 28752
rect 10988 28736 11004 28752
rect 11020 28736 11036 28752
rect 11052 28736 11068 28752
rect 11084 28736 11100 28752
rect 11116 28736 11132 28752
rect 11148 28736 11164 28752
rect 11180 28736 11196 28752
rect 11212 28736 11228 28752
rect 11244 28736 11260 28752
rect 11276 28736 11292 28752
rect 11308 28736 11324 28752
rect 11340 28736 11356 28752
rect 11372 28736 11388 28752
rect 11404 28736 11420 28752
rect 11436 28736 11452 28752
rect 11468 28736 11484 28752
rect 11500 28736 11516 28752
rect 11532 28736 11548 28752
rect 11564 28736 11580 28752
rect 11596 28736 11612 28752
rect 11628 28736 11644 28752
rect 11660 28736 11676 28752
rect 11692 28736 11708 28752
rect 11724 28736 11740 28752
rect 10060 28704 10076 28720
rect 10092 28704 10108 28720
rect 10124 28704 10140 28720
rect 10156 28704 10172 28720
rect 10188 28704 10204 28720
rect 10220 28704 10236 28720
rect 10252 28704 10268 28720
rect 10284 28704 10300 28720
rect 10316 28704 10332 28720
rect 10348 28704 10364 28720
rect 10380 28704 10396 28720
rect 10412 28704 10428 28720
rect 10444 28704 10460 28720
rect 10476 28704 10492 28720
rect 10508 28704 10524 28720
rect 10540 28704 10556 28720
rect 10572 28704 10588 28720
rect 10604 28704 10620 28720
rect 10636 28704 10652 28720
rect 10668 28704 10684 28720
rect 10700 28704 10716 28720
rect 10732 28704 10748 28720
rect 10764 28704 10780 28720
rect 10796 28704 10812 28720
rect 10828 28704 10844 28720
rect 10860 28704 10876 28720
rect 10892 28704 10908 28720
rect 10924 28704 10940 28720
rect 10956 28704 10972 28720
rect 10988 28704 11004 28720
rect 11020 28704 11036 28720
rect 11052 28704 11068 28720
rect 11084 28704 11100 28720
rect 11116 28704 11132 28720
rect 11148 28704 11164 28720
rect 11180 28704 11196 28720
rect 11212 28704 11228 28720
rect 11244 28704 11260 28720
rect 11276 28704 11292 28720
rect 11308 28704 11324 28720
rect 11340 28704 11356 28720
rect 11372 28704 11388 28720
rect 11404 28704 11420 28720
rect 11436 28704 11452 28720
rect 11468 28704 11484 28720
rect 11500 28704 11516 28720
rect 11532 28704 11548 28720
rect 11564 28704 11580 28720
rect 11596 28704 11612 28720
rect 11628 28704 11644 28720
rect 11660 28704 11676 28720
rect 11692 28704 11708 28720
rect 11724 28704 11740 28720
rect 10060 28672 10076 28688
rect 10092 28672 10108 28688
rect 10124 28672 10140 28688
rect 10156 28672 10172 28688
rect 10188 28672 10204 28688
rect 10220 28672 10236 28688
rect 10252 28672 10268 28688
rect 10284 28672 10300 28688
rect 10316 28672 10332 28688
rect 10348 28672 10364 28688
rect 10380 28672 10396 28688
rect 10412 28672 10428 28688
rect 10444 28672 10460 28688
rect 10476 28672 10492 28688
rect 10508 28672 10524 28688
rect 10540 28672 10556 28688
rect 10572 28672 10588 28688
rect 10604 28672 10620 28688
rect 10636 28672 10652 28688
rect 10668 28672 10684 28688
rect 10700 28672 10716 28688
rect 10732 28672 10748 28688
rect 10764 28672 10780 28688
rect 10796 28672 10812 28688
rect 10828 28672 10844 28688
rect 10860 28672 10876 28688
rect 10892 28672 10908 28688
rect 10924 28672 10940 28688
rect 10956 28672 10972 28688
rect 10988 28672 11004 28688
rect 11020 28672 11036 28688
rect 11052 28672 11068 28688
rect 11084 28672 11100 28688
rect 11116 28672 11132 28688
rect 11148 28672 11164 28688
rect 11180 28672 11196 28688
rect 11212 28672 11228 28688
rect 11244 28672 11260 28688
rect 11276 28672 11292 28688
rect 11308 28672 11324 28688
rect 11340 28672 11356 28688
rect 11372 28672 11388 28688
rect 11404 28672 11420 28688
rect 11436 28672 11452 28688
rect 11468 28672 11484 28688
rect 11500 28672 11516 28688
rect 11532 28672 11548 28688
rect 11564 28672 11580 28688
rect 11596 28672 11612 28688
rect 11628 28672 11644 28688
rect 11660 28672 11676 28688
rect 11692 28672 11708 28688
rect 11724 28672 11740 28688
rect 10060 28640 10076 28656
rect 10092 28640 10108 28656
rect 10124 28640 10140 28656
rect 10156 28640 10172 28656
rect 10188 28640 10204 28656
rect 10220 28640 10236 28656
rect 10252 28640 10268 28656
rect 10284 28640 10300 28656
rect 10316 28640 10332 28656
rect 10348 28640 10364 28656
rect 10380 28640 10396 28656
rect 10412 28640 10428 28656
rect 10444 28640 10460 28656
rect 10476 28640 10492 28656
rect 10508 28640 10524 28656
rect 10540 28640 10556 28656
rect 10572 28640 10588 28656
rect 10604 28640 10620 28656
rect 10636 28640 10652 28656
rect 10668 28640 10684 28656
rect 10700 28640 10716 28656
rect 10732 28640 10748 28656
rect 10764 28640 10780 28656
rect 10796 28640 10812 28656
rect 10828 28640 10844 28656
rect 10860 28640 10876 28656
rect 10892 28640 10908 28656
rect 10924 28640 10940 28656
rect 10956 28640 10972 28656
rect 10988 28640 11004 28656
rect 11020 28640 11036 28656
rect 11052 28640 11068 28656
rect 11084 28640 11100 28656
rect 11116 28640 11132 28656
rect 11148 28640 11164 28656
rect 11180 28640 11196 28656
rect 11212 28640 11228 28656
rect 11244 28640 11260 28656
rect 11276 28640 11292 28656
rect 11308 28640 11324 28656
rect 11340 28640 11356 28656
rect 11372 28640 11388 28656
rect 11404 28640 11420 28656
rect 11436 28640 11452 28656
rect 11468 28640 11484 28656
rect 11500 28640 11516 28656
rect 11532 28640 11548 28656
rect 11564 28640 11580 28656
rect 11596 28640 11612 28656
rect 11628 28640 11644 28656
rect 11660 28640 11676 28656
rect 11692 28640 11708 28656
rect 11724 28640 11740 28656
rect 10060 28608 10076 28624
rect 10092 28608 10108 28624
rect 10124 28608 10140 28624
rect 10156 28608 10172 28624
rect 10188 28608 10204 28624
rect 10220 28608 10236 28624
rect 10252 28608 10268 28624
rect 10284 28608 10300 28624
rect 10316 28608 10332 28624
rect 10348 28608 10364 28624
rect 10380 28608 10396 28624
rect 10412 28608 10428 28624
rect 10444 28608 10460 28624
rect 10476 28608 10492 28624
rect 10508 28608 10524 28624
rect 10540 28608 10556 28624
rect 10572 28608 10588 28624
rect 10604 28608 10620 28624
rect 10636 28608 10652 28624
rect 10668 28608 10684 28624
rect 10700 28608 10716 28624
rect 10732 28608 10748 28624
rect 10764 28608 10780 28624
rect 10796 28608 10812 28624
rect 10828 28608 10844 28624
rect 10860 28608 10876 28624
rect 10892 28608 10908 28624
rect 10924 28608 10940 28624
rect 10956 28608 10972 28624
rect 10988 28608 11004 28624
rect 11020 28608 11036 28624
rect 11052 28608 11068 28624
rect 11084 28608 11100 28624
rect 11116 28608 11132 28624
rect 11148 28608 11164 28624
rect 11180 28608 11196 28624
rect 11212 28608 11228 28624
rect 11244 28608 11260 28624
rect 11276 28608 11292 28624
rect 11308 28608 11324 28624
rect 11340 28608 11356 28624
rect 11372 28608 11388 28624
rect 11404 28608 11420 28624
rect 11436 28608 11452 28624
rect 11468 28608 11484 28624
rect 11500 28608 11516 28624
rect 11532 28608 11548 28624
rect 11564 28608 11580 28624
rect 11596 28608 11612 28624
rect 11628 28608 11644 28624
rect 11660 28608 11676 28624
rect 11692 28608 11708 28624
rect 11724 28608 11740 28624
rect 10060 28576 10076 28592
rect 10092 28576 10108 28592
rect 10124 28576 10140 28592
rect 10156 28576 10172 28592
rect 10188 28576 10204 28592
rect 10220 28576 10236 28592
rect 10252 28576 10268 28592
rect 10284 28576 10300 28592
rect 10316 28576 10332 28592
rect 10348 28576 10364 28592
rect 10380 28576 10396 28592
rect 10412 28576 10428 28592
rect 10444 28576 10460 28592
rect 10476 28576 10492 28592
rect 10508 28576 10524 28592
rect 10540 28576 10556 28592
rect 10572 28576 10588 28592
rect 10604 28576 10620 28592
rect 10636 28576 10652 28592
rect 10668 28576 10684 28592
rect 10700 28576 10716 28592
rect 10732 28576 10748 28592
rect 10764 28576 10780 28592
rect 10796 28576 10812 28592
rect 10828 28576 10844 28592
rect 10860 28576 10876 28592
rect 10892 28576 10908 28592
rect 10924 28576 10940 28592
rect 10956 28576 10972 28592
rect 10988 28576 11004 28592
rect 11020 28576 11036 28592
rect 11052 28576 11068 28592
rect 11084 28576 11100 28592
rect 11116 28576 11132 28592
rect 11148 28576 11164 28592
rect 11180 28576 11196 28592
rect 11212 28576 11228 28592
rect 11244 28576 11260 28592
rect 11276 28576 11292 28592
rect 11308 28576 11324 28592
rect 11340 28576 11356 28592
rect 11372 28576 11388 28592
rect 11404 28576 11420 28592
rect 11436 28576 11452 28592
rect 11468 28576 11484 28592
rect 11500 28576 11516 28592
rect 11532 28576 11548 28592
rect 11564 28576 11580 28592
rect 11596 28576 11612 28592
rect 11628 28576 11644 28592
rect 11660 28576 11676 28592
rect 11692 28576 11708 28592
rect 11724 28576 11740 28592
rect 10060 28544 10076 28560
rect 10092 28544 10108 28560
rect 10124 28544 10140 28560
rect 10156 28544 10172 28560
rect 10188 28544 10204 28560
rect 10220 28544 10236 28560
rect 10252 28544 10268 28560
rect 10284 28544 10300 28560
rect 10316 28544 10332 28560
rect 10348 28544 10364 28560
rect 10380 28544 10396 28560
rect 10412 28544 10428 28560
rect 10444 28544 10460 28560
rect 10476 28544 10492 28560
rect 10508 28544 10524 28560
rect 10540 28544 10556 28560
rect 10572 28544 10588 28560
rect 10604 28544 10620 28560
rect 10636 28544 10652 28560
rect 10668 28544 10684 28560
rect 10700 28544 10716 28560
rect 10732 28544 10748 28560
rect 10764 28544 10780 28560
rect 10796 28544 10812 28560
rect 10828 28544 10844 28560
rect 10860 28544 10876 28560
rect 10892 28544 10908 28560
rect 10924 28544 10940 28560
rect 10956 28544 10972 28560
rect 10988 28544 11004 28560
rect 11020 28544 11036 28560
rect 11052 28544 11068 28560
rect 11084 28544 11100 28560
rect 11116 28544 11132 28560
rect 11148 28544 11164 28560
rect 11180 28544 11196 28560
rect 11212 28544 11228 28560
rect 11244 28544 11260 28560
rect 11276 28544 11292 28560
rect 11308 28544 11324 28560
rect 11340 28544 11356 28560
rect 11372 28544 11388 28560
rect 11404 28544 11420 28560
rect 11436 28544 11452 28560
rect 11468 28544 11484 28560
rect 11500 28544 11516 28560
rect 11532 28544 11548 28560
rect 11564 28544 11580 28560
rect 11596 28544 11612 28560
rect 11628 28544 11644 28560
rect 11660 28544 11676 28560
rect 11692 28544 11708 28560
rect 11724 28544 11740 28560
rect 10060 28512 10076 28528
rect 10092 28512 10108 28528
rect 10124 28512 10140 28528
rect 10156 28512 10172 28528
rect 10188 28512 10204 28528
rect 10220 28512 10236 28528
rect 10252 28512 10268 28528
rect 10284 28512 10300 28528
rect 10316 28512 10332 28528
rect 10348 28512 10364 28528
rect 10380 28512 10396 28528
rect 10412 28512 10428 28528
rect 10444 28512 10460 28528
rect 10476 28512 10492 28528
rect 10508 28512 10524 28528
rect 10540 28512 10556 28528
rect 10572 28512 10588 28528
rect 10604 28512 10620 28528
rect 10636 28512 10652 28528
rect 10668 28512 10684 28528
rect 10700 28512 10716 28528
rect 10732 28512 10748 28528
rect 10764 28512 10780 28528
rect 10796 28512 10812 28528
rect 10828 28512 10844 28528
rect 10860 28512 10876 28528
rect 10892 28512 10908 28528
rect 10924 28512 10940 28528
rect 10956 28512 10972 28528
rect 10988 28512 11004 28528
rect 11020 28512 11036 28528
rect 11052 28512 11068 28528
rect 11084 28512 11100 28528
rect 11116 28512 11132 28528
rect 11148 28512 11164 28528
rect 11180 28512 11196 28528
rect 11212 28512 11228 28528
rect 11244 28512 11260 28528
rect 11276 28512 11292 28528
rect 11308 28512 11324 28528
rect 11340 28512 11356 28528
rect 11372 28512 11388 28528
rect 11404 28512 11420 28528
rect 11436 28512 11452 28528
rect 11468 28512 11484 28528
rect 11500 28512 11516 28528
rect 11532 28512 11548 28528
rect 11564 28512 11580 28528
rect 11596 28512 11612 28528
rect 11628 28512 11644 28528
rect 11660 28512 11676 28528
rect 11692 28512 11708 28528
rect 11724 28512 11740 28528
rect 9260 27668 9276 27684
rect 9292 27668 9308 27684
rect 9324 27668 9340 27684
rect 9356 27668 9372 27684
rect 9388 27668 9404 27684
rect 9420 27668 9436 27684
rect 9452 27668 9468 27684
rect 9484 27668 9500 27684
rect 9516 27668 9532 27684
rect 9548 27668 9564 27684
rect 9580 27668 9596 27684
rect 9612 27668 9628 27684
rect 9644 27668 9660 27684
rect 9260 27636 9276 27652
rect 9292 27636 9308 27652
rect 9324 27636 9340 27652
rect 9356 27636 9372 27652
rect 9388 27636 9404 27652
rect 9420 27636 9436 27652
rect 9452 27636 9468 27652
rect 9484 27636 9500 27652
rect 9516 27636 9532 27652
rect 9548 27636 9564 27652
rect 9580 27636 9596 27652
rect 9612 27636 9628 27652
rect 9644 27636 9660 27652
rect 9260 27604 9276 27620
rect 9292 27604 9308 27620
rect 9324 27604 9340 27620
rect 9356 27604 9372 27620
rect 9388 27604 9404 27620
rect 9420 27604 9436 27620
rect 9452 27604 9468 27620
rect 9484 27604 9500 27620
rect 9516 27604 9532 27620
rect 9548 27604 9564 27620
rect 9580 27604 9596 27620
rect 9612 27604 9628 27620
rect 9644 27604 9660 27620
rect 9260 27572 9276 27588
rect 9292 27572 9308 27588
rect 9324 27572 9340 27588
rect 9356 27572 9372 27588
rect 9388 27572 9404 27588
rect 9420 27572 9436 27588
rect 9452 27572 9468 27588
rect 9484 27572 9500 27588
rect 9516 27572 9532 27588
rect 9548 27572 9564 27588
rect 9580 27572 9596 27588
rect 9612 27572 9628 27588
rect 9644 27572 9660 27588
rect 9260 27540 9276 27556
rect 9292 27540 9308 27556
rect 9324 27540 9340 27556
rect 9356 27540 9372 27556
rect 9388 27540 9404 27556
rect 9420 27540 9436 27556
rect 9452 27540 9468 27556
rect 9484 27540 9500 27556
rect 9516 27540 9532 27556
rect 9548 27540 9564 27556
rect 9580 27540 9596 27556
rect 9612 27540 9628 27556
rect 9644 27540 9660 27556
rect 9260 27508 9276 27524
rect 9292 27508 9308 27524
rect 9324 27508 9340 27524
rect 9356 27508 9372 27524
rect 9388 27508 9404 27524
rect 9420 27508 9436 27524
rect 9452 27508 9468 27524
rect 9484 27508 9500 27524
rect 9516 27508 9532 27524
rect 9548 27508 9564 27524
rect 9580 27508 9596 27524
rect 9612 27508 9628 27524
rect 9644 27508 9660 27524
rect 9260 27476 9276 27492
rect 9292 27476 9308 27492
rect 9324 27476 9340 27492
rect 9356 27476 9372 27492
rect 9388 27476 9404 27492
rect 9420 27476 9436 27492
rect 9452 27476 9468 27492
rect 9484 27476 9500 27492
rect 9516 27476 9532 27492
rect 9548 27476 9564 27492
rect 9580 27476 9596 27492
rect 9612 27476 9628 27492
rect 9644 27476 9660 27492
rect 9260 27444 9276 27460
rect 9292 27444 9308 27460
rect 9324 27444 9340 27460
rect 9356 27444 9372 27460
rect 9388 27444 9404 27460
rect 9420 27444 9436 27460
rect 9452 27444 9468 27460
rect 9484 27444 9500 27460
rect 9516 27444 9532 27460
rect 9548 27444 9564 27460
rect 9580 27444 9596 27460
rect 9612 27444 9628 27460
rect 9644 27444 9660 27460
rect 9260 27412 9276 27428
rect 9292 27412 9308 27428
rect 9324 27412 9340 27428
rect 9356 27412 9372 27428
rect 9388 27412 9404 27428
rect 9420 27412 9436 27428
rect 9452 27412 9468 27428
rect 9484 27412 9500 27428
rect 9516 27412 9532 27428
rect 9548 27412 9564 27428
rect 9580 27412 9596 27428
rect 9612 27412 9628 27428
rect 9644 27412 9660 27428
rect 9260 27380 9276 27396
rect 9292 27380 9308 27396
rect 9324 27380 9340 27396
rect 9356 27380 9372 27396
rect 9388 27380 9404 27396
rect 9420 27380 9436 27396
rect 9452 27380 9468 27396
rect 9484 27380 9500 27396
rect 9516 27380 9532 27396
rect 9548 27380 9564 27396
rect 9580 27380 9596 27396
rect 9612 27380 9628 27396
rect 9644 27380 9660 27396
rect 9260 27348 9276 27364
rect 9292 27348 9308 27364
rect 9324 27348 9340 27364
rect 9356 27348 9372 27364
rect 9388 27348 9404 27364
rect 9420 27348 9436 27364
rect 9452 27348 9468 27364
rect 9484 27348 9500 27364
rect 9516 27348 9532 27364
rect 9548 27348 9564 27364
rect 9580 27348 9596 27364
rect 9612 27348 9628 27364
rect 9644 27348 9660 27364
rect 9260 27316 9276 27332
rect 9292 27316 9308 27332
rect 9324 27316 9340 27332
rect 9356 27316 9372 27332
rect 9388 27316 9404 27332
rect 9420 27316 9436 27332
rect 9452 27316 9468 27332
rect 9484 27316 9500 27332
rect 9516 27316 9532 27332
rect 9548 27316 9564 27332
rect 9580 27316 9596 27332
rect 9612 27316 9628 27332
rect 9644 27316 9660 27332
rect 9260 27284 9276 27300
rect 9292 27284 9308 27300
rect 9324 27284 9340 27300
rect 9356 27284 9372 27300
rect 9388 27284 9404 27300
rect 9420 27284 9436 27300
rect 9452 27284 9468 27300
rect 9484 27284 9500 27300
rect 9516 27284 9532 27300
rect 9548 27284 9564 27300
rect 9580 27284 9596 27300
rect 9612 27284 9628 27300
rect 9644 27284 9660 27300
rect 9260 27252 9276 27268
rect 9292 27252 9308 27268
rect 9324 27252 9340 27268
rect 9356 27252 9372 27268
rect 9388 27252 9404 27268
rect 9420 27252 9436 27268
rect 9452 27252 9468 27268
rect 9484 27252 9500 27268
rect 9516 27252 9532 27268
rect 9548 27252 9564 27268
rect 9580 27252 9596 27268
rect 9612 27252 9628 27268
rect 9644 27252 9660 27268
rect 9260 27220 9276 27236
rect 9292 27220 9308 27236
rect 9324 27220 9340 27236
rect 9356 27220 9372 27236
rect 9388 27220 9404 27236
rect 9420 27220 9436 27236
rect 9452 27220 9468 27236
rect 9484 27220 9500 27236
rect 9516 27220 9532 27236
rect 9548 27220 9564 27236
rect 9580 27220 9596 27236
rect 9612 27220 9628 27236
rect 9644 27220 9660 27236
rect 9260 27188 9276 27204
rect 9292 27188 9308 27204
rect 9324 27188 9340 27204
rect 9356 27188 9372 27204
rect 9388 27188 9404 27204
rect 9420 27188 9436 27204
rect 9452 27188 9468 27204
rect 9484 27188 9500 27204
rect 9516 27188 9532 27204
rect 9548 27188 9564 27204
rect 9580 27188 9596 27204
rect 9612 27188 9628 27204
rect 9644 27188 9660 27204
rect 9260 27156 9276 27172
rect 9292 27156 9308 27172
rect 9324 27156 9340 27172
rect 9356 27156 9372 27172
rect 9388 27156 9404 27172
rect 9420 27156 9436 27172
rect 9452 27156 9468 27172
rect 9484 27156 9500 27172
rect 9516 27156 9532 27172
rect 9548 27156 9564 27172
rect 9580 27156 9596 27172
rect 9612 27156 9628 27172
rect 9644 27156 9660 27172
rect 9260 27124 9276 27140
rect 9292 27124 9308 27140
rect 9324 27124 9340 27140
rect 9356 27124 9372 27140
rect 9388 27124 9404 27140
rect 9420 27124 9436 27140
rect 9452 27124 9468 27140
rect 9484 27124 9500 27140
rect 9516 27124 9532 27140
rect 9548 27124 9564 27140
rect 9580 27124 9596 27140
rect 9612 27124 9628 27140
rect 9644 27124 9660 27140
rect 9260 27092 9276 27108
rect 9292 27092 9308 27108
rect 9324 27092 9340 27108
rect 9356 27092 9372 27108
rect 9388 27092 9404 27108
rect 9420 27092 9436 27108
rect 9452 27092 9468 27108
rect 9484 27092 9500 27108
rect 9516 27092 9532 27108
rect 9548 27092 9564 27108
rect 9580 27092 9596 27108
rect 9612 27092 9628 27108
rect 9644 27092 9660 27108
rect 9260 27060 9276 27076
rect 9292 27060 9308 27076
rect 9324 27060 9340 27076
rect 9356 27060 9372 27076
rect 9388 27060 9404 27076
rect 9420 27060 9436 27076
rect 9452 27060 9468 27076
rect 9484 27060 9500 27076
rect 9516 27060 9532 27076
rect 9548 27060 9564 27076
rect 9580 27060 9596 27076
rect 9612 27060 9628 27076
rect 9644 27060 9660 27076
rect 9260 27028 9276 27044
rect 9292 27028 9308 27044
rect 9324 27028 9340 27044
rect 9356 27028 9372 27044
rect 9388 27028 9404 27044
rect 9420 27028 9436 27044
rect 9452 27028 9468 27044
rect 9484 27028 9500 27044
rect 9516 27028 9532 27044
rect 9548 27028 9564 27044
rect 9580 27028 9596 27044
rect 9612 27028 9628 27044
rect 9644 27028 9660 27044
rect 9260 26996 9276 27012
rect 9292 26996 9308 27012
rect 9324 26996 9340 27012
rect 9356 26996 9372 27012
rect 9388 26996 9404 27012
rect 9420 26996 9436 27012
rect 9452 26996 9468 27012
rect 9484 26996 9500 27012
rect 9516 26996 9532 27012
rect 9548 26996 9564 27012
rect 9580 26996 9596 27012
rect 9612 26996 9628 27012
rect 9644 26996 9660 27012
rect 9260 26964 9276 26980
rect 9292 26964 9308 26980
rect 9324 26964 9340 26980
rect 9356 26964 9372 26980
rect 9388 26964 9404 26980
rect 9420 26964 9436 26980
rect 9452 26964 9468 26980
rect 9484 26964 9500 26980
rect 9516 26964 9532 26980
rect 9548 26964 9564 26980
rect 9580 26964 9596 26980
rect 9612 26964 9628 26980
rect 9644 26964 9660 26980
rect 9260 26932 9276 26948
rect 9292 26932 9308 26948
rect 9324 26932 9340 26948
rect 9356 26932 9372 26948
rect 9388 26932 9404 26948
rect 9420 26932 9436 26948
rect 9452 26932 9468 26948
rect 9484 26932 9500 26948
rect 9516 26932 9532 26948
rect 9548 26932 9564 26948
rect 9580 26932 9596 26948
rect 9612 26932 9628 26948
rect 9644 26932 9660 26948
rect 9260 26900 9276 26916
rect 9292 26900 9308 26916
rect 9324 26900 9340 26916
rect 9356 26900 9372 26916
rect 9388 26900 9404 26916
rect 9420 26900 9436 26916
rect 9452 26900 9468 26916
rect 9484 26900 9500 26916
rect 9516 26900 9532 26916
rect 9548 26900 9564 26916
rect 9580 26900 9596 26916
rect 9612 26900 9628 26916
rect 9644 26900 9660 26916
rect 9260 26868 9276 26884
rect 9292 26868 9308 26884
rect 9324 26868 9340 26884
rect 9356 26868 9372 26884
rect 9388 26868 9404 26884
rect 9420 26868 9436 26884
rect 9452 26868 9468 26884
rect 9484 26868 9500 26884
rect 9516 26868 9532 26884
rect 9548 26868 9564 26884
rect 9580 26868 9596 26884
rect 9612 26868 9628 26884
rect 9644 26868 9660 26884
rect 9260 26836 9276 26852
rect 9292 26836 9308 26852
rect 9324 26836 9340 26852
rect 9356 26836 9372 26852
rect 9388 26836 9404 26852
rect 9420 26836 9436 26852
rect 9452 26836 9468 26852
rect 9484 26836 9500 26852
rect 9516 26836 9532 26852
rect 9548 26836 9564 26852
rect 9580 26836 9596 26852
rect 9612 26836 9628 26852
rect 9644 26836 9660 26852
rect 9260 26804 9276 26820
rect 9292 26804 9308 26820
rect 9324 26804 9340 26820
rect 9356 26804 9372 26820
rect 9388 26804 9404 26820
rect 9420 26804 9436 26820
rect 9452 26804 9468 26820
rect 9484 26804 9500 26820
rect 9516 26804 9532 26820
rect 9548 26804 9564 26820
rect 9580 26804 9596 26820
rect 9612 26804 9628 26820
rect 9644 26804 9660 26820
rect 9260 26772 9276 26788
rect 9292 26772 9308 26788
rect 9324 26772 9340 26788
rect 9356 26772 9372 26788
rect 9388 26772 9404 26788
rect 9420 26772 9436 26788
rect 9452 26772 9468 26788
rect 9484 26772 9500 26788
rect 9516 26772 9532 26788
rect 9548 26772 9564 26788
rect 9580 26772 9596 26788
rect 9612 26772 9628 26788
rect 9644 26772 9660 26788
rect 9260 26740 9276 26756
rect 9292 26740 9308 26756
rect 9324 26740 9340 26756
rect 9356 26740 9372 26756
rect 9388 26740 9404 26756
rect 9420 26740 9436 26756
rect 9452 26740 9468 26756
rect 9484 26740 9500 26756
rect 9516 26740 9532 26756
rect 9548 26740 9564 26756
rect 9580 26740 9596 26756
rect 9612 26740 9628 26756
rect 9644 26740 9660 26756
rect 9260 26708 9276 26724
rect 9292 26708 9308 26724
rect 9324 26708 9340 26724
rect 9356 26708 9372 26724
rect 9388 26708 9404 26724
rect 9420 26708 9436 26724
rect 9452 26708 9468 26724
rect 9484 26708 9500 26724
rect 9516 26708 9532 26724
rect 9548 26708 9564 26724
rect 9580 26708 9596 26724
rect 9612 26708 9628 26724
rect 9644 26708 9660 26724
rect 9260 26676 9276 26692
rect 9292 26676 9308 26692
rect 9324 26676 9340 26692
rect 9356 26676 9372 26692
rect 9388 26676 9404 26692
rect 9420 26676 9436 26692
rect 9452 26676 9468 26692
rect 9484 26676 9500 26692
rect 9516 26676 9532 26692
rect 9548 26676 9564 26692
rect 9580 26676 9596 26692
rect 9612 26676 9628 26692
rect 9644 26676 9660 26692
rect 9260 26644 9276 26660
rect 9292 26644 9308 26660
rect 9324 26644 9340 26660
rect 9356 26644 9372 26660
rect 9388 26644 9404 26660
rect 9420 26644 9436 26660
rect 9452 26644 9468 26660
rect 9484 26644 9500 26660
rect 9516 26644 9532 26660
rect 9548 26644 9564 26660
rect 9580 26644 9596 26660
rect 9612 26644 9628 26660
rect 9644 26644 9660 26660
rect 9260 26612 9276 26628
rect 9292 26612 9308 26628
rect 9324 26612 9340 26628
rect 9356 26612 9372 26628
rect 9388 26612 9404 26628
rect 9420 26612 9436 26628
rect 9452 26612 9468 26628
rect 9484 26612 9500 26628
rect 9516 26612 9532 26628
rect 9548 26612 9564 26628
rect 9580 26612 9596 26628
rect 9612 26612 9628 26628
rect 9644 26612 9660 26628
rect 9260 26580 9276 26596
rect 9292 26580 9308 26596
rect 9324 26580 9340 26596
rect 9356 26580 9372 26596
rect 9388 26580 9404 26596
rect 9420 26580 9436 26596
rect 9452 26580 9468 26596
rect 9484 26580 9500 26596
rect 9516 26580 9532 26596
rect 9548 26580 9564 26596
rect 9580 26580 9596 26596
rect 9612 26580 9628 26596
rect 9644 26580 9660 26596
rect 9260 26548 9276 26564
rect 9292 26548 9308 26564
rect 9324 26548 9340 26564
rect 9356 26548 9372 26564
rect 9388 26548 9404 26564
rect 9420 26548 9436 26564
rect 9452 26548 9468 26564
rect 9484 26548 9500 26564
rect 9516 26548 9532 26564
rect 9548 26548 9564 26564
rect 9580 26548 9596 26564
rect 9612 26548 9628 26564
rect 9644 26548 9660 26564
rect 9260 26516 9276 26532
rect 9292 26516 9308 26532
rect 9324 26516 9340 26532
rect 9356 26516 9372 26532
rect 9388 26516 9404 26532
rect 9420 26516 9436 26532
rect 9452 26516 9468 26532
rect 9484 26516 9500 26532
rect 9516 26516 9532 26532
rect 9548 26516 9564 26532
rect 9580 26516 9596 26532
rect 9612 26516 9628 26532
rect 9644 26516 9660 26532
<< metal2 >>
rect 10040 29020 11760 29180
rect 10041 29008 11759 29020
rect 10041 28992 10060 29008
rect 10076 28992 10092 29008
rect 10108 28992 10124 29008
rect 10140 28992 10156 29008
rect 10172 28992 10188 29008
rect 10204 28992 10220 29008
rect 10236 28992 10252 29008
rect 10268 28992 10284 29008
rect 10300 28992 10316 29008
rect 10332 28992 10348 29008
rect 10364 28992 10380 29008
rect 10396 28992 10412 29008
rect 10428 28992 10444 29008
rect 10460 28992 10476 29008
rect 10492 28992 10508 29008
rect 10524 28992 10540 29008
rect 10556 28992 10572 29008
rect 10588 28992 10604 29008
rect 10620 28992 10636 29008
rect 10652 28992 10668 29008
rect 10684 28992 10700 29008
rect 10716 28992 10732 29008
rect 10748 28992 10764 29008
rect 10780 28992 10796 29008
rect 10812 28992 10828 29008
rect 10844 28992 10860 29008
rect 10876 28992 10892 29008
rect 10908 28992 10924 29008
rect 10940 28992 10956 29008
rect 10972 28992 10988 29008
rect 11004 28992 11020 29008
rect 11036 28992 11052 29008
rect 11068 28992 11084 29008
rect 11100 28992 11116 29008
rect 11132 28992 11148 29008
rect 11164 28992 11180 29008
rect 11196 28992 11212 29008
rect 11228 28992 11244 29008
rect 11260 28992 11276 29008
rect 11292 28992 11308 29008
rect 11324 28992 11340 29008
rect 11356 28992 11372 29008
rect 11388 28992 11404 29008
rect 11420 28992 11436 29008
rect 11452 28992 11468 29008
rect 11484 28992 11500 29008
rect 11516 28992 11532 29008
rect 11548 28992 11564 29008
rect 11580 28992 11596 29008
rect 11612 28992 11628 29008
rect 11644 28992 11660 29008
rect 11676 28992 11692 29008
rect 11708 28992 11724 29008
rect 11740 28992 11759 29008
rect 10041 28976 11759 28992
rect 10041 28960 10060 28976
rect 10076 28960 10092 28976
rect 10108 28960 10124 28976
rect 10140 28960 10156 28976
rect 10172 28960 10188 28976
rect 10204 28960 10220 28976
rect 10236 28960 10252 28976
rect 10268 28960 10284 28976
rect 10300 28960 10316 28976
rect 10332 28960 10348 28976
rect 10364 28960 10380 28976
rect 10396 28960 10412 28976
rect 10428 28960 10444 28976
rect 10460 28960 10476 28976
rect 10492 28960 10508 28976
rect 10524 28960 10540 28976
rect 10556 28960 10572 28976
rect 10588 28960 10604 28976
rect 10620 28960 10636 28976
rect 10652 28960 10668 28976
rect 10684 28960 10700 28976
rect 10716 28960 10732 28976
rect 10748 28960 10764 28976
rect 10780 28960 10796 28976
rect 10812 28960 10828 28976
rect 10844 28960 10860 28976
rect 10876 28960 10892 28976
rect 10908 28960 10924 28976
rect 10940 28960 10956 28976
rect 10972 28960 10988 28976
rect 11004 28960 11020 28976
rect 11036 28960 11052 28976
rect 11068 28960 11084 28976
rect 11100 28960 11116 28976
rect 11132 28960 11148 28976
rect 11164 28960 11180 28976
rect 11196 28960 11212 28976
rect 11228 28960 11244 28976
rect 11260 28960 11276 28976
rect 11292 28960 11308 28976
rect 11324 28960 11340 28976
rect 11356 28960 11372 28976
rect 11388 28960 11404 28976
rect 11420 28960 11436 28976
rect 11452 28960 11468 28976
rect 11484 28960 11500 28976
rect 11516 28960 11532 28976
rect 11548 28960 11564 28976
rect 11580 28960 11596 28976
rect 11612 28960 11628 28976
rect 11644 28960 11660 28976
rect 11676 28960 11692 28976
rect 11708 28960 11724 28976
rect 11740 28960 11759 28976
rect 10041 28944 11759 28960
rect 10041 28928 10060 28944
rect 10076 28928 10092 28944
rect 10108 28928 10124 28944
rect 10140 28928 10156 28944
rect 10172 28928 10188 28944
rect 10204 28928 10220 28944
rect 10236 28928 10252 28944
rect 10268 28928 10284 28944
rect 10300 28928 10316 28944
rect 10332 28928 10348 28944
rect 10364 28928 10380 28944
rect 10396 28928 10412 28944
rect 10428 28928 10444 28944
rect 10460 28928 10476 28944
rect 10492 28928 10508 28944
rect 10524 28928 10540 28944
rect 10556 28928 10572 28944
rect 10588 28928 10604 28944
rect 10620 28928 10636 28944
rect 10652 28928 10668 28944
rect 10684 28928 10700 28944
rect 10716 28928 10732 28944
rect 10748 28928 10764 28944
rect 10780 28928 10796 28944
rect 10812 28928 10828 28944
rect 10844 28928 10860 28944
rect 10876 28928 10892 28944
rect 10908 28928 10924 28944
rect 10940 28928 10956 28944
rect 10972 28928 10988 28944
rect 11004 28928 11020 28944
rect 11036 28928 11052 28944
rect 11068 28928 11084 28944
rect 11100 28928 11116 28944
rect 11132 28928 11148 28944
rect 11164 28928 11180 28944
rect 11196 28928 11212 28944
rect 11228 28928 11244 28944
rect 11260 28928 11276 28944
rect 11292 28928 11308 28944
rect 11324 28928 11340 28944
rect 11356 28928 11372 28944
rect 11388 28928 11404 28944
rect 11420 28928 11436 28944
rect 11452 28928 11468 28944
rect 11484 28928 11500 28944
rect 11516 28928 11532 28944
rect 11548 28928 11564 28944
rect 11580 28928 11596 28944
rect 11612 28928 11628 28944
rect 11644 28928 11660 28944
rect 11676 28928 11692 28944
rect 11708 28928 11724 28944
rect 11740 28928 11759 28944
rect 10041 28912 11759 28928
rect 10041 28896 10060 28912
rect 10076 28896 10092 28912
rect 10108 28896 10124 28912
rect 10140 28896 10156 28912
rect 10172 28896 10188 28912
rect 10204 28896 10220 28912
rect 10236 28896 10252 28912
rect 10268 28896 10284 28912
rect 10300 28896 10316 28912
rect 10332 28896 10348 28912
rect 10364 28896 10380 28912
rect 10396 28896 10412 28912
rect 10428 28896 10444 28912
rect 10460 28896 10476 28912
rect 10492 28896 10508 28912
rect 10524 28896 10540 28912
rect 10556 28896 10572 28912
rect 10588 28896 10604 28912
rect 10620 28896 10636 28912
rect 10652 28896 10668 28912
rect 10684 28896 10700 28912
rect 10716 28896 10732 28912
rect 10748 28896 10764 28912
rect 10780 28896 10796 28912
rect 10812 28896 10828 28912
rect 10844 28896 10860 28912
rect 10876 28896 10892 28912
rect 10908 28896 10924 28912
rect 10940 28896 10956 28912
rect 10972 28896 10988 28912
rect 11004 28896 11020 28912
rect 11036 28896 11052 28912
rect 11068 28896 11084 28912
rect 11100 28896 11116 28912
rect 11132 28896 11148 28912
rect 11164 28896 11180 28912
rect 11196 28896 11212 28912
rect 11228 28896 11244 28912
rect 11260 28896 11276 28912
rect 11292 28896 11308 28912
rect 11324 28896 11340 28912
rect 11356 28896 11372 28912
rect 11388 28896 11404 28912
rect 11420 28896 11436 28912
rect 11452 28896 11468 28912
rect 11484 28896 11500 28912
rect 11516 28896 11532 28912
rect 11548 28896 11564 28912
rect 11580 28896 11596 28912
rect 11612 28896 11628 28912
rect 11644 28896 11660 28912
rect 11676 28896 11692 28912
rect 11708 28896 11724 28912
rect 11740 28896 11759 28912
rect 10041 28880 11759 28896
rect 10041 28864 10060 28880
rect 10076 28864 10092 28880
rect 10108 28864 10124 28880
rect 10140 28864 10156 28880
rect 10172 28864 10188 28880
rect 10204 28864 10220 28880
rect 10236 28864 10252 28880
rect 10268 28864 10284 28880
rect 10300 28864 10316 28880
rect 10332 28864 10348 28880
rect 10364 28864 10380 28880
rect 10396 28864 10412 28880
rect 10428 28864 10444 28880
rect 10460 28864 10476 28880
rect 10492 28864 10508 28880
rect 10524 28864 10540 28880
rect 10556 28864 10572 28880
rect 10588 28864 10604 28880
rect 10620 28864 10636 28880
rect 10652 28864 10668 28880
rect 10684 28864 10700 28880
rect 10716 28864 10732 28880
rect 10748 28864 10764 28880
rect 10780 28864 10796 28880
rect 10812 28864 10828 28880
rect 10844 28864 10860 28880
rect 10876 28864 10892 28880
rect 10908 28864 10924 28880
rect 10940 28864 10956 28880
rect 10972 28864 10988 28880
rect 11004 28864 11020 28880
rect 11036 28864 11052 28880
rect 11068 28864 11084 28880
rect 11100 28864 11116 28880
rect 11132 28864 11148 28880
rect 11164 28864 11180 28880
rect 11196 28864 11212 28880
rect 11228 28864 11244 28880
rect 11260 28864 11276 28880
rect 11292 28864 11308 28880
rect 11324 28864 11340 28880
rect 11356 28864 11372 28880
rect 11388 28864 11404 28880
rect 11420 28864 11436 28880
rect 11452 28864 11468 28880
rect 11484 28864 11500 28880
rect 11516 28864 11532 28880
rect 11548 28864 11564 28880
rect 11580 28864 11596 28880
rect 11612 28864 11628 28880
rect 11644 28864 11660 28880
rect 11676 28864 11692 28880
rect 11708 28864 11724 28880
rect 11740 28864 11759 28880
rect 10041 28848 11759 28864
rect 10041 28832 10060 28848
rect 10076 28832 10092 28848
rect 10108 28832 10124 28848
rect 10140 28832 10156 28848
rect 10172 28832 10188 28848
rect 10204 28832 10220 28848
rect 10236 28832 10252 28848
rect 10268 28832 10284 28848
rect 10300 28832 10316 28848
rect 10332 28832 10348 28848
rect 10364 28832 10380 28848
rect 10396 28832 10412 28848
rect 10428 28832 10444 28848
rect 10460 28832 10476 28848
rect 10492 28832 10508 28848
rect 10524 28832 10540 28848
rect 10556 28832 10572 28848
rect 10588 28832 10604 28848
rect 10620 28832 10636 28848
rect 10652 28832 10668 28848
rect 10684 28832 10700 28848
rect 10716 28832 10732 28848
rect 10748 28832 10764 28848
rect 10780 28832 10796 28848
rect 10812 28832 10828 28848
rect 10844 28832 10860 28848
rect 10876 28832 10892 28848
rect 10908 28832 10924 28848
rect 10940 28832 10956 28848
rect 10972 28832 10988 28848
rect 11004 28832 11020 28848
rect 11036 28832 11052 28848
rect 11068 28832 11084 28848
rect 11100 28832 11116 28848
rect 11132 28832 11148 28848
rect 11164 28832 11180 28848
rect 11196 28832 11212 28848
rect 11228 28832 11244 28848
rect 11260 28832 11276 28848
rect 11292 28832 11308 28848
rect 11324 28832 11340 28848
rect 11356 28832 11372 28848
rect 11388 28832 11404 28848
rect 11420 28832 11436 28848
rect 11452 28832 11468 28848
rect 11484 28832 11500 28848
rect 11516 28832 11532 28848
rect 11548 28832 11564 28848
rect 11580 28832 11596 28848
rect 11612 28832 11628 28848
rect 11644 28832 11660 28848
rect 11676 28832 11692 28848
rect 11708 28832 11724 28848
rect 11740 28832 11759 28848
rect 10041 28816 11759 28832
rect 10041 28800 10060 28816
rect 10076 28800 10092 28816
rect 10108 28800 10124 28816
rect 10140 28800 10156 28816
rect 10172 28800 10188 28816
rect 10204 28800 10220 28816
rect 10236 28800 10252 28816
rect 10268 28800 10284 28816
rect 10300 28800 10316 28816
rect 10332 28800 10348 28816
rect 10364 28800 10380 28816
rect 10396 28800 10412 28816
rect 10428 28800 10444 28816
rect 10460 28800 10476 28816
rect 10492 28800 10508 28816
rect 10524 28800 10540 28816
rect 10556 28800 10572 28816
rect 10588 28800 10604 28816
rect 10620 28800 10636 28816
rect 10652 28800 10668 28816
rect 10684 28800 10700 28816
rect 10716 28800 10732 28816
rect 10748 28800 10764 28816
rect 10780 28800 10796 28816
rect 10812 28800 10828 28816
rect 10844 28800 10860 28816
rect 10876 28800 10892 28816
rect 10908 28800 10924 28816
rect 10940 28800 10956 28816
rect 10972 28800 10988 28816
rect 11004 28800 11020 28816
rect 11036 28800 11052 28816
rect 11068 28800 11084 28816
rect 11100 28800 11116 28816
rect 11132 28800 11148 28816
rect 11164 28800 11180 28816
rect 11196 28800 11212 28816
rect 11228 28800 11244 28816
rect 11260 28800 11276 28816
rect 11292 28800 11308 28816
rect 11324 28800 11340 28816
rect 11356 28800 11372 28816
rect 11388 28800 11404 28816
rect 11420 28800 11436 28816
rect 11452 28800 11468 28816
rect 11484 28800 11500 28816
rect 11516 28800 11532 28816
rect 11548 28800 11564 28816
rect 11580 28800 11596 28816
rect 11612 28800 11628 28816
rect 11644 28800 11660 28816
rect 11676 28800 11692 28816
rect 11708 28800 11724 28816
rect 11740 28800 11759 28816
rect 10041 28784 11759 28800
rect 10041 28768 10060 28784
rect 10076 28768 10092 28784
rect 10108 28768 10124 28784
rect 10140 28768 10156 28784
rect 10172 28768 10188 28784
rect 10204 28768 10220 28784
rect 10236 28768 10252 28784
rect 10268 28768 10284 28784
rect 10300 28768 10316 28784
rect 10332 28768 10348 28784
rect 10364 28768 10380 28784
rect 10396 28768 10412 28784
rect 10428 28768 10444 28784
rect 10460 28768 10476 28784
rect 10492 28768 10508 28784
rect 10524 28768 10540 28784
rect 10556 28768 10572 28784
rect 10588 28768 10604 28784
rect 10620 28768 10636 28784
rect 10652 28768 10668 28784
rect 10684 28768 10700 28784
rect 10716 28768 10732 28784
rect 10748 28768 10764 28784
rect 10780 28768 10796 28784
rect 10812 28768 10828 28784
rect 10844 28768 10860 28784
rect 10876 28768 10892 28784
rect 10908 28768 10924 28784
rect 10940 28768 10956 28784
rect 10972 28768 10988 28784
rect 11004 28768 11020 28784
rect 11036 28768 11052 28784
rect 11068 28768 11084 28784
rect 11100 28768 11116 28784
rect 11132 28768 11148 28784
rect 11164 28768 11180 28784
rect 11196 28768 11212 28784
rect 11228 28768 11244 28784
rect 11260 28768 11276 28784
rect 11292 28768 11308 28784
rect 11324 28768 11340 28784
rect 11356 28768 11372 28784
rect 11388 28768 11404 28784
rect 11420 28768 11436 28784
rect 11452 28768 11468 28784
rect 11484 28768 11500 28784
rect 11516 28768 11532 28784
rect 11548 28768 11564 28784
rect 11580 28768 11596 28784
rect 11612 28768 11628 28784
rect 11644 28768 11660 28784
rect 11676 28768 11692 28784
rect 11708 28768 11724 28784
rect 11740 28768 11759 28784
rect 10041 28752 11759 28768
rect 10041 28736 10060 28752
rect 10076 28736 10092 28752
rect 10108 28736 10124 28752
rect 10140 28736 10156 28752
rect 10172 28736 10188 28752
rect 10204 28736 10220 28752
rect 10236 28736 10252 28752
rect 10268 28736 10284 28752
rect 10300 28736 10316 28752
rect 10332 28736 10348 28752
rect 10364 28736 10380 28752
rect 10396 28736 10412 28752
rect 10428 28736 10444 28752
rect 10460 28736 10476 28752
rect 10492 28736 10508 28752
rect 10524 28736 10540 28752
rect 10556 28736 10572 28752
rect 10588 28736 10604 28752
rect 10620 28736 10636 28752
rect 10652 28736 10668 28752
rect 10684 28736 10700 28752
rect 10716 28736 10732 28752
rect 10748 28736 10764 28752
rect 10780 28736 10796 28752
rect 10812 28736 10828 28752
rect 10844 28736 10860 28752
rect 10876 28736 10892 28752
rect 10908 28736 10924 28752
rect 10940 28736 10956 28752
rect 10972 28736 10988 28752
rect 11004 28736 11020 28752
rect 11036 28736 11052 28752
rect 11068 28736 11084 28752
rect 11100 28736 11116 28752
rect 11132 28736 11148 28752
rect 11164 28736 11180 28752
rect 11196 28736 11212 28752
rect 11228 28736 11244 28752
rect 11260 28736 11276 28752
rect 11292 28736 11308 28752
rect 11324 28736 11340 28752
rect 11356 28736 11372 28752
rect 11388 28736 11404 28752
rect 11420 28736 11436 28752
rect 11452 28736 11468 28752
rect 11484 28736 11500 28752
rect 11516 28736 11532 28752
rect 11548 28736 11564 28752
rect 11580 28736 11596 28752
rect 11612 28736 11628 28752
rect 11644 28736 11660 28752
rect 11676 28736 11692 28752
rect 11708 28736 11724 28752
rect 11740 28736 11759 28752
rect 10041 28720 11759 28736
rect 10041 28704 10060 28720
rect 10076 28704 10092 28720
rect 10108 28704 10124 28720
rect 10140 28704 10156 28720
rect 10172 28704 10188 28720
rect 10204 28704 10220 28720
rect 10236 28704 10252 28720
rect 10268 28704 10284 28720
rect 10300 28704 10316 28720
rect 10332 28704 10348 28720
rect 10364 28704 10380 28720
rect 10396 28704 10412 28720
rect 10428 28704 10444 28720
rect 10460 28704 10476 28720
rect 10492 28704 10508 28720
rect 10524 28704 10540 28720
rect 10556 28704 10572 28720
rect 10588 28704 10604 28720
rect 10620 28704 10636 28720
rect 10652 28704 10668 28720
rect 10684 28704 10700 28720
rect 10716 28704 10732 28720
rect 10748 28704 10764 28720
rect 10780 28704 10796 28720
rect 10812 28704 10828 28720
rect 10844 28704 10860 28720
rect 10876 28704 10892 28720
rect 10908 28704 10924 28720
rect 10940 28704 10956 28720
rect 10972 28704 10988 28720
rect 11004 28704 11020 28720
rect 11036 28704 11052 28720
rect 11068 28704 11084 28720
rect 11100 28704 11116 28720
rect 11132 28704 11148 28720
rect 11164 28704 11180 28720
rect 11196 28704 11212 28720
rect 11228 28704 11244 28720
rect 11260 28704 11276 28720
rect 11292 28704 11308 28720
rect 11324 28704 11340 28720
rect 11356 28704 11372 28720
rect 11388 28704 11404 28720
rect 11420 28704 11436 28720
rect 11452 28704 11468 28720
rect 11484 28704 11500 28720
rect 11516 28704 11532 28720
rect 11548 28704 11564 28720
rect 11580 28704 11596 28720
rect 11612 28704 11628 28720
rect 11644 28704 11660 28720
rect 11676 28704 11692 28720
rect 11708 28704 11724 28720
rect 11740 28704 11759 28720
rect 10041 28688 11759 28704
rect 10041 28672 10060 28688
rect 10076 28672 10092 28688
rect 10108 28672 10124 28688
rect 10140 28672 10156 28688
rect 10172 28672 10188 28688
rect 10204 28672 10220 28688
rect 10236 28672 10252 28688
rect 10268 28672 10284 28688
rect 10300 28672 10316 28688
rect 10332 28672 10348 28688
rect 10364 28672 10380 28688
rect 10396 28672 10412 28688
rect 10428 28672 10444 28688
rect 10460 28672 10476 28688
rect 10492 28672 10508 28688
rect 10524 28672 10540 28688
rect 10556 28672 10572 28688
rect 10588 28672 10604 28688
rect 10620 28672 10636 28688
rect 10652 28672 10668 28688
rect 10684 28672 10700 28688
rect 10716 28672 10732 28688
rect 10748 28672 10764 28688
rect 10780 28672 10796 28688
rect 10812 28672 10828 28688
rect 10844 28672 10860 28688
rect 10876 28672 10892 28688
rect 10908 28672 10924 28688
rect 10940 28672 10956 28688
rect 10972 28672 10988 28688
rect 11004 28672 11020 28688
rect 11036 28672 11052 28688
rect 11068 28672 11084 28688
rect 11100 28672 11116 28688
rect 11132 28672 11148 28688
rect 11164 28672 11180 28688
rect 11196 28672 11212 28688
rect 11228 28672 11244 28688
rect 11260 28672 11276 28688
rect 11292 28672 11308 28688
rect 11324 28672 11340 28688
rect 11356 28672 11372 28688
rect 11388 28672 11404 28688
rect 11420 28672 11436 28688
rect 11452 28672 11468 28688
rect 11484 28672 11500 28688
rect 11516 28672 11532 28688
rect 11548 28672 11564 28688
rect 11580 28672 11596 28688
rect 11612 28672 11628 28688
rect 11644 28672 11660 28688
rect 11676 28672 11692 28688
rect 11708 28672 11724 28688
rect 11740 28672 11759 28688
rect 10041 28656 11759 28672
rect 10041 28640 10060 28656
rect 10076 28640 10092 28656
rect 10108 28640 10124 28656
rect 10140 28640 10156 28656
rect 10172 28640 10188 28656
rect 10204 28640 10220 28656
rect 10236 28640 10252 28656
rect 10268 28640 10284 28656
rect 10300 28640 10316 28656
rect 10332 28640 10348 28656
rect 10364 28640 10380 28656
rect 10396 28640 10412 28656
rect 10428 28640 10444 28656
rect 10460 28640 10476 28656
rect 10492 28640 10508 28656
rect 10524 28640 10540 28656
rect 10556 28640 10572 28656
rect 10588 28640 10604 28656
rect 10620 28640 10636 28656
rect 10652 28640 10668 28656
rect 10684 28640 10700 28656
rect 10716 28640 10732 28656
rect 10748 28640 10764 28656
rect 10780 28640 10796 28656
rect 10812 28640 10828 28656
rect 10844 28640 10860 28656
rect 10876 28640 10892 28656
rect 10908 28640 10924 28656
rect 10940 28640 10956 28656
rect 10972 28640 10988 28656
rect 11004 28640 11020 28656
rect 11036 28640 11052 28656
rect 11068 28640 11084 28656
rect 11100 28640 11116 28656
rect 11132 28640 11148 28656
rect 11164 28640 11180 28656
rect 11196 28640 11212 28656
rect 11228 28640 11244 28656
rect 11260 28640 11276 28656
rect 11292 28640 11308 28656
rect 11324 28640 11340 28656
rect 11356 28640 11372 28656
rect 11388 28640 11404 28656
rect 11420 28640 11436 28656
rect 11452 28640 11468 28656
rect 11484 28640 11500 28656
rect 11516 28640 11532 28656
rect 11548 28640 11564 28656
rect 11580 28640 11596 28656
rect 11612 28640 11628 28656
rect 11644 28640 11660 28656
rect 11676 28640 11692 28656
rect 11708 28640 11724 28656
rect 11740 28640 11759 28656
rect 10041 28624 11759 28640
rect 10041 28608 10060 28624
rect 10076 28608 10092 28624
rect 10108 28608 10124 28624
rect 10140 28608 10156 28624
rect 10172 28608 10188 28624
rect 10204 28608 10220 28624
rect 10236 28608 10252 28624
rect 10268 28608 10284 28624
rect 10300 28608 10316 28624
rect 10332 28608 10348 28624
rect 10364 28608 10380 28624
rect 10396 28608 10412 28624
rect 10428 28608 10444 28624
rect 10460 28608 10476 28624
rect 10492 28608 10508 28624
rect 10524 28608 10540 28624
rect 10556 28608 10572 28624
rect 10588 28608 10604 28624
rect 10620 28608 10636 28624
rect 10652 28608 10668 28624
rect 10684 28608 10700 28624
rect 10716 28608 10732 28624
rect 10748 28608 10764 28624
rect 10780 28608 10796 28624
rect 10812 28608 10828 28624
rect 10844 28608 10860 28624
rect 10876 28608 10892 28624
rect 10908 28608 10924 28624
rect 10940 28608 10956 28624
rect 10972 28608 10988 28624
rect 11004 28608 11020 28624
rect 11036 28608 11052 28624
rect 11068 28608 11084 28624
rect 11100 28608 11116 28624
rect 11132 28608 11148 28624
rect 11164 28608 11180 28624
rect 11196 28608 11212 28624
rect 11228 28608 11244 28624
rect 11260 28608 11276 28624
rect 11292 28608 11308 28624
rect 11324 28608 11340 28624
rect 11356 28608 11372 28624
rect 11388 28608 11404 28624
rect 11420 28608 11436 28624
rect 11452 28608 11468 28624
rect 11484 28608 11500 28624
rect 11516 28608 11532 28624
rect 11548 28608 11564 28624
rect 11580 28608 11596 28624
rect 11612 28608 11628 28624
rect 11644 28608 11660 28624
rect 11676 28608 11692 28624
rect 11708 28608 11724 28624
rect 11740 28608 11759 28624
rect 10041 28592 11759 28608
rect 10041 28576 10060 28592
rect 10076 28576 10092 28592
rect 10108 28576 10124 28592
rect 10140 28576 10156 28592
rect 10172 28576 10188 28592
rect 10204 28576 10220 28592
rect 10236 28576 10252 28592
rect 10268 28576 10284 28592
rect 10300 28576 10316 28592
rect 10332 28576 10348 28592
rect 10364 28576 10380 28592
rect 10396 28576 10412 28592
rect 10428 28576 10444 28592
rect 10460 28576 10476 28592
rect 10492 28576 10508 28592
rect 10524 28576 10540 28592
rect 10556 28576 10572 28592
rect 10588 28576 10604 28592
rect 10620 28576 10636 28592
rect 10652 28576 10668 28592
rect 10684 28576 10700 28592
rect 10716 28576 10732 28592
rect 10748 28576 10764 28592
rect 10780 28576 10796 28592
rect 10812 28576 10828 28592
rect 10844 28576 10860 28592
rect 10876 28576 10892 28592
rect 10908 28576 10924 28592
rect 10940 28576 10956 28592
rect 10972 28576 10988 28592
rect 11004 28576 11020 28592
rect 11036 28576 11052 28592
rect 11068 28576 11084 28592
rect 11100 28576 11116 28592
rect 11132 28576 11148 28592
rect 11164 28576 11180 28592
rect 11196 28576 11212 28592
rect 11228 28576 11244 28592
rect 11260 28576 11276 28592
rect 11292 28576 11308 28592
rect 11324 28576 11340 28592
rect 11356 28576 11372 28592
rect 11388 28576 11404 28592
rect 11420 28576 11436 28592
rect 11452 28576 11468 28592
rect 11484 28576 11500 28592
rect 11516 28576 11532 28592
rect 11548 28576 11564 28592
rect 11580 28576 11596 28592
rect 11612 28576 11628 28592
rect 11644 28576 11660 28592
rect 11676 28576 11692 28592
rect 11708 28576 11724 28592
rect 11740 28576 11759 28592
rect 10041 28560 11759 28576
rect 10041 28544 10060 28560
rect 10076 28544 10092 28560
rect 10108 28544 10124 28560
rect 10140 28544 10156 28560
rect 10172 28544 10188 28560
rect 10204 28544 10220 28560
rect 10236 28544 10252 28560
rect 10268 28544 10284 28560
rect 10300 28544 10316 28560
rect 10332 28544 10348 28560
rect 10364 28544 10380 28560
rect 10396 28544 10412 28560
rect 10428 28544 10444 28560
rect 10460 28544 10476 28560
rect 10492 28544 10508 28560
rect 10524 28544 10540 28560
rect 10556 28544 10572 28560
rect 10588 28544 10604 28560
rect 10620 28544 10636 28560
rect 10652 28544 10668 28560
rect 10684 28544 10700 28560
rect 10716 28544 10732 28560
rect 10748 28544 10764 28560
rect 10780 28544 10796 28560
rect 10812 28544 10828 28560
rect 10844 28544 10860 28560
rect 10876 28544 10892 28560
rect 10908 28544 10924 28560
rect 10940 28544 10956 28560
rect 10972 28544 10988 28560
rect 11004 28544 11020 28560
rect 11036 28544 11052 28560
rect 11068 28544 11084 28560
rect 11100 28544 11116 28560
rect 11132 28544 11148 28560
rect 11164 28544 11180 28560
rect 11196 28544 11212 28560
rect 11228 28544 11244 28560
rect 11260 28544 11276 28560
rect 11292 28544 11308 28560
rect 11324 28544 11340 28560
rect 11356 28544 11372 28560
rect 11388 28544 11404 28560
rect 11420 28544 11436 28560
rect 11452 28544 11468 28560
rect 11484 28544 11500 28560
rect 11516 28544 11532 28560
rect 11548 28544 11564 28560
rect 11580 28544 11596 28560
rect 11612 28544 11628 28560
rect 11644 28544 11660 28560
rect 11676 28544 11692 28560
rect 11708 28544 11724 28560
rect 11740 28544 11759 28560
rect 10041 28528 11759 28544
rect 10041 28512 10060 28528
rect 10076 28512 10092 28528
rect 10108 28512 10124 28528
rect 10140 28512 10156 28528
rect 10172 28512 10188 28528
rect 10204 28512 10220 28528
rect 10236 28512 10252 28528
rect 10268 28512 10284 28528
rect 10300 28512 10316 28528
rect 10332 28512 10348 28528
rect 10364 28512 10380 28528
rect 10396 28512 10412 28528
rect 10428 28512 10444 28528
rect 10460 28512 10476 28528
rect 10492 28512 10508 28528
rect 10524 28512 10540 28528
rect 10556 28512 10572 28528
rect 10588 28512 10604 28528
rect 10620 28512 10636 28528
rect 10652 28512 10668 28528
rect 10684 28512 10700 28528
rect 10716 28512 10732 28528
rect 10748 28512 10764 28528
rect 10780 28512 10796 28528
rect 10812 28512 10828 28528
rect 10844 28512 10860 28528
rect 10876 28512 10892 28528
rect 10908 28512 10924 28528
rect 10940 28512 10956 28528
rect 10972 28512 10988 28528
rect 11004 28512 11020 28528
rect 11036 28512 11052 28528
rect 11068 28512 11084 28528
rect 11100 28512 11116 28528
rect 11132 28512 11148 28528
rect 11164 28512 11180 28528
rect 11196 28512 11212 28528
rect 11228 28512 11244 28528
rect 11260 28512 11276 28528
rect 11292 28512 11308 28528
rect 11324 28512 11340 28528
rect 11356 28512 11372 28528
rect 11388 28512 11404 28528
rect 11420 28512 11436 28528
rect 11452 28512 11468 28528
rect 11484 28512 11500 28528
rect 11516 28512 11532 28528
rect 11548 28512 11564 28528
rect 11580 28512 11596 28528
rect 11612 28512 11628 28528
rect 11644 28512 11660 28528
rect 11676 28512 11692 28528
rect 11708 28512 11724 28528
rect 11740 28512 11759 28528
rect 10041 28501 11759 28512
rect 8820 27699 9240 27700
rect 8820 27684 9679 27699
rect 8820 27668 9260 27684
rect 9276 27668 9292 27684
rect 9308 27668 9324 27684
rect 9340 27668 9356 27684
rect 9372 27668 9388 27684
rect 9404 27668 9420 27684
rect 9436 27668 9452 27684
rect 9468 27668 9484 27684
rect 9500 27668 9516 27684
rect 9532 27668 9548 27684
rect 9564 27668 9580 27684
rect 9596 27668 9612 27684
rect 9628 27668 9644 27684
rect 9660 27668 9679 27684
rect 8820 27652 9679 27668
rect 8820 27636 9260 27652
rect 9276 27636 9292 27652
rect 9308 27636 9324 27652
rect 9340 27636 9356 27652
rect 9372 27636 9388 27652
rect 9404 27636 9420 27652
rect 9436 27636 9452 27652
rect 9468 27636 9484 27652
rect 9500 27636 9516 27652
rect 9532 27636 9548 27652
rect 9564 27636 9580 27652
rect 9596 27636 9612 27652
rect 9628 27636 9644 27652
rect 9660 27636 9679 27652
rect 8820 27620 9679 27636
rect 8820 27604 9260 27620
rect 9276 27604 9292 27620
rect 9308 27604 9324 27620
rect 9340 27604 9356 27620
rect 9372 27604 9388 27620
rect 9404 27604 9420 27620
rect 9436 27604 9452 27620
rect 9468 27604 9484 27620
rect 9500 27604 9516 27620
rect 9532 27604 9548 27620
rect 9564 27604 9580 27620
rect 9596 27604 9612 27620
rect 9628 27604 9644 27620
rect 9660 27604 9679 27620
rect 8820 27588 9679 27604
rect 8820 27572 9260 27588
rect 9276 27572 9292 27588
rect 9308 27572 9324 27588
rect 9340 27572 9356 27588
rect 9372 27572 9388 27588
rect 9404 27572 9420 27588
rect 9436 27572 9452 27588
rect 9468 27572 9484 27588
rect 9500 27572 9516 27588
rect 9532 27572 9548 27588
rect 9564 27572 9580 27588
rect 9596 27572 9612 27588
rect 9628 27572 9644 27588
rect 9660 27572 9679 27588
rect 8820 27556 9679 27572
rect 8820 27540 9260 27556
rect 9276 27540 9292 27556
rect 9308 27540 9324 27556
rect 9340 27540 9356 27556
rect 9372 27540 9388 27556
rect 9404 27540 9420 27556
rect 9436 27540 9452 27556
rect 9468 27540 9484 27556
rect 9500 27540 9516 27556
rect 9532 27540 9548 27556
rect 9564 27540 9580 27556
rect 9596 27540 9612 27556
rect 9628 27540 9644 27556
rect 9660 27540 9679 27556
rect 8820 27524 9679 27540
rect 8820 27508 9260 27524
rect 9276 27508 9292 27524
rect 9308 27508 9324 27524
rect 9340 27508 9356 27524
rect 9372 27508 9388 27524
rect 9404 27508 9420 27524
rect 9436 27508 9452 27524
rect 9468 27508 9484 27524
rect 9500 27508 9516 27524
rect 9532 27508 9548 27524
rect 9564 27508 9580 27524
rect 9596 27508 9612 27524
rect 9628 27508 9644 27524
rect 9660 27508 9679 27524
rect 8820 27492 9679 27508
rect 8820 27476 9260 27492
rect 9276 27476 9292 27492
rect 9308 27476 9324 27492
rect 9340 27476 9356 27492
rect 9372 27476 9388 27492
rect 9404 27476 9420 27492
rect 9436 27476 9452 27492
rect 9468 27476 9484 27492
rect 9500 27476 9516 27492
rect 9532 27476 9548 27492
rect 9564 27476 9580 27492
rect 9596 27476 9612 27492
rect 9628 27476 9644 27492
rect 9660 27476 9679 27492
rect 8820 27460 9679 27476
rect 8820 27444 9260 27460
rect 9276 27444 9292 27460
rect 9308 27444 9324 27460
rect 9340 27444 9356 27460
rect 9372 27444 9388 27460
rect 9404 27444 9420 27460
rect 9436 27444 9452 27460
rect 9468 27444 9484 27460
rect 9500 27444 9516 27460
rect 9532 27444 9548 27460
rect 9564 27444 9580 27460
rect 9596 27444 9612 27460
rect 9628 27444 9644 27460
rect 9660 27444 9679 27460
rect 8820 27428 9679 27444
rect 8820 27412 9260 27428
rect 9276 27412 9292 27428
rect 9308 27412 9324 27428
rect 9340 27412 9356 27428
rect 9372 27412 9388 27428
rect 9404 27412 9420 27428
rect 9436 27412 9452 27428
rect 9468 27412 9484 27428
rect 9500 27412 9516 27428
rect 9532 27412 9548 27428
rect 9564 27412 9580 27428
rect 9596 27412 9612 27428
rect 9628 27412 9644 27428
rect 9660 27412 9679 27428
rect 8820 27396 9679 27412
rect 8820 27380 9260 27396
rect 9276 27380 9292 27396
rect 9308 27380 9324 27396
rect 9340 27380 9356 27396
rect 9372 27380 9388 27396
rect 9404 27380 9420 27396
rect 9436 27380 9452 27396
rect 9468 27380 9484 27396
rect 9500 27380 9516 27396
rect 9532 27380 9548 27396
rect 9564 27380 9580 27396
rect 9596 27380 9612 27396
rect 9628 27380 9644 27396
rect 9660 27380 9679 27396
rect 8820 27364 9679 27380
rect 8820 27348 9260 27364
rect 9276 27348 9292 27364
rect 9308 27348 9324 27364
rect 9340 27348 9356 27364
rect 9372 27348 9388 27364
rect 9404 27348 9420 27364
rect 9436 27348 9452 27364
rect 9468 27348 9484 27364
rect 9500 27348 9516 27364
rect 9532 27348 9548 27364
rect 9564 27348 9580 27364
rect 9596 27348 9612 27364
rect 9628 27348 9644 27364
rect 9660 27348 9679 27364
rect 8820 27332 9679 27348
rect 8820 27316 9260 27332
rect 9276 27316 9292 27332
rect 9308 27316 9324 27332
rect 9340 27316 9356 27332
rect 9372 27316 9388 27332
rect 9404 27316 9420 27332
rect 9436 27316 9452 27332
rect 9468 27316 9484 27332
rect 9500 27316 9516 27332
rect 9532 27316 9548 27332
rect 9564 27316 9580 27332
rect 9596 27316 9612 27332
rect 9628 27316 9644 27332
rect 9660 27316 9679 27332
rect 8820 27300 9679 27316
rect 8820 27284 9260 27300
rect 9276 27284 9292 27300
rect 9308 27284 9324 27300
rect 9340 27284 9356 27300
rect 9372 27284 9388 27300
rect 9404 27284 9420 27300
rect 9436 27284 9452 27300
rect 9468 27284 9484 27300
rect 9500 27284 9516 27300
rect 9532 27284 9548 27300
rect 9564 27284 9580 27300
rect 9596 27284 9612 27300
rect 9628 27284 9644 27300
rect 9660 27284 9679 27300
rect 8820 27268 9679 27284
rect 8820 27252 9260 27268
rect 9276 27252 9292 27268
rect 9308 27252 9324 27268
rect 9340 27252 9356 27268
rect 9372 27252 9388 27268
rect 9404 27252 9420 27268
rect 9436 27252 9452 27268
rect 9468 27252 9484 27268
rect 9500 27252 9516 27268
rect 9532 27252 9548 27268
rect 9564 27252 9580 27268
rect 9596 27252 9612 27268
rect 9628 27252 9644 27268
rect 9660 27252 9679 27268
rect 8820 27236 9679 27252
rect 8820 27220 9260 27236
rect 9276 27220 9292 27236
rect 9308 27220 9324 27236
rect 9340 27220 9356 27236
rect 9372 27220 9388 27236
rect 9404 27220 9420 27236
rect 9436 27220 9452 27236
rect 9468 27220 9484 27236
rect 9500 27220 9516 27236
rect 9532 27220 9548 27236
rect 9564 27220 9580 27236
rect 9596 27220 9612 27236
rect 9628 27220 9644 27236
rect 9660 27220 9679 27236
rect 8820 27204 9679 27220
rect 8820 27188 9260 27204
rect 9276 27188 9292 27204
rect 9308 27188 9324 27204
rect 9340 27188 9356 27204
rect 9372 27188 9388 27204
rect 9404 27188 9420 27204
rect 9436 27188 9452 27204
rect 9468 27188 9484 27204
rect 9500 27188 9516 27204
rect 9532 27188 9548 27204
rect 9564 27188 9580 27204
rect 9596 27188 9612 27204
rect 9628 27188 9644 27204
rect 9660 27188 9679 27204
rect 8820 27172 9679 27188
rect 8820 27156 9260 27172
rect 9276 27156 9292 27172
rect 9308 27156 9324 27172
rect 9340 27156 9356 27172
rect 9372 27156 9388 27172
rect 9404 27156 9420 27172
rect 9436 27156 9452 27172
rect 9468 27156 9484 27172
rect 9500 27156 9516 27172
rect 9532 27156 9548 27172
rect 9564 27156 9580 27172
rect 9596 27156 9612 27172
rect 9628 27156 9644 27172
rect 9660 27156 9679 27172
rect 8820 27140 9679 27156
rect 8820 27124 9260 27140
rect 9276 27124 9292 27140
rect 9308 27124 9324 27140
rect 9340 27124 9356 27140
rect 9372 27124 9388 27140
rect 9404 27124 9420 27140
rect 9436 27124 9452 27140
rect 9468 27124 9484 27140
rect 9500 27124 9516 27140
rect 9532 27124 9548 27140
rect 9564 27124 9580 27140
rect 9596 27124 9612 27140
rect 9628 27124 9644 27140
rect 9660 27124 9679 27140
rect 8820 27108 9679 27124
rect 8820 27092 9260 27108
rect 9276 27092 9292 27108
rect 9308 27092 9324 27108
rect 9340 27092 9356 27108
rect 9372 27092 9388 27108
rect 9404 27092 9420 27108
rect 9436 27092 9452 27108
rect 9468 27092 9484 27108
rect 9500 27092 9516 27108
rect 9532 27092 9548 27108
rect 9564 27092 9580 27108
rect 9596 27092 9612 27108
rect 9628 27092 9644 27108
rect 9660 27092 9679 27108
rect 8820 27076 9679 27092
rect 8820 27060 9260 27076
rect 9276 27060 9292 27076
rect 9308 27060 9324 27076
rect 9340 27060 9356 27076
rect 9372 27060 9388 27076
rect 9404 27060 9420 27076
rect 9436 27060 9452 27076
rect 9468 27060 9484 27076
rect 9500 27060 9516 27076
rect 9532 27060 9548 27076
rect 9564 27060 9580 27076
rect 9596 27060 9612 27076
rect 9628 27060 9644 27076
rect 9660 27060 9679 27076
rect 8820 27044 9679 27060
rect 8820 27028 9260 27044
rect 9276 27028 9292 27044
rect 9308 27028 9324 27044
rect 9340 27028 9356 27044
rect 9372 27028 9388 27044
rect 9404 27028 9420 27044
rect 9436 27028 9452 27044
rect 9468 27028 9484 27044
rect 9500 27028 9516 27044
rect 9532 27028 9548 27044
rect 9564 27028 9580 27044
rect 9596 27028 9612 27044
rect 9628 27028 9644 27044
rect 9660 27028 9679 27044
rect 8820 27012 9679 27028
rect 8820 26996 9260 27012
rect 9276 26996 9292 27012
rect 9308 26996 9324 27012
rect 9340 26996 9356 27012
rect 9372 26996 9388 27012
rect 9404 26996 9420 27012
rect 9436 26996 9452 27012
rect 9468 26996 9484 27012
rect 9500 26996 9516 27012
rect 9532 26996 9548 27012
rect 9564 26996 9580 27012
rect 9596 26996 9612 27012
rect 9628 26996 9644 27012
rect 9660 26996 9679 27012
rect 8820 26980 9679 26996
rect 8820 26964 9260 26980
rect 9276 26964 9292 26980
rect 9308 26964 9324 26980
rect 9340 26964 9356 26980
rect 9372 26964 9388 26980
rect 9404 26964 9420 26980
rect 9436 26964 9452 26980
rect 9468 26964 9484 26980
rect 9500 26964 9516 26980
rect 9532 26964 9548 26980
rect 9564 26964 9580 26980
rect 9596 26964 9612 26980
rect 9628 26964 9644 26980
rect 9660 26964 9679 26980
rect 8820 26948 9679 26964
rect 8820 26932 9260 26948
rect 9276 26932 9292 26948
rect 9308 26932 9324 26948
rect 9340 26932 9356 26948
rect 9372 26932 9388 26948
rect 9404 26932 9420 26948
rect 9436 26932 9452 26948
rect 9468 26932 9484 26948
rect 9500 26932 9516 26948
rect 9532 26932 9548 26948
rect 9564 26932 9580 26948
rect 9596 26932 9612 26948
rect 9628 26932 9644 26948
rect 9660 26932 9679 26948
rect 8820 26916 9679 26932
rect 8820 26900 9260 26916
rect 9276 26900 9292 26916
rect 9308 26900 9324 26916
rect 9340 26900 9356 26916
rect 9372 26900 9388 26916
rect 9404 26900 9420 26916
rect 9436 26900 9452 26916
rect 9468 26900 9484 26916
rect 9500 26900 9516 26916
rect 9532 26900 9548 26916
rect 9564 26900 9580 26916
rect 9596 26900 9612 26916
rect 9628 26900 9644 26916
rect 9660 26900 9679 26916
rect 8820 26884 9679 26900
rect 8820 26868 9260 26884
rect 9276 26868 9292 26884
rect 9308 26868 9324 26884
rect 9340 26868 9356 26884
rect 9372 26868 9388 26884
rect 9404 26868 9420 26884
rect 9436 26868 9452 26884
rect 9468 26868 9484 26884
rect 9500 26868 9516 26884
rect 9532 26868 9548 26884
rect 9564 26868 9580 26884
rect 9596 26868 9612 26884
rect 9628 26868 9644 26884
rect 9660 26868 9679 26884
rect 8820 26852 9679 26868
rect 8820 26836 9260 26852
rect 9276 26836 9292 26852
rect 9308 26836 9324 26852
rect 9340 26836 9356 26852
rect 9372 26836 9388 26852
rect 9404 26836 9420 26852
rect 9436 26836 9452 26852
rect 9468 26836 9484 26852
rect 9500 26836 9516 26852
rect 9532 26836 9548 26852
rect 9564 26836 9580 26852
rect 9596 26836 9612 26852
rect 9628 26836 9644 26852
rect 9660 26836 9679 26852
rect 8820 26820 9679 26836
rect 8820 26804 9260 26820
rect 9276 26804 9292 26820
rect 9308 26804 9324 26820
rect 9340 26804 9356 26820
rect 9372 26804 9388 26820
rect 9404 26804 9420 26820
rect 9436 26804 9452 26820
rect 9468 26804 9484 26820
rect 9500 26804 9516 26820
rect 9532 26804 9548 26820
rect 9564 26804 9580 26820
rect 9596 26804 9612 26820
rect 9628 26804 9644 26820
rect 9660 26804 9679 26820
rect 8820 26788 9679 26804
rect 8820 26772 9260 26788
rect 9276 26772 9292 26788
rect 9308 26772 9324 26788
rect 9340 26772 9356 26788
rect 9372 26772 9388 26788
rect 9404 26772 9420 26788
rect 9436 26772 9452 26788
rect 9468 26772 9484 26788
rect 9500 26772 9516 26788
rect 9532 26772 9548 26788
rect 9564 26772 9580 26788
rect 9596 26772 9612 26788
rect 9628 26772 9644 26788
rect 9660 26772 9679 26788
rect 8820 26756 9679 26772
rect 8820 26740 9260 26756
rect 9276 26740 9292 26756
rect 9308 26740 9324 26756
rect 9340 26740 9356 26756
rect 9372 26740 9388 26756
rect 9404 26740 9420 26756
rect 9436 26740 9452 26756
rect 9468 26740 9484 26756
rect 9500 26740 9516 26756
rect 9532 26740 9548 26756
rect 9564 26740 9580 26756
rect 9596 26740 9612 26756
rect 9628 26740 9644 26756
rect 9660 26740 9679 26756
rect 8820 26724 9679 26740
rect 8820 26708 9260 26724
rect 9276 26708 9292 26724
rect 9308 26708 9324 26724
rect 9340 26708 9356 26724
rect 9372 26708 9388 26724
rect 9404 26708 9420 26724
rect 9436 26708 9452 26724
rect 9468 26708 9484 26724
rect 9500 26708 9516 26724
rect 9532 26708 9548 26724
rect 9564 26708 9580 26724
rect 9596 26708 9612 26724
rect 9628 26708 9644 26724
rect 9660 26708 9679 26724
rect 8820 26692 9679 26708
rect 8820 26676 9260 26692
rect 9276 26676 9292 26692
rect 9308 26676 9324 26692
rect 9340 26676 9356 26692
rect 9372 26676 9388 26692
rect 9404 26676 9420 26692
rect 9436 26676 9452 26692
rect 9468 26676 9484 26692
rect 9500 26676 9516 26692
rect 9532 26676 9548 26692
rect 9564 26676 9580 26692
rect 9596 26676 9612 26692
rect 9628 26676 9644 26692
rect 9660 26676 9679 26692
rect 8820 26660 9679 26676
rect 8820 26644 9260 26660
rect 9276 26644 9292 26660
rect 9308 26644 9324 26660
rect 9340 26644 9356 26660
rect 9372 26644 9388 26660
rect 9404 26644 9420 26660
rect 9436 26644 9452 26660
rect 9468 26644 9484 26660
rect 9500 26644 9516 26660
rect 9532 26644 9548 26660
rect 9564 26644 9580 26660
rect 9596 26644 9612 26660
rect 9628 26644 9644 26660
rect 9660 26644 9679 26660
rect 8820 26628 9679 26644
rect 8820 26612 9260 26628
rect 9276 26612 9292 26628
rect 9308 26612 9324 26628
rect 9340 26612 9356 26628
rect 9372 26612 9388 26628
rect 9404 26612 9420 26628
rect 9436 26612 9452 26628
rect 9468 26612 9484 26628
rect 9500 26612 9516 26628
rect 9532 26612 9548 26628
rect 9564 26612 9580 26628
rect 9596 26612 9612 26628
rect 9628 26612 9644 26628
rect 9660 26612 9679 26628
rect 12480 26720 12580 29180
rect 15180 26920 15280 29180
rect 17880 27281 17980 29180
rect 17880 27280 18179 27281
rect 17881 27254 18179 27280
rect 17881 27238 17894 27254
rect 17910 27238 17926 27254
rect 17942 27238 17958 27254
rect 17974 27238 17990 27254
rect 18006 27238 18022 27254
rect 18038 27238 18054 27254
rect 18070 27238 18086 27254
rect 18102 27238 18118 27254
rect 18134 27238 18150 27254
rect 18166 27238 18179 27254
rect 17881 27222 18179 27238
rect 17881 27206 17894 27222
rect 17910 27206 17926 27222
rect 17942 27206 17958 27222
rect 17974 27206 17990 27222
rect 18006 27206 18022 27222
rect 18038 27206 18054 27222
rect 18070 27206 18086 27222
rect 18102 27206 18118 27222
rect 18134 27206 18150 27222
rect 18166 27206 18179 27222
rect 17881 27181 18179 27206
rect 20580 27080 20680 29180
rect 25440 28400 25540 29180
rect 28140 28400 28240 29180
rect 25320 28300 25540 28400
rect 26020 28320 28240 28400
rect 24301 27254 24599 27279
rect 24301 27238 24314 27254
rect 24330 27238 24346 27254
rect 24362 27238 24378 27254
rect 24394 27238 24410 27254
rect 24426 27238 24442 27254
rect 24458 27238 24474 27254
rect 24490 27238 24506 27254
rect 24522 27238 24538 27254
rect 24554 27238 24570 27254
rect 24586 27238 24599 27254
rect 24301 27222 24599 27238
rect 24301 27206 24314 27222
rect 24330 27206 24346 27222
rect 24362 27206 24378 27222
rect 24394 27206 24410 27222
rect 24426 27206 24442 27222
rect 24458 27206 24474 27222
rect 24490 27206 24506 27222
rect 24522 27206 24538 27222
rect 24554 27206 24570 27222
rect 24586 27206 24599 27222
rect 24301 27180 24599 27206
rect 24301 27179 24600 27180
rect 20580 27000 24460 27080
rect 15180 26820 24320 26920
rect 12480 26620 17580 26720
rect 8820 26596 9679 26612
rect 8820 26580 9260 26596
rect 9276 26580 9292 26596
rect 9308 26580 9324 26596
rect 9340 26580 9356 26596
rect 9372 26580 9388 26596
rect 9404 26580 9420 26596
rect 9436 26580 9452 26596
rect 9468 26580 9484 26596
rect 9500 26580 9516 26596
rect 9532 26580 9548 26596
rect 9564 26580 9580 26596
rect 9596 26580 9612 26596
rect 9628 26580 9644 26596
rect 9660 26580 9679 26596
rect 8820 26564 9679 26580
rect 8820 26548 9260 26564
rect 9276 26548 9292 26564
rect 9308 26548 9324 26564
rect 9340 26548 9356 26564
rect 9372 26548 9388 26564
rect 9404 26548 9420 26564
rect 9436 26548 9452 26564
rect 9468 26548 9484 26564
rect 9500 26548 9516 26564
rect 9532 26548 9548 26564
rect 9564 26548 9580 26564
rect 9596 26548 9612 26564
rect 9628 26548 9644 26564
rect 9660 26548 9679 26564
rect 8820 26532 9679 26548
rect 8820 26516 9260 26532
rect 9276 26516 9292 26532
rect 9308 26516 9324 26532
rect 9340 26516 9356 26532
rect 9372 26516 9388 26532
rect 9404 26516 9420 26532
rect 9436 26516 9452 26532
rect 9468 26516 9484 26532
rect 9500 26516 9516 26532
rect 9532 26516 9548 26532
rect 9564 26516 9580 26532
rect 9596 26516 9612 26532
rect 9628 26516 9644 26532
rect 9660 26516 9679 26532
rect 8820 26501 9679 26516
rect 8820 26500 9240 26501
rect 17480 26400 17580 26620
rect 24240 26380 24320 26820
rect 24380 26380 24460 27000
rect 24520 26380 24600 27179
rect 25320 26340 25420 28300
rect 26020 26380 26100 28320
rect 27720 28160 29180 28240
rect 10101 25484 10179 25499
rect 10101 25468 10116 25484
rect 10132 25468 10148 25484
rect 10164 25468 10179 25484
rect 10101 25452 10179 25468
rect 10101 25436 10116 25452
rect 10132 25436 10148 25452
rect 10164 25436 10179 25452
rect 10101 25420 10179 25436
rect 9941 25324 10019 25339
rect 9941 25308 9956 25324
rect 9972 25308 9988 25324
rect 10004 25308 10019 25324
rect 9941 25292 10019 25308
rect 9941 25276 9956 25292
rect 9972 25276 9988 25292
rect 10004 25276 10019 25292
rect 9941 25260 10019 25276
rect 9781 25164 9859 25179
rect 9781 25148 9796 25164
rect 9812 25148 9828 25164
rect 9844 25148 9859 25164
rect 9781 25132 9859 25148
rect 9781 25116 9796 25132
rect 9812 25116 9828 25132
rect 9844 25116 9859 25132
rect 9781 25100 9859 25116
rect 9621 24464 9699 24479
rect 9621 24448 9636 24464
rect 9652 24448 9668 24464
rect 9684 24448 9699 24464
rect 9621 24432 9699 24448
rect 9621 24416 9636 24432
rect 9652 24416 9668 24432
rect 9684 24416 9699 24432
rect 9621 24400 9699 24416
rect 8820 23379 8960 23380
rect 8820 23354 9099 23379
rect 8820 23338 8974 23354
rect 8990 23338 9006 23354
rect 9022 23338 9038 23354
rect 9054 23338 9070 23354
rect 9086 23338 9099 23354
rect 8820 23322 9099 23338
rect 8820 23306 8974 23322
rect 8990 23306 9006 23322
rect 9022 23306 9038 23322
rect 9054 23306 9070 23322
rect 9086 23306 9099 23322
rect 8820 23290 9099 23306
rect 8820 23274 8974 23290
rect 8990 23274 9006 23290
rect 9022 23274 9038 23290
rect 9054 23274 9070 23290
rect 9086 23274 9099 23290
rect 8820 23258 9099 23274
rect 8820 23242 8974 23258
rect 8990 23242 9006 23258
rect 9022 23242 9038 23258
rect 9054 23242 9070 23258
rect 9086 23242 9099 23258
rect 8820 23240 9099 23242
rect 8959 23226 9099 23240
rect 8959 23210 8974 23226
rect 8990 23210 9006 23226
rect 9022 23210 9038 23226
rect 9054 23210 9070 23226
rect 9086 23210 9099 23226
rect 8959 23194 9099 23210
rect 8959 23178 8974 23194
rect 8990 23178 9006 23194
rect 9022 23178 9038 23194
rect 9054 23178 9070 23194
rect 9086 23178 9099 23194
rect 8959 23162 9099 23178
rect 8959 23146 8974 23162
rect 8990 23146 9006 23162
rect 9022 23146 9038 23162
rect 9054 23146 9070 23162
rect 9086 23146 9099 23162
rect 8959 23130 9099 23146
rect 8959 23114 8974 23130
rect 8990 23114 9006 23130
rect 9022 23114 9038 23130
rect 9054 23114 9070 23130
rect 9086 23114 9099 23130
rect 8959 23098 9099 23114
rect 8959 23082 8974 23098
rect 8990 23082 9006 23098
rect 9022 23082 9038 23098
rect 9054 23082 9070 23098
rect 9086 23082 9099 23098
rect 8959 23066 9099 23082
rect 8959 23050 8974 23066
rect 8990 23050 9006 23066
rect 9022 23050 9038 23066
rect 9054 23050 9070 23066
rect 9086 23050 9099 23066
rect 8959 23034 9099 23050
rect 8959 23018 8974 23034
rect 8990 23018 9006 23034
rect 9022 23018 9038 23034
rect 9054 23018 9070 23034
rect 9086 23018 9099 23034
rect 8959 23002 9099 23018
rect 8959 22986 8974 23002
rect 8990 22986 9006 23002
rect 9022 22986 9038 23002
rect 9054 22986 9070 23002
rect 9086 22986 9099 23002
rect 8959 22961 9099 22986
rect 8820 20679 9240 20680
rect 8820 20654 9379 20679
rect 8820 20638 9254 20654
rect 9270 20638 9286 20654
rect 9302 20638 9318 20654
rect 9334 20638 9350 20654
rect 9366 20638 9379 20654
rect 8820 20622 9379 20638
rect 8820 20606 9254 20622
rect 9270 20606 9286 20622
rect 9302 20606 9318 20622
rect 9334 20606 9350 20622
rect 9366 20606 9379 20622
rect 8820 20590 9379 20606
rect 8820 20574 9254 20590
rect 9270 20574 9286 20590
rect 9302 20574 9318 20590
rect 9334 20574 9350 20590
rect 9366 20574 9379 20590
rect 8820 20558 9379 20574
rect 8820 20542 9254 20558
rect 9270 20542 9286 20558
rect 9302 20542 9318 20558
rect 9334 20542 9350 20558
rect 9366 20542 9379 20558
rect 8820 20540 9379 20542
rect 9239 20526 9379 20540
rect 9239 20510 9254 20526
rect 9270 20510 9286 20526
rect 9302 20510 9318 20526
rect 9334 20510 9350 20526
rect 9366 20510 9379 20526
rect 9239 20494 9379 20510
rect 9239 20478 9254 20494
rect 9270 20478 9286 20494
rect 9302 20478 9318 20494
rect 9334 20478 9350 20494
rect 9366 20478 9379 20494
rect 9239 20462 9379 20478
rect 9239 20446 9254 20462
rect 9270 20446 9286 20462
rect 9302 20446 9318 20462
rect 9334 20446 9350 20462
rect 9366 20446 9379 20462
rect 9239 20430 9379 20446
rect 9239 20414 9254 20430
rect 9270 20414 9286 20430
rect 9302 20414 9318 20430
rect 9334 20414 9350 20430
rect 9366 20414 9379 20430
rect 9239 20398 9379 20414
rect 9239 20382 9254 20398
rect 9270 20382 9286 20398
rect 9302 20382 9318 20398
rect 9334 20382 9350 20398
rect 9366 20382 9379 20398
rect 9239 20366 9379 20382
rect 9239 20350 9254 20366
rect 9270 20350 9286 20366
rect 9302 20350 9318 20366
rect 9334 20350 9350 20366
rect 9366 20350 9379 20366
rect 9239 20334 9379 20350
rect 9239 20318 9254 20334
rect 9270 20318 9286 20334
rect 9302 20318 9318 20334
rect 9334 20318 9350 20334
rect 9366 20318 9379 20334
rect 9239 20302 9379 20318
rect 9239 20286 9254 20302
rect 9270 20286 9286 20302
rect 9302 20286 9318 20302
rect 9334 20286 9350 20302
rect 9366 20286 9379 20302
rect 9239 20261 9379 20286
rect 9620 17960 9700 24400
rect 8820 17880 9700 17960
rect 9780 15260 9860 25100
rect 8820 15180 9860 15260
rect 9940 12560 10020 25260
rect 8820 12480 10020 12560
rect 10100 9840 10180 25420
rect 27720 16720 27800 28160
rect 27880 25460 29180 25540
rect 27880 18160 27960 25460
rect 28041 23018 28119 23039
rect 28041 23002 28056 23018
rect 28072 23002 28088 23018
rect 28104 23002 28119 23018
rect 28041 22986 28119 23002
rect 28041 22970 28056 22986
rect 28072 22970 28088 22986
rect 28104 22970 28119 22986
rect 28041 22954 28119 22970
rect 28041 22938 28056 22954
rect 28072 22938 28088 22954
rect 28104 22938 28119 22954
rect 28041 22922 28119 22938
rect 28041 22906 28056 22922
rect 28072 22906 28088 22922
rect 28104 22906 28119 22922
rect 28041 22890 28119 22906
rect 28041 22874 28056 22890
rect 28072 22874 28088 22890
rect 28104 22874 28119 22890
rect 28041 22858 28119 22874
rect 28041 22842 28056 22858
rect 28072 22842 28088 22858
rect 28104 22842 28119 22858
rect 28041 22820 28119 22842
rect 28040 22740 29180 22820
rect 28421 20284 28501 20299
rect 28421 20268 28436 20284
rect 28452 20268 28468 20284
rect 28484 20268 28501 20284
rect 28421 20252 28501 20268
rect 28421 20236 28436 20252
rect 28452 20236 28468 20252
rect 28484 20236 28501 20252
rect 28421 20220 28501 20236
rect 28421 20204 28436 20220
rect 28452 20204 28468 20220
rect 28484 20204 28501 20220
rect 28421 20188 28501 20204
rect 28421 20172 28436 20188
rect 28452 20172 28468 20188
rect 28484 20172 28501 20188
rect 28421 20156 28501 20172
rect 28421 20140 28436 20156
rect 28452 20140 28468 20156
rect 28484 20140 28501 20156
rect 28421 20124 29180 20140
rect 28421 20108 28436 20124
rect 28452 20108 28468 20124
rect 28484 20108 29180 20124
rect 28421 20092 29180 20108
rect 28421 20076 28436 20092
rect 28452 20076 28468 20092
rect 28484 20076 29180 20092
rect 28421 20061 29180 20076
rect 28500 20060 29180 20061
rect 27881 18144 27959 18160
rect 27881 18128 27896 18144
rect 27912 18128 27928 18144
rect 27944 18128 27959 18144
rect 27881 18112 27959 18128
rect 27881 18096 27896 18112
rect 27912 18096 27928 18112
rect 27944 18096 27959 18112
rect 27881 18080 27959 18096
rect 27881 18064 27896 18080
rect 27912 18064 27928 18080
rect 27944 18064 27959 18080
rect 27881 18048 27959 18064
rect 27881 18032 27896 18048
rect 27912 18032 27928 18048
rect 27944 18032 27959 18048
rect 27881 18016 27959 18032
rect 27881 18000 27896 18016
rect 27912 18000 27928 18016
rect 27944 18000 27959 18016
rect 27881 17984 27959 18000
rect 27881 17968 27896 17984
rect 27912 17968 27928 17984
rect 27944 17968 27959 17984
rect 27881 17952 27959 17968
rect 27881 17936 27896 17952
rect 27912 17936 27928 17952
rect 27944 17936 27959 17952
rect 27881 17921 27959 17936
rect 28581 17584 28661 17599
rect 28581 17568 28596 17584
rect 28612 17568 28628 17584
rect 28644 17568 28661 17584
rect 28581 17552 28661 17568
rect 28581 17536 28596 17552
rect 28612 17536 28628 17552
rect 28644 17536 28661 17552
rect 28581 17520 28661 17536
rect 28581 17504 28596 17520
rect 28612 17504 28628 17520
rect 28644 17504 28661 17520
rect 28581 17488 28661 17504
rect 28581 17472 28596 17488
rect 28612 17472 28628 17488
rect 28644 17472 28661 17488
rect 28581 17456 28661 17472
rect 28581 17440 28596 17456
rect 28612 17440 28628 17456
rect 28644 17440 28661 17456
rect 28581 17424 29180 17440
rect 28581 17408 28596 17424
rect 28612 17408 28628 17424
rect 28644 17408 29180 17424
rect 28581 17392 29180 17408
rect 28581 17376 28596 17392
rect 28612 17376 28628 17392
rect 28644 17376 29180 17392
rect 28581 17361 29180 17376
rect 28660 17360 29180 17361
rect 27721 16704 27799 16720
rect 27721 16688 27736 16704
rect 27752 16688 27768 16704
rect 27784 16688 27799 16704
rect 27721 16672 27799 16688
rect 27721 16656 27736 16672
rect 27752 16656 27768 16672
rect 27784 16656 27799 16672
rect 27721 16640 27799 16656
rect 27721 16624 27736 16640
rect 27752 16624 27768 16640
rect 27784 16624 27799 16640
rect 27721 16608 27799 16624
rect 27721 16592 27736 16608
rect 27752 16592 27768 16608
rect 27784 16592 27799 16608
rect 27721 16576 27799 16592
rect 27721 16560 27736 16576
rect 27752 16560 27768 16576
rect 27784 16560 27799 16576
rect 27721 16544 27799 16560
rect 27721 16528 27736 16544
rect 27752 16528 27768 16544
rect 27784 16528 27799 16544
rect 27721 16512 27799 16528
rect 27721 16496 27736 16512
rect 27752 16496 27768 16512
rect 27784 16496 27799 16512
rect 27721 16481 27799 16496
rect 28741 14884 28821 14899
rect 28741 14868 28756 14884
rect 28772 14868 28788 14884
rect 28804 14868 28821 14884
rect 28741 14852 28821 14868
rect 28741 14836 28756 14852
rect 28772 14836 28788 14852
rect 28804 14836 28821 14852
rect 28741 14820 28821 14836
rect 28741 14804 28756 14820
rect 28772 14804 28788 14820
rect 28804 14804 28821 14820
rect 28741 14788 28821 14804
rect 28741 14772 28756 14788
rect 28772 14772 28788 14788
rect 28804 14772 28821 14788
rect 28741 14756 28821 14772
rect 28741 14740 28756 14756
rect 28772 14740 28788 14756
rect 28804 14740 28821 14756
rect 28741 14724 29180 14740
rect 28741 14708 28756 14724
rect 28772 14708 28788 14724
rect 28804 14708 29180 14724
rect 28741 14692 29180 14708
rect 28741 14676 28756 14692
rect 28772 14676 28788 14692
rect 28804 14676 29180 14692
rect 28741 14661 29180 14676
rect 28820 14660 29180 14661
rect 28901 12184 28981 12199
rect 28901 12168 28916 12184
rect 28932 12168 28948 12184
rect 28964 12168 28981 12184
rect 28901 12152 28981 12168
rect 28901 12136 28916 12152
rect 28932 12136 28948 12152
rect 28964 12136 28981 12152
rect 28901 12120 28981 12136
rect 28901 12104 28916 12120
rect 28932 12104 28948 12120
rect 28964 12104 28981 12120
rect 28901 12088 28981 12104
rect 28901 12072 28916 12088
rect 28932 12072 28948 12088
rect 28964 12072 28981 12088
rect 28901 12056 28981 12072
rect 28901 12040 28916 12056
rect 28932 12040 28948 12056
rect 28964 12040 28981 12056
rect 28901 12024 29180 12040
rect 28901 12008 28916 12024
rect 28932 12008 28948 12024
rect 28964 12008 29180 12024
rect 28901 11992 29180 12008
rect 28901 11976 28916 11992
rect 28932 11976 28948 11992
rect 28964 11976 29180 11992
rect 28901 11961 29180 11976
rect 28980 11960 29180 11961
rect 11750 10550 11830 11780
rect 11890 10770 11950 11780
rect 12000 11740 12160 11780
rect 12060 10980 12160 11740
rect 12780 11180 12880 11780
rect 20280 11380 20380 11780
rect 22740 11580 22840 11780
rect 22740 11480 25540 11580
rect 20280 11280 22840 11380
rect 12780 11080 20140 11180
rect 12060 10880 17440 10980
rect 11890 10660 14740 10770
rect 11750 10440 12040 10550
rect 8820 9760 10180 9840
rect 11940 8820 12040 10440
rect 14640 8820 14740 10660
rect 17340 8820 17440 10880
rect 20040 8820 20140 11080
rect 22740 8820 22840 11280
rect 25440 8820 25540 11480
rect 25960 9200 26060 11780
rect 25960 9100 28240 9200
rect 28140 8820 28240 9100
<< m3contact >>
rect 17894 27238 17910 27254
rect 17926 27238 17942 27254
rect 17958 27238 17974 27254
rect 17990 27238 18006 27254
rect 18022 27238 18038 27254
rect 18054 27238 18070 27254
rect 18086 27238 18102 27254
rect 18118 27238 18134 27254
rect 18150 27238 18166 27254
rect 17894 27206 17910 27222
rect 17926 27206 17942 27222
rect 17958 27206 17974 27222
rect 17990 27206 18006 27222
rect 18022 27206 18038 27222
rect 18054 27206 18070 27222
rect 18086 27206 18102 27222
rect 18118 27206 18134 27222
rect 18150 27206 18166 27222
rect 24314 27238 24330 27254
rect 24346 27238 24362 27254
rect 24378 27238 24394 27254
rect 24410 27238 24426 27254
rect 24442 27238 24458 27254
rect 24474 27238 24490 27254
rect 24506 27238 24522 27254
rect 24538 27238 24554 27254
rect 24570 27238 24586 27254
rect 24314 27206 24330 27222
rect 24346 27206 24362 27222
rect 24378 27206 24394 27222
rect 24410 27206 24426 27222
rect 24442 27206 24458 27222
rect 24474 27206 24490 27222
rect 24506 27206 24522 27222
rect 24538 27206 24554 27222
rect 24570 27206 24586 27222
rect 10116 25468 10132 25484
rect 10148 25468 10164 25484
rect 10116 25436 10132 25452
rect 10148 25436 10164 25452
rect 9956 25308 9972 25324
rect 9988 25308 10004 25324
rect 9956 25276 9972 25292
rect 9988 25276 10004 25292
rect 9796 25148 9812 25164
rect 9828 25148 9844 25164
rect 9796 25116 9812 25132
rect 9828 25116 9844 25132
rect 9636 24448 9652 24464
rect 9668 24448 9684 24464
rect 9636 24416 9652 24432
rect 9668 24416 9684 24432
rect 8974 23338 8990 23354
rect 9006 23338 9022 23354
rect 9038 23338 9054 23354
rect 9070 23338 9086 23354
rect 8974 23306 8990 23322
rect 9006 23306 9022 23322
rect 9038 23306 9054 23322
rect 9070 23306 9086 23322
rect 8974 23274 8990 23290
rect 9006 23274 9022 23290
rect 9038 23274 9054 23290
rect 9070 23274 9086 23290
rect 8974 23242 8990 23258
rect 9006 23242 9022 23258
rect 9038 23242 9054 23258
rect 9070 23242 9086 23258
rect 8974 23210 8990 23226
rect 9006 23210 9022 23226
rect 9038 23210 9054 23226
rect 9070 23210 9086 23226
rect 8974 23178 8990 23194
rect 9006 23178 9022 23194
rect 9038 23178 9054 23194
rect 9070 23178 9086 23194
rect 8974 23146 8990 23162
rect 9006 23146 9022 23162
rect 9038 23146 9054 23162
rect 9070 23146 9086 23162
rect 8974 23114 8990 23130
rect 9006 23114 9022 23130
rect 9038 23114 9054 23130
rect 9070 23114 9086 23130
rect 8974 23082 8990 23098
rect 9006 23082 9022 23098
rect 9038 23082 9054 23098
rect 9070 23082 9086 23098
rect 8974 23050 8990 23066
rect 9006 23050 9022 23066
rect 9038 23050 9054 23066
rect 9070 23050 9086 23066
rect 8974 23018 8990 23034
rect 9006 23018 9022 23034
rect 9038 23018 9054 23034
rect 9070 23018 9086 23034
rect 8974 22986 8990 23002
rect 9006 22986 9022 23002
rect 9038 22986 9054 23002
rect 9070 22986 9086 23002
rect 9254 20638 9270 20654
rect 9286 20638 9302 20654
rect 9318 20638 9334 20654
rect 9350 20638 9366 20654
rect 9254 20606 9270 20622
rect 9286 20606 9302 20622
rect 9318 20606 9334 20622
rect 9350 20606 9366 20622
rect 9254 20574 9270 20590
rect 9286 20574 9302 20590
rect 9318 20574 9334 20590
rect 9350 20574 9366 20590
rect 9254 20542 9270 20558
rect 9286 20542 9302 20558
rect 9318 20542 9334 20558
rect 9350 20542 9366 20558
rect 9254 20510 9270 20526
rect 9286 20510 9302 20526
rect 9318 20510 9334 20526
rect 9350 20510 9366 20526
rect 9254 20478 9270 20494
rect 9286 20478 9302 20494
rect 9318 20478 9334 20494
rect 9350 20478 9366 20494
rect 9254 20446 9270 20462
rect 9286 20446 9302 20462
rect 9318 20446 9334 20462
rect 9350 20446 9366 20462
rect 9254 20414 9270 20430
rect 9286 20414 9302 20430
rect 9318 20414 9334 20430
rect 9350 20414 9366 20430
rect 9254 20382 9270 20398
rect 9286 20382 9302 20398
rect 9318 20382 9334 20398
rect 9350 20382 9366 20398
rect 9254 20350 9270 20366
rect 9286 20350 9302 20366
rect 9318 20350 9334 20366
rect 9350 20350 9366 20366
rect 9254 20318 9270 20334
rect 9286 20318 9302 20334
rect 9318 20318 9334 20334
rect 9350 20318 9366 20334
rect 9254 20286 9270 20302
rect 9286 20286 9302 20302
rect 9318 20286 9334 20302
rect 9350 20286 9366 20302
rect 28056 23002 28072 23018
rect 28088 23002 28104 23018
rect 28056 22970 28072 22986
rect 28088 22970 28104 22986
rect 28056 22938 28072 22954
rect 28088 22938 28104 22954
rect 28056 22906 28072 22922
rect 28088 22906 28104 22922
rect 28056 22874 28072 22890
rect 28088 22874 28104 22890
rect 28056 22842 28072 22858
rect 28088 22842 28104 22858
rect 28436 20268 28452 20284
rect 28468 20268 28484 20284
rect 28436 20236 28452 20252
rect 28468 20236 28484 20252
rect 28436 20204 28452 20220
rect 28468 20204 28484 20220
rect 28436 20172 28452 20188
rect 28468 20172 28484 20188
rect 28436 20140 28452 20156
rect 28468 20140 28484 20156
rect 28436 20108 28452 20124
rect 28468 20108 28484 20124
rect 28436 20076 28452 20092
rect 28468 20076 28484 20092
rect 27896 18128 27912 18144
rect 27928 18128 27944 18144
rect 27896 18096 27912 18112
rect 27928 18096 27944 18112
rect 27896 18064 27912 18080
rect 27928 18064 27944 18080
rect 27896 18032 27912 18048
rect 27928 18032 27944 18048
rect 27896 18000 27912 18016
rect 27928 18000 27944 18016
rect 27896 17968 27912 17984
rect 27928 17968 27944 17984
rect 27896 17936 27912 17952
rect 27928 17936 27944 17952
rect 28596 17568 28612 17584
rect 28628 17568 28644 17584
rect 28596 17536 28612 17552
rect 28628 17536 28644 17552
rect 28596 17504 28612 17520
rect 28628 17504 28644 17520
rect 28596 17472 28612 17488
rect 28628 17472 28644 17488
rect 28596 17440 28612 17456
rect 28628 17440 28644 17456
rect 28596 17408 28612 17424
rect 28628 17408 28644 17424
rect 28596 17376 28612 17392
rect 28628 17376 28644 17392
rect 27736 16688 27752 16704
rect 27768 16688 27784 16704
rect 27736 16656 27752 16672
rect 27768 16656 27784 16672
rect 27736 16624 27752 16640
rect 27768 16624 27784 16640
rect 27736 16592 27752 16608
rect 27768 16592 27784 16608
rect 27736 16560 27752 16576
rect 27768 16560 27784 16576
rect 27736 16528 27752 16544
rect 27768 16528 27784 16544
rect 27736 16496 27752 16512
rect 27768 16496 27784 16512
rect 28756 14868 28772 14884
rect 28788 14868 28804 14884
rect 28756 14836 28772 14852
rect 28788 14836 28804 14852
rect 28756 14804 28772 14820
rect 28788 14804 28804 14820
rect 28756 14772 28772 14788
rect 28788 14772 28804 14788
rect 28756 14740 28772 14756
rect 28788 14740 28804 14756
rect 28756 14708 28772 14724
rect 28788 14708 28804 14724
rect 28756 14676 28772 14692
rect 28788 14676 28804 14692
rect 28916 12168 28932 12184
rect 28948 12168 28964 12184
rect 28916 12136 28932 12152
rect 28948 12136 28964 12152
rect 28916 12104 28932 12120
rect 28948 12104 28964 12120
rect 28916 12072 28932 12088
rect 28948 12072 28964 12088
rect 28916 12040 28932 12056
rect 28948 12040 28964 12056
rect 28916 12008 28932 12024
rect 28948 12008 28964 12024
rect 28916 11976 28932 11992
rect 28948 11976 28964 11992
<< metal3 >>
rect 18180 27279 24300 27280
rect 17881 27254 24599 27279
rect 17881 27238 17894 27254
rect 17910 27238 17926 27254
rect 17942 27238 17958 27254
rect 17974 27238 17990 27254
rect 18006 27238 18022 27254
rect 18038 27238 18054 27254
rect 18070 27238 18086 27254
rect 18102 27238 18118 27254
rect 18134 27238 18150 27254
rect 18166 27238 24314 27254
rect 24330 27238 24346 27254
rect 24362 27238 24378 27254
rect 24394 27238 24410 27254
rect 24426 27238 24442 27254
rect 24458 27238 24474 27254
rect 24490 27238 24506 27254
rect 24522 27238 24538 27254
rect 24554 27238 24570 27254
rect 24586 27238 24599 27254
rect 17881 27222 24599 27238
rect 17881 27206 17894 27222
rect 17910 27206 17926 27222
rect 17942 27206 17958 27222
rect 17974 27206 17990 27222
rect 18006 27206 18022 27222
rect 18038 27206 18054 27222
rect 18070 27206 18086 27222
rect 18102 27206 18118 27222
rect 18134 27206 18150 27222
rect 18166 27206 24314 27222
rect 24330 27206 24346 27222
rect 24362 27206 24378 27222
rect 24394 27206 24410 27222
rect 24426 27206 24442 27222
rect 24458 27206 24474 27222
rect 24490 27206 24506 27222
rect 24522 27206 24538 27222
rect 24554 27206 24570 27222
rect 24586 27206 24599 27222
rect 17881 27181 24599 27206
rect 18180 27180 24300 27181
rect 26740 26200 28980 26280
rect 26740 26060 28820 26140
rect 26740 25920 28660 26000
rect 26740 25780 28500 25860
rect 10180 25499 11280 25500
rect 10101 25484 11280 25499
rect 10101 25468 10116 25484
rect 10132 25468 10148 25484
rect 10164 25468 11280 25484
rect 10101 25452 11280 25468
rect 10101 25436 10116 25452
rect 10132 25436 10148 25452
rect 10164 25436 11280 25452
rect 10101 25421 11280 25436
rect 10180 25420 11280 25421
rect 10020 25339 11280 25340
rect 9941 25324 11280 25339
rect 9941 25308 9956 25324
rect 9972 25308 9988 25324
rect 10004 25308 11280 25324
rect 9941 25292 11280 25308
rect 9941 25276 9956 25292
rect 9972 25276 9988 25292
rect 10004 25276 11280 25292
rect 9941 25261 11280 25276
rect 10020 25260 11280 25261
rect 9860 25179 11280 25180
rect 9781 25164 11280 25179
rect 9781 25148 9796 25164
rect 9812 25148 9828 25164
rect 9844 25148 11280 25164
rect 9781 25132 11280 25148
rect 9781 25116 9796 25132
rect 9812 25116 9828 25132
rect 9844 25116 11280 25132
rect 9781 25101 11280 25116
rect 9860 25100 11280 25101
rect 9700 24479 11280 24480
rect 9621 24464 11280 24479
rect 9621 24448 9636 24464
rect 9652 24448 9668 24464
rect 9684 24448 11280 24464
rect 9621 24432 11280 24448
rect 9621 24416 9636 24432
rect 9652 24416 9668 24432
rect 9684 24416 11280 24432
rect 9621 24401 11280 24416
rect 9700 24400 11280 24401
rect 8961 23354 9099 23379
rect 8961 23338 8974 23354
rect 8990 23338 9006 23354
rect 9022 23338 9038 23354
rect 9054 23338 9070 23354
rect 9086 23338 9099 23354
rect 8961 23322 9099 23338
rect 8961 23306 8974 23322
rect 8990 23306 9006 23322
rect 9022 23306 9038 23322
rect 9054 23306 9070 23322
rect 9086 23306 9099 23322
rect 8961 23290 9099 23306
rect 8961 23274 8974 23290
rect 8990 23274 9006 23290
rect 9022 23274 9038 23290
rect 9054 23274 9070 23290
rect 9086 23274 9099 23290
rect 8961 23258 9099 23274
rect 8961 23242 8974 23258
rect 8990 23242 9006 23258
rect 9022 23242 9038 23258
rect 9054 23242 9070 23258
rect 9086 23242 9099 23258
rect 8961 23226 9099 23242
rect 8961 23210 8974 23226
rect 8990 23210 9006 23226
rect 9022 23210 9038 23226
rect 9054 23210 9070 23226
rect 9086 23210 9099 23226
rect 8961 23194 9099 23210
rect 8961 23178 8974 23194
rect 8990 23178 9006 23194
rect 9022 23178 9038 23194
rect 9054 23178 9070 23194
rect 9086 23178 9099 23194
rect 8961 23162 9099 23178
rect 8961 23146 8974 23162
rect 8990 23146 9006 23162
rect 9022 23146 9038 23162
rect 9054 23146 9070 23162
rect 9086 23146 9099 23162
rect 8961 23130 9099 23146
rect 8961 23114 8974 23130
rect 8990 23114 9006 23130
rect 9022 23114 9038 23130
rect 9054 23114 9070 23130
rect 9086 23114 9099 23130
rect 8961 23098 9099 23114
rect 8961 23082 8974 23098
rect 8990 23082 9006 23098
rect 9022 23082 9038 23098
rect 9054 23082 9070 23098
rect 9086 23082 9099 23098
rect 8961 23066 9099 23082
rect 8961 23050 8974 23066
rect 8990 23050 9006 23066
rect 9022 23050 9038 23066
rect 9054 23050 9070 23066
rect 9086 23050 9099 23066
rect 8961 23034 9099 23050
rect 8961 23018 8974 23034
rect 8990 23018 9006 23034
rect 9022 23018 9038 23034
rect 9054 23018 9070 23034
rect 9086 23018 9099 23034
rect 8961 23002 9099 23018
rect 8961 22986 8974 23002
rect 8990 22986 9006 23002
rect 9022 22986 9038 23002
rect 9054 22986 9070 23002
rect 9086 22986 9099 23002
rect 8961 22960 9099 22986
rect 26740 23039 28040 23040
rect 26740 23018 28119 23039
rect 26740 23002 28056 23018
rect 28072 23002 28088 23018
rect 28104 23002 28119 23018
rect 26740 22986 28119 23002
rect 26740 22970 28056 22986
rect 28072 22970 28088 22986
rect 28104 22970 28119 22986
rect 26740 22960 28119 22970
rect 8960 18760 9100 22960
rect 28040 22954 28119 22960
rect 28040 22938 28056 22954
rect 28072 22938 28088 22954
rect 28104 22938 28119 22954
rect 28040 22922 28119 22938
rect 28040 22906 28056 22922
rect 28072 22906 28088 22922
rect 28104 22906 28119 22922
rect 28040 22890 28119 22906
rect 28040 22874 28056 22890
rect 28072 22874 28088 22890
rect 28104 22874 28119 22890
rect 28040 22858 28119 22874
rect 28040 22842 28056 22858
rect 28072 22842 28088 22858
rect 28104 22842 28119 22858
rect 28040 22821 28119 22842
rect 9241 20654 9379 20679
rect 9241 20638 9254 20654
rect 9270 20638 9286 20654
rect 9302 20638 9318 20654
rect 9334 20638 9350 20654
rect 9366 20638 9379 20654
rect 9241 20622 9379 20638
rect 9241 20606 9254 20622
rect 9270 20606 9286 20622
rect 9302 20606 9318 20622
rect 9334 20606 9350 20622
rect 9366 20606 9379 20622
rect 9241 20590 9379 20606
rect 9241 20574 9254 20590
rect 9270 20574 9286 20590
rect 9302 20574 9318 20590
rect 9334 20574 9350 20590
rect 9366 20574 9379 20590
rect 9241 20558 9379 20574
rect 9241 20542 9254 20558
rect 9270 20542 9286 20558
rect 9302 20542 9318 20558
rect 9334 20542 9350 20558
rect 9366 20542 9379 20558
rect 9241 20526 9379 20542
rect 9241 20510 9254 20526
rect 9270 20510 9286 20526
rect 9302 20510 9318 20526
rect 9334 20510 9350 20526
rect 9366 20510 9379 20526
rect 9241 20494 9379 20510
rect 9241 20478 9254 20494
rect 9270 20478 9286 20494
rect 9302 20478 9318 20494
rect 9334 20478 9350 20494
rect 9366 20478 9379 20494
rect 9241 20462 9379 20478
rect 9241 20446 9254 20462
rect 9270 20446 9286 20462
rect 9302 20446 9318 20462
rect 9334 20446 9350 20462
rect 9366 20446 9379 20462
rect 9241 20430 9379 20446
rect 9241 20414 9254 20430
rect 9270 20414 9286 20430
rect 9302 20414 9318 20430
rect 9334 20414 9350 20430
rect 9366 20414 9379 20430
rect 9241 20398 9379 20414
rect 9241 20382 9254 20398
rect 9270 20382 9286 20398
rect 9302 20382 9318 20398
rect 9334 20382 9350 20398
rect 9366 20382 9379 20398
rect 9241 20366 9379 20382
rect 9241 20350 9254 20366
rect 9270 20350 9286 20366
rect 9302 20350 9318 20366
rect 9334 20350 9350 20366
rect 9366 20350 9379 20366
rect 9241 20334 9379 20350
rect 9241 20318 9254 20334
rect 9270 20318 9286 20334
rect 9302 20318 9318 20334
rect 9334 20318 9350 20334
rect 9366 20318 9379 20334
rect 9241 20302 9379 20318
rect 9241 20286 9254 20302
rect 9270 20286 9286 20302
rect 9302 20286 9318 20302
rect 9334 20286 9350 20302
rect 9366 20286 9379 20302
rect 28420 20300 28500 25780
rect 9241 20260 9379 20286
rect 28421 20284 28499 20300
rect 28421 20268 28436 20284
rect 28452 20268 28468 20284
rect 28484 20268 28499 20284
rect 9240 19040 9380 20260
rect 28421 20252 28499 20268
rect 28421 20236 28436 20252
rect 28452 20236 28468 20252
rect 28484 20236 28499 20252
rect 28421 20220 28499 20236
rect 28421 20204 28436 20220
rect 28452 20204 28468 20220
rect 28484 20204 28499 20220
rect 28421 20188 28499 20204
rect 28421 20172 28436 20188
rect 28452 20172 28468 20188
rect 28484 20172 28499 20188
rect 28421 20156 28499 20172
rect 28421 20140 28436 20156
rect 28452 20140 28468 20156
rect 28484 20140 28499 20156
rect 28421 20124 28499 20140
rect 28421 20108 28436 20124
rect 28452 20108 28468 20124
rect 28484 20108 28499 20124
rect 28421 20092 28499 20108
rect 28421 20076 28436 20092
rect 28452 20076 28468 20092
rect 28484 20076 28499 20092
rect 28421 20061 28499 20076
rect 9240 18900 11300 19040
rect 11160 18820 11300 18900
rect 8960 18620 11300 18760
rect 27880 18144 27959 18159
rect 27880 18128 27896 18144
rect 27912 18128 27928 18144
rect 27944 18128 27959 18144
rect 27880 18112 27959 18128
rect 27880 18096 27896 18112
rect 27912 18096 27928 18112
rect 27944 18096 27959 18112
rect 27880 18080 27959 18096
rect 27880 18064 27896 18080
rect 27912 18064 27928 18080
rect 27944 18064 27959 18080
rect 27880 18048 27959 18064
rect 27880 18032 27896 18048
rect 27912 18032 27928 18048
rect 27944 18032 27959 18048
rect 27880 18016 27959 18032
rect 27880 18000 27896 18016
rect 27912 18000 27928 18016
rect 27944 18000 27959 18016
rect 26740 17984 27959 18000
rect 26740 17968 27896 17984
rect 27912 17968 27928 17984
rect 27944 17968 27959 17984
rect 26740 17952 27959 17968
rect 26740 17936 27896 17952
rect 27912 17936 27928 17952
rect 27944 17936 27959 17952
rect 26740 17921 27959 17936
rect 26740 17920 27880 17921
rect 28580 17600 28660 25920
rect 28581 17584 28659 17600
rect 28581 17568 28596 17584
rect 28612 17568 28628 17584
rect 28644 17568 28659 17584
rect 28581 17552 28659 17568
rect 28581 17536 28596 17552
rect 28612 17536 28628 17552
rect 28644 17536 28659 17552
rect 28581 17520 28659 17536
rect 28581 17504 28596 17520
rect 28612 17504 28628 17520
rect 28644 17504 28659 17520
rect 28581 17488 28659 17504
rect 28581 17472 28596 17488
rect 28612 17472 28628 17488
rect 28644 17472 28659 17488
rect 28581 17456 28659 17472
rect 28581 17440 28596 17456
rect 28612 17440 28628 17456
rect 28644 17440 28659 17456
rect 28581 17424 28659 17440
rect 28581 17408 28596 17424
rect 28612 17408 28628 17424
rect 28644 17408 28659 17424
rect 28581 17392 28659 17408
rect 28581 17376 28596 17392
rect 28612 17376 28628 17392
rect 28644 17376 28659 17392
rect 28581 17361 28659 17376
rect 27720 16704 27799 16719
rect 27720 16688 27736 16704
rect 27752 16688 27768 16704
rect 27784 16688 27799 16704
rect 27720 16672 27799 16688
rect 27720 16656 27736 16672
rect 27752 16656 27768 16672
rect 27784 16656 27799 16672
rect 27720 16640 27799 16656
rect 27720 16624 27736 16640
rect 27752 16624 27768 16640
rect 27784 16624 27799 16640
rect 27720 16608 27799 16624
rect 27720 16592 27736 16608
rect 27752 16592 27768 16608
rect 27784 16592 27799 16608
rect 27720 16576 27799 16592
rect 27720 16560 27736 16576
rect 27752 16560 27768 16576
rect 27784 16560 27799 16576
rect 26740 16544 27799 16560
rect 26740 16528 27736 16544
rect 27752 16528 27768 16544
rect 27784 16528 27799 16544
rect 26740 16512 27799 16528
rect 26740 16496 27736 16512
rect 27752 16496 27768 16512
rect 27784 16496 27799 16512
rect 26740 16481 27799 16496
rect 26740 16480 27720 16481
rect 28740 14900 28820 26060
rect 28741 14884 28819 14900
rect 28741 14868 28756 14884
rect 28772 14868 28788 14884
rect 28804 14868 28819 14884
rect 28741 14852 28819 14868
rect 28741 14836 28756 14852
rect 28772 14836 28788 14852
rect 28804 14836 28819 14852
rect 28741 14820 28819 14836
rect 28741 14804 28756 14820
rect 28772 14804 28788 14820
rect 28804 14804 28819 14820
rect 28741 14788 28819 14804
rect 28741 14772 28756 14788
rect 28772 14772 28788 14788
rect 28804 14772 28819 14788
rect 28741 14756 28819 14772
rect 28741 14740 28756 14756
rect 28772 14740 28788 14756
rect 28804 14740 28819 14756
rect 28741 14724 28819 14740
rect 28741 14708 28756 14724
rect 28772 14708 28788 14724
rect 28804 14708 28819 14724
rect 28741 14692 28819 14708
rect 28741 14676 28756 14692
rect 28772 14676 28788 14692
rect 28804 14676 28819 14692
rect 28741 14661 28819 14676
rect 28900 12200 28980 26200
rect 28901 12184 28979 12200
rect 28901 12168 28916 12184
rect 28932 12168 28948 12184
rect 28964 12168 28979 12184
rect 28901 12152 28979 12168
rect 28901 12136 28916 12152
rect 28932 12136 28948 12152
rect 28964 12136 28979 12152
rect 28901 12120 28979 12136
rect 28901 12104 28916 12120
rect 28932 12104 28948 12120
rect 28964 12104 28979 12120
rect 28901 12088 28979 12104
rect 28901 12072 28916 12088
rect 28932 12072 28948 12088
rect 28964 12072 28979 12088
rect 28901 12056 28979 12072
rect 28901 12040 28916 12056
rect 28932 12040 28948 12056
rect 28964 12040 28979 12056
rect 28901 12024 28979 12040
rect 28901 12008 28916 12024
rect 28932 12008 28948 12024
rect 28964 12008 28979 12024
rect 28901 11992 28979 12008
rect 28901 11976 28916 11992
rect 28932 11976 28948 11992
rect 28964 11976 28979 11992
rect 28901 11961 28979 11976
<< end >>
