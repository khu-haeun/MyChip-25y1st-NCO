/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module nco(
    inout vdd,
    inout gnd,
    output [11:0] Dout,
    input En,
    input [19:0] FCW,
    output Vld,
    input clk,
    input selSign,
    input selXY
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire \genblk1[0].u_ce.Vld_bF$buf4  ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire [1:0] \a[5]  ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire \genblk1[2].u_ce.Vld_bF$buf0  ;
wire [1:0] \genblk1[2].u_ce.Y_  ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _7004_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire \u_ot.ISreg_bF$buf3  ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire [1:0] \genblk1[5].u_ce.Yin0  ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _7042_ ;
wire _6833__bF$buf0 ;
wire _6833__bF$buf1 ;
wire _6833__bF$buf2 ;
wire _6833__bF$buf3 ;
wire _6833__bF$buf4 ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6771_ ;
wire _6351_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf1  ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf2  ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire [1:0] \genblk1[2].u_ce.Xin1  ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire \genblk1[0].u_ce.Vld_bF$buf1  ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7001_ ;
wire [11:0] \u_pa.Atmp  ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire \u_ot.ISreg_bF$buf0  ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire \genblk1[2].u_ce.ISout  ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire [11:0] \genblk1[5].u_ce.Xcalc  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6956_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _1834__bF$buf0 ;
wire _1834__bF$buf1 ;
wire _1834__bF$buf2 ;
wire _1834__bF$buf3 ;
wire _1834__bF$buf4 ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf2  ;
wire _4925_ ;
wire _4505_ ;
wire \genblk1[5].u_ce.Vld_bF$buf2  ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _3524__bF$buf0 ;
wire _3524__bF$buf1 ;
wire _3524__bF$buf2 ;
wire _3524__bF$buf3 ;
wire _3524__bF$buf4 ;
wire _3524__bF$buf5 ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5151__bF$buf0 ;
wire _5151__bF$buf1 ;
wire _5151__bF$buf2 ;
wire _5151__bF$buf3 ;
wire _5748_ ;
wire _5151__bF$buf4 ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _197_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf1  ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire \u_ot.ISreg  ;
wire _6821_ ;
wire _6401_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire [11:0] \u_ot.Xcalc  ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire [1:0] \genblk1[0].u_ce.Ain1  ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire [1:0] \genblk1[3].u_ce.Y_  ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf2  ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _7033_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf3  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire [11:4] \genblk1[0].u_ce.Yin12b  ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire [1:0] \genblk1[1].u_ce.Xin0  ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire [11:0] _7071_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _158__bF$buf0 ;
wire _158__bF$buf1 ;
wire _158__bF$buf2 ;
wire _158__bF$buf3 ;
wire _158__bF$buf4 ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire [11:4] \genblk1[2].u_ce.Yin12b  ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire \genblk1[2].u_ce.Vld  ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _7068_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire [11:4] \genblk1[4].u_ce.Yin12b  ;
wire _1054_ ;
wire _385_ ;
wire [1:0] \a[0]  ;
wire _2679_ ;
wire _2259_ ;
wire [1:0] \genblk1[3].u_ce.Yin1  ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire [1:0] \genblk1[6].u_ce.Ain0  ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire [11:4] \u_ot.Yin12b  ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire [11:4] \genblk1[6].u_ce.Yin12b  ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _4348__bF$buf0 ;
wire _4348__bF$buf1 ;
wire _4348__bF$buf2 ;
wire _4348__bF$buf3 ;
wire _4348__bF$buf4 ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _6912_ ;
wire _2832_ ;
wire _2412_ ;
wire [11:0] \genblk1[7].u_ce.Ycalc  ;
wire _3617_ ;
wire _6089_ ;
wire _7030_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf0  ;
wire _6721_ ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire En_bF$buf0 ;
wire En_bF$buf1 ;
wire En_bF$buf2 ;
wire En_bF$buf3 ;
wire En_bF$buf4 ;
wire _5704_ ;
wire \genblk1[3].u_ce.Vld_bF$buf2  ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _973__bF$buf0 ;
wire _973__bF$buf1 ;
wire _973__bF$buf2 ;
wire _973__bF$buf3 ;
wire _973__bF$buf4 ;
wire _6718_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf1  ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _7065_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire [11:0] \genblk1[2].u_ce.Xcalc  ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire \genblk1[7].u_ce.Vld  ;
wire _896_ ;
wire _476_ ;
wire [5:0] \genblk1[1].u_ce.LoadCtl  ;
wire _3711_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf2  ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire [1:0] \genblk1[6].u_ce.Xin1  ;
wire _5683_ ;
wire _5263_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf3  ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _6812_ ;
wire _2732_ ;
wire _2312_ ;
wire \genblk1[1].u_ce.Vld_bF$buf3  ;
wire _3937_ ;
wire _3517_ ;
wire [1:1] \a[7]  ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire [1:0] \genblk1[4].u_ce.Y_  ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _39_ ;
wire _6906_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _7024_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _2649__bF$buf0 ;
wire _2649__bF$buf1 ;
wire _2649__bF$buf2 ;
wire _2649__bF$buf3 ;
wire _2649__bF$buf4 ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire \genblk1[6].u_ce.ISout  ;
wire _3649_ ;
wire _3229_ ;
wire _7062_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire [1:0] \genblk1[2].u_ce.Yin0  ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _172__bF$buf0 ;
wire _172__bF$buf1 ;
wire _172__bF$buf2 ;
wire _172__bF$buf3 ;
wire _172__bF$buf4 ;
wire _2958_ ;
wire _172__bF$buf5 ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire [5:0] \u_pa.RdyCtl  ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf0  ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _7059_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _2672__bF$buf0 ;
wire _2672__bF$buf1 ;
wire _2672__bF$buf2 ;
wire _2672__bF$buf3 ;
wire _2672__bF$buf4 ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire selXY ;
wire _4625_ ;
wire _4205_ ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire \genblk1[1].u_ce.Vld_bF$buf0  ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire selSign ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf3  ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _6903_ ;
wire _4090_ ;
wire _4362__bF$buf0 ;
wire _2823_ ;
wire _4362__bF$buf1 ;
wire _2403_ ;
wire _4362__bF$buf2 ;
wire _4362__bF$buf3 ;
wire _4362__bF$buf4 ;
wire _4362__bF$buf5 ;
wire _5295_ ;
wire _3608_ ;
wire _7021_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf2  ;
wire _5601_ ;
wire [1:0] \genblk1[4].u_ce.Ain1  ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire [11:0] \genblk1[4].u_ce.Ycalc  ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf3  ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire [1:0] \genblk1[5].u_ce.Xin0  ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire [11:0] \genblk1[5].u_ce.Acalc  ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7056_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire \genblk1[0].u_ce.Vld  ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf0  ;
wire \genblk1[6].u_ce.Vld_bF$buf1  ;
wire [1:0] \genblk1[7].u_ce.Yin1  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _6900_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire [1:0] \u_ot.Yin1  ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _6803_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf0  ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire [1:0] \genblk1[5].u_ce.Y_  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _7053_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire [11:4] \genblk1[1].u_ce.Yin12b  ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \u_ot.LoadCtl_6_bF$buf4  ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf3  ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire \genblk1[4].u_ce.Vld_bF$buf2  ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire \genblk1[3].u_ce.ISout  ;
wire _4713_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire [11:0] \genblk1[6].u_ce.Xcalc  ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire En ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf2  ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire [1:0] \a[2]  ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire \genblk1[5].u_ce.Vld  ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire _2088_ ;
wire _5174__bF$buf0 ;
wire _5174__bF$buf1 ;
wire _5174__bF$buf2 ;
wire _5174__bF$buf3 ;
wire _5174__bF$buf4 ;
wire [1:0] \genblk1[0].u_ce.Yin1  ;
wire \genblk1[0].u_ce.Rdy_bF$buf2  ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire [1:0] \genblk1[3].u_ce.Ain0  ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire [1:0] \genblk1[0].u_ce.X_  ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf3  ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _7012_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf4  ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _7050_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire \u_ot.LoadCtl_6_bF$buf1  ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf0  ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire [5:0] \genblk1[3].u_ce.LoadCtl  ;
wire _690_ ;
wire _270_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _6929_ ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire [1:0] \genblk1[6].u_ce.Yin0  ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _7047_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire [11:0] \genblk1[1].u_ce.Ycalc  ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _3487__bF$buf0 ;
wire _3487__bF$buf1 ;
wire _3487__bF$buf2 ;
wire _3487__bF$buf3 ;
wire _3487__bF$buf4 ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf0  ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf1  ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _1679_ ;
wire _1259_ ;
wire [1:0] \genblk1[3].u_ce.Xin1  ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _6603_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire \genblk1[2].u_ce.Vld_bF$buf2  ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire [11:4] \genblk1[6].u_ce.Ain12b  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire [1:0] \genblk1[6].u_ce.Y_  ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _7044_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _6773_ ;
wire _6353_ ;
wire _2693_ ;
wire _2273_ ;
wire _996__bF$buf0 ;
wire _996__bF$buf1 ;
wire _996__bF$buf2 ;
wire _996__bF$buf3 ;
wire _3898_ ;
wire _996__bF$buf4 ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf3  ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire [11:0] Dout ;
wire _5909_ ;
wire _3096_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf4  ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire \genblk1[0].u_ce.ISout  ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire \genblk1[0].u_ce.Vld_bF$buf3  ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire [11:0] \genblk1[3].u_ce.Xcalc  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire [1:0] \genblk1[1].u_ce.X_  ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7003_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire \u_ot.ISreg_bF$buf2  ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _7041_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf0  ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire [1:0] \genblk1[1].u_ce.Ain1  ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf1  ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire \genblk1[7].u_ce.ISout  ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire [1:0] \genblk1[2].u_ce.Xin0  ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire \genblk1[0].u_ce.Vld_bF$buf0  ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf4  ;
wire _4927_ ;
wire _4507_ ;
wire \genblk1[5].u_ce.Vld_bF$buf4  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7000_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire [7:0] \genblk1  ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire [1:0] \genblk1[4].u_ce.Yin1  ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire \genblk1[3].u_ce.Vld  ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _199_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf3  ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _6823_ ;
wire _6403_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire [1:0] \genblk1[7].u_ce.Y_  ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire [11:0] \genblk1[5].u_ce.Ycalc  ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf1  ;
wire _4924_ ;
wire _4504_ ;
wire \genblk1[5].u_ce.Vld_bF$buf1  ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire [11:1] \genblk1[6].u_ce.Acalc  ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _1810__bF$buf0 ;
wire _1810__bF$buf1 ;
wire _1810__bF$buf2 ;
wire _1810__bF$buf3 ;
wire _1810__bF$buf4 ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire [5:0] \genblk1[0].u_ce.LoadCtl  ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _196_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf0  ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire [1:0] \a[4]  ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire [19:0] \u_pa.acc_reg  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire [1:0] \genblk1[2].u_ce.X_  ;
wire [1:0] \genblk1[7].u_ce.Xin1  ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire [1:0] \genblk1[0].u_ce.Ain0  ;
wire _1188_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf1  ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire [5:0] \genblk1[5].u_ce.LoadCtl  ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _6914_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire [11:0] \genblk1[0].u_ce.Xcalc  ;
wire _7032_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf2  ;
wire _6723_ ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire [1:0] \u_ot.Xin1  ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _7070_ ;
wire _5803_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _2686__bF$buf0 ;
wire _2686__bF$buf1 ;
wire _2686__bF$buf2 ;
wire _2686__bF$buf3 ;
wire _2686__bF$buf4 ;
wire _2686__bF$buf5 ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire \genblk1[3].u_ce.Vld_bF$buf4  ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf3  ;
wire _5744_ ;
wire _5324_ ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _7067_ ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire [1:0] \genblk1[3].u_ce.Yin0  ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire clk_bF$buf76 ;
wire _134__bF$buf0 ;
wire clk_bF$buf77 ;
wire _134__bF$buf1 ;
wire clk_bF$buf78 ;
wire _134__bF$buf2 ;
wire _134__bF$buf3 ;
wire _134__bF$buf4 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire [11:4] \genblk1[1].u_ce.Ain12b  ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire \genblk1[4].u_ce.ISout  ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [11:4] \genblk1[3].u_ce.Ain12b  ;
wire _1185_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire [11:0] \genblk1[7].u_ce.Xcalc  ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _6911_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire [1:0] \genblk1[0].u_ce.Xin1  ;
wire [11:4] \genblk1[5].u_ce.Ain12b  ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire \genblk1[0].u_ce.ISin  ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _4324__bF$buf0 ;
wire _4324__bF$buf1 ;
wire _4324__bF$buf2 ;
wire _4324__bF$buf3 ;
wire _4324__bF$buf4 ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire [11:11] \genblk1[7].u_ce.Ain12b  ;
wire _5703_ ;
wire \genblk1[3].u_ce.Vld_bF$buf1  ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _5949__bF$buf0 ;
wire _5949__bF$buf1 ;
wire _5949__bF$buf2 ;
wire _5949__bF$buf3 ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire [19:0] FCW ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf0  ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _7064_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire [1:0] \genblk1[5].u_ce.Ain1  ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf1  ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire [1:0] \genblk1[6].u_ce.Xin0  ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf2  ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire [11:0] \genblk1[2].u_ce.Ycalc  ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire [11:4] \genblk1[7].u_ce.Xin12b  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire [11:0] \genblk1[3].u_ce.Acalc  ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _2731_ ;
wire _2311_ ;
wire \genblk1[1].u_ce.Vld_bF$buf2  ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire [1:0] \genblk1[3].u_ce.X_  ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _3510__bF$buf0 ;
wire _3510__bF$buf1 ;
wire _3510__bF$buf2 ;
wire _3510__bF$buf3 ;
wire _3510__bF$buf4 ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7023_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire \genblk1[1].u_ce.Vld  ;
wire _6714_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _7061_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _7058_ ;
wire _2193_ ;
wire \genblk1[0].u_ce.Rdy  ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _5829_ ;
wire _5409_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf2  ;
wire \genblk1[6].u_ce.Vld_bF$buf3  ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _6902_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7020_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire \genblk1[1].u_ce.ISout  ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire [1:0] \genblk1[1].u_ce.Yin1  ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf1  ;
wire _4239_ ;
wire _5600_ ;
wire [1:0] \genblk1[4].u_ce.Ain0  ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire [11:0] \genblk1[4].u_ce.Xcalc  ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf2  ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _7055_ ;
wire _2190_ ;
wire _3395_ ;
wire _5963__bF$buf0 ;
wire _5963__bF$buf1 ;
wire _5963__bF$buf2 ;
wire _5963__bF$buf3 ;
wire _5963__bF$buf4 ;
wire _5963__bF$buf5 ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _4621_ ;
wire _4201_ ;
wire [5:0] \genblk1[2].u_ce.LoadCtl  ;
wire _5826_ ;
wire _5406_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire \genblk1[4].u_ce.Vld_bF$buf4  ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire \genblk1[6].u_ce.Vld_bF$buf0  ;
wire _1649_ ;
wire _1229_ ;
wire [1:0] \genblk1[7].u_ce.Yin0  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire [5:0] \genblk1[7].u_ce.LoadCtl  ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire [1:0] \u_ot.Yin0  ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf4  ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire [1:0] \a[6]  ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire [1:0] \genblk1[4].u_ce.X_  ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7014_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire [1:0] \genblk1[4].u_ce.Xin1  ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire [11:0] \genblk1[0].u_ce.Acalc  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _7052_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \u_ot.LoadCtl_6_bF$buf3  ;
wire _3677_ ;
wire _3257_ ;
wire _5823_ ;
wire _5403_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf2  ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire \genblk1[4].u_ce.Vld_bF$buf1  ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire [11:4] \genblk1[0].u_ce.Ain12b  ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _7049_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf1  ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire [11:4] \genblk1[2].u_ce.Ain12b  ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire [11:0] \genblk1[6].u_ce.Ycalc  ;
wire [1:0] \genblk1[0].u_ce.Yin0  ;
wire \genblk1[0].u_ce.Rdy_bF$buf1  ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf2  ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire [11:4] \genblk1[4].u_ce.Ain12b  ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _7011_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf3  ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _5150__bF$buf0 ;
wire _5150__bF$buf1 ;
wire _5150__bF$buf2 ;
wire _5150__bF$buf3 ;
wire _5150__bF$buf4 ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1848__bF$buf0 ;
wire _1848__bF$buf1 ;
wire _1848__bF$buf2 ;
wire _1848__bF$buf3 ;
wire _1848__bF$buf4 ;
wire _1848__bF$buf5 ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire \u_ot.LoadCtl_6_bF$buf0  ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire \genblk1[2].u_ce.Vld_bF$buf4  ;
wire [11:4] \genblk1[2].u_ce.Xin12b  ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _5723_ ;
wire _5303_ ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _6562__bF$buf0 ;
wire _6562__bF$buf1 ;
wire _6562__bF$buf2 ;
wire _6562__bF$buf3 ;
wire _6562__bF$buf4 ;
wire [11:0] \genblk1[1].u_ce.Xcalc  ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7046_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire [11:4] \genblk1[4].u_ce.Xin12b  ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire Vld ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire [1:0] \genblk1[2].u_ce.Ain1  ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire _3098_ ;
wire [11:4] \genblk1[6].u_ce.Xin12b  ;
wire _5664_ ;
wire _5244_ ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf0  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _1678_ ;
wire _1258_ ;
wire [1:0] \genblk1[3].u_ce.Xin0  ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire \genblk1[2].u_ce.Vld_bF$buf1  ;
wire [1:0] \genblk1[5].u_ce.X_  ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire \u_ot.ISreg_bF$buf4  ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire [1:0] \genblk1[5].u_ce.Yin1  ;
wire _2425_ ;
wire _2005_ ;
wire _7043_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf2  ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf3  ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire [1:0] \a[1]  ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _972__bF$buf0 ;
wire _972__bF$buf1 ;
wire _972__bF$buf2 ;
wire _972__bF$buf3 ;
wire _972__bF$buf4 ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6998_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire \genblk1[0].u_ce.Vld_bF$buf2  ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7002_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [11:0] \genblk1[3].u_ce.Ycalc  ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire \u_ot.ISreg_bF$buf1  ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7040_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire [11:0] \genblk1[4].u_ce.Acalc  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire [5:0] \genblk1[4].u_ce.LoadCtl  ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire [1:0] \genblk1[1].u_ce.Ain0  ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf0  ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _2648__bF$buf0 ;
wire _4641_ ;
wire _2648__bF$buf1 ;
wire _4221_ ;
wire _2648__bF$buf2 ;
wire _2648__bF$buf3 ;
wire _2648__bF$buf4 ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf3  ;
wire _4926_ ;
wire _4506_ ;
wire \genblk1[5].u_ce.Vld_bF$buf3  ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire [1:0] \genblk1[4].u_ce.Yin0  ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _198_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf2  ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire [1:0] \genblk1[6].u_ce.X_  ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire [11:0] \u_ot.Ycalc  ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf3  ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _7034_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf4  ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire [1:0] \genblk1[1].u_ce.Xin1  ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf0  ;
wire _4923_ ;
wire _4503_ ;
wire \genblk1[5].u_ce.Vld_bF$buf0  ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _7069_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire [1:0] \genblk1[6].u_ce.Ain1  ;
wire _5784_ ;
wire _5364_ ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire [1:0] \genblk1[7].u_ce.Xin0  ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf0  ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _6913_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _7031_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf1  ;
wire _6722_ ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire [1:0] \u_ot.Xin0  ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire [11:4] \genblk1[1].u_ce.Xin12b  ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire [11:0] \genblk1[0].u_ce.Ycalc  ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire [11:4] \genblk1[3].u_ce.Xin12b  ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire \genblk1[3].u_ce.Vld_bF$buf3  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire [11:0] \genblk1[1].u_ce.Acalc  ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf2  ;
wire _5743_ ;
wire _5323_ ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _7066_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire [11:4] \genblk1[5].u_ce.Xin12b  ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf3  ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf4  ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _6910_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire [1:0] \genblk1[0].u_ce.Xin0  ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire \genblk1[1].u_ce.Vld_bF$buf4  ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire [1:0] \genblk1[7].u_ce.X_  ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire \genblk1[3].u_ce.Vld_bF$buf0  ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _7063_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire [1:0] \genblk1[2].u_ce.Yin1  ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _5605_ ;
wire [1:0] \genblk1[5].u_ce.Ain0  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _5188__bF$buf0 ;
wire _5188__bF$buf1 ;
wire _5188__bF$buf2 ;
wire _5188__bF$buf3 ;
wire _5188__bF$buf4 ;
wire _5188__bF$buf5 ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf0  ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _5925__bF$buf0 ;
wire _5925__bF$buf1 ;
wire _5925__bF$buf2 ;
wire _1848_ ;
wire _5925__bF$buf3 ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf1  ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire [1:0] \a[3]  ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _3486__bF$buf0 ;
wire _3486__bF$buf1 ;
wire _6598_ ;
wire _3486__bF$buf2 ;
wire _6178_ ;
wire _3486__bF$buf3 ;
wire _3486__bF$buf4 ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire \genblk1[1].u_ce.Vld_bF$buf1  ;
wire _3935_ ;
wire _3515_ ;
wire [5:0] \genblk1[6].u_ce.LoadCtl  ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _1598_ ;
wire _1178_ ;
wire [1:0] \genblk1[0].u_ce.Y_  ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _6904_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7022_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _7060_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire \genblk1[6].u_ce.Vld  ;
wire _6751_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf3  ;
wire _5602_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf4  ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1811__bF$buf0 ;
wire _1811__bF$buf1 ;
wire _1811__bF$buf2 ;
wire _1811__bF$buf3 ;
wire _1811__bF$buf4 ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire _1845_ ;
wire [1:0] \genblk1[5].u_ce.Xin1  ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _7057_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf1  ;
wire \genblk1[6].u_ce.Vld_bF$buf2  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _6901_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [1:0] \genblk1[1].u_ce.Yin0  ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf0  ;
wire _4238_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _6613_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf1  ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _135__bF$buf0 ;
wire _135__bF$buf1 ;
wire _135__bF$buf2 ;
wire _135__bF$buf3 ;
wire _135__bF$buf4 ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _7054_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _1010__bF$buf0 ;
wire _1010__bF$buf1 ;
wire _1010__bF$buf2 ;
wire _1010__bF$buf3 ;
wire _847_ ;
wire _1010__bF$buf4 ;
wire _427_ ;
wire _1010__bF$buf5 ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _2283_ ;
wire [6:0] \u_ot.LoadCtl  ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf4  ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire \genblk1[4].u_ce.Vld_bF$buf3  ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf3  ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _4325__bF$buf0 ;
wire _4325__bF$buf1 ;
wire _4325__bF$buf2 ;
wire _4325__bF$buf3 ;
wire _4325__bF$buf4 ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf3  ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire [1:0] \genblk1[3].u_ce.Ain1  ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire [1:0] \genblk1[1].u_ce.Y_  ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire [11:4] \genblk1[0].u_ce.Xin12b  ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _7013_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire [1:0] \genblk1[4].u_ce.Xin0  ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _7051_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \u_ot.LoadCtl_6_bF$buf2  ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf1  ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire \genblk1[4].u_ce.Vld_bF$buf0  ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _1645_ ;
wire _1225_ ;
wire [1:0] \genblk1[6].u_ce.Yin1  ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _7048_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire [11:4] \genblk1[3].u_ce.Yin12b  ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf0  ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire [11:4] \u_ot.Xin12b  ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf0  ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire [11:4] \genblk1[5].u_ce.Yin12b  ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf1  ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7010_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf2  ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire [11:4] \genblk1[7].u_ce.Yin12b  ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire \genblk1[5].u_ce.ISout  ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire \genblk1[2].u_ce.Vld_bF$buf3  ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire _5926__bF$buf0 ;
wire _5926__bF$buf1 ;
wire _5926__bF$buf2 ;
wire _5926__bF$buf3 ;
wire _5926__bF$buf4 ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7045_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire \genblk1[4].u_ce.Vld  ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire [1:0] \genblk1[2].u_ce.Ain0  ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire [11:0] \genblk1[2].u_ce.Acalc  ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;

DFFPOSX1 _11689_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.LoadCtl [4])
);

NAND3X1 _11269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3873_),
    .B(_3894_),
    .C(_3877_),
    .Y(_3908_)
);

FILL FILL_1__13772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12765_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5112_),
    .B(_5115_),
    .C(_5109_),
    .Y(_5116_)
);

FILL FILL_0__12345_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4755_),
    .B(_4756_),
    .Y(_4763_)
);

DFFPOSX1 _9837_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[2].u_ce.LoadCtl [0])
);

AND2X2 _9417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2212_),
    .B(_2227_),
    .Y(_2229_)
);

FILL FILL_1__8794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14137_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [11]),
    .Y(_6202_)
);

OAI21X1 _13415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5832_),
    .B(_5804_),
    .C(_5095_),
    .Y(_5088_)
);

FILL FILL_0__14911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7484_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2389_),
    .Y(_2391_)
);

AOI21X1 _9170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1979_),
    .B(_1976_),
    .C(_1971_),
    .Y(_1992_)
);

FILL FILL_0__10831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10411_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_807_),
    .C(_73_),
    .Y(_66_)
);

FILL FILL_2__13630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9648_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4436_),
    .B(_4453_),
    .C(_4435_),
    .Y(_4467_)
);

FILL FILL_0__9210_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_7010_)
);

FILL FILL_0__14088_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6654_),
    .B(_6662_),
    .Y(_6666_)
);

FILL FILL_1__7645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13408_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3019_),
    .B(_3020_),
    .C(_2694_),
    .Y(_3021_)
);

DFFPOSX1 _8861_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_859_),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.Xcalc [8])
);

OR2X2 _8441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(_1340_),
    .Y(_1341_)
);

OAI21X1 _8021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(\genblk1[1].u_ce.Ycalc [8]),
    .C(_924_),
    .Y(_941_)
);

NOR2X1 _11498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4112_),
    .B(_4098_),
    .Y(_4123_)
);

NAND3X1 _11078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf3),
    .B(_3725_),
    .C(_3724_),
    .Y(_3726_)
);

FILL FILL_1__13581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12154_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .Y(_2443_)
);

INVX1 _9226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2046_)
);

FILL FILL_1__8183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13779_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6019_),
    .B(_6017_),
    .C(_5997_),
    .Y(_5838_)
);

FILL FILL_0__13359_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain0 [0]),
    .Y(_5680_)
);

FILL FILL_0__14720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7059_),
    .B(_7060_),
    .Y(_6788_)
);

NAND3X1 _14429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6714_),
    .B(_6712_),
    .C(_6689_),
    .Y(_6715_)
);

NOR2X1 _14009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6364_),
    .B(_6368_),
    .Y(_6369_)
);

FILL FILL_0__7293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10220_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(gnd),
    .S(_685_),
    .Y(_687_)
);

FILL FILL_0__8498_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3433_)
);

FILL FILL_0__8078_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf3),
    .B(_3073_),
    .C(_3070_),
    .Y(_3074_)
);

FILL FILL_1__12852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11425_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [5]),
    .Y(_4287_)
);

FILL FILL_0__11005_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14182_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5858_),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.Xcalc [10])
);

DFFPOSX1 _8917_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.LoadCtl [4])
);

FILL FILL_1__7874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x86550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13217_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5386_)
);

FILL FILL_1__8659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9600_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1555_),
    .C(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .Y(_1557_)
);

OAI21X1 _8250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(_1156_),
    .C(_1157_),
    .Y(_1158_)
);

BUFX2 BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert121 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf4 )
);

FILL FILL_2__7103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13390_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert123 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert124 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert126 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 )
);

FILL FILL_2__11769_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 )
);

FILL FILL_2__11349_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert128 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 )
);

FILL FILL_0__12383_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 )
);

FILL FILL_2__12710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7769_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[3].u_ce.Ycalc [0]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Ycalc [2]),
    .Y(_2623_)
);

FILL FILL_0__7349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .B(_2232_),
    .C(_1848__bF$buf2),
    .Y(_2265_)
);

NAND3X1 _9035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf1),
    .B(_1826_),
    .C(_1863_),
    .Y(_1864_)
);

FILL FILL_1__11703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14595_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6238_)
);

FILL FILL_0__13588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13168_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13453_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5053_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Acalc [1])
);

INVX1 _13033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5499_)
);

FILL FILL_1__9197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10095_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6877_),
    .Y(_6885_)
);

NAND2X1 _14238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(\u_ot.Xcalc [7]),
    .Y(_6552_)
);

FILL FILL_2__8481_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7941_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Acalc [0])
);

AOI21X1 _7521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(_506_),
    .C(_180_),
    .Y(_507_)
);

OAI21X1 _7101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_105_),
    .C(_106_),
    .Y(_107_)
);

AOI21X1 _10998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3610_),
    .B(_3487__bF$buf2),
    .C(_3631_),
    .Y(_3649_)
);

NOR2X1 _10578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3283_),
    .B(_3288_),
    .Y(_3289_)
);

NAND3X1 _10158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2889_),
    .C(_2886_),
    .Y(_2892_)
);

FILL FILL_1__12661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_1584_),
    .Y(_1609_)
);

NAND3X1 _8306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1211_),
    .C(_1210_),
    .Y(_1212_)
);

FILL FILL_1__7683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12859_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf0),
    .B(_5166_),
    .C(_5203_),
    .Y(_5204_)
);

FILL FILL_0__12439_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4851_),
    .B(_4850_),
    .C(_4843_),
    .Y(_4214_)
);

FILL FILL_0__12019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10793_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6248_),
    .B(_6031_),
    .Y(_6292_)
);

NOR2X1 _13509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[7].u_ce.LoadCtl [1]),
    .Y(_5892_)
);

FILL FILL_2__11998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_2475_),
    .C(_2476_),
    .Y(_1713_)
);

OR2X2 _9264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2082_),
    .B(_2078_),
    .Y(_2083_)
);

FILL FILL_1__11932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10505_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6055_),
    .B(_6054_),
    .Y(_6056_)
);

FILL FILL_0__13397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5716_),
    .B(_5707_),
    .C(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .Y(_5717_)
);

FILL FILL_1__12717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9304_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14887_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6778_),
    .CLK(clk_bF$buf50),
    .Q(\u_pa.acc_reg [11])
);

OAI21X1 _14467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6731_),
    .B(_6740_),
    .C(_6742_),
    .Y(_6521_)
);

AOI21X1 _14047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6404_),
    .B(_6403_),
    .C(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6405_)
);

FILL FILL_1__7739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(_241_),
    .C(_172__bF$buf3),
    .Y(_722_)
);

INVX1 _7330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_324_)
);

NOR2X1 _10387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3096_),
    .B(_3086_),
    .Y(_3111_)
);

FILL FILL_1__12890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11043_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1786_),
    .C(_1787_),
    .Y(_1788_)
);

NAND2X1 _8535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1424_),
    .B(_1427_),
    .Y(_1431_)
);

MUX2X1 _8115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .S(vdd),
    .Y(_1030_)
);

FILL FILL_1__7492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13255_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5422_),
    .B(_5418_),
    .Y(_5423_)
);

FILL FILL_0__12668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12248_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4854_),
    .C(_4268_),
    .Y(_4261_)
);

NAND2X1 _12113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4625_),
    .B(_4430_),
    .Y(_4670_)
);

FILL FILL_1__8697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6078_),
    .B(_6080_),
    .C(_6108_),
    .Y(_6109_)
);

INVX1 _13318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5769_),
    .Y(_5770_)
);

FILL FILL_1_CLKBUF1_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2299_),
    .B(_2300_),
    .Y(_2301_)
);

INVX1 _9073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .Y(_1900_)
);

FILL FILL_1__11741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13491_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5091_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Ain1 [0])
);

FILL FILL_0_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5534_),
    .Y(_5535_)
);

FILL FILL_0_BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_774_),
    .Y(_775_)
);

FILL FILL_1__12946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11519_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4373_),
    .C(_4374_),
    .Y(_4375_)
);

FILL FILL_0__9113_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6919_),
    .B(_6916_),
    .Y(_6921_)
);

OAI21X1 _14276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf2),
    .B(_6580_),
    .C(_6581_),
    .Y(_6491_)
);

FILL FILL_1__7548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14318_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2927_),
    .Y(_2928_)
);

FILL FILL_2__10658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11272_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1636_),
    .B(_923_),
    .Y(_1641_)
);

NAND2X1 _8344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .B(_1162_),
    .Y(_1248_)
);

FILL FILL_2__7617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12897_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5239_),
    .Y(_5240_)
);

FILL FILL_0__12477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12057_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4878_),
    .B(_4883_),
    .Y(_4886_)
);

INVX1 _9969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2711_),
    .Y(_2712_)
);

OR2X2 _9549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2353_)
);

NAND3X1 _9129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1922_),
    .B(_1939_),
    .C(_1921_),
    .Y(_1953_)
);

FILL FILL_1__8086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6312_),
    .B(_6316_),
    .Y(_6328_)
);

INVX8 _13547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_5926_)
);

AND2X2 _13127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5582_),
    .Y(_5589_)
);

FILL FILL_0__14623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10123_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_572_),
    .Y(_597_)
);

FILL FILL_1__12755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11328_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11613_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3353_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Ycalc [1])
);

AND2X2 _14085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6429_),
    .B(_6440_),
    .Y(_6441_)
);

FILL FILL_1__7777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5262_),
    .B(_5279_),
    .C(_5261_),
    .Y(_5293_)
);

FILL FILL257250x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9503_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(gnd),
    .Y(_1823_)
);

NAND2X1 _8573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1073_),
    .B(_1466_),
    .Y(_1467_)
);

OAI21X1 _8153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1065_),
    .C(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_1066_)
);

FILL FILL_1__10821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13293_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf4),
    .B(_5458_),
    .C(_5447_),
    .Y(_5459_)
);

DFFPOSX1 _12571_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4225_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [10])
);

FILL FILL_0__12286_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4575_),
    .C(_4705_),
    .Y(_4706_)
);

DFFPOSX1 _9778_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1690_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Xcalc [1])
);

NAND2X1 _9358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [10]),
    .Y(_2172_)
);

FILL FILL_1__11606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14078_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6139_),
    .B(_6145_),
    .C(_6142_),
    .Y(_6146_)
);

OAI21X1 _13356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Xin12b [9]),
    .Y(_5803_)
);

FILL FILL_2__13818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10352_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Xin12b [9]),
    .Y(_806_)
);

INVX1 _7424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .Y(_414_)
);

FILL FILL_1__12984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11557_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4410_),
    .Y(_4411_)
);

FILL FILL_2__9169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11137_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf3),
    .B(_4051_),
    .C(_3524__bF$buf2),
    .Y(_4052_)
);

INVX1 _11002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3651_),
    .Y(_3653_)
);

NAND2X1 _8629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1508_),
    .B(_1517_),
    .Y(_1519_)
);

NAND2X1 _8209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf4),
    .B(_1029_),
    .Y(_1119_)
);

FILL FILL_1__7586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13349_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [5]),
    .Y(_5113_)
);

OAI21X1 _12207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4721_),
    .B(_4704_),
    .C(_4759_),
    .Y(_4760_)
);

FILL FILL_1__14710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9312_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_984_),
    .B(_1281_),
    .Y(_1284_)
);

FILL FILL_1__10630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14908_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(_4921_),
    .Y(_4922_)
);

FILL FILL_0__12095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12422_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2105_),
    .C(_2387_),
    .Y(_2388_)
);

OAI21X1 _9167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .B(_1988_),
    .C(_1989_),
    .Y(_1990_)
);

FILL FILL_1__11835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10408_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _13585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5963_)
);

OAI21X1 _13165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5602_),
    .B(_5599_),
    .C(_5188__bF$buf2),
    .Y(_5625_)
);

FILL FILL_2__13627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10161_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_631_),
    .C(_619_),
    .Y(_22_)
);

OAI21X1 _7233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_207_),
    .C(_220_),
    .Y(_231_)
);

FILL FILL_1__12793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11366_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11651_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3391_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xin12b [8])
);

OAI21X1 _11231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3788_),
    .C(_3871_),
    .Y(_3872_)
);

DFFPOSX1 _8858_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_856_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[1].u_ce.Xcalc [5])
);

NAND2X1 _8438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1079_),
    .B(_1286_),
    .Y(_1338_)
);

AOI22X1 _8018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.Acalc [1]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Acalc [3]),
    .Y(_939_)
);

FILL FILL_1__7395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5324_),
    .B(_5328_),
    .C(_5329_),
    .Y(_5330_)
);

OAI22X1 _12436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4284_),
    .B(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .C(_4973_),
    .D(_4972_),
    .Y(_4224_)
);

INVX1 _12016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4576_),
    .Y(_4577_)
);

FILL FILL_0__13932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9121_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1081_),
    .B(_1072_),
    .C(_1010__bF$buf1),
    .Y(_1102_)
);

FILL FILL_0__14717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7884_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2190_),
    .Y(_2209_)
);

FILL FILL_1__11224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8651_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3571_),
    .B(_3573_),
    .C(_3559_),
    .Y(_3577_)
);

FILL FILL_0__8231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10637_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3212_),
    .B(_3216_),
    .Y(_3218_)
);

FILL FILL_0__10217_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5824_)
);

FILL FILL_2__9610_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_676_),
    .C(_681_),
    .Y(_684_)
);

FILL FILL_2__13856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9436_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [9]),
    .Y(_4284_)
);

FILL FILL_0__9016_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6802_),
    .B(_6834_),
    .Y(_6764_)
);

DFFPOSX1 _14179_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5855_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [7])
);

FILL FILL_0__10390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8812_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_827_)
);

OAI21X1 _7462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_171_),
    .C(_449_),
    .Y(_450_)
);

AOI21X1 _10099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2834_),
    .B(_2818_),
    .C(_2830_),
    .Y(_2835_)
);

FILL FILL256650x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11595_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4447_)
);

FILL FILL_0__11175_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4086_),
    .Y(_4087_)
);

NOR2X1 _11040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3689_),
    .B(_3673_),
    .Y(_3690_)
);

FILL FILL_2__11922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(_1552_),
    .Y(_1554_)
);

AND2X2 _8247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .B(_1109_),
    .Y(_1155_)
);

FILL FILL_1__10915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13387_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Xcalc [1]),
    .C(_5146_),
    .D(_5109_),
    .Y(_5147_)
);

OAI21X1 _12245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4795_),
    .C(_4775_),
    .Y(_4796_)
);

FILL FILL_2__12707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9350_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_7027_)
);

FILL FILL_0__14106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8040_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10731_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2557_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xin12b [4])
);

FILL FILL_0__10446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10026_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .B(_3035_),
    .Y(_3038_)
);

DFFPOSX1 _7938_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [9])
);

OAI21X1 _7518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_474_),
    .C(_172__bF$buf0),
    .Y(_504_)
);

FILL FILL_2__13665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9665_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4462_),
    .B(_4444_),
    .C(_4500_),
    .Y(_4501_)
);

FILL FILL_0__9245_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4138_),
    .Y(_4139_)
);

FILL FILL_1__8621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8201_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [0]),
    .B(_158__bF$buf4),
    .Y(_668_)
);

FILL FILL_1__14804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_267_),
    .C(_265_),
    .Y(_268_)
);

FILL FILL_1__9406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8896_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_894_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[1].u_ce.Yin12b [5])
);

FILL FILL_0_CLKBUF1_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1352_),
    .C(_1365_),
    .Y(_1374_)
);

FILL FILL_0_CLKBUF1_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _8056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_972_)
);

FILL FILL_0_CLKBUF1_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5276_),
    .C(_5342_),
    .Y(_5366_)
);

NAND2X1 _12474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_5000_),
    .Y(_5002_)
);

FILL FILL_0__12189_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [0]),
    .B(_4348__bF$buf0),
    .Y(_4613_)
);

FILL FILL_2__12936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf0),
    .B(_6051_),
    .C(_6052_),
    .Y(_6053_)
);

NAND2X1 _13259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5708_),
    .B(_5712_),
    .Y(_5714_)
);

FILL FILL_0__14755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14335_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6850_),
    .B(_6849_),
    .Y(_6851_)
);

DFFPOSX1 _14200_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5876_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Yin12b [6])
);

FILL FILL_1__11262_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf0),
    .B(_3515_),
    .Y(_3613_)
);

FILL FILL_0__10675_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2678_),
    .C(_2648__bF$buf4),
    .Y(_3253_)
);

FILL FILL_0__10255_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2855_),
    .Y(_2856_)
);

OAI21X1 _7747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_718_),
    .C(_709_),
    .Y(_29_)
);

AOI21X1 _7327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_304_),
    .C(_316_),
    .Y(_321_)
);

FILL FILL_2__13894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9474_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(\genblk1[5].u_ce.Xcalc [9]),
    .C(_4276_),
    .Y(_4318_)
);

FILL FILL_0__9054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .B(_3961_),
    .Y(_3962_)
);

FILL FILL_0__12821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14613_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _7080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_88_)
);

FILL FILL_0__13606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11120_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_)
);

FILL FILL_1__10953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7138_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4812_),
    .B(_4831_),
    .C(_4362__bF$buf2),
    .Y(_4832_)
);

FILL FILL_2__12745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8325_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13488_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5088_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain12b [7])
);

OAI21X1 _13068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5401_),
    .C(_5531_),
    .Y(_5532_)
);

FILL FILL_0__14564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10064_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7976_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_60_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin0 [1])
);

NAND2X1 _7556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf0),
    .B(_459_),
    .Y(_540_)
);

OAI21X1 _7136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_136_),
    .C(_137_),
    .Y(_138_)
);

FILL FILL_1__12696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12276_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4536_),
    .B(_4510_),
    .C(_4535_),
    .Y(_4537_)
);

FILL FILL_0__9283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11269_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_4166_)
);

NAND2X1 _11134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3778_),
    .Y(_3779_)
);

FILL FILL_0__12630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14068_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2486_),
    .Y(_2488_)
);

INVX1 _12759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5236_),
    .Y(_5237_)
);

NAND2X1 _12339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .B(_4883_),
    .Y(_4884_)
);

FILL FILL_1__14842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13835_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf1),
    .B(_6071_),
    .C(_6072_),
    .Y(_6073_)
);

FILL FILL_0__13415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9024_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1009_)
);

FILL FILL_1__10342_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14905_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6796_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.Atmp [9])
);

FILL FILL_2__7787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf3),
    .B(_4649_),
    .C(_4642_),
    .Y(_4650_)
);

FILL FILL_2__12974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x201750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf3),
    .B(_2111_),
    .Y(_2116_)
);

FILL FILL_1__11967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8554_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3478_),
    .B(_3435_),
    .C(_3483_),
    .Y(\genblk1[4].u_ce.X_ [1])
);

FILL FILL_0__8134_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3127_),
    .B(_3126_),
    .C(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3128_)
);

NAND2X1 _13297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [6]),
    .B(_5749_),
    .Y(_5750_)
);

FILL FILL_2__9933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10620_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_172__bF$buf5),
    .Y(_755_)
);

NAND3X1 _7365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .B(_357_),
    .C(_356_),
    .Y(_358_)
);

FILL FILL_1__12085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11498_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_4354_)
);

FILL FILL_0__9092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11078_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3994_),
    .B(_3992_),
    .Y(_3998_)
);

FILL FILL_1__10818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7825_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2668_),
    .Y(_2674_)
);

FILL FILL_0__7405_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2298_),
    .B(_2317_),
    .C(_1848__bF$buf0),
    .Y(_2318_)
);

NAND2X1 _12988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5451_),
    .Y(_5456_)
);

DFFPOSX1 _12568_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4222_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [7])
);

AOI22X1 _12148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4348__bF$buf2),
    .C(_4703_),
    .D(_4346_),
    .Y(_4206_)
);

FILL FILL_1__14651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x111750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert111 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert112 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert114 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert116 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert118 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert119 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14429_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6929_),
    .B(_6919_),
    .Y(_6937_)
);

FILL FILL_0__14009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8363_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[2].u_ce.X_ [1]),
    .Y(_3330_)
);

FILL FILL_0__10349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf3),
    .B(_2941_),
    .C(_2944_),
    .Y(_2945_)
);

FILL FILL_0__11710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9568_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4406_),
    .B(_4407_),
    .Y(_4408_)
);

FILL FILL_0__9148_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4048_),
    .Y(_4049_)
);

FILL FILL_1__13922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8104_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_575_),
    .C(_576_),
    .Y(_577_)
);

FILL FILL_1__14707_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_173_),
    .C(_174_),
    .Y(_175_)
);

OAI21X1 _11592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4185_),
    .B(_4155_),
    .C(_4186_),
    .Y(_3415_)
);

OAI21X1 _11172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3795_),
    .C(_3815_),
    .Y(_3816_)
);

FILL FILL_1__9729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1645_),
    .C(_1661_),
    .Y(_891_)
);

OAI21X1 _8379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_984_),
    .B(_1281_),
    .C(_994_),
    .Y(_1282_)
);

FILL FILL_1__10627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7634_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [1]),
    .B(_2475_),
    .Y(_2508_)
);

FILL FILL_0__7214_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf2),
    .B(_2135_),
    .C(_2128_),
    .Y(_2136_)
);

FILL FILL_1__13099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5273_)
);

INVX1 _12377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4918_),
    .Y(_4919_)
);

FILL FILL_1__14460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14658_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14523_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6511_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Ycalc [11])
);

FILL FILL_0__14238_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6047_),
    .B(_6455_),
    .C(_6456_),
    .Y(_5860_)
);

FILL FILL_2__12172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8592_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(gnd),
    .C(_3487__bF$buf4),
    .Y(_3520_)
);

FILL FILL_0__8172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10158_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3152_),
    .B(_3163_),
    .Y(_3164_)
);

AOI21X1 _10023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2761_),
    .B(_2758_),
    .C(_2747_),
    .Y(_2763_)
);

FILL FILL_2__10905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9377_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11648_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3388_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [11])
);

NAND2X1 _11228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3868_),
    .Y(_3869_)
);

FILL FILL_1__13731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9118_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf0),
    .B(_1001_),
    .Y(_1099_)
);

FILL FILL_1__10856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7443_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4366_),
    .B(_4737_),
    .C(_4733_),
    .Y(_4740_)
);

FILL FILL_2__8822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8648_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3573_),
    .B(_3571_),
    .Y(_3574_)
);

FILL FILL_0__8228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14467_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6972_)
);

FILL FILL_0__14047_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6627_),
    .C(_6630_),
    .Y(_6631_)
);

FILL FILL_1__7604_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert390 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert391 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

FILL FILL_1__11394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [6]),
    .B(_3321_),
    .Y(_3351_)
);

FILL FILL_0__10387_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2980_),
    .B(_2981_),
    .Y(_2982_)
);

FILL FILL_1__8809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9360_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_810_),
    .C(_825_),
    .Y(_55_)
);

NAND2X1 _7459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_447_)
);

FILL FILL_2__13186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(_1641_),
    .C(_1672_),
    .Y(_901_)
);

OAI21X1 _8400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1281_),
    .C(_1301_),
    .Y(_1302_)
);

FILL FILL_1__12179_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4421_),
    .B(_4438_),
    .C(_4439_),
    .Y(_4444_)
);

FILL FILL_0__9186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _11457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3449_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_4082_),
    .D(_4084_),
    .Y(_3382_)
);

NAND3X1 _11037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(_3685_),
    .C(_3686_),
    .Y(_3687_)
);

FILL FILL_1__13960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12113_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .Y(_2405_)
);

FILL FILL_1__8982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x136950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13738_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(\genblk1[7].u_ce.Xin12b [5]),
    .S(vdd),
    .Y(_5981_)
);

FILL FILL_0__13318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10245_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7023_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(_7024_),
    .Y(_6783_)
);

FILL FILL_0__7672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8037_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10728_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2554_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xin12b [9])
);

INVX1 _10308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3035_)
);

FILL FILL_1__12811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14276_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [4]),
    .Y(_6804_)
);

NAND2X1 _14141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .B(_6463_),
    .Y(_6479_)
);

FILL FILL_1__7833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14603_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3197_),
    .B(_3190_),
    .C(_3195_),
    .Y(_3198_)
);

FILL FILL_0__10196_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2796_),
    .Y(_2799_)
);

FILL FILL_1__8618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10103_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_662_),
    .Y(_665_)
);

OR2X2 _7268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_263_),
    .Y(_265_)
);

FILL FILL256950x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11686_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.LoadCtl [1])
);

OAI21X1 _11266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3904_),
    .B(_3905_),
    .C(_3508_),
    .Y(_3906_)
);

FILL FILL_2__11308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7728_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9834_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1746_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Ain1 [1])
);

FILL FILL_0__7308_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_2223_),
    .C(_2219_),
    .Y(_2226_)
);

FILL FILL_1__8791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13547_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [11]),
    .B(_5949__bF$buf3),
    .Y(_6199_)
);

FILL FILL_0__13127_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [6]),
    .B(_5804_),
    .Y(_5834_)
);

FILL FILL_1__9996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10054_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6838_),
    .B(_6841_),
    .C(_6839_),
    .Y(_6848_)
);

FILL FILL_0__7481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12686_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [6]),
    .B(_807_),
    .Y(_837_)
);

FILL FILL_1__11259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8686_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3608_),
    .C(_3609_),
    .Y(_3610_)
);

FILL FILL_0__8266_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3228_),
    .B(_3242_),
    .C(_3240_),
    .Y(_3250_)
);

OAI21X1 _10117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2822_),
    .B(_2826_),
    .C(_2821_),
    .Y(_2853_)
);

FILL FILL_1__12620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7006_),
    .B(_7005_),
    .Y(_7007_)
);

FILL FILL_0__14085_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6654_),
    .B(_6662_),
    .Y(_6663_)
);

FILL FILL_1__7642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12818_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2997_),
    .B(_2988_),
    .C(_2686__bF$buf3),
    .Y(_3018_)
);

FILL FILL_1__8427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf0),
    .B(_483_),
    .C(_474_),
    .Y(_484_)
);

INVX4 _7077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .Y(_85_)
);

AOI21X1 _11495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4117_),
    .B(_4053_),
    .C(\genblk1[4].u_ce.Ain12b [8]),
    .Y(_4120_)
);

NOR3X1 _11075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .B(_3702_),
    .C(_3675_),
    .Y(_3723_)
);

FILL FILL_0__12991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7537_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1830_),
    .Y(_2440_)
);

FILL FILL_0__7117_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(_2042_),
    .C(_2040_),
    .Y(_2043_)
);

FILL FILL_1__8180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13776_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6015_),
    .B(_6016_),
    .C(_5951_),
    .Y(_6017_)
);

FILL FILL_0__13356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5677_),
    .B(_5676_),
    .C(_5669_),
    .Y(_5052_)
);

FILL FILL_1__9385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7057_),
    .B(_7058_),
    .Y(_6787_)
);

NAND2X1 _14426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(\u_ot.Yin12b [10]),
    .Y(_6712_)
);

NAND3X1 _14006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6341_),
    .B(_6365_),
    .C(_6340_),
    .Y(_6366_)
);

FILL FILL_0__7290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert100 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert101 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert102 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert103 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert104 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert105 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert106 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert107 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8075_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10766_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.LoadCtl [5])
);

AOI21X1 _10346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf1),
    .B(_3030_),
    .C(_3052_),
    .Y(_3071_)
);

FILL FILL_2__10808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11002_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8914_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.LoadCtl [1])
);

FILL FILL_1__7871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13214_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5328_),
    .B(_5382_),
    .C(_5380_),
    .Y(_5383_)
);

FILL FILL_0__12627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7766_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [6]),
    .B(_2603_),
    .Y(_2620_)
);

FILL FILL_0__7346_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2174_),
    .C(_2261_),
    .Y(_2262_)
);

OAI21X1 _9032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1859_),
    .C(_1860_),
    .Y(_1861_)
);

FILL FILL_1__11700_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4466_),
    .C(_4646_),
    .Y(_4647_)
);

FILL FILL_2__8725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256050x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13585_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6235_),
    .B(_6230_),
    .C(_6214_),
    .Y(_5848_)
);

FILL FILL_0__13165_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13450_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5050_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [9])
);

NAND2X1 _13030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5451_),
    .B(_5256_),
    .Y(_5496_)
);

FILL FILL_1__9194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10092_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [5]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf1),
    .Y(_6883_)
);

NAND2X1 _14235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [6]),
    .Y(_6550_)
);

FILL FILL_1__7507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11297_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [6]),
    .Y(_3646_)
);

AOI21X1 _10575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3285_),
    .B(_3250_),
    .C(_3284_),
    .Y(_3286_)
);

INVX1 _10155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2887_),
    .Y(_2889_)
);

FILL FILL_0__11231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13089_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1539_),
    .C(\genblk1[1].u_ce.Ain12b [8]),
    .Y(_1606_)
);

NOR3X1 _8303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(_1188_),
    .C(_1161_),
    .Y(_1209_)
);

FILL FILL_1__7680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12856_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5199_),
    .C(_5200_),
    .Y(_5201_)
);

FILL FILL_0__12436_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4848_),
    .B(_4847_),
    .Y(_4849_)
);

FILL FILL_0__12016_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2646_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_2671_),
    .Y(_2514_)
);

OAI21X1 _9508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2233_),
    .C(_2261_),
    .Y(_2315_)
);

FILL FILL_1__8465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14228_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6288_),
    .B(_6245_),
    .S(vdd),
    .Y(_6289_)
);

NOR2X1 _13506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .B(\genblk1[7].u_ce.LoadCtl [3]),
    .Y(_5889_)
);

FILL FILL_2__11575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7575_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1762_),
    .B(_1768_),
    .Y(_2474_)
);

FILL FILL_0__7155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2056_),
    .C(_2035_),
    .Y(_2080_)
);

FILL FILL_0__10922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14599_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14884_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6775_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [8])
);

OAI21X1 _14464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Xin1 [0]),
    .Y(_6741_)
);

AOI21X1 _14044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6401_),
    .B(_6399_),
    .C(_6394_),
    .Y(_6402_)
);

FILL FILL_1__7736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2687_),
    .B(_3106_),
    .C(_3107_),
    .Y(_3108_)
);

FILL FILL_2__10846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11040_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(_1784_),
    .Y(\genblk1[2].u_ce.Y_ [0])
);

NAND2X1 _8532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1427_),
    .Y(_1428_)
);

MUX2X1 _8112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .S(vdd),
    .Y(_1027_)
);

OAI21X1 _11589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf4),
    .B(_4151_),
    .C(_4184_),
    .Y(_3414_)
);

NAND3X1 _11169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf1),
    .B(_3812_),
    .C(_3790_),
    .Y(_3813_)
);

FILL FILL_1__13672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13252_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5393_),
    .B(_5396_),
    .C(_5375_),
    .Y(_5420_)
);

FILL FILL_0__12665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12245_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_4267_)
);

NAND2X1 _12110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4623_),
    .Y(_4667_)
);

OAI21X1 _9737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1847_),
    .C(_2506_),
    .Y(_1736_)
);

OAI21X1 _9317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1952_),
    .C(_2132_),
    .Y(_2133_)
);

FILL FILL_1__8694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14037_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [7]),
    .Y(_6106_)
);

NOR2X1 _13315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5170_),
    .Y(_5767_)
);

FILL FILL_1_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7384_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2215_),
    .C(_2261_),
    .Y(_2298_)
);

INVX1 _9070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .Y(_1897_)
);

FILL FILL_2__8763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10311_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_736_),
    .C(_770_),
    .Y(_772_)
);

FILL FILL_2__13530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4370_),
    .C(_4371_),
    .Y(_4372_)
);

FILL FILL_0__9110_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6918_)
);

OR2X2 _14273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6577_),
    .B(\u_ot.Xin1 [1]),
    .Y(_6579_)
);

FILL FILL_1__7545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13308_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_2925_)
);

NAND2X1 _8761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1637_),
    .Y(_1639_)
);

AOI22X1 _8341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_940_),
    .B(_996__bF$buf4),
    .C(_1245_),
    .D(_1068_),
    .Y(_849_)
);

OAI21X1 _11398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4025_),
    .B(_4027_),
    .C(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4030_)
);

FILL FILL_1__13061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12054_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .B(_2705_),
    .S(_2648__bF$buf3),
    .Y(_2709_)
);

OAI21X1 _9546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(_2338_),
    .C(_1848__bF$buf3),
    .Y(_2350_)
);

AOI22X1 _9126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1781_),
    .B(_1834__bF$buf3),
    .C(_1950_),
    .D(_1906_),
    .Y(_1681_)
);

FILL FILL_1__8083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13679_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5912_),
    .B(_5949__bF$buf0),
    .C(_6325_),
    .D(_5947_),
    .Y(_5852_)
);

INVX1 _13544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [0]),
    .Y(_5923_)
);

FILL FILL_0__13259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5547_),
    .B(_5530_),
    .C(_5585_),
    .Y(_5586_)
);

FILL FILL_0__14620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10186_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6962_),
    .Y(_6969_)
);

INVX1 _14329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [10]),
    .Y(_6628_)
);

FILL FILL_0__7193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_592_),
    .C(_593_),
    .Y(_594_)
);

FILL FILL_0__8398_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [1]),
    .Y(_3349_)
);

AOI21X1 _10249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2975_),
    .B(_2978_),
    .C(_2697_),
    .Y(_2979_)
);

FILL FILL_1__12752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11325_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[4] [1]),
    .Y(_3431_)
);

NOR2X1 _14082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6431_),
    .B(_6433_),
    .Y(_6438_)
);

OAI21X1 _8817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf5),
    .B(_1637_),
    .C(_1670_),
    .Y(_900_)
);

FILL FILL_1__7774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13117_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5121_),
    .B(_5174__bF$buf2),
    .C(_5290_),
    .D(_5246_),
    .Y(_5033_)
);

FILL FILL_1__8979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9500_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1820_)
);

OR2X2 _8570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1462_),
    .B(_1461_),
    .Y(_1464_)
);

OAI21X1 _8150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1057_),
    .B(_1059_),
    .C(_1045_),
    .Y(_1063_)
);

FILL FILL_1__13290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7669_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9775_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1687_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Ycalc [10])
);

FILL FILL_0__7249_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834__bF$buf4),
    .B(_2169_),
    .C(_2148_),
    .Y(_1691_)
);

FILL FILL_1__11603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14075_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6118_),
    .B(_6114_),
    .Y(_6143_)
);

FILL FILL_0__13068_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5801_)
);

FILL FILL_2__13815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12808_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [6]),
    .Y(_6801_)
);

INVX1 _14138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6477_)
);

FILL FILL257250x237750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8381_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_804_)
);

INVX1 _7421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_411_)
);

AOI21X1 _10898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3554_),
    .B(_3553_),
    .C(_3512_),
    .Y(_3555_)
);

NAND2X1 _10478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .B(_3195_),
    .Y(_3196_)
);

OAI21X1 _10058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf2),
    .B(_2794_),
    .C(_2795_),
    .Y(_2796_)
);

FILL FILL_1__12981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11134_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(_1513_),
    .C(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1516_)
);

NAND2X1 _8206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1116_)
);

FILL FILL_1__7583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12759_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [9]),
    .Y(_5110_)
);

FILL FILL_0__12339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4756_),
    .B(_4755_),
    .Y(_4757_)
);

FILL FILL_0__13700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6194_),
    .B(_6196_),
    .C(_6018_),
    .Y(_6197_)
);

INVX1 _13409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [1]),
    .Y(_5832_)
);

FILL FILL_2__11898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [4]),
    .B(_1834__bF$buf2),
    .Y(_2385_)
);

OAI21X1 _9164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_1930_),
    .C(_1986_),
    .Y(_1987_)
);

FILL FILL_1__11832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10405_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf1),
    .B(_5959_),
    .C(_5958_),
    .Y(_5960_)
);

FILL FILL_0__13297_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5621_),
    .C(_5601_),
    .Y(_5622_)
);

FILL FILL257250x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9204_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7003_),
    .B(_6977_),
    .Y(_7004_)
);

OAI21X1 _14367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6543_),
    .B(\u_ot.LoadCtl_6_bF$buf4 ),
    .C(_6660_),
    .Y(_6503_)
);

FILL FILL_1__7639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_629_),
    .Y(_630_)
);

OAI21X1 _7230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_226_),
    .C(_206_),
    .Y(_3_)
);

NAND2X1 _10287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2971_),
    .B(_2754_),
    .Y(_3015_)
);

FILL FILL_1__12790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11363_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8855_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_853_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Xcalc [2])
);

OAI21X1 _8435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1208_),
    .C(_1334_),
    .Y(_1335_)
);

NAND2X1 _8015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [7]),
    .B(_927_),
    .Y(_936_)
);

FILL FILL_1__7392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12988_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5288_),
    .B(_5270_),
    .C(_5326_),
    .Y(_5327_)
);

FILL FILL_0__12148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4970_),
    .B(_4969_),
    .Y(_4971_)
);

OAI21X1 _12013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4300_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4574_),
    .Y(_4200_)
);

FILL FILL_1__8597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5998_),
    .B(_6013_),
    .Y(_6014_)
);

NOR2X1 _13218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5674_),
    .B(_5673_),
    .Y(_5675_)
);

FILL FILL_0__14714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_2205_),
    .C(_2204_),
    .Y(_2206_)
);

FILL FILL_1__11221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10214_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5271_),
    .B(_5807_),
    .C(_5822_),
    .Y(_5077_)
);

NAND2X1 _7706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_681_),
    .Y(_682_)
);

FILL FILL_1__12846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4282_)
);

FILL FILL_0__9013_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [0]),
    .B(En_bF$buf3),
    .Y(_6761_)
);

DFFPOSX1 _14176_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5852_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [4])
);

FILL FILL_1__7868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14218_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5379_),
    .B(_5351_),
    .Y(_5380_)
);

NAND3X1 _10096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2803_),
    .C(_2831_),
    .Y(_2832_)
);

FILL FILL_2__10558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11172_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1510_),
    .C(_1550_),
    .Y(_1551_)
);

AOI22X1 _8244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1132_),
    .B(_996__bF$buf4),
    .C(_1152_),
    .D(_1068_),
    .Y(_845_)
);

FILL FILL_1__10912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12797_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(\genblk1[6].u_ce.Xcalc [9]),
    .C(_5106_),
    .Y(_5144_)
);

FILL FILL_0__12377_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4793_)
);

OAI21X1 _9869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(\genblk1[3].u_ce.Ycalc [8]),
    .C(_2600_),
    .Y(_2617_)
);

NAND2X1 _9449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2237_),
    .Y(_2259_)
);

OAI21X1 _9029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1856_),
    .C(_1857_),
    .Y(_1858_)
);

FILL FILL257550x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14589_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6231_),
    .B(_6232_),
    .Y(_6233_)
);

DFFPOSX1 _13447_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5047_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [6])
);

NAND2X1 _13027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5449_),
    .Y(_5493_)
);

FILL FILL_0__14103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10023_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7935_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.Xcalc [6])
);

NAND2X1 _7515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_240_),
    .Y(_501_)
);

FILL FILL_1__12655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9662_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4494_),
    .B(_4497_),
    .Y(_4498_)
);

FILL FILL_0__9242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11228_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [10]),
    .B(_3510__bF$buf2),
    .Y(_4136_)
);

FILL FILL_1__7677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14447_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5196_),
    .C(_5197_),
    .Y(_5198_)
);

FILL FILL_1__14801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8893_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_891_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[1].u_ce.Yin12b [6])
);

NAND2X1 _8473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(_1370_),
    .Y(_1372_)
);

FILL FILL_0_CLKBUF1_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(_921_),
    .C(_969_),
    .Y(\genblk1[1].u_ce.X_ [1])
);

FILL FILL_0_CLKBUF1_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13193_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5362_),
    .B(_5336_),
    .C(_5361_),
    .Y(_5363_)
);

FILL FILL_0__12186_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4282_),
    .B(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_5000_)
);

OAI21X1 _12051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4607_),
    .B(_4610_),
    .C(_4417_),
    .Y(_4611_)
);

FILL FILL_2__12513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_2464_),
    .C(_2467_),
    .Y(_2472_)
);

NAND3X1 _9258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2035_),
    .B(_2057_),
    .C(_2043_),
    .Y(_2077_)
);

FILL FILL_1__11926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_5999_),
    .Y(_6050_)
);

OAI21X1 _13256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_5711_)
);

FILL FILL_2__13718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10252_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_704_),
    .C(_703_),
    .Y(_717_)
);

NAND3X1 _7324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_289_),
    .C(_317_),
    .Y(_318_)
);

FILL FILL_1__12884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9471_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4315_),
    .B(_4314_),
    .Y(\genblk1[5].u_ce.X_ [0])
);

FILL FILL_0__11457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11037_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .Y(_3959_)
);

OAI21X1 _8949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1764_),
    .B(_1781_),
    .C(_1782_),
    .Y(_1783_)
);

NAND3X1 _8529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf1),
    .B(_1424_),
    .C(_1421_),
    .Y(_1425_)
);

MUX2X1 _8109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .B(_1020_),
    .S(_973__bF$buf4),
    .Y(_1024_)
);

FILL FILL_1__7486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5375_),
    .B(_5397_),
    .C(_5383_),
    .Y(_5417_)
);

OAI21X1 _12527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4911_),
    .B(_5000_),
    .C(_4265_),
    .Y(_4258_)
);

NAND2X1 _12107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4633_),
    .B(_4650_),
    .Y(_4664_)
);

FILL FILL_1__14610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9212_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1188_),
    .C(_1187_),
    .Y(_1189_)
);

FILL FILL_1__10950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7555_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4747_),
    .C(_4775_),
    .Y(_4829_)
);

FILL FILL_2__12322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [9]),
    .B(_1834__bF$buf4),
    .Y(_2295_)
);

NAND2X1 _9067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1892_),
    .B(_1893_),
    .Y(_1894_)
);

FILL FILL_1__11735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10308_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13485_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5085_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Ain12b [8])
);

AOI22X1 _13065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5142_),
    .B(_5174__bF$buf3),
    .C(_5529_),
    .D(_5172_),
    .Y(_5044_)
);

FILL FILL_2__9701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10061_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7973_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_57_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin1 [0])
);

NAND2X1 _7553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_525_),
    .Y(_537_)
);

INVX8 _7133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_135_)
);

FILL FILL_1__12693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12273_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [8]),
    .Y(_4534_)
);

FILL FILL_2__9298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9280_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_4162_),
    .C(_4164_),
    .Y(_3396_)
);

FILL FILL_0__11266_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3776_)
);

NOR2X1 _8758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1635_),
    .B(_1636_),
    .Y(_1637_)
);

OAI21X1 _8338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .B(_1185_),
    .C(_1238_),
    .Y(_1243_)
);

FILL FILL_1__7295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13058_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5232_),
    .B(_5233_),
    .Y(_5234_)
);

INVX1 _12336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4880_),
    .Y(_4881_)
);

FILL FILL_0__13832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9021_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(vdd),
    .C(_973__bF$buf4),
    .Y(_1006_)
);

DFFPOSX1 _14902_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6793_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [6])
);

FILL FILL_0__14617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7784_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2112_),
    .Y(_2113_)
);

FILL FILL_1__11964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8551_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.Xcalc [5]),
    .C(_3441_),
    .D(\genblk1[4].u_ce.Xcalc [7]),
    .Y(_3481_)
);

FILL FILL_0__8131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10117_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3124_),
    .B(_3122_),
    .C(_3117_),
    .Y(_3125_)
);

NAND2X1 _13294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5746_),
    .Y(_5747_)
);

FILL FILL_2__9510_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(_587_),
    .C(_590_),
    .Y(_591_)
);

FILL FILL_2__13756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4187_),
    .B(_3435_),
    .C(_3429_),
    .Y(_3422_)
);

OAI21X1 _14499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6565_),
    .C(_6759_),
    .Y(_6536_)
);

OR2X2 _14079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6433_),
    .B(_6431_),
    .Y(_6435_)
);

FILL FILL_0__10290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8712_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_749_),
    .Y(_752_)
);

NAND3X1 _7362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_354_),
    .C(_351_),
    .Y(_355_)
);

FILL FILL_1__12082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11495_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(\genblk1[5].u_ce.Xin12b [6]),
    .S(vdd),
    .Y(_4351_)
);

FILL FILL_0__11075_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3992_),
    .B(_3994_),
    .Y(_3995_)
);

FILL FILL_1__9917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11822_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1815_),
    .C(_1816_),
    .Y(_1817_)
);

INVX1 _8567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .Y(_1461_)
);

OR2X2 _8147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1059_),
    .B(_1057_),
    .Y(_1060_)
);

FILL FILL_1__10815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5452_),
    .Y(_5453_)
);

DFFPOSX1 _12565_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4219_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [4])
);

OR2X2 _12145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4700_),
    .B(_4685_),
    .Y(_4701_)
);

FILL FILL_0__13641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14426_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6934_)
);

FILL FILL_0__14006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8360_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_2597_),
    .C(_3328_),
    .Y(_2560_)
);

FILL FILL_0__10346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .Y(_2942_)
);

OAI21X1 _7838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_799_),
    .C(_801_),
    .Y(_38_)
);

NAND2X1 _7418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [11]),
    .B(_158__bF$buf1),
    .Y(_408_)
);

FILL FILL_2__13985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9565_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4403_),
    .B(_4404_),
    .Y(_4405_)
);

FILL FILL_0__9145_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _11416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3432_),
    .B(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .C(_4044_),
    .D(_4046_),
    .Y(_3379_)
);

FILL FILL_0__12912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8101_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_530_),
    .Y(_574_)
);

FILL FILL_1__14704_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _7171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_172_)
);

FILL FILL_1__9726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9306_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1660_)
);

NAND2X1 _8376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1271_),
    .Y(_1279_)
);

FILL FILL_1__10624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5247_),
    .B(_5264_),
    .C(_5265_),
    .Y(_5270_)
);

OR2X2 _12374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4915_),
    .B(_4911_),
    .Y(_4916_)
);

FILL FILL_0__12089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8416_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6319_),
    .B(_6320_),
    .C(_5930_),
    .Y(_6359_)
);

AOI21X1 _13579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5956_),
    .B(_5935_),
    .C(_5926__bF$buf4),
    .Y(_5957_)
);

INVX1 _13159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5619_)
);

FILL FILL_0__14655_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14520_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6508_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Ycalc [8])
);

FILL FILL_0__14235_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5889_),
    .B(_5892_),
    .Y(_6454_)
);

FILL FILL_1__11582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10995_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(_3516_),
    .Y(_3517_)
);

FILL FILL_0__10575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3154_),
    .B(_3156_),
    .Y(_3161_)
);

INVX1 _10020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .Y(_2760_)
);

NAND3X1 _7647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(_625_),
    .C(_626_),
    .Y(_627_)
);

AOI21X1 _7227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_225_),
    .C(_160_),
    .Y(_226_)
);

FILL FILL_2__13794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9374_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11645_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3385_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[4].u_ce.Acalc [8])
);

AOI21X1 _11225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3846_),
    .B(_3861_),
    .C(_3859_),
    .Y(_3866_)
);

FILL FILL_0__12721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11020_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1094_),
    .C(_1095_),
    .Y(_1096_)
);

FILL FILL_1__10853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4731_),
    .B(_4736_),
    .Y(_4737_)
);

FILL FILL_2__12645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8645_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3570_),
    .B(_3567_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3571_)
);

FILL FILL_0__8225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(_5804_),
    .Y(_5821_)
);

FILL FILL_0__14464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8806_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(_807_),
    .Y(_824_)
);

OAI21X1 _7456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_439_),
    .C(_423_),
    .Y(_13_)
);

FILL FILL_1__12176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11589_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4441_),
    .B(_4422_),
    .C(_4350_),
    .Y(_4442_)
);

FILL FILL_0__9183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4072_),
    .Y(_4082_)
);

NAND3X1 _11034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3674_),
    .B(_3680_),
    .C(_3683_),
    .Y(_3684_)
);

FILL FILL_0__12950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10909_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2401_),
    .B(_2397_),
    .Y(_2402_)
);

NAND2X1 _12659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5141_),
    .B(_5140_),
    .Y(\genblk1[6].u_ce.X_ [0])
);

OAI21X1 _12239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4755_),
    .B(_4785_),
    .C(_4781_),
    .Y(_4790_)
);

FILL FILL_1__14742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13735_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5977_),
    .B(_5970_),
    .S(_5925__bF$buf2),
    .Y(_5978_)
);

FILL FILL_0__13315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10242_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7010_),
    .B(_7011_),
    .C(_7021_),
    .Y(_7022_)
);

FILL FILL_2__7687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12034_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [8]),
    .Y(_2020_)
);

FILL FILL_1__11867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x111750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8034_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10725_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2551_),
    .CLK(clk_bF$buf50),
    .Q(\genblk1[3].u_ce.Xin12b [10])
);

OAI21X1 _10305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2990_),
    .C(_3031_),
    .Y(_3032_)
);

OAI21X1 _13197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5573_),
    .C(_5601_),
    .Y(_5655_)
);

FILL FILL_0__11801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10520_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_135__bF$buf4),
    .C(_154_),
    .Y(_662_)
);

OAI21X1 _7265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf3),
    .B(_260_),
    .C(_261_),
    .Y(_262_)
);

DFFPOSX1 _11683_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3423_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[4].u_ce.Ain0 [0])
);

FILL FILL_0__11398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .B(_3901_),
    .Y(_3903_)
);

FILL FILL_0__7725_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9831_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1743_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Ain12b [4])
);

FILL FILL_0__7305_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2222_),
    .Y(_2223_)
);

INVX1 _12888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [8]),
    .Y(_5360_)
);

OAI21X1 _12468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4992_),
    .B(_4997_),
    .C(_4998_),
    .Y(_4231_)
);

INVX1 _12048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4607_),
    .Y(_4608_)
);

FILL FILL_1__14131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6842_),
    .B(_6845_),
    .Y(_6846_)
);

FILL FILL_2__7496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8683_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3607_)
);

FILL FILL_0__8263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10669_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [6]),
    .B(_2672__bF$buf1),
    .Y(_3247_)
);

FILL FILL_0__10249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2846_),
    .B(_2849_),
    .Y(_2850_)
);

FILL FILL256950x93750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9468_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(_4311_),
    .C(_4312_),
    .Y(_4313_)
);

FILL FILL_0__9048_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3911_),
    .B(_3940_),
    .C(_3913_),
    .Y(_3956_)
);

FILL FILL_1__13822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14607_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_480_),
    .Y(_481_)
);

NOR2X1 _7074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_81_),
    .Y(_82_)
);

INVX1 _11492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4117_)
);

INVX1 _11072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3710_),
    .Y(_3720_)
);

FILL FILL_1__9629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11534_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1583_),
    .Y(_1584_)
);

INVX1 _8279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1186_)
);

FILL FILL_1__10947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7534_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2428_),
    .B(_2436_),
    .C(_1834__bF$buf1),
    .Y(_2438_)
);

FILL FILL_0__7114_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2039_),
    .B(_2011_),
    .Y(_2040_)
);

MUX2X1 _12697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(\genblk1[6].u_ce.Xin12b [6]),
    .S(gnd),
    .Y(_5177_)
);

NOR2X1 _12277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4804_),
    .Y(_4826_)
);

FILL FILL_1__14780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14558_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7046_),
    .B(_7047_),
    .C(_7056_),
    .D(_7053_),
    .Y(_6786_)
);

FILL FILL_0__14138_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [11]),
    .B(_6635_),
    .Y(_6709_)
);

NOR2X1 _14003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6358_),
    .B(_6362_),
    .Y(_6363_)
);

FILL FILL257250x187350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10478_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10763_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.LoadCtl [2])
);

FILL FILL_0__10058_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3049_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3068_),
    .Y(_2532_)
);

FILL FILL_2__10805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13277_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8911_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_909_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Ain0 [0])
);

FILL FILL_0__9697_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4531_),
    .Y(_4532_)
);

FILL FILL_0__9277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4162_),
    .Y(_4163_)
);

OAI21X1 _11128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3771_),
    .B(_3773_),
    .C(_3582_),
    .Y(_3774_)
);

FILL FILL_1__13631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(_1002_),
    .Y(_1003_)
);

FILL FILL_1__10336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7343_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4512_),
    .C(_4643_),
    .Y(_4644_)
);

FILL FILL_2__8722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8548_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [3]),
    .Y(_3478_)
);

FILL FILL_0__8128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14367_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6879_),
    .B(_6876_),
    .Y(_6880_)
);

NAND2X1 _14232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [5]),
    .Y(_6548_)
);

FILL FILL_1__7504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3642_),
    .B(_3627_),
    .C(_3579_),
    .Y(_3644_)
);

NOR2X1 _10572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3282_),
    .B(_3281_),
    .Y(_3283_)
);

FILL FILL_0__10287_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2885_),
    .Y(_2886_)
);

FILL FILL_1__8709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9260_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_749_),
    .Y(_750_)
);

NOR2X1 _7359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_323_),
    .Y(_352_)
);

FILL FILL_2__13086_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1602_),
    .Y(_1603_)
);

INVX1 _8300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .Y(_1206_)
);

FILL FILL_1__12499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12079_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _11777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4348_)
);

FILL FILL_0__9086_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3991_),
    .Y(_3992_)
);

FILL FILL_1__13860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2668_),
    .C(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .Y(_2669_)
);

NOR2X1 _9505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2290_),
    .Y(_2312_)
);

FILL FILL_1__8462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14225_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6285_),
    .Y(_6286_)
);

FILL FILL_0__13638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5885_),
    .Y(_5886_)
);

FILL FILL_1__9667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10145_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833__bF$buf1),
    .B(_6931_),
    .Y(_6932_)
);

FILL FILL_0__7572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert100 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert101 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert102 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert103 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert104 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert105 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert106 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert107 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8357_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_3327_)
);

NAND2X1 _10208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2939_)
);

FILL FILL_1__12711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14596_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14881_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6772_),
    .CLK(clk_bF$buf50),
    .Q(\u_pa.acc_reg [5])
);

NAND2X1 _14461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [5]),
    .B(_6737_),
    .Y(_6739_)
);

NAND3X1 _14041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf0),
    .B(_6398_),
    .C(_6395_),
    .Y(_6399_)
);

FILL FILL_1__7733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(_3101_),
    .C(_3104_),
    .Y(_3105_)
);

FILL FILL_1__8938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10003_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_570_),
    .Y(_571_)
);

NAND3X1 _7168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf2),
    .B(_168_),
    .C(_167_),
    .Y(_169_)
);

NAND2X1 _11586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [0]),
    .B(_4151_),
    .Y(_4183_)
);

NAND2X1 _11166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf0),
    .B(_3809_),
    .Y(_3810_)
);

FILL FILL_0__12662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7628_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Y_ [0]),
    .Y(_2505_)
);

FILL FILL_0__7208_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1998_),
    .C(_2129_),
    .Y(_2130_)
);

FILL FILL_1__8691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13867_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6103_),
    .B(_6099_),
    .C(_5951_),
    .Y(_6104_)
);

FILL FILL_0__13027_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5756_),
    .B(_5764_),
    .Y(_5765_)
);

FILL FILL_1__9896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10374_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14517_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6505_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Ycalc [5])
);

FILL FILL_0__7381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11999_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_767_),
    .Y(_769_)
);

FILL FILL_1__11579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8586_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .B(\genblk1[4].u_ce.Xin12b [4]),
    .S(gnd),
    .Y(_3514_)
);

FILL FILL_0__8166_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3156_),
    .B(_3154_),
    .Y(_3158_)
);

OAI21X1 _10017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf0),
    .B(_2753_),
    .C(_2756_),
    .Y(_2757_)
);

FILL FILL_1__12940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6912_),
    .B(_6909_),
    .C(_6914_),
    .Y(_6915_)
);

OAI21X1 _14270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf4),
    .B(_6575_),
    .C(_6576_),
    .Y(_6490_)
);

FILL FILL_1__7542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x122550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [11]),
    .B(_2672__bF$buf3),
    .Y(_2922_)
);

FILL FILL_1__8747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10232_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_375_),
    .C(_387_),
    .Y(_388_)
);

AND2X2 _11395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4026_),
    .B(_4024_),
    .Y(_4027_)
);

FILL FILL_2__11857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7857_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .S(vdd),
    .Y(_2706_)
);

FILL FILL_0__7437_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_2347_)
);

NAND2X1 _9123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1947_),
    .B(_1944_),
    .Y(_1948_)
);

FILL FILL_1__8080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14263_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6305_),
    .B(_6322_),
    .Y(_6323_)
);

FILL FILL_0__13676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13256_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5918_),
    .B(_5919_),
    .C(_5920_),
    .Y(_5921_)
);

NAND2X1 _13121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5582_),
    .B(_5581_),
    .Y(_5583_)
);

FILL FILL_1__9285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10183_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6962_),
    .B(_6965_),
    .Y(_6967_)
);

NOR2X1 _14326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .Y(_6625_)
);

FILL FILL_0__7190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8395_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [0]),
    .Y(_3347_)
);

MUX2X1 _10246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2971_),
    .B(_2968_),
    .S(_2649__bF$buf1),
    .Y(_2976_)
);

FILL FILL_0__11742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [0]),
    .B(_1637_),
    .Y(_1669_)
);

FILL FILL_1__7771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12947_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5287_),
    .B(_5284_),
    .Y(_5288_)
);

FILL FILL_0__12527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7666_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9772_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1684_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Ycalc [7])
);

FILL FILL_0__7246_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2166_),
    .B(_2149_),
    .Y(_2167_)
);

FILL FILL_1__11600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14072_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6114_),
    .B(_6118_),
    .Y(_6140_)
);

OAI21X1 _13350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5340_),
    .B(_5796_),
    .C(_5798_),
    .Y(_5060_)
);

FILL FILL_0__13065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12805_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14555_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6536_),
    .CLK(clk_bF$buf51),
    .Q(\u_ot.ISreg )
);

INVX1 _14135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6475_)
);

FILL FILL_1__7827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x198150 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3550_),
    .B(_3551_),
    .Y(_3552_)
);

NAND2X1 _10475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3192_),
    .B(_3191_),
    .Y(_3193_)
);

INVX1 _10055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .Y(_2793_)
);

FILL FILL_0__11971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11131_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1510_),
    .Y(_1513_)
);

OAI21X1 _8203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1110_),
    .B(_1092_),
    .C(_1109_),
    .Y(_1113_)
);

FILL FILL_1__7580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12756_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5107_)
);

FILL FILL_0__12336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4750_),
    .B(_4753_),
    .Y(_4754_)
);

DFFPOSX1 _9828_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1740_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Ain12b [9])
);

NOR2X1 _9408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2175_),
    .Y(_2220_)
);

FILL FILL_1__8785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14128_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6188_),
    .B(_6184_),
    .Y(_6194_)
);

INVX1 _13406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [0]),
    .Y(_5830_)
);

FILL FILL_2__11475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7475_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2382_),
    .B(_2373_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2383_)
);

NAND2X1 _9161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1980_),
    .B(_1983_),
    .Y(_1984_)
);

FILL FILL_0__10822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14499_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6957_),
    .B(_7000_),
    .Y(_7001_)
);

FILL FILL_0__14079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin1 [1]),
    .B(_6657_),
    .Y(_6658_)
);

FILL FILL_1__7636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13819_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3011_),
    .B(_2968_),
    .S(vdd),
    .Y(_3012_)
);

FILL FILL_0__11780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11360_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8852_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_850_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Ycalc [11])
);

OAI21X1 _8432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1327_),
    .B(_1311_),
    .C(_1325_),
    .Y(_1332_)
);

OAI21X1 _8012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [11]),
    .C(_924_),
    .Y(_933_)
);

AOI22X1 _11489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4103_),
    .B(_3510__bF$buf0),
    .C(_4113_),
    .D(_4114_),
    .Y(_3384_)
);

AND2X2 _11069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3656_),
    .B(_3659_),
    .Y(_3717_)
);

FILL FILL_1__13992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12985_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5320_),
    .B(_5323_),
    .Y(_5324_)
);

FILL FILL_0__12145_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4964_),
    .B(_4959_),
    .C(_4957_),
    .Y(_4968_)
);

AND2X2 _12010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4559_),
    .B(_4571_),
    .Y(_4572_)
);

NAND2X1 _9637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2429_),
    .B(_2432_),
    .Y(_2435_)
);

OAI21X1 _9217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2023_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_)
);

FILL FILL_1__8594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x93750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin1 [0]),
    .B(_6006_),
    .C(_6009_),
    .Y(_6011_)
);

NAND2X1 _13215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf2),
    .B(_5659_),
    .Y(_5672_)
);

FILL FILL_0__14711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(_2202_),
    .C(_2200_),
    .Y(_2203_)
);

FILL FILL_2_BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12489_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_677_),
    .Y(_679_)
);

FILL FILL_2__13010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9448_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(\genblk1[5].u_ce.LoadCtl [3]),
    .Y(_4279_)
);

FILL FILL_0__11416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9010_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _14593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .Y(_6833_)
);

DFFPOSX1 _14173_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5849_),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.Xcalc [1])
);

DFFPOSX1 _8908_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_906_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Ain12b [5])
);

FILL FILL_1__7865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5363_),
    .B(_5376_),
    .C(_5377_),
    .Y(_5378_)
);

FILL FILL_1_BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [7]),
    .Y(_2829_)
);

INVX1 _8661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [4]),
    .Y(_1548_)
);

NAND2X1 _8241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1149_),
    .Y(_1150_)
);

NOR2X1 _11298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf1),
    .B(_3763_),
    .Y(_3936_)
);

FILL FILL_1__13381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12374_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.Acalc [1]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Acalc [3]),
    .Y(_2615_)
);

OAI21X1 _9446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2256_),
    .Y(_1695_)
);

MUX2X1 _9026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1854_),
    .B(_1851_),
    .S(_1811__bF$buf4),
    .Y(_1855_)
);

FILL FILL_0__8701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13579_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .B(_6229_),
    .Y(_6230_)
);

FILL FILL_0__13159_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13444_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5044_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Xcalc [3])
);

NAND2X1 _13024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .B(_5476_),
    .Y(_5490_)
);

FILL FILL_2__13906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10086_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6877_)
);

NAND2X1 _14229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(\u_ot.Xcalc [4]),
    .Y(_6546_)
);

FILL FILL_0__7093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12298_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7932_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [3])
);

MUX2X1 _7512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .B(_454_),
    .S(gnd),
    .Y(_498_)
);

INVX1 _10989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3640_),
    .Y(_3641_)
);

FILL FILL_0__8298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [8]),
    .B(_3215_),
    .C(_3279_),
    .Y(_3280_)
);

AOI21X1 _10149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2881_),
    .B(_2869_),
    .C(_2882_),
    .Y(_2883_)
);

FILL FILL_1__12652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9677_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf0),
    .B(_4491_),
    .C(_4486_),
    .Y(_4495_)
);

FILL FILL_2__9257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11225_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4130_),
    .B(_4133_),
    .Y(_4134_)
);

AOI22X1 _8717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1589_),
    .B(_996__bF$buf3),
    .C(_1599_),
    .D(_1600_),
    .Y(_870_)
);

FILL FILL_1__7674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x237750 (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5194_),
    .B(_5191_),
    .S(_5151__bF$buf3),
    .Y(_5195_)
);

FILL FILL_1__8459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9400_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8890_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_888_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[1].u_ce.Yin12b [11])
);

NAND2X1 _8470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1368_),
    .Y(_1369_)
);

AOI22X1 _8050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.Xcalc [5]),
    .C(_927_),
    .D(\genblk1[1].u_ce.Xcalc [7]),
    .Y(_967_)
);

FILL FILL_1__13190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7569_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_2464_),
    .C(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2470_)
);

FILL FILL_0__7149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2069_),
    .B(_2073_),
    .Y(_2074_)
);

FILL FILL_1__11923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [10]),
    .Y(_6047_)
);

INVX1 _13253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain1 [1]),
    .Y(_5708_)
);

FILL FILL_2__13715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9715_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14878_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6769_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [2])
);

NAND3X1 _14458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [2]),
    .B(_6718_),
    .C(_6736_),
    .Y(_6737_)
);

INVX1 _14038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6309_),
    .Y(_6396_)
);

FILL FILL_2__8281_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_713_),
    .B(_710_),
    .Y(_714_)
);

INVX1 _7321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [7]),
    .Y(_315_)
);

OAI21X1 _10798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3456_),
    .B(_3459_),
    .C(_3444_),
    .Y(_3460_)
);

INVX1 _10378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3100_),
    .Y(_3102_)
);

FILL FILL_1__12881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11034_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_1778_),
    .C(_1779_),
    .Y(_1780_)
);

NOR2X1 _8526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf3),
    .B(_1249_),
    .Y(_1422_)
);

INVX1 _8106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .Y(_1021_)
);

FILL FILL_1__7483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13246_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5409_),
    .B(_5413_),
    .Y(_5414_)
);

FILL FILL_0__12659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [0]),
    .B(_5000_),
    .Y(_4264_)
);

OAI21X1 _12104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348__bF$buf0),
    .B(_4661_),
    .C(_4635_),
    .Y(_4204_)
);

FILL FILL_0__13600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8268_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6100_),
    .B(_6079_),
    .Y(_6101_)
);

INVX1 _13309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5761_),
    .Y(_5762_)
);

FILL FILL_0__14805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2290_),
    .Y(_2293_)
);

NAND2X1 _9064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1889_),
    .B(_1890_),
    .Y(_1891_)
);

FILL FILL_1__11732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13197_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13482_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5082_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin0 [1])
);

OR2X2 _13062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .B(_5511_),
    .Y(_5527_)
);

FILL FILL_2__13944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9104_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6911_),
    .B(_6868_),
    .C(_6877_),
    .Y(_6912_)
);

OAI21X1 _14267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6573_),
    .C(_6570_),
    .Y(_6574_)
);

FILL FILL_1__7539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14309_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7970_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_54_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin12b [7])
);

AOI22X1 _7550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_158__bF$buf0),
    .C(_534_),
    .D(_156_),
    .Y(_17_)
);

INVX1 _7130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [0]),
    .Y(_132_)
);

OAI21X1 _10187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2917_),
    .B(_2919_),
    .C(_2741_),
    .Y(_2920_)
);

FILL FILL_1__12690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11263_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996__bF$buf2),
    .B(_1634_),
    .C(_1633_),
    .Y(_874_)
);

AOI21X1 _8335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .B(_1238_),
    .C(_1236_),
    .Y(_1240_)
);

FILL FILL_1__7292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12888_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5229_),
    .B(_5230_),
    .Y(_5231_)
);

FILL FILL_0__12468_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain1 [0]),
    .B(_4877_),
    .Y(_4878_)
);

FILL FILL_0__12048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6316_),
    .C(_6311_),
    .Y(_6320_)
);

NOR2X1 _13538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Xcalc [11]),
    .Y(_5918_)
);

NAND2X1 _13118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(_5579_),
    .Y(_5580_)
);

FILL FILL257250x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7187_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_2110_)
);

FILL FILL_1__11961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10114_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5741_),
    .B(_5726_),
    .C(_5743_),
    .Y(_5744_)
);

INVX1 _7606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .Y(_588_)
);

FILL FILL_1__12746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_3428_)
);

NAND2X1 _14496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.Y_ [1]),
    .Y(_6758_)
);

OR2X2 _14076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6395_),
    .B(_6397_),
    .Y(_6432_)
);

FILL FILL_1__7768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14118_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5279_),
    .B(_5280_),
    .Y(_5285_)
);

FILL FILL_2__10458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1812_),
    .C(_1813_),
    .Y(_1814_)
);

NOR2X1 _8564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1455_),
    .B(_1440_),
    .Y(_1458_)
);

AOI21X1 _8144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .B(_1053_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1057_)
);

FILL FILL_1__10812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5450_)
);

FILL FILL_0__12697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12277_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12562_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4216_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Acalc [1])
);

INVX1 _12142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4697_),
    .Y(_4698_)
);

DFFPOSX1 _9769_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1681_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Ycalc [4])
);

INVX1 _9349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .Y(_2164_)
);

FILL FILL_0__8604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6099_),
    .B(_6127_),
    .Y(_6137_)
);

NAND2X1 _13347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5796_),
    .Y(_5797_)
);

FILL FILL_0__14843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10343_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_799_),
    .Y(_800_)
);

OAI21X1 _7415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .B(_405_),
    .C(_227_),
    .Y(_406_)
);

FILL FILL_2__13982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11548_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _11833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4401_),
    .B(_4352_),
    .C(_4400_),
    .D(_4344_),
    .Y(_4402_)
);

FILL FILL_0__9142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4043_),
    .B(_4036_),
    .Y(_4044_)
);

FILL FILL_1__7997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14347_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5103_),
    .Y(_5104_)
);

FILL FILL_1__14701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9303_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1658_)
);

AND2X2 _8373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(_1275_),
    .Y(_1276_)
);

FILL FILL_1__10621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13093_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5267_),
    .B(_5248_),
    .C(_5176_),
    .Y(_5268_)
);

OAI21X1 _12371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(_4344_),
    .Y(_4913_)
);

FILL FILL_0__12086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12413_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2735_),
    .C(_2721_),
    .Y(_2739_)
);

NAND2X1 _9578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2374_),
    .B(_2378_),
    .Y(_2380_)
);

NAND3X1 _9158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf4),
    .B(_1977_),
    .C(_1972_),
    .Y(_1981_)
);

FILL FILL_1__11826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(_6355_),
    .Y(_6356_)
);

MUX2X1 _13576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5953_),
    .B(_5952_),
    .S(_5926__bF$buf2),
    .Y(_5954_)
);

OAI21X1 _13156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5611_),
    .C(_5607_),
    .Y(_5616_)
);

FILL FILL_2__13618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10152_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .B(_604_),
    .C(_172__bF$buf0),
    .Y(_624_)
);

NOR2X1 _7224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_222_),
    .Y(_223_)
);

FILL FILL_1__12784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11357_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11642_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3382_),
    .CLK(clk_bF$buf38),
    .Q(\genblk1[4].u_ce.Acalc [5])
);

NAND2X1 _11222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3847_),
    .B(_3862_),
    .Y(_3864_)
);

DFFPOSX1 _8849_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_847_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Ycalc [8])
);

NOR2X1 _8429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1328_),
    .Y(_1330_)
);

AOI22X1 _8009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Acalc [0]),
    .C(_929_),
    .D(_930_),
    .Y(_931_)
);

FILL FILL_1__7386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf5),
    .B(_5317_),
    .C(_5312_),
    .Y(_5321_)
);

NAND2X1 _12427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4959_),
    .B(_4964_),
    .Y(_4966_)
);

OAI21X1 _12007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4561_),
    .C(_4563_),
    .Y(_4569_)
);

FILL FILL_0__13923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9112_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1093_)
);

FILL FILL_1__10850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7455_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4692_),
    .B(_4689_),
    .Y(_4734_)
);

FILL FILL_2__12222_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .B(_2197_),
    .Y(_2200_)
);

FILL FILL_1__11215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8642_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3565_),
    .Y(_3568_)
);

FILL FILL_0__8222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10208_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5800_),
    .C(_5819_),
    .Y(_5074_)
);

FILL FILL_2__9601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_803_),
    .C(_822_),
    .Y(_52_)
);

NAND2X1 _7453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_441_),
    .Y(_442_)
);

FILL FILL_1__12173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11586_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4437_),
    .B(_4434_),
    .C(_4423_),
    .Y(_4439_)
);

FILL FILL_2__9198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11166_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4073_),
    .B(_4077_),
    .Y(_4079_)
);

INVX1 _11031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .Y(_3681_)
);

AOI21X1 _8658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1535_),
    .B(_1544_),
    .C(_1545_),
    .Y(_1546_)
);

AOI21X1 _8238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1103_),
    .B(_1105_),
    .C(_1093_),
    .Y(_1147_)
);

FILL FILL_1__7195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5137_),
    .C(_5138_),
    .Y(_5139_)
);

INVX1 _12236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4785_),
    .Y(_4788_)
);

FILL FILL_0__13732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9341_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7005_),
    .B(_7006_),
    .Y(_7019_)
);

FILL FILL_2__7684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12031_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .Y(_2018_)
);

FILL FILL_1__11864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8451_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10722_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2548_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Acalc [9])
);

FILL FILL_0__8031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10017_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_3029_)
);

NOR2X1 _13194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5630_),
    .Y(_5652_)
);

FILL FILL_2__9410_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7929_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xcalc [0])
);

INVX1 _7509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_495_)
);

FILL FILL_2__13656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9656_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4472_),
    .B(_4467_),
    .C(_4362__bF$buf0),
    .Y(_4492_)
);

FILL FILL_0__9236_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf4),
    .B(\genblk1[4].u_ce.Ain12b [9]),
    .Y(_4131_)
);

NAND2X1 _14399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6673_),
    .B(_6687_),
    .Y(_6688_)
);

FILL FILL_0__10190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8612_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .B(_659_),
    .Y(_660_)
);

NAND2X1 _7262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf3),
    .B(_208_),
    .Y(_259_)
);

FILL FILL_0__11395_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11680_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3420_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[4].u_ce.Ain12b [5])
);

AOI21X1 _11260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3895_),
    .B(_3899_),
    .C(_3528_),
    .Y(_3900_)
);

FILL FILL_2__11722_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8887_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_885_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Xin0 [0])
);

OR2X2 _8467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1358_),
    .Y(_1366_)
);

INVX1 _8047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [3]),
    .Y(_964_)
);

FILL FILL_0__7722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13187_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5357_),
    .Y(_5358_)
);

OAI21X1 _12465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4995_),
    .B(_4993_),
    .C(_4996_),
    .Y(_4230_)
);

NAND2X1 _12045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4604_),
    .B(_4580_),
    .Y(_4605_)
);

FILL FILL_0__13961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6840_),
    .B(_6841_),
    .Y(_6843_)
);

FILL FILL_2__12260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert390 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert391 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8698_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3584_),
    .B(_3603_),
    .C(_3604_),
    .Y(_3605_)
);

FILL FILL_0__8260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10666_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3243_),
    .B(_3234_),
    .Y(_3245_)
);

FILL FILL_0__10246_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf2),
    .B(_2843_),
    .C(_2837_),
    .Y(_2847_)
);

AOI21X1 _7738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(gnd),
    .C(_172__bF$buf5),
    .Y(_711_)
);

AOI21X1 _7318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_308_),
    .C(_160_),
    .Y(_313_)
);

FILL FILL_2__13885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9465_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4308_),
    .C(_4309_),
    .Y(_4310_)
);

FILL FILL_0__9045_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3919_),
    .B(_3947_),
    .Y(_3953_)
);

FILL FILL_0__12812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14604_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf2),
    .B(_476_),
    .C(_477_),
    .Y(_478_)
);

FILL FILL_1__9626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9206_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(_1579_),
    .Y(_1581_)
);

OAI21X1 _8276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1174_),
    .C(_1173_),
    .Y(_1183_)
);

FILL FILL_1__10944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10104_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf3 )
);

FILL FILL_0__7531_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf2 )
);

FILL FILL_0__7111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7129_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf0 )
);

INVX8 _12694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .Y(_5174_)
);

INVX1 _12274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [10]),
    .Y(_4823_)
);

FILL FILL_2__12736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [2]),
    .B(_5949__bF$buf2),
    .Y(_6263_)
);

DFFPOSX1 _13479_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5079_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin1 [0])
);

INVX1 _13059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5523_),
    .Y(_5524_)
);

AOI21X1 _14840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7034_),
    .B(_7038_),
    .C(_7036_),
    .Y(_7054_)
);

FILL FILL_0__14135_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [11]),
    .B(_6562__bF$buf3),
    .Y(_6706_)
);

NOR2X1 _14000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6359_),
    .B(_6339_),
    .Y(_6360_)
);

FILL FILL_1__11482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10895_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10760_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2586_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[3].u_ce.Ain0 [1])
);

FILL FILL_0__10475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10055_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3065_),
    .B(_3050_),
    .Y(_3066_)
);

DFFPOSX1 _7967_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_51_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin12b [8])
);

OR2X2 _7547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_531_),
    .Y(_532_)
);

OAI21X1 _7127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_128_),
    .C(_129_),
    .Y(_130_)
);

FILL FILL_2__13694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9694_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4498_),
    .B(_4502_),
    .C(_4497_),
    .Y(_4529_)
);

FILL FILL_0__9274_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(_4159_),
    .Y(_4161_)
);

NOR3X1 _11125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3761_),
    .B(_3770_),
    .C(_3754_),
    .Y(_3771_)
);

FILL FILL_0__12621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11760_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .B(\genblk1[1].u_ce.Xin12b [4]),
    .S(vdd),
    .Y(_1000_)
);

FILL FILL_1__10333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7340_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4640_),
    .B(_4638_),
    .S(_4325__bF$buf2),
    .Y(_4641_)
);

FILL FILL_2__12965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8545_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3472_),
    .B(_3475_),
    .C(_3444_),
    .Y(_3476_)
);

FILL FILL_0__8125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5736_),
    .B(_5740_),
    .Y(_5741_)
);

FILL FILL_2__9924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10611_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .Y(_747_)
);

OR2X2 _7356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_327_),
    .Y(_349_)
);

FILL FILL_1__12496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11489_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4345_),
    .Y(_4346_)
);

FILL FILL_0__9083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3979_),
    .B(_3981_),
    .C(_3988_),
    .Y(_3989_)
);

FILL FILL_0__12850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7816_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .B(_2664_),
    .Y(_2666_)
);

INVX1 _9502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [10]),
    .Y(_2309_)
);

NAND3X1 _12979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf2),
    .B(_5443_),
    .C(_5446_),
    .Y(_5447_)
);

DFFPOSX1 _12559_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4213_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [10])
);

OR2X2 _12139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4694_),
    .B(_4693_),
    .Y(_4695_)
);

FILL FILL_1__14642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13635_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6283_),
    .B(_6282_),
    .C(_6018_),
    .Y(_6284_)
);

FILL FILL_0__13215_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13500_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[6].u_ce.LoadCtl [5])
);

FILL FILL_1__9664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10142_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6925_),
    .B(_6928_),
    .Y(_6929_)
);

FILL FILL256650x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12774_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .B(_1920_),
    .C(_1909_),
    .Y(_1925_)
);

FILL FILL_1__11767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8354_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .B(_3324_),
    .C(_3325_),
    .Y(_2557_)
);

NAND2X1 _10205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2936_),
    .Y(_2526_)
);

NOR2X1 _13097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518_),
    .B(_5515_),
    .Y(_5560_)
);

FILL FILL_0__11701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10420_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_529_),
    .C(_139_),
    .Y(_568_)
);

AOI21X1 _7165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_144_),
    .C(_135__bF$buf4),
    .Y(_166_)
);

FILL FILL_0__11298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3485_),
    .C(_4181_),
    .Y(_3411_)
);

INVX1 _11163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3806_),
    .Y(_3807_)
);

FILL FILL_1__10618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7625_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .B(_1759_),
    .C(_2503_),
    .Y(_1733_)
);

FILL FILL_0__7205_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2124_),
    .S(_1811__bF$buf2),
    .Y(_2127_)
);

AOI21X1 _12788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5263_),
    .B(_5260_),
    .C(_5249_),
    .Y(_5265_)
);

OAI21X1 _12368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4906_),
    .B(_4907_),
    .C(_4904_),
    .Y(_4910_)
);

FILL FILL_1__14451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14649_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14514_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6502_),
    .CLK(clk_bF$buf9),
    .Q(\u_ot.Ycalc [2])
);

FILL FILL_0__14229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8583_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [1]),
    .B(_3510__bF$buf3),
    .Y(_3511_)
);

FILL FILL_0__8163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10149_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3118_),
    .B(_3120_),
    .Y(_3155_)
);

NOR2X1 _10014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2649__bF$buf0),
    .Y(_2754_)
);

FILL FILL_2__9962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9368_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11639_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3379_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [2])
);

NAND3X1 _11219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3532_),
    .B(_3858_),
    .C(_3857_),
    .Y(_3861_)
);

FILL FILL_1__13722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x187350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8324_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .Y(_385_)
);

AOI21X1 _11392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(vdd),
    .C(_4023_),
    .Y(_4024_)
);

FILL FILL_1__9949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11434_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [11]),
    .B(_996__bF$buf1),
    .Y(_1491_)
);

OAI21X1 _8179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1070_),
    .B(_1089_),
    .C(_1090_),
    .Y(_1091_)
);

FILL FILL_1__10847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7854_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .S(vdd),
    .Y(_2703_)
);

FILL FILL_0__7434_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834__bF$buf2),
    .B(_2343_),
    .C(_2344_),
    .Y(_1701_)
);

NOR2X1 _9120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1940_),
    .Y(_1945_)
);

DFFPOSX1 _12597_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4251_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Ain12b [10])
);

OAI21X1 _12177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf3),
    .B(_4729_),
    .C(_4730_),
    .Y(_4731_)
);

FILL FILL_2__8813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14458_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6964_)
);

FILL FILL_0__14038_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6618_),
    .B(_6562__bF$buf2),
    .C(_6621_),
    .D(_6622_),
    .Y(_6497_)
);

FILL FILL_1__11385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8392_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3303_),
    .B(_3313_),
    .C(_3345_),
    .Y(_2575_)
);

FILL FILL_0__10378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf1),
    .B(_2969_),
    .C(_2972_),
    .Y(_2973_)
);

FILL FILL_2__13177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_971_),
    .C(_1667_),
    .Y(_897_)
);

FILL FILL_0__9597_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .Y(_4436_)
);

FILL FILL_0__9177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4075_),
    .B(_3524__bF$buf2),
    .Y(_4076_)
);

INVX1 _11028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3677_),
    .Y(_3678_)
);

FILL FILL_1__13951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8028_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10719_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2545_),
    .CLK(clk_bF$buf73),
    .Q(\genblk1[3].u_ce.Acalc [6])
);

FILL FILL_1__9091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14687_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14552_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [3]),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.LoadCtl [4])
);

FILL FILL_0__14267_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6176_),
    .B(_6455_),
    .C(_6473_),
    .Y(_5872_)
);

FILL FILL_1__7824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11194_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3548_),
    .B(_3540_),
    .C(_3523_),
    .Y(_3549_)
);

FILL FILL_0__10187_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3189_),
    .B(_3187_),
    .Y(_3190_)
);

INVX1 _10052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_2790_)
);

FILL FILL_1__8609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9160_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_656_),
    .Y(_657_)
);

INVX1 _7259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_256_)
);

AOI21X1 _8620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(gnd),
    .C(_1509_),
    .Y(_1510_)
);

AOI21X1 _8200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(_1110_),
    .C(_998_),
    .Y(_1111_)
);

FILL FILL_1__12399_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11677_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3417_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[4].u_ce.Ain12b [6])
);

NAND3X1 _11257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3834_),
    .B(_3896_),
    .C(_3837_),
    .Y(_3897_)
);

FILL FILL_1__13760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7719_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9825_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1737_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Ain12b [10])
);

OAI21X1 _9405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf3),
    .B(_2215_),
    .C(_2216_),
    .Y(_2217_)
);

FILL FILL_1__8782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13958_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6159_),
    .B(_6168_),
    .C(_6190_),
    .Y(_6191_)
);

FILL FILL_0__13538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13118_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5788_),
    .B(_5796_),
    .C(_5828_),
    .Y(_5083_)
);

FILL FILL_1__9987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10045_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6839_),
    .Y(_6840_)
);

FILL FILL_0__7892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8677_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3601_),
    .Y(_3602_)
);

FILL FILL_0__8257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3241_),
    .B(_3240_),
    .Y(_3242_)
);

OAI21X1 _10108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .B(_2810_),
    .C(_2686__bF$buf2),
    .Y(_2844_)
);

FILL FILL_2__9636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14496_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6993_),
    .B(_6997_),
    .C(_6998_),
    .Y(_6782_)
);

FILL FILL_0__14076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6655_),
    .C(_6653_),
    .Y(_6656_)
);

FILL FILL_1__7633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12809_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3008_),
    .Y(_3009_)
);

FILL FILL_1__8838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8418_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_370_),
    .Y(_475_)
);

NAND2X1 _11486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4111_),
    .B(_4110_),
    .Y(_4112_)
);

AOI22X1 _11066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3696_),
    .B(_3510__bF$buf1),
    .C(_3714_),
    .D(_3694_),
    .Y(_3361_)
);

FILL FILL_2__11948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7528_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2431_),
    .Y(_2432_)
);

FILL FILL_0__7108_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2031_),
    .B(_2034_),
    .Y(_2035_)
);

FILL FILL_1__8591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13767_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5941_),
    .B(_5978_),
    .C(_5963__bF$buf4),
    .Y(_6008_)
);

FILL FILL_0__13347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [11]),
    .B(_5174__bF$buf4),
    .Y(_5669_)
);

FILL FILL_1__9376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_7051_)
);

NAND2X1 _14417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6702_),
    .B(_6703_),
    .Y(_6704_)
);

FILL FILL_2_BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11899_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_675_),
    .B(_673_),
    .Y(_676_)
);

FILL FILL_1__11479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8066_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10757_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2583_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Ain1 [0])
);

INVX1 _10337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3062_),
    .Y(_3063_)
);

FILL FILL_1__12840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256050x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6827_),
    .B(_6830_),
    .Y(_6831_)
);

DFFPOSX1 _14170_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5846_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Ycalc [10])
);

DFFPOSX1 _8905_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_903_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Ain12b [6])
);

FILL FILL_1__7862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5371_),
    .B(_5374_),
    .Y(_5375_)
);

FILL FILL_0__12618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2822_),
    .C(_2674_),
    .Y(_2827_)
);

FILL FILL_1__8647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10132_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_291_),
    .C(_230_),
    .Y(_293_)
);

FILL FILL256650x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [7]),
    .Y(_3933_)
);

FILL FILL_2__11757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7757_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [7]),
    .B(_2603_),
    .Y(_2612_)
);

FILL FILL_0__7337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2249_),
    .B(_2253_),
    .Y(_2254_)
);

INVX1 _9023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1852_)
);

FILL FILL_1__14583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13996_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6226_),
    .B(_6224_),
    .S(_5926__bF$buf4),
    .Y(_6227_)
);

FILL FILL_0__13576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13156_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13441_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5041_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Xcalc [0])
);

FILL FILL256650x150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174__bF$buf3),
    .B(_5487_),
    .C(_5461_),
    .Y(_5042_)
);

FILL FILL_1__9185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10083_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [4]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf1),
    .Y(_6875_)
);

NAND2X1 _14226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(\u_ot.Xcalc [3]),
    .Y(_6544_)
);

FILL FILL_0__7090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11288_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3636_),
    .C(_3637_),
    .Y(_3638_)
);

FILL FILL_0__8295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [8]),
    .B(_2672__bF$buf3),
    .Y(_3277_)
);

NAND3X1 _10146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2846_),
    .B(_2849_),
    .C(_2879_),
    .Y(_2880_)
);

FILL FILL_2__9674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11222_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1597_),
    .B(_1596_),
    .Y(_1598_)
);

FILL FILL_1__7671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12847_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5192_)
);

FILL FILL_0__12427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12007_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2662_),
    .B(_2659_),
    .S(_2649__bF$buf4),
    .Y(_2663_)
);

FILL FILL_1__8456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x198150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14219_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6280_),
    .B(_6279_),
    .Y(_6281_)
);

FILL FILL_2__7320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7566_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .B(_1848__bF$buf1),
    .Y(_2467_)
);

FILL FILL_0__7146_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_1848__bF$buf5),
    .Y(_2071_)
);

FILL FILL_1__11920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13385_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6020_),
    .B(_5949__bF$buf1),
    .C(_6044_),
    .D(_6021_),
    .Y(_5839_)
);

NOR2X1 _13250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [3]),
    .B(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .Y(_5705_)
);

FILL FILL_1__12705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9712_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14875_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6766_),
    .CLK(clk_bF$buf72),
    .Q(\genblk1[0].u_ce.Rdy )
);

NAND2X1 _14455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [7]),
    .B(_6733_),
    .Y(_6735_)
);

AOI21X1 _14035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6392_),
    .B(_6368_),
    .C(_6391_),
    .Y(_6393_)
);

FILL FILL_1__7727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11097_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [4]),
    .Y(_3457_)
);

INVX1 _10375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3098_),
    .Y(_3099_)
);

FILL FILL_0__11871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11031_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .B(_1776_),
    .Y(\a[3] [1])
);

INVX1 _8523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [7]),
    .Y(_1419_)
);

INVX1 _8103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1018_)
);

FILL FILL_1__7480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12656_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5405_),
    .B(_5188__bF$buf1),
    .Y(_5411_)
);

FILL FILL_0__12236_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5023_),
    .B(_4997_),
    .C(_5027_),
    .Y(_4255_)
);

NAND2X1 _12101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4636_),
    .B(_4658_),
    .Y(_4659_)
);

NAND2X1 _9728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2486_),
    .Y(_2502_)
);

OAI21X1 _9308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1909_),
    .C(_2123_),
    .Y(_2124_)
);

FILL FILL_1__8685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14028_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .B(_6096_),
    .C(_6097_),
    .Y(_6098_)
);

OR2X2 _13306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5683_),
    .B(_5188__bF$buf4),
    .Y(_5759_)
);

FILL FILL_0__14802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7375_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2288_),
    .C(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2290_)
);

OAI22X1 _9061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1887_),
    .B(_1838_),
    .C(_1886_),
    .D(_1830_),
    .Y(_1888_)
);

FILL FILL_2__8334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14399_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .B(_6890_),
    .C(_6908_),
    .Y(_6909_)
);

OAI21X1 _14264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .C(\u_ot.ISreg_bF$buf2 ),
    .Y(_6571_)
);

FILL FILL_1__7536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13719_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2911_),
    .B(_2907_),
    .Y(_2917_)
);

FILL FILL_0__11260_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1632_),
    .B(_1631_),
    .C(_1622_),
    .Y(_873_)
);

AOI21X1 _8332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1212_),
    .B(_1214_),
    .C(_1208_),
    .Y(_1237_)
);

NAND2X1 _11389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [1]),
    .B(_3510__bF$buf2),
    .Y(_4021_)
);

FILL FILL_1__13892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12885_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _12750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5227_),
    .B(_5178_),
    .C(_5226_),
    .D(_5170_),
    .Y(_5228_)
);

FILL FILL_0__12465_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4354_),
    .B(_4325__bF$buf3),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4875_)
);

FILL FILL_0__12045_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2699_),
    .B(_2696_),
    .S(_2649__bF$buf2),
    .Y(_2700_)
);

NAND2X1 _9537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2341_),
    .Y(_2342_)
);

NOR2X1 _9117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1910_),
    .Y(_1942_)
);

FILL FILL_1__8494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6316_),
    .C(_6312_),
    .Y(_6317_)
);

FILL FILL_0_BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[7].u_ce.Xcalc [0]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Xcalc [2]),
    .Y(_5916_)
);

FILL FILL_0_BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5536_),
    .B(_5557_),
    .C(_5561_),
    .Y(_5577_)
);

FILL FILL_0_BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7184_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf0),
    .B(_2103_),
    .C(_2106_),
    .Y(_2107_)
);

FILL FILL_2__8983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12389_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .Y(_585_)
);

FILL FILL_0__8389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11316_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4062_),
    .B(_4162_),
    .C(_3426_),
    .Y(_3419_)
);

OAI21X1 _14493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6749_),
    .B(_6740_),
    .C(_6756_),
    .Y(_6533_)
);

OAI21X1 _14073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6393_),
    .B(_6428_),
    .C(_6426_),
    .Y(_6429_)
);

OAI21X1 _8808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1666_)
);

FILL FILL_1__7765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13108_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5259_),
    .B(_5250_),
    .Y(_5282_)
);

FILL FILL257250x244950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9911_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _8981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_1811_)
);

OAI21X1 _8561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1455_),
    .B(_1440_),
    .C(_994_),
    .Y(_1456_)
);

INVX1 _8141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1054_)
);

AOI21X1 _11198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3836_),
    .B(_3838_),
    .C(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3841_)
);

FILL FILL_2__7834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12274_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9766_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1678_),
    .CLK(clk_bF$buf9),
    .Q(\genblk1[2].u_ce.ISout )
);

AOI21X1 _9346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2113_),
    .C(_2139_),
    .Y(_2161_)
);

FILL FILL_0__8601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13899_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6106_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6134_),
    .Y(_5843_)
);

FILL FILL_0__13059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [5]),
    .B(_5105_),
    .Y(_5794_)
);

FILL FILL_2__13806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9088_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14549_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [0]),
    .CLK(clk_bF$buf38),
    .Q(\u_ot.LoadCtl [1])
);

NAND2X1 _14129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.X_ [1]),
    .Y(_6472_)
);

FILL FILL_2__8372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [5]),
    .B(_85_),
    .Y(_797_)
);

AND2X2 _7412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_393_),
    .Y(_403_)
);

MUX2X1 _10889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3545_),
    .B(_3544_),
    .S(_3487__bF$buf3),
    .Y(_3546_)
);

FILL FILL_0__8198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3186_),
    .Y(_3187_)
);

OAI21X1 _10049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2786_),
    .C(_2787_),
    .Y(_2788_)
);

FILL FILL_1__12972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11545_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4398_),
    .B(_4351_),
    .S(gnd),
    .Y(_4399_)
);

FILL FILL_2__9157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11125_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4039_),
    .B(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_4041_)
);

NAND2X1 _8617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [1]),
    .B(_996__bF$buf3),
    .Y(_1507_)
);

FILL FILL_1__7574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13337_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12615_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Vld )
);

FILL FILL_1__8779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9300_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1637_),
    .Y(_1656_)
);

OAI21X1 _8370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1093_),
    .C(_1272_),
    .Y(_1273_)
);

FILL FILL_1__13090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7889_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2735_),
    .B(_2733_),
    .Y(_2736_)
);

FILL FILL_0__7469_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_2377_)
);

OAI21X1 _9155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1958_),
    .B(_1953_),
    .C(_1848__bF$buf4),
    .Y(_1978_)
);

FILL FILL_1__11823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14295_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6350_),
    .Y(_6353_)
);

NOR2X1 _13573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5945_),
    .Y(_5951_)
);

FILL FILL_0__13288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5611_),
    .Y(_5614_)
);

FILL FILL_2__13615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9615_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6989_),
    .B(_6995_),
    .Y(_6996_)
);

OR2X2 _14358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6652_),
    .B(_6651_),
    .Y(_6653_)
);

FILL FILL_2__8181_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_620_),
    .Y(_621_)
);

NAND3X1 _7221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .B(_215_),
    .C(_218_),
    .Y(_220_)
);

DFFPOSX1 _10698_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2524_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Ycalc [9])
);

OAI21X1 _10278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3006_),
    .B(_3005_),
    .C(_2741_),
    .Y(_3007_)
);

FILL FILL_1__12781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11354_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8846_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_844_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Ycalc [5])
);

AOI21X1 _8426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1322_),
    .B(_1324_),
    .C(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1327_)
);

AOI22X1 _8006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.Acalc [4]),
    .C(_927_),
    .D(\genblk1[1].u_ce.Acalc [6]),
    .Y(_928_)
);

FILL FILL_1__7383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12979_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5298_),
    .B(_5293_),
    .C(_5188__bF$buf5),
    .Y(_5318_)
);

FILL FILL_0__12139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4924_),
    .B(_4919_),
    .C(_4961_),
    .Y(_4963_)
);

OAI21X1 _12004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4561_),
    .C(_4565_),
    .Y(_4566_)
);

FILL FILL_0__13920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8168_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5986_),
    .B(_5961_),
    .C(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_6005_)
);

NOR2X1 _13209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5665_),
    .B(_5654_),
    .Y(_5667_)
);

FILL FILL_0__14705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7278_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .Y(_2197_)
);

FILL FILL_2_BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11212_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3561_),
    .C(_3564_),
    .Y(_3565_)
);

FILL FILL_0__10625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13097_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5816_),
    .B(_5800_),
    .C(_5817_),
    .Y(_5073_)
);

FILL FILL_2__13844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9004_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [18]),
    .Y(_6828_)
);

DFFPOSX1 _14167_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5843_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Ycalc [7])
);

FILL FILL_1__7859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8800_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_803_),
    .C(_820_),
    .Y(_51_)
);

NOR2X1 _7450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .B(_438_),
    .Y(_439_)
);

NOR2X1 _10087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2823_),
    .B(_2802_),
    .Y(_2824_)
);

FILL FILL_1__12170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11910_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1542_),
    .Y(_1543_)
);

NAND2X1 _8235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1140_),
    .Y(_1144_)
);

FILL FILL_1__7192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12788_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5134_),
    .C(_5135_),
    .Y(_5136_)
);

FILL FILL_0__12368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4781_),
    .B(_4784_),
    .Y(_4785_)
);

FILL FILL_1__8397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6086_),
    .C(_6223_),
    .Y(_6224_)
);

DFFPOSX1 _13438_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5038_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [9])
);

NAND2X1 _13018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .B(_5484_),
    .Y(_5485_)
);

FILL FILL257250x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .B(_1988_),
    .C(_1983_),
    .Y(_2015_)
);

FILL FILL_1__11861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10014_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [10]),
    .Y(_5649_)
);

DFFPOSX1 _7926_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[0].u_ce.Ycalc [9])
);

OAI21X1 _7506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .B(_491_),
    .C(_227_),
    .Y(_493_)
);

FILL FILL_2__13653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9653_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf1),
    .B(_4487_),
    .C(_4488_),
    .Y(_4489_)
);

FILL FILL_0__9233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11219_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4128_),
    .Y(_4129_)
);

OAI21X1 _14396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6551_),
    .B(\u_ot.LoadCtl_6_bF$buf1 ),
    .C(_6685_),
    .Y(_6507_)
);

FILL FILL_1__7668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14018_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5189_)
);

FILL FILL_2__10358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11392_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8884_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_882_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Xin12b [5])
);

NOR2X1 _8464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1341_),
    .B(_1360_),
    .Y(_1363_)
);

OAI21X1 _8044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_958_),
    .B(_961_),
    .C(_930_),
    .Y(_962_)
);

FILL FILL_2__7737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13184_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5324_),
    .B(_5328_),
    .C(_5323_),
    .Y(_5355_)
);

FILL FILL_0__12177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4992_),
    .B(_4993_),
    .C(_4994_),
    .Y(_4229_)
);

NAND2X1 _12042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .B(_4601_),
    .Y(_4602_)
);

FILL FILL_2__12924_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2450_),
    .B(_2463_),
    .C(_2461_),
    .Y(_2464_)
);

OAI21X1 _9249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2066_),
    .C(_2067_),
    .Y(_2068_)
);

FILL FILL_1__11917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6039_),
    .B(_6041_),
    .Y(_6042_)
);

NAND2X1 _13247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5701_),
    .Y(_5702_)
);

FILL FILL_0__14743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10243_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_708_),
    .Y(_28_)
);

NOR2X1 _7315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_288_),
    .Y(_310_)
);

FILL FILL_2__13882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11448_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4307_),
    .B(_4306_),
    .Y(\genblk1[5].u_ce.Y_ [1])
);

FILL FILL_0__9042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11028_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .B(_3950_),
    .C(_3507_),
    .Y(_3951_)
);

FILL FILL_1__7897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14247_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5404_),
    .B(_5406_),
    .C(_5407_),
    .Y(_5408_)
);

OAI21X1 _12518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Ain12b [9]),
    .Y(_5026_)
);

FILL FILL_1__14601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9203_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1577_),
    .B(_1537_),
    .Y(_1578_)
);

OAI21X1 _8273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1176_),
    .C(_1180_),
    .Y(_1181_)
);

FILL FILL_1__10941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10101_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925_),
    .Y(_5925__bF$buf2)
);

FILL FILL_2__7546_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925_),
    .Y(_5925__bF$buf1)
);

BUFX2 BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925_),
    .Y(_5925__bF$buf0)
);

BUFX2 BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf5)
);

BUFX2 BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf4)
);

BUFX2 BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf3)
);

BUFX2 BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf2)
);

BUFX2 BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf1)
);

BUFX2 BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963_),
    .Y(_5963__bF$buf0)
);

INVX2 _12691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5171_),
    .Y(_5172_)
);

BUFX2 BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 )
);

AND2X2 _12271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4811_),
    .B(_4820_),
    .Y(_4821_)
);

FILL FILL_2__12733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12313_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.Xcalc [5]),
    .C(_2603_),
    .D(\genblk1[3].u_ce.Xcalc [7]),
    .Y(_2643_)
);

AOI21X1 _9478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .B(_2284_),
    .C(_2279_),
    .Y(_2287_)
);

MUX2X1 _9058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1837_),
    .S(vdd),
    .Y(_1885_)
);

FILL FILL_1__11726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8313_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6259_),
    .B(_6237_),
    .Y(_6261_)
);

DFFPOSX1 _13476_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5076_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [7])
);

OR2X2 _13056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5520_),
    .B(_5519_),
    .Y(_5521_)
);

FILL FILL_2__13518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10052_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7964_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_48_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin0 [1])
);

OAI21X1 _7544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_525_),
    .C(_520_),
    .Y(_529_)
);

NOR2X1 _7124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Xcalc [11]),
    .Y(_127_)
);

FILL FILL_1__12684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9691_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4522_),
    .B(_4525_),
    .Y(_4526_)
);

FILL FILL_0__9271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3444_),
    .B(_3441_),
    .Y(_4159_)
);

NAND2X1 _11122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .B(_3747_),
    .Y(_3768_)
);

NAND2X1 _8749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1628_),
    .B(_1629_),
    .Y(_1630_)
);

NAND2X1 _8329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(_1233_),
    .Y(_1234_)
);

FILL FILL_1__7286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13049_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5224_),
    .B(_5177_),
    .S(vdd),
    .Y(_5225_)
);

OAI21X1 _12327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4870_),
    .B(_4872_),
    .C(_4859_),
    .Y(_4216_)
);

FILL FILL_1__14830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9012_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [1]),
    .B(_996__bF$buf0),
    .Y(_997_)
);

FILL FILL_1__10330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7355_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4423_),
    .C(_4637_),
    .Y(_4638_)
);

FILL FILL_2__12962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12122_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_2104_)
);

FILL FILL_1_CLKBUF1_insert390 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert391 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8542_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [4]),
    .Y(_3473_)
);

FILL FILL_0__8122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10108_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .B(_5738_),
    .Y(_5739_)
);

FILL FILL_2__9921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [6]),
    .B(_743_),
    .Y(_744_)
);

NOR2X1 _7353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_336_),
    .Y(_346_)
);

FILL FILL_1__12493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11486_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4342_),
    .Y(_4343_)
);

FILL FILL_0__9080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11066_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3979_),
    .Y(_3986_)
);

FILL FILL_1__9908_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [0]),
    .Y(_1808_)
);

OAI21X1 _8558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1452_),
    .C(_1440_),
    .Y(_1453_)
);

AOI21X1 _8138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1047_),
    .C(_1050_),
    .Y(_1051_)
);

FILL FILL_1__7095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13278_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_5444_)
);

DFFPOSX1 _12556_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4210_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xcalc [7])
);

NAND2X1 _12136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4690_),
    .B(_4691_),
    .Y(_4692_)
);

FILL FILL_0__13632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14417_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[9]),
    .Y(_6926_)
);

FILL FILL_2__7584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12351_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .Y(_1922_)
);

FILL FILL_1__11764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8351_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_3321_),
    .C(_3323_),
    .Y(_2556_)
);

FILL FILL_0__10337_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .B(_2917_),
    .C(_2923_),
    .Y(_2934_)
);

OAI21X1 _13094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf1),
    .B(_5555_),
    .C(_5556_),
    .Y(_5557_)
);

FILL FILL_2__9310_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [11]),
    .B(_158__bF$buf2),
    .Y(_795_)
);

AOI21X1 _7409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_377_),
    .C(_399_),
    .Y(_400_)
);

FILL FILL_2__13556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [2]),
    .B(_4348__bF$buf4),
    .Y(_4396_)
);

FILL FILL_0__9136_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(vdd),
    .Y(_4038_)
);

FILL FILL_1__13910_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [6]),
    .B(_6562__bF$buf1),
    .Y(_6602_)
);

FILL FILL_0__12903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(_564_),
    .Y(_565_)
);

MUX2X1 _7162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_161_),
    .S(_135__bF$buf3),
    .Y(_163_)
);

OAI21X1 _11580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_4180_)
);

FILL FILL_0__11295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf2),
    .B(_3803_),
    .Y(_3804_)
);

FILL FILL_1__9717_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1021_),
    .C(_1654_),
    .Y(_886_)
);

NAND2X1 _8367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1270_)
);

FILL FILL_1__10615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13087_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5259_),
    .Y(_5262_)
);

AND2X2 _12365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4907_),
    .B(_4906_),
    .Y(_4908_)
);

FILL FILL_0__13861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14226_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14511_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6499_),
    .CLK(clk_bF$buf4),
    .Q(\u_ot.Xcalc [11])
);

FILL FILL_2__7393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3503_),
    .B(_3505_),
    .C(_3508_),
    .Y(_3509_)
);

FILL FILL_0__8160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10146_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3116_),
    .B(_3151_),
    .C(_3149_),
    .Y(_3152_)
);

OAI21X1 _10011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2749_),
    .C(_2750_),
    .Y(_2751_)
);

OAI22X1 _7638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_618_),
    .D(_616_),
    .Y(_21_)
);

OAI21X1 _7218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_187_),
    .C(_172__bF$buf1),
    .Y(_217_)
);

FILL FILL_2__13365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9365_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11636_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3376_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [11])
);

OAI21X1 _11216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3851_),
    .B(_3854_),
    .C(_3856_),
    .Y(_3858_)
);

FILL FILL_0__12712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8321_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_369_),
    .C(_227_),
    .Y(_383_)
);

FILL FILL_0__13917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9106_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1487_),
    .B(_1476_),
    .Y(_1489_)
);

INVX1 _8176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .Y(_1088_)
);

FILL FILL_1__10844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7431_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12594_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4248_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin1 [1])
);

NOR2X1 _12174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4601_),
    .Y(_4728_)
);

FILL FILL_2__8810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8636_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .S(gnd),
    .Y(_3562_)
);

FILL FILL_0__8216_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6161_),
    .B(_6167_),
    .C(_6165_),
    .Y(_6168_)
);

OAI21X1 _13379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5427_),
    .B(_5796_),
    .C(_5815_),
    .Y(_5072_)
);

FILL FILL_0__14455_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6958_),
    .B(_6960_),
    .Y(_6961_)
);

FILL FILL_0__14035_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6610_),
    .C(_6613_),
    .Y(_6620_)
);

FILL FILL_1__11382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10795_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[2].u_ce.Y_ [1]),
    .Y(_3344_)
);

FILL FILL_0__10375_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2970_)
);

OAI21X1 _7867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_411_),
    .B(_799_),
    .C(_818_),
    .Y(_50_)
);

MUX2X1 _7447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_433_),
    .S(_135__bF$buf2),
    .Y(_436_)
);

FILL FILL_2__13594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9594_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf2),
    .B(_4429_),
    .C(_4432_),
    .Y(_4433_)
);

FILL FILL_0__9174_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [5]),
    .Y(_4073_)
);

NAND3X1 _11025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3637_),
    .B(_3653_),
    .C(_3636_),
    .Y(_3675_)
);

FILL FILL_0__12941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8025_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10716_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2542_),
    .CLK(clk_bF$buf4),
    .Q(\genblk1[3].u_ce.Acalc [3])
);

AND2X2 _13188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5637_),
    .B(_5646_),
    .Y(_5647_)
);

FILL FILL_0__14684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10511_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .Y(_654_)
);

AOI22X1 _7256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_158__bF$buf1),
    .C(_253_),
    .D(_230_),
    .Y(_4_)
);

FILL FILL_1__12396_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11674_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3414_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Ain12b [11])
);

FILL FILL_0__11389_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .Y(_3894_)
);

FILL FILL_0__12750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7716_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9822_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1734_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Yin1 [1])
);

NOR2X1 _9402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf1),
    .B(_2087_),
    .Y(_2214_)
);

NAND2X1 _12879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5348_),
    .B(_5351_),
    .Y(_5352_)
);

INVX1 _12459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [0]),
    .Y(_4992_)
);

INVX1 _12039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4587_),
    .Y(_4599_)
);

FILL FILL_1__14122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13955_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [10]),
    .B(_6182_),
    .C(_6187_),
    .Y(_6188_)
);

FILL FILL_0__13535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13115_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5827_)
);

FILL FILL_1__9984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10042_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6835_),
    .B(_6836_),
    .C(_6837_),
    .Y(_6767_)
);

FILL FILL_2__12674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8674_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3597_),
    .C(_3598_),
    .Y(_3599_)
);

FILL FILL_0__8254_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3236_),
    .B(_3238_),
    .Y(_3239_)
);

OAI21X1 _10105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2753_),
    .C(_2840_),
    .Y(_2841_)
);

FILL FILL_0__11601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10320_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [2]),
    .B(_158__bF$buf3),
    .Y(_472_)
);

FILL FILL_0__11198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4105_),
    .B(_4108_),
    .Y(_4109_)
);

INVX1 _11063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3711_),
    .Y(_3712_)
);

FILL FILL_2__11525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7525_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .Y(_2429_)
);

FILL FILL_0__7105_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_2029_),
    .C(_2025_),
    .Y(_2032_)
);

INVX1 _12688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5168_),
    .Y(_5169_)
);

NAND2X1 _12268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4815_),
    .B(_4816_),
    .Y(_4818_)
);

FILL FILL_1__14771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10271_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7036_),
    .Y(_7048_)
);

FILL FILL_0__14129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(\u_ot.Yin12b [10]),
    .C(_6700_),
    .Y(_6701_)
);

FILL FILL_2__7296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8063_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10754_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2580_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Ain12b [7])
);

FILL FILL_0__10469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .B(_3059_),
    .C(_2686__bF$buf5),
    .Y(_3060_)
);

FILL FILL_2__9862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11410_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8902_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_900_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Ain12b [11])
);

FILL FILL_0__9688_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf0),
    .B(_4519_),
    .C(_4513_),
    .Y(_4523_)
);

FILL FILL_0__9268_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [1]),
    .Y(_4157_)
);

NAND2X1 _11119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3762_),
    .B(_3764_),
    .Y(_3765_)
);

FILL FILL_1__13622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5369_),
    .C(_5365_),
    .Y(_5372_)
);

FILL FILL_1_BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14407_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_289_),
    .Y(_290_)
);

OAI21X1 _11292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .B(_3924_),
    .C(_3579_),
    .Y(_3931_)
);

FILL FILL_1__9849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1395_),
    .Y(_1396_)
);

OAI21X1 _8079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_989_),
    .B(_991_),
    .C(_994_),
    .Y(_995_)
);

FILL FILL_1__10327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7754_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [11]),
    .C(_2600_),
    .Y(_2609_)
);

FILL FILL_0__7334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2250_),
    .C(_2225_),
    .Y(_2251_)
);

INVX1 _9020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1849_)
);

OAI21X1 _12497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5011_),
    .B(_4997_),
    .C(_5014_),
    .Y(_4244_)
);

NAND2X1 _12077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [1]),
    .B(_4348__bF$buf0),
    .Y(_4635_)
);

FILL FILL_2__8713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14358_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6869_),
    .B(_6868_),
    .Y(_6872_)
);

NAND2X1 _14223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [2]),
    .Y(_6542_)
);

FILL FILL_1__7915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf3),
    .B(_3634_),
    .C(_3629_),
    .Y(_3635_)
);

FILL FILL_0__8292_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3274_),
    .Y(_3275_)
);

FILL FILL_0__10278_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2830_),
    .B(_2846_),
    .Y(_2877_)
);

FILL FILL_2__13077_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .Y(_1595_)
);

FILL FILL_0__9497_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4339_),
    .B(_4332_),
    .S(_4324__bF$buf0),
    .Y(_4340_)
);

FILL FILL_0__9077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982_),
    .B(_3973_),
    .C(_3508_),
    .Y(_3984_)
);

FILL FILL_1__13851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12004_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .Y(_2660_)
);

FILL FILL_1__8453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13629_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(_6277_),
    .C(_6275_),
    .Y(_6278_)
);

FILL FILL_0__13209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(_3321_),
    .Y(_3322_)
);

FILL FILL_1__12702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9307_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14872_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6763_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [3])
);

FILL FILL_0__14587_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [3]),
    .B(_6720_),
    .Y(_6733_)
);

AOI22X1 _14032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6372_),
    .B(_5949__bF$buf0),
    .C(_6390_),
    .D(_6387_),
    .Y(_5855_)
);

FILL FILL_1__7724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11094_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [10]),
    .Y(_3454_)
);

FILL FILL_0__10087_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3079_),
    .Y(_3096_)
);

FILL FILL_1__8929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10834_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _7999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .Y(_921_)
);

FILL FILL_2__9060_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .Y(_562_)
);

NOR2X1 _7159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_154_),
    .Y(_160_)
);

OAI21X1 _8940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1764_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1775_)
);

OAI21X1 _8520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1410_),
    .C(_1065_),
    .Y(_1417_)
);

NAND2X1 _8100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_1015_)
);

FILL FILL_1__12299_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4557_),
    .B(_4545_),
    .C(_4558_),
    .Y(_4559_)
);

OAI21X1 _11577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3628_),
    .B(_4162_),
    .C(_4178_),
    .Y(_3408_)
);

NAND2X1 _11157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3801_)
);

FILL FILL_1__13660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_2483_),
    .C(_2500_),
    .Y(_1730_)
);

NAND2X1 _9305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [1]),
    .B(_1834__bF$buf0),
    .Y(_2121_)
);

FILL FILL_1__8682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13858_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6086_),
    .B(_6091_),
    .C(_6094_),
    .Y(_6095_)
);

FILL FILL_0__13018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5750_),
    .B(_5754_),
    .Y(_5756_)
);

FILL FILL_1__9887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10365_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14508_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6496_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Xcalc [8])
);

FILL FILL_0__7792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8577_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf0),
    .B(_3487__bF$buf3),
    .Y(_3506_)
);

FILL FILL_0__8157_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3143_),
    .C(_3148_),
    .Y(_3149_)
);

NAND3X1 _10008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2709_),
    .C(_2727_),
    .Y(_2748_)
);

FILL FILL_1__12931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14396_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6906_)
);

NAND2X1 _14261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [1]),
    .B(_6562__bF$buf2),
    .Y(_6569_)
);

FILL FILL_1__7533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12709_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2882_),
    .B(_2891_),
    .C(_2913_),
    .Y(_2914_)
);

FILL FILL_1__8738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8318_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .B(_379_),
    .C(_378_),
    .Y(_380_)
);

FILL FILL256350x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4015_),
    .B(_4018_),
    .Y(_4019_)
);

FILL FILL_2__11848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7848_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .Y(_2697_)
);

FILL FILL_0__7428_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(_2338_),
    .C(\genblk1[2].u_ce.Ain0 [0]),
    .Y(_2339_)
);

INVX2 _9114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1938_),
    .Y(_1939_)
);

FILL FILL_1__8491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13667_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6294_),
    .B(_6313_),
    .C(_5963__bF$buf2),
    .Y(_6314_)
);

FILL FILL_0_BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13247_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [6]),
    .B(_5891_),
    .Y(_5913_)
);

NAND2X1 _13112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5573_),
    .Y(_5574_)
);

FILL FILL_0_BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x216150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10174_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6935_),
    .B(_6941_),
    .C(_6950_),
    .Y(_6958_)
);

OAI21X1 _14317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf1),
    .B(_6616_),
    .C(_6617_),
    .Y(_6496_)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11799_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .Y(_582_)
);

FILL FILL_1__11379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8386_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3335_),
    .B(_2597_),
    .C(_3342_),
    .Y(_2572_)
);

NAND2X1 _10237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_2967_)
);

FILL FILL_1__12740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11313_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Yin1 [0]),
    .Y(_6755_)
);

AOI21X1 _14070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6420_),
    .C(_6425_),
    .Y(_6426_)
);

OAI21X1 _8805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1114_),
    .B(_1648_),
    .C(_1664_),
    .Y(_894_)
);

FILL FILL_1__7762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12938_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5278_),
    .Y(_5279_)
);

FILL FILL_0__12518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10032_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .Y(_198_)
);

FILL FILL257250x126150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3837_),
    .C(_3834_),
    .Y(_3838_)
);

FILL FILL_0__12691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7657_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2359_),
    .C(_1755_),
    .Y(_1748_)
);

FILL FILL_0__7237_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(gnd),
    .C(_2157_),
    .Y(_2158_)
);

FILL FILL_1__14483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13896_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf1),
    .B(_6018_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_6132_)
);

FILL FILL_0__13056_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [11]),
    .B(_5174__bF$buf0),
    .Y(_5792_)
);

FILL FILL_1__9085_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14546_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6534_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Yin0 [0])
);

OAI21X1 _14126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6461_),
    .B(_5887_),
    .C(_6470_),
    .Y(_5869_)
);

FILL FILL_1__7818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11188_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3542_),
    .B(_3541_),
    .S(_3487__bF$buf3),
    .Y(_3543_)
);

FILL FILL_0__8195_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3177_),
    .Y(_3184_)
);

OAI21X1 _10046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2783_),
    .B(_2784_),
    .C(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2785_)
);

FILL FILL_0__11962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11122_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1504_),
    .Y(_1505_)
);

FILL FILL_1__7571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12747_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12612_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.LoadCtl [3])
);

FILL FILL_0__12327_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9819_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1731_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Yin12b [4])
);

FILL FILL_1__8776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14119_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6179_),
    .Y(_6185_)
);

FILL FILL_2__11886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7886_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2732_),
    .B(_2729_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2733_)
);

FILL FILL_0__7466_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_2374_)
);

OAI21X1 _9152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf4),
    .B(_1973_),
    .C(_1974_),
    .Y(_1975_)
);

FILL FILL_1__11820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14292_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6269_),
    .C(_6349_),
    .Y(_6350_)
);

OAI21X1 _13570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5923_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_5948_),
    .Y(_5835_)
);

FILL FILL_0__13285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5607_),
    .B(_5610_),
    .Y(_5611_)
);

FILL FILL_0__9612_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6988_),
    .B(_6992_),
    .C(_6984_),
    .Y(_6993_)
);

OAI21X1 _14355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6539_),
    .B(\u_ot.LoadCtl_6_bF$buf3 ),
    .C(_6650_),
    .Y(_6501_)
);

FILL FILL_1__7627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14817_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10695_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2521_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [6])
);

NOR2X1 _10275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3003_),
    .B(_3002_),
    .Y(_3004_)
);

FILL FILL_0__11771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11351_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8843_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_841_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Ycalc [2])
);

OAI21X1 _8423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1323_),
    .C(_1320_),
    .Y(_1324_)
);

OAI21X1 _8003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(\genblk1[1].u_ce.Acalc [8]),
    .C(_924_),
    .Y(_925_)
);

FILL FILL_1__7380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12976_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf4),
    .B(_5313_),
    .C(_5314_),
    .Y(_5315_)
);

OAI21X1 _12421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4934_),
    .B(_4950_),
    .C(_4948_),
    .Y(_4960_)
);

FILL FILL_0__12136_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4470_),
    .C(_4516_),
    .Y(_4563_)
);

OAI21X1 _9628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2426_),
    .C(_2409_),
    .Y(_1707_)
);

INVX1 _9208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .Y(_2029_)
);

FILL FILL_1__8585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5925__bF$buf0),
    .Y(_6002_)
);

OAI21X1 _13206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5663_),
    .B(_5662_),
    .C(_5272_),
    .Y(_5664_)
);

FILL FILL_0__14702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2152_),
    .C(_2193_),
    .Y(_2194_)
);

FILL FILL_2__8234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14299_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [0]),
    .B(_6824_),
    .C(_6825_),
    .Y(\a[0] [1])
);

DFFPOSX1 _14164_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5840_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[7].u_ce.Ycalc [4])
);

FILL FILL_1__7856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .B(_2819_),
    .C(_2820_),
    .Y(_2821_)
);

FILL FILL_2__10546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11160_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_1539_),
    .C(_1538_),
    .Y(_1540_)
);

NAND2X1 _8232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1140_),
    .Y(_1141_)
);

FILL FILL_1__10900_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3920_),
    .B(_3902_),
    .C(_3900_),
    .Y(_3928_)
);

FILL FILL_2__7505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12785_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5133_),
    .B(_5132_),
    .Y(\genblk1[6].u_ce.Y_ [1])
);

FILL FILL_0__12365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf1),
    .B(_4778_),
    .C(_4773_),
    .Y(_4782_)
);

AOI22X1 _9857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.Acalc [0]),
    .C(_2605_),
    .D(_2606_),
    .Y(_2607_)
);

NOR2X1 _9437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .B(_2247_),
    .Y(_2248_)
);

OAI22X1 _9017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(_1845_),
    .C(_1810__bF$buf1),
    .D(_1839_),
    .Y(_1846_)
);

FILL FILL_1__8394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x244950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .B(_6219_),
    .C(_6220_),
    .D(\genblk1[7].u_ce.Yin0 [1]),
    .Y(_6221_)
);

DFFPOSX1 _13435_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5035_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [6])
);

INVX1 _13015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5481_),
    .Y(_5482_)
);

FILL FILL_1__9599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7084_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_2011_),
    .Y(_2012_)
);

FILL FILL_0__10851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12289_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7923_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[0].u_ce.Ycalc [6])
);

NOR2X1 _7503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_488_),
    .Y(_490_)
);

FILL FILL_0__8289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9650_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4453_),
    .B(_4475_),
    .C(_4456_),
    .Y(_4486_)
);

FILL FILL_0__9230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11216_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4125_),
    .B(_4069_),
    .C(_4124_),
    .Y(_4126_)
);

NAND2X1 _14393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(\u_ot.Yin12b [6]),
    .Y(_6683_)
);

NAND2X1 _8708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf4),
    .B(_1509_),
    .Y(_1592_)
);

FILL FILL_1__7665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13008_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _12706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .B(_5185_),
    .C(_5150__bF$buf3),
    .D(_5179_),
    .Y(_5186_)
);

DFFPOSX1 _8881_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_879_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Xin12b [6])
);

NAND3X1 _8461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1320_),
    .B(_1281_),
    .C(_1298_),
    .Y(_1360_)
);

INVX1 _8041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [4]),
    .Y(_959_)
);

NAND2X1 _11098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3737_),
    .B(_3744_),
    .Y(_3745_)
);

FILL FILL_2__7734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12501_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_2442_),
    .C(_2456_),
    .Y(_2461_)
);

NAND3X1 _9246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2051_),
    .B(_2063_),
    .C(_2047_),
    .Y(_2065_)
);

FILL FILL_1__11914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13799_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6024_),
    .B(_6035_),
    .C(_6038_),
    .Y(_6039_)
);

FILL FILL_0__13379_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5698_),
    .B(vdd),
    .S(_5697_),
    .Y(_5699_)
);

FILL FILL_2__13706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9706_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14869_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6760_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [0])
);

INVX1 _14449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.X_ [1]),
    .Y(_6731_)
);

NOR2X1 _14029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6373_),
    .B(_6363_),
    .Y(_6388_)
);

FILL FILL_2__8272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_705_),
    .Y(_706_)
);

NAND3X1 _7312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .B(_305_),
    .C(_306_),
    .Y(_307_)
);

OAI21X1 _10789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .B(_3451_),
    .C(_3444_),
    .Y(_3452_)
);

FILL FILL_0__8098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .B(_3093_),
    .Y(_3094_)
);

FILL FILL_1__12872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11445_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(_4303_),
    .C(_4304_),
    .Y(_4305_)
);

FILL FILL_2__9057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11025_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3934_),
    .B(_3924_),
    .C(_3947_),
    .Y(_3948_)
);

AOI21X1 _8937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1770_),
    .C(_1771_),
    .Y(_1772_)
);

AOI21X1 _8517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1406_),
    .B(_1388_),
    .C(_1386_),
    .Y(_1414_)
);

FILL FILL_1__7894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13237_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5391_),
    .B(_5403_),
    .C(_5387_),
    .Y(_5405_)
);

OAI21X1 _12515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Ain12b [8]),
    .Y(_5024_)
);

FILL FILL256050x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9200_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .Y(_1575_)
);

OAI21X1 _8270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1174_),
    .B(_1177_),
    .C(_1065_),
    .Y(_1178_)
);

BUFX2 BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf5)
);

BUFX2 BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf4)
);

BUFX2 BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf3)
);

BUFX2 BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf2)
);

BUFX2 BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf1)
);

BUFX2 BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .Y(_3524__bF$buf0)
);

FILL FILL_2__12310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7789_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [3]),
    .Y(_2640_)
);

FILL FILL_0__7369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf0),
    .B(_2283_),
    .C(_2280_),
    .Y(_2284_)
);

NAND2X1 _9055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [2]),
    .B(_1834__bF$buf1),
    .Y(_1882_)
);

FILL FILL_1__11723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8310_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5974_),
    .B(_6255_),
    .C(_6252_),
    .Y(_6258_)
);

FILL FILL_0__13188_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13473_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5073_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin12b [8])
);

NAND2X1 _13053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5516_),
    .B(_5517_),
    .Y(_5518_)
);

FILL FILL_2__13935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9515_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [7]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf1),
    .Y(_6904_)
);

INVX1 _14258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin0 [1]),
    .Y(_6566_)
);

FILL FILL257250x230550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8081_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7961_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_45_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin1 [0])
);

OAI21X1 _7541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_525_),
    .C(_521_),
    .Y(_526_)
);

AOI22X1 _7121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.Xcalc [0]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Xcalc [2]),
    .Y(_125_)
);

AND2X2 _10598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3302_),
    .B(_3306_),
    .Y(_3307_)
);

NAND3X1 _10178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .B(_2905_),
    .C(_2910_),
    .Y(_2911_)
);

FILL FILL_1__12681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11254_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .Y(_1627_)
);

NAND2X1 _8326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1223_),
    .B(_1230_),
    .Y(_1231_)
);

FILL FILL_1__7283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12879_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [2]),
    .B(_5174__bF$buf1),
    .Y(_5222_)
);

FILL FILL_0__12459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4860_),
    .B(_4869_),
    .Y(_4870_)
);

FILL FILL_0__12039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8068_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6227_),
    .C(_6310_),
    .Y(_6311_)
);

OAI21X1 _13529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Xcalc [10]),
    .C(_5889_),
    .Y(_5910_)
);

INVX1 _13109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [6]),
    .Y(_5571_)
);

FILL FILL_0__14605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2101_)
);

FILL FILL_1__11952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10945_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [8]),
    .Y(_3470_)
);

FILL FILL_0__10525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10105_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5735_),
    .Y(_5736_)
);

FILL FILL_2__13744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9324_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6737_),
    .C(_6753_),
    .Y(_6530_)
);

OAI21X1 _14067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6423_),
    .B(_6422_),
    .C(_6410_),
    .Y(_5857_)
);

FILL FILL_1__7759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8700_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_740_),
    .Y(_741_)
);

OAI21X1 _7350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_343_),
    .Y(_8_)
);

FILL FILL_1__12490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11810_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1803_),
    .B(_1804_),
    .C(_1805_),
    .Y(_1806_)
);

NAND3X1 _8555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf3),
    .B(_1444_),
    .C(_1442_),
    .Y(_1450_)
);

MUX2X1 _8135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .S(vdd),
    .Y(_1048_)
);

FILL FILL_1__7092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12688_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5441_)
);

DFFPOSX1 _12553_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4207_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [4])
);

FILL FILL_0__12268_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf3),
    .B(_4688_),
    .Y(_4689_)
);

FILL FILL_1__8297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6128_),
    .B(_6112_),
    .Y(_6129_)
);

NAND2X1 _13338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5788_),
    .Y(_5789_)
);

FILL FILL_0__14834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14414_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf2),
    .B(_1915_),
    .C(_1918_),
    .Y(_1919_)
);

FILL FILL_1__11761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5427_),
    .Y(_5554_)
);

AND2X2 _7826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_792_),
    .Y(_793_)
);

NAND3X1 _7406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .B(_391_),
    .C(_396_),
    .Y(_397_)
);

FILL FILL_2__13973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11539_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.ISout ),
    .Y(_4394_)
);

FILL FILL_0__9133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11119_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4035_)
);

NAND2X1 _14296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(_6596_),
    .Y(_6599_)
);

FILL FILL_0__12900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14758_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12609_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .CLK(clk_bF$buf47),
    .Q(\genblk1[5].u_ce.LoadCtl [0])
);

FILL FILL_2__10678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9714_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.X_ [0]),
    .Y(_1653_)
);

NOR2X1 _8364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1002_),
    .Y(_1267_)
);

FILL FILL_1__10612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13084_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf2),
    .B(_5255_),
    .C(_5258_),
    .Y(_5259_)
);

FILL FILL_0__12497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12077_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4900_),
    .B(_4903_),
    .Y(_4905_)
);

FILL FILL_2__12824_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .Y(_2730_)
);

NOR2X1 _9569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [3]),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2371_)
);

NAND3X1 _9149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1961_),
    .C(_1942_),
    .Y(_1972_)
);

FILL FILL_1__11817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6312_),
    .B(_6333_),
    .C(_6316_),
    .Y(_6347_)
);

OAI21X1 _13567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5945_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_5946_)
);

NAND3X1 _13147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf2),
    .B(_5604_),
    .C(_5599_),
    .Y(_5608_)
);

FILL FILL_0__14643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10143_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .Y(_616_)
);

AOI21X1 _7215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_170_),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_214_)
);

FILL FILL_2__13782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11348_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11633_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3373_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [8])
);

OR2X2 _11213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3851_),
    .B(_3854_),
    .Y(_3855_)
);

FILL FILL_1__7797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5279_),
    .B(_5301_),
    .C(_5282_),
    .Y(_5312_)
);

INVX1 _12418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4956_),
    .Y(_4957_)
);

FILL FILL_0__13914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9103_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1484_),
    .C(_1094_),
    .Y(_1486_)
);

OAI21X1 _8173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1083_),
    .C(_1084_),
    .Y(_1085_)
);

FILL FILL_1__10841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7446_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12591_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4245_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Yin12b [4])
);

INVX1 _12171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [5]),
    .Y(_4725_)
);

FILL FILL_2__12633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12213_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9798_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1710_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Acalc [9])
);

NAND2X1 _9378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2191_)
);

FILL FILL_1__11206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8633_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3504_),
    .B(_3551_),
    .C(_3549_),
    .Y(_3559_)
);

FILL FILL_0__8213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf3),
    .B(_6164_),
    .C(_6163_),
    .Y(_6165_)
);

NAND2X1 _13376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5796_),
    .Y(_5814_)
);

FILL FILL_0__14452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_799_),
    .Y(_817_)
);

OAI21X1 _7444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_295_),
    .C(_432_),
    .Y(_433_)
);

FILL FILL_2__13591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11577_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4325__bF$buf2),
    .Y(_4430_)
);

FILL FILL_0__9171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11157_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4068_),
    .B(_4069_),
    .C(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Y(_4071_)
);

OAI21X1 _11022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(_3670_),
    .C(_3671_),
    .Y(_3672_)
);

NOR2X1 _8649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_973__bF$buf3),
    .Y(_1537_)
);

NAND3X1 _8229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf2),
    .B(_1137_),
    .C(_1134_),
    .Y(_1138_)
);

FILL FILL_1__7186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5129_),
    .C(_5130_),
    .Y(_5131_)
);

OAI21X1 _12227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4752_),
    .B(_4746_),
    .C(_4362__bF$buf1),
    .Y(_4779_)
);

FILL FILL_1__14730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12022_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf4),
    .B(_2005_),
    .C(_1999_),
    .Y(_2009_)
);

FILL FILL_1__11855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8022_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10713_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2539_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Acalc [0])
);

FILL FILL_0__10428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10008_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5641_),
    .B(_5642_),
    .Y(_5644_)
);

FILL FILL_2__13227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9647_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4303_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4483_),
    .Y(_4196_)
);

FILL FILL_0__9227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8603_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_651_),
    .Y(_652_)
);

NAND2X1 _7253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_250_),
    .Y(_251_)
);

FILL FILL_1__12393_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11671_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3411_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Yin0 [0])
);

FILL FILL_0__11386_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf1),
    .B(_3849_),
    .C(_3890_),
    .Y(_3891_)
);

DFFPOSX1 _8878_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_876_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[1].u_ce.Xin12b [11])
);

NAND2X1 _8458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1356_),
    .Y(_1357_)
);

INVX1 _8038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [8]),
    .Y(_956_)
);

FILL FILL_0__7713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf5),
    .B(_5345_),
    .C(_5339_),
    .Y(_5349_)
);

OAI21X1 _12456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4446_),
    .B(_4989_),
    .C(_4990_),
    .Y(_4227_)
);

OR2X2 _12036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4596_),
    .B(_4592_),
    .Y(_4597_)
);

FILL FILL_0__13952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14317_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [0]),
    .Y(_6835_)
);

FILL FILL_2__7484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8671_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf3),
    .B(_3595_),
    .C(_3586_),
    .Y(_3596_)
);

FILL FILL_2__8269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10657_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2942_),
    .B(_2755_),
    .C(_2686__bF$buf0),
    .Y(_3236_)
);

FILL FILL_0__10237_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2838_)
);

FILL FILL_2__9210_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_702_),
    .Y(_703_)
);

NAND3X1 _7309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_300_),
    .C(_303_),
    .Y(_304_)
);

FILL FILL_2__13036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9456_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4300_),
    .C(_4301_),
    .Y(_4302_)
);

FILL FILL_0__9036_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .B(_3941_),
    .Y(_3945_)
);

FILL FILL_1__13810_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14199_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5875_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Yin12b [9])
);

FILL FILL_0__12803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8412_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_468_),
    .B(_446_),
    .Y(_470_)
);

FILL FILL_0__11195_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf4),
    .B(_4023_),
    .Y(_4106_)
);

OAI21X1 _11060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3704_),
    .C(_3702_),
    .Y(_3709_)
);

FILL FILL_1__9617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11522_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .Y(_1572_)
);

INVX1 _8267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1174_),
    .Y(_1175_)
);

FILL FILL_1__10935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10515_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949_),
    .Y(_5949__bF$buf3)
);

FILL FILL_0__7522_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949_),
    .Y(_5949__bF$buf2)
);

FILL FILL_0__7102_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949_),
    .Y(_5949__bF$buf1)
);

BUFX2 BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949_),
    .Y(_5949__bF$buf0)
);

BUFX2 BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf5)
);

BUFX2 BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf4)
);

BUFX2 BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf3)
);

BUFX2 BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf2)
);

BUFX2 BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf1)
);

MUX2X1 _12685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5165_),
    .B(_5158_),
    .S(_5150__bF$buf0),
    .Y(_5166_)
);

BUFX2 BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .Y(_4362__bF$buf0)
);

NAND2X1 _12265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4813_),
    .B(_4814_),
    .Y(_4815_)
);

FILL FILL_0__13761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9370_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7044_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(_7045_),
    .Y(_6785_)
);

FILL FILL_0__14126_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6673_),
    .B(_6687_),
    .Y(_6698_)
);

FILL FILL_2__7293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10466_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10751_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2577_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Ain12b [8])
);

FILL FILL_0__10046_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf5),
    .B(_3056_),
    .C(_3051_),
    .Y(_3057_)
);

DFFPOSX1 _7958_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_42_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xin12b [7])
);

OAI21X1 _7538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_522_),
    .C(_172__bF$buf4),
    .Y(_523_)
);

NAND2X1 _7118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [6]),
    .B(_89_),
    .Y(_122_)
);

FILL FILL_2__13265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9685_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4489_),
    .B(_4486_),
    .C(_4362__bF$buf0),
    .Y(_4520_)
);

FILL FILL_0__9265_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4150_),
    .B(_3437_),
    .Y(_4155_)
);

NAND2X1 _11116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .B(_3676_),
    .Y(_3762_)
);

FILL FILL_1__8641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_283_),
    .C(_286_),
    .Y(_287_)
);

FILL FILL_0__13817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9006_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [6]),
    .Y(_1393_)
);

NAND2X1 _8076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf1),
    .B(_973__bF$buf3),
    .Y(_992_)
);

FILL FILL_1__10324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7331_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .B(_4997_),
    .Y(_5013_)
);

OAI21X1 _12074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf3),
    .B(_4632_),
    .C(_4621_),
    .Y(_4633_)
);

FILL FILL_2__8710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8536_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3464_),
    .B(_3467_),
    .C(_3444_),
    .Y(_3468_)
);

FILL FILL_0__8116_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf1),
    .B(_5982_),
    .Y(_6072_)
);

OR2X2 _13279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5732_),
    .B(_5728_),
    .Y(_5733_)
);

FILL FILL_0__14775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6869_)
);

NAND2X1 _14220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [1]),
    .Y(_6540_)
);

FILL FILL_1__7912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11282_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3589_),
    .B(_3487__bF$buf2),
    .C(_3631_),
    .Y(_3632_)
);

INVX1 _10560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3271_),
    .Y(_3272_)
);

FILL FILL_0__10275_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2861_),
    .B(_2874_),
    .C(_2674_),
    .Y(_2875_)
);

OAI21X1 _7767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .B(_717_),
    .C(_737_),
    .Y(_738_)
);

OAI21X1 _7347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf5),
    .B(_227_),
    .C(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Y(_341_)
);

FILL FILL_2__13074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9494_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(vdd),
    .Y(_4337_)
);

FILL FILL_0__9074_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3587_),
    .B(_3980_),
    .Y(_3981_)
);

FILL FILL_2__11807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7807_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2657_)
);

FILL FILL_1__8450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14633_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf2),
    .B(_6274_),
    .C(_6265_),
    .Y(_6275_)
);

FILL FILL_0__13626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8345_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Xin12b [9]),
    .Y(_3320_)
);

INVX1 _13088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [5]),
    .Y(_5551_)
);

FILL FILL_2__9724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10411_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [2]),
    .Y(_918_)
);

OAI21X1 _7576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_478_),
    .C(_558_),
    .Y(_559_)
);

OAI21X1 _7156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_157_),
    .Y(_0_)
);

FILL FILL_1__12296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4522_),
    .B(_4525_),
    .C(_4555_),
    .Y(_4556_)
);

NAND2X1 _11574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4162_),
    .Y(_4177_)
);

FILL FILL_0__11289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3498_),
    .B(_3795_),
    .Y(_3798_)
);

FILL FILL_0__12650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7616_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .B(_2483_),
    .Y(_2499_)
);

OAI21X1 _9302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf2),
    .B(_2118_),
    .C(_2107_),
    .Y(_2119_)
);

NOR2X1 _12779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5151__bF$buf3),
    .Y(_5256_)
);

OAI21X1 _12359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4619_),
    .C(_4901_),
    .Y(_4902_)
);

FILL FILL_1__14862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x194550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13855_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6090_),
    .Y(_6092_)
);

FILL FILL_0__13015_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5752_),
    .Y(_5753_)
);

FILL FILL_1__9884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10362_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14505_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6493_),
    .CLK(clk_bF$buf9),
    .Q(\u_ot.Xcalc [5])
);

FILL FILL_1__11987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8574_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3485_),
    .B(_3502_),
    .Y(_3503_)
);

FILL FILL_0__8154_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .B(_3145_),
    .C(_3133_),
    .Y(_2536_)
);

OAI21X1 _10005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2721_),
    .C(_2734_),
    .Y(_2745_)
);

FILL FILL_0__11921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14918_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_376_),
    .C(_374_),
    .Y(_377_)
);

FILL FILL_0__11098_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain0 [0]),
    .Y(_4016_)
);

FILL FILL_2__11425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7845_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2694_)
);

FILL FILL_0__7425_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2335_),
    .B(_2331_),
    .C(_1832_),
    .Y(_2337_)
);

OAI21X1 _9111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf4),
    .B(_1934_),
    .C(_1935_),
    .Y(_1936_)
);

DFFPOSX1 _12588_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4242_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin12b [9])
);

NAND2X1 _12168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4721_),
    .B(_4704_),
    .Y(_4723_)
);

FILL FILL_1__14671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14449_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [12]),
    .B(_6833__bF$buf3),
    .Y(_6955_)
);

FILL FILL_0__14029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6610_),
    .B(_6613_),
    .Y(_6615_)
);

FILL FILL_2__7196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8383_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_3341_)
);

FILL FILL_0__10369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2685_),
    .C(_2963_),
    .Y(_2964_)
);

FILL FILL_0__11730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11310_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1648_),
    .Y(_1663_)
);

FILL FILL_0__9588_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4425_),
    .C(_4426_),
    .Y(_4427_)
);

FILL FILL_0__9168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4067_),
    .B(_4066_),
    .Y(_4068_)
);

AND2X2 _11019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3620_),
    .B(_3623_),
    .Y(_3669_)
);

FILL FILL_1__13942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12935_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf2),
    .B(_5274_),
    .C(_5275_),
    .Y(_5276_)
);

FILL FILL_0__12515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x237750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14307_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_191_),
    .S(_134__bF$buf1),
    .Y(_195_)
);

INVX1 _11192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3834_),
    .Y(_3835_)
);

FILL FILL_1__9749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11234_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1300_),
    .B(_1289_),
    .S(gnd),
    .Y(_1301_)
);

FILL FILL_1__10647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10227_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf23)
);

FILL FILL_0__7654_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf22)
);

NAND2X1 _9760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[2] [0]),
    .Y(_1754_)
);

FILL FILL_0__7234_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf21)
);

NAND2X1 _9340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_2102_),
    .Y(_2155_)
);

CLKBUF1 CLKBUF1_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf18)
);

NOR2X1 _12397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4937_),
    .B(_4928_),
    .Y(_4938_)
);

FILL FILL_2__8613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14678_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14543_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6531_),
    .CLK(clk_bF$buf51),
    .Q(\u_ot.Yin12b [5])
);

FILL FILL_0__14258_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_6469_)
);

FILL FILL257250x180150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11185_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf2),
    .B(_3502_),
    .C(_3539_),
    .Y(_3540_)
);

FILL FILL_0__8192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10598_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [0]),
    .B(_2672__bF$buf1),
    .Y(_3182_)
);

FILL FILL_0__10178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2769_),
    .B(_2781_),
    .C(_2779_),
    .Y(_2782_)
);

FILL FILL257250x147750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain0 [0]),
    .Y(_1502_)
);

FILL FILL_0__9397_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11668_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3408_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Yin12b [5])
);

OAI21X1 _11248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3883_),
    .B(_3866_),
    .C(_3879_),
    .Y(_3888_)
);

FILL FILL_1__13751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12324_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9816_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1728_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Yin12b [9])
);

FILL FILL_1__8773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13949_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6177_),
    .Y(_6182_)
);

FILL FILL_0__13529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8668_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_3593_)
);

FILL FILL_0__8248_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3233_),
    .B(_3232_),
    .C(_3223_),
    .Y(_2543_)
);

FILL FILL_2__9627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14487_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6989_),
    .Y(_6990_)
);

FILL FILL_0__14067_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [1]),
    .Y(_6648_)
);

FILL FILL_1__7624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13807_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10692_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2518_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [3])
);

NAND3X1 _10272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(_3000_),
    .C(_2998_),
    .Y(_3001_)
);

FILL FILL_1__8829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_803_),
    .C(_836_),
    .Y(_64_)
);

NAND3X1 _7479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_464_),
    .C(_461_),
    .Y(_467_)
);

DFFPOSX1 _8840_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_838_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Ycalc [0])
);

INVX1 _8420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1320_),
    .Y(_1321_)
);

FILL FILL_1__12199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [10]),
    .Y(_922_)
);

OAI21X1 _11897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4444_),
    .B(_4462_),
    .C(_4463_),
    .Y(_4464_)
);

INVX1 _11477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [7]),
    .Y(_4103_)
);

OAI21X1 _11057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3704_),
    .C(_3705_),
    .Y(_3706_)
);

FILL FILL_1__13980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .B(_2414_),
    .Y(_2424_)
);

OAI21X1 _9205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1936_),
    .C(_2002_),
    .Y(_2026_)
);

FILL FILL_1__8582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13758_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .B(\genblk1[7].u_ce.Xin12b [8]),
    .S(vdd),
    .Y(_5999_)
);

FILL FILL_0__13338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [10]),
    .B(_5659_),
    .C(_5660_),
    .Y(_5661_)
);

FILL FILL_1__9367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7036_),
    .B(_7037_),
    .C(_7042_),
    .Y(_7043_)
);

OR2X2 _14408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .B(_6694_),
    .Y(_6696_)
);

FILL FILL_2_BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8057_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10748_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2574_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin0 [1])
);

NAND2X1 _10328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf1),
    .B(_2973_),
    .Y(_3054_)
);

FILL FILL_1__12831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [1]),
    .B(_6822_),
    .Y(_6823_)
);

DFFPOSX1 _14161_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5837_),
    .CLK(clk_bF$buf47),
    .Q(\genblk1[7].u_ce.ISout )
);

FILL FILL_1__7853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2809_),
    .B(_2814_),
    .C(_2817_),
    .Y(_2818_)
);

FILL FILL_1__8638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _7288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_262_),
    .C(_234_),
    .Y(_284_)
);

AND2X2 _11286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .B(_3918_),
    .Y(_3925_)
);

FILL FILL_2__11748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7748_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.Acalc [4]),
    .C(_2603_),
    .D(\genblk1[3].u_ce.Acalc [6]),
    .Y(_2604_)
);

FILL FILL_0__7328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2244_),
    .B(_2224_),
    .Y(_2245_)
);

NAND3X1 _9014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .B(_1840_),
    .C(_1811__bF$buf0),
    .Y(_1843_)
);

FILL FILL_1__8391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13987_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6217_),
    .Y(_6218_)
);

FILL FILL_0__13567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13147_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13432_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5032_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Ycalc [3])
);

MUX2X1 _13012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .B(_5467_),
    .S(vdd),
    .Y(_5479_)
);

FILL FILL_1__9596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x126150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10074_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6865_),
    .B(_6849_),
    .C(_6857_),
    .Y(_6866_)
);

NAND2X1 _14217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [0]),
    .B(selXY_bF$buf0),
    .Y(_6538_)
);

FILL FILL_0__7081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12286_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7920_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Ycalc [3])
);

FILL FILL_1__11699_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(_486_),
    .C(_484_),
    .Y(_487_)
);

FILL FILL_1__11279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3598_),
    .B(_3615_),
    .C(_3597_),
    .Y(_3629_)
);

FILL FILL_0__8286_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3185_),
    .B(_2686__bF$buf1),
    .Y(_3269_)
);

NAND3X1 _10137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .B(_2871_),
    .C(_2870_),
    .Y(_2872_)
);

FILL FILL_1__12640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6676_),
    .B(_6673_),
    .C(_6666_),
    .Y(_6680_)
);

INVX1 _8705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [7]),
    .Y(_1589_)
);

FILL FILL_1__7662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12838_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .B(_5180_),
    .C(_5151__bF$buf1),
    .Y(_5183_)
);

FILL FILL_0__12418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10772_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(\genblk1[0].u_ce.Ycalc [8]),
    .C(_86_),
    .Y(_103_)
);

NAND2X1 _13908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6270_),
    .B(_6271_),
    .Y(_6272_)
);

NAND2X1 _11095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf3),
    .B(_3741_),
    .Y(_3742_)
);

FILL FILL_2__11977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7557_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_2454_),
    .C(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2459_)
);

FILL FILL_0__7137_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1973_),
    .C(_2002_),
    .Y(_2062_)
);

FILL FILL_1__11911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13796_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6025_),
    .Y(_6036_)
);

FILL FILL_0__13376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5695_),
    .B(_5688_),
    .C(_5693_),
    .Y(_5696_)
);

FILL FILL_2__13703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [11]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .Y(_7069_)
);

NAND2X1 _14446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6728_),
    .B(_6720_),
    .Y(_6729_)
);

NAND3X1 _14026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5964_),
    .B(_6383_),
    .C(_6384_),
    .Y(_6385_)
);

FILL FILL_1__7718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11088_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [5]),
    .Y(_3449_)
);

FILL FILL_0__8095_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3028_),
    .B(_3089_),
    .C(_3090_),
    .Y(_3091_)
);

FILL FILL_0__11862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11022_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1756_),
    .B(_1759_),
    .C(_1769_),
    .Y(\a[3] [0])
);

AND2X2 _8514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1404_),
    .Y(_1411_)
);

FILL FILL_1__7891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12647_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5313_),
    .C(_5342_),
    .Y(_5402_)
);

FILL FILL_0__12227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [1]),
    .B(_4989_),
    .Y(_5022_)
);

INVX1 _9719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [1]),
    .Y(_2497_)
);

FILL FILL_1__8676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf0),
    .B(_6000_),
    .Y(_6089_)
);

FILL FILL_2__11786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7786_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2634_),
    .B(_2637_),
    .C(_2606_),
    .Y(_2638_)
);

FILL FILL_0__7366_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2194_),
    .Y(_2281_)
);

INVX1 _9052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.ISout ),
    .Y(_1880_)
);

FILL FILL_1__11720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11300_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_6234_),
    .C(_6254_),
    .Y(_6255_)
);

FILL FILL_0__13185_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13470_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5070_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin0 [1])
);

NOR2X1 _13050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf1),
    .B(_5514_),
    .Y(_5515_)
);

FILL FILL_2__13932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6899_),
    .B(_6900_),
    .Y(_6901_)
);

OAI21X1 _14255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6561_),
    .B(_6562__bF$buf4),
    .C(_6563_),
    .Y(_6488_)
);

FILL FILL_1__7527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14717_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3303_),
    .Y(_3304_)
);

INVX1 _10175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2902_),
    .Y(_2908_)
);

FILL FILL_2__10637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11251_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_1618_),
    .C(_1607_),
    .Y(_1624_)
);

NAND2X1 _8323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf3),
    .B(_1227_),
    .Y(_1228_)
);

FILL FILL_1__7280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12876_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.ISout ),
    .Y(_5220_)
);

FILL FILL_0__12456_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4866_),
    .B(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4867_)
);

FILL FILL_0__12036_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_2691_)
);

AOI21X1 _9528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2319_),
    .B(_1848__bF$buf5),
    .C(_2090_),
    .Y(_2334_)
);

NAND2X1 _9108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_1933_)
);

FILL FILL_1__8485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6307_),
    .Y(_6308_)
);

FILL FILL_0_BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[7].u_ce.Ycalc [1]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Ycalc [3]),
    .Y(_5908_)
);

FILL FILL_0_BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .B(_5567_),
    .Y(_5569_)
);

FILL FILL_0_BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7175_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2084_),
    .B(_2098_),
    .Y(_1688_)
);

FILL FILL_2__8974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11307_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [7]),
    .B(_6733_),
    .Y(_6752_)
);

NAND2X1 _14064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6418_),
    .B(_6420_),
    .Y(_6421_)
);

FILL FILL_1__7756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9902_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Xcalc [11]),
    .Y(_1803_)
);

OAI21X1 _8552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1424_),
    .B(_1421_),
    .C(_1010__bF$buf1),
    .Y(_1447_)
);

AOI21X1 _8132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_990_),
    .B(_1037_),
    .C(_1035_),
    .Y(_1045_)
);

FILL FILL_1__10800_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3787_),
    .B(_3592_),
    .Y(_3832_)
);

FILL FILL_2__7825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13272_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5424_),
    .B(_5438_),
    .Y(_5040_)
);

FILL FILL_0__12685_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12550_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4204_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [1])
);

FILL FILL_0__12265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [10]),
    .Y(_4686_)
);

OAI21X1 _9757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_1759_),
    .C(_1752_),
    .Y(_1745_)
);

OAI21X1 _9337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .C(_2151_),
    .Y(_2152_)
);

FILL FILL_1__8294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14057_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .B(_6124_),
    .C(_6125_),
    .Y(_6126_)
);

INVX1 _13335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5785_),
    .Y(_5786_)
);

FILL FILL_0__14831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1811__bF$buf3),
    .Y(_1916_)
);

FILL FILL_0__10331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12189_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_789_),
    .Y(_790_)
);

INVX1 _7403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .Y(_394_)
);

FILL FILL_2__13970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11536_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4390_),
    .B(_4342_),
    .Y(_4392_)
);

FILL FILL_2__9148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11116_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4022_),
    .B(_4031_),
    .Y(_4033_)
);

NAND2X1 _14293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6595_),
    .B(_6586_),
    .Y(_6596_)
);

OAI21X1 _8608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1499_),
    .B(_1498_),
    .C(_1491_),
    .Y(_862_)
);

FILL FILL_1__7565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13328_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12606_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4260_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Ain1 [1])
);

FILL FILL_2__10675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9711_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1640_),
    .B(_921_),
    .C(_1651_),
    .Y(_883_)
);

OAI21X1 _8361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1262_),
    .C(_1263_),
    .Y(_1264_)
);

FILL FILL_2__7634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12401_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2723_),
    .C(_2726_),
    .Y(_2727_)
);

NAND2X1 _9566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2367_),
    .B(_2360_),
    .Y(_2369_)
);

OAI21X1 _9146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1789_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_1969_),
    .Y(_1682_)
);

FILL FILL_1__11814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6343_),
    .B(_6344_),
    .C(_5947_),
    .Y(_6345_)
);

FILL FILL_0__13699_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5924_),
    .B(_5941_),
    .Y(_5943_)
);

FILL FILL_0__13279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5578_),
    .B(_5572_),
    .C(_5188__bF$buf3),
    .Y(_5605_)
);

FILL FILL_2__13606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9606_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6986_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(_6987_),
    .Y(_6781_)
);

OAI21X1 _14349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .B(_6537_),
    .C(_6645_),
    .Y(_6500_)
);

FILL FILL_0__10980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10140_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_609_),
    .Y(_613_)
);

NAND2X1 _7212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_134__bF$buf1),
    .Y(_211_)
);

DFFPOSX1 _10689_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2515_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Ycalc [1])
);

NAND3X1 _10269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf3),
    .B(_2997_),
    .C(_2988_),
    .Y(_2998_)
);

FILL FILL_1__12772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11345_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11630_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3370_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [5])
);

NAND2X1 _11210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3593_),
    .B(_3800_),
    .Y(_3852_)
);

OAI21X1 _8837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1502_),
    .C(_916_),
    .Y(_909_)
);

NAND2X1 _8417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(_1078_),
    .Y(_1318_)
);

FILL FILL_1__7794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x230550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5129_),
    .B(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .C(_5309_),
    .Y(_5034_)
);

NOR2X1 _12415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4344_),
    .Y(_4954_)
);

FILL FILL_0__13911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9100_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [10]),
    .B(_1481_),
    .C(_1482_),
    .Y(_1483_)
);

NAND3X1 _8170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf1),
    .B(_1081_),
    .C(_1072_),
    .Y(_1082_)
);

FILL FILL_2__7863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9795_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1707_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Acalc [6])
);

FILL FILL_0__7269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2188_),
    .B(_2187_),
    .Y(_2189_)
);

FILL FILL_1__11203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8648_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(\genblk1[3].u_ce.ISout ),
    .Y(_3557_)
);

FILL FILL_0__8210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6118_),
    .B(_6141_),
    .C(_6114_),
    .Y(_6162_)
);

FILL FILL_0__13088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5162_),
    .C(_5812_),
    .Y(_5069_)
);

FILL FILL_2__13835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [3]),
    .B(_6817_),
    .C(_6819_),
    .Y(_6820_)
);

OAI21X1 _14158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf5),
    .B(_6455_),
    .C(_6487_),
    .Y(_5884_)
);

OAI21X1 _7861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_146_),
    .C(_815_),
    .Y(_47_)
);

AOI22X1 _7441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .B(_428_),
    .C(_429_),
    .D(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_430_)
);

OAI21X1 _10498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf4),
    .B(_3213_),
    .C(_2686__bF$buf1),
    .Y(_3214_)
);

INVX1 _10078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .Y(_2815_)
);

FILL FILL_1__12161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1526_),
    .B(_1531_),
    .Y(_1534_)
);

AOI21X1 _8226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_973__bF$buf0),
    .C(_1117_),
    .Y(_1135_)
);

FILL FILL_1__7183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12779_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5126_),
    .C(_5127_),
    .Y(_5128_)
);

FILL FILL_0__12359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4688_),
    .C(_4775_),
    .Y(_4776_)
);

FILL FILL_0__13720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6215_)
);

DFFPOSX1 _13429_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5029_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Ycalc [1])
);

OAI21X1 _13009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf1),
    .B(_5475_),
    .C(_5468_),
    .Y(_5476_)
);

FILL FILL_2__7672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .B(_1972_),
    .C(_1848__bF$buf4),
    .Y(_2006_)
);

FILL FILL_1__11852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10425_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10710_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2536_),
    .CLK(clk_bF$buf34),
    .Q(\genblk1[3].u_ce.Xcalc [9])
);

FILL FILL_0__10005_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5639_),
    .B(_5640_),
    .Y(_5641_)
);

DFFPOSX1 _7917_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ycalc [1])
);

FILL FILL_2__13644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9644_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4465_),
    .B(_4480_),
    .Y(_4481_)
);

FILL FILL_0__9224_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6676_),
    .B(_6677_),
    .Y(_6678_)
);

FILL FILL_1__7659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8600_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_645_),
    .Y(_649_)
);

NAND3X1 _7250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_244_),
    .C(_247_),
    .Y(_248_)
);

FILL FILL_1__12390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11710_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8875_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_873_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[1].u_ce.Acalc [10])
);

OAI21X1 _8455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1223_),
    .C(_1353_),
    .Y(_1354_)
);

OAI21X1 _8035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(_953_),
    .C(_930_),
    .Y(_954_)
);

FILL FILL_0__7710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13175_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .B(_5312_),
    .C(_5188__bF$buf5),
    .Y(_5346_)
);

FILL FILL_0__12168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4276_),
    .B(_4282_),
    .Y(_4988_)
);

NAND3X1 _12033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4567_),
    .B(_4570_),
    .C(_4549_),
    .Y(_4594_)
);

FILL FILL_2__12915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11908_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5973_),
    .B(_6032_),
    .C(_6031_),
    .D(_5969_),
    .Y(_6033_)
);

NAND2X1 _13238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .B(_5693_),
    .Y(_5694_)
);

FILL FILL_0__14734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10234_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf2),
    .B(_699_),
    .C(_172__bF$buf5),
    .Y(_700_)
);

INVX1 _7306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .Y(_301_)
);

FILL FILL_2__13873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11439_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4299_),
    .B(_4298_),
    .Y(\genblk1[5].u_ce.Y_ [0])
);

FILL FILL_0__9033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3940_),
    .B(_3941_),
    .Y(_3942_)
);

DFFPOSX1 _14196_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5872_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Yin12b [10])
);

FILL FILL_0__12800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14658_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5399_),
    .B(_5398_),
    .C(_5246_),
    .Y(_5400_)
);

OAI21X1 _12509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4361_),
    .C(_5020_),
    .Y(_4250_)
);

FILL FILL_2__10998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9614_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1569_),
    .Y(_1570_)
);

NAND2X1 _8264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(_1168_),
    .Y(_1172_)
);

FILL FILL_1__10932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10512_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf3)
);

BUFX2 BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf2)
);

FILL FILL_2__7117_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf1)
);

BUFX2 BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf0)
);

BUFX2 BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .Y(_1834__bF$buf4)
);

BUFX2 BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .Y(_1834__bF$buf3)
);

BUFX2 BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .Y(_1834__bF$buf2)
);

BUFX2 BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .Y(_1834__bF$buf1)
);

BUFX2 BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .Y(_1834__bF$buf0)
);

NAND2X1 _12682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(gnd),
    .Y(_5163_)
);

FILL FILL_0__12397_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_134__bF$buf4)
);

OAI21X1 _12262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4729_),
    .C(_4775_),
    .Y(_4812_)
);

FILL FILL_2__12724_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [4]),
    .Y(_2635_)
);

AOI21X1 _9469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2277_),
    .B(_2253_),
    .C(_2276_),
    .Y(_2278_)
);

OR2X2 _9049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(_1828_),
    .Y(_1878_)
);

FILL FILL_1__11717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf2),
    .B(_6251_),
    .C(_6229_),
    .Y(_6252_)
);

DFFPOSX1 _13467_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5067_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin1 [0])
);

NAND2X1 _13047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [10]),
    .Y(_5512_)
);

FILL FILL_0__14123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10043_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7955_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_39_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin12b [8])
);

OAI21X1 _7535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_436_),
    .C(_519_),
    .Y(_520_)
);

OAI21X1 _7115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Xcalc [10]),
    .C(_86_),
    .Y(_119_)
);

FILL FILL_2__13682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9682_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4429_),
    .C(_4516_),
    .Y(_4517_)
);

FILL FILL_0__9262_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4151_),
    .Y(_4153_)
);

FILL FILL_0__11248_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3454_),
    .B(_3510__bF$buf1),
    .C(_3759_),
    .D(_3582_),
    .Y(_3363_)
);

FILL FILL_1__7697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5216_),
    .B(_5168_),
    .Y(_5218_)
);

OAI21X1 _12318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4619_),
    .B(_4852_),
    .C(_4362__bF$buf4),
    .Y(_4864_)
);

FILL FILL_1__14821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9003_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1374_),
    .B(_1389_),
    .Y(_1391_)
);

NOR2X1 _8073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_988_),
    .Y(_989_)
);

FILL FILL_1__10321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7346_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [1]),
    .Y(_5011_)
);

NAND2X1 _12071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf2),
    .B(_4625_),
    .Y(_4630_)
);

FILL FILL_2__12953_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .B(_2483_),
    .C(_2485_),
    .Y(_1718_)
);

AOI21X1 _9278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2081_),
    .B(_2079_),
    .C(_2085_),
    .Y(_2096_)
);

FILL FILL_1__11946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8533_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [5]),
    .Y(_3465_)
);

FILL FILL_0__8113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6069_)
);

OAI21X1 _13276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(_5170_),
    .Y(_5730_)
);

FILL FILL_2__9912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10272_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_734_),
    .Y(_735_)
);

NOR2X1 _7344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_337_),
    .B(_321_),
    .Y(_338_)
);

FILL FILL_1__12484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11477_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4334_)
);

FILL FILL_0__9071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11057_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3976_),
    .B(_3975_),
    .Y(_3978_)
);

AOI22X1 _8969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Xcalc [0]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Xcalc [2]),
    .Y(_1801_)
);

OAI21X1 _8549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1443_),
    .C(_1423_),
    .Y(_1444_)
);

NAND2X1 _8129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .B(\genblk1[0].u_ce.ISout ),
    .Y(_1043_)
);

FILL FILL_1__7086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2654_)
);

FILL FILL_1__13689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13269_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5421_),
    .B(_5419_),
    .C(_5425_),
    .Y(_5436_)
);

DFFPOSX1 _12547_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4201_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Ycalc [10])
);

OAI21X1 _12127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348__bF$buf0),
    .B(_4683_),
    .C(_4662_),
    .Y(_4205_)
);

FILL FILL_1__14630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12762_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1911_),
    .C(_1912_),
    .Y(_1913_)
);

FILL FILL_1__11755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8342_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3318_)
);

FILL FILL_0__10328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5547_),
    .B(_5530_),
    .Y(_5549_)
);

FILL FILL_2__13127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9547_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4361_),
    .B(_4378_),
    .C(_4386_),
    .Y(_4389_)
);

FILL FILL_0__9127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8503_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7993_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[0].u_ce.LoadCtl [4])
);

NAND3X1 _7573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_542_),
    .C(_525_),
    .Y(_556_)
);

OAI21X1 _7153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_154_),
    .C(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_155_)
);

FILL FILL_1__12293_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4506_),
    .B(_4522_),
    .Y(_4553_)
);

OAI21X1 _11571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4171_),
    .B(_4159_),
    .C(_4175_),
    .Y(_3405_)
);

FILL FILL_0__11286_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3498_),
    .B(_3795_),
    .C(_3508_),
    .Y(_3796_)
);

FILL FILL_1__9708_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1648_),
    .Y(_1650_)
);

NAND2X1 _8358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [0]),
    .B(_996__bF$buf4),
    .Y(_1261_)
);

FILL FILL_1__10606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5251_),
    .C(_5252_),
    .Y(_5253_)
);

NAND2X1 _12356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [4]),
    .B(_4348__bF$buf3),
    .Y(_4899_)
);

FILL FILL_0__13852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14217_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14502_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6490_),
    .CLK(clk_bF$buf46),
    .Q(\u_ot.Xcalc [2])
);

FILL FILL_2__7384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8589_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3498_),
    .C(_3499_),
    .Y(_3500_)
);

FILL FILL_0__8151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10137_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3141_),
    .B(_3143_),
    .Y(_3144_)
);

OAI21X1 _10002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2742_),
    .B(_2740_),
    .C(_2720_),
    .Y(_2517_)
);

FILL FILL_2__9950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9110_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .B(_609_),
    .Y(_610_)
);

MUX2X1 _7209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(\genblk1[0].u_ce.Xin12b [8]),
    .S(gnd),
    .Y(_208_)
);

FILL FILL257550x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9356_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11627_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3367_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xcalc [2])
);

OAI21X1 _11207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3722_),
    .C(_3848_),
    .Y(_3849_)
);

FILL FILL_1__13710_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [5]),
    .B(_5888_),
    .Y(_6453_)
);

FILL FILL_0__12703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14915_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_373_),
    .C(_372_),
    .Y(_374_)
);

FILL FILL_0__13908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11095_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4013_),
    .B(_4012_),
    .C(_4005_),
    .Y(_3376_)
);

FILL FILL_1__9937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11422_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1479_),
    .C(_1010__bF$buf3),
    .Y(_1480_)
);

NOR2X1 _8167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_1079_)
);

FILL FILL_1__10835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7422_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12585_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4239_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Yin12b [10])
);

NAND3X1 _12165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4329_),
    .B(_4719_),
    .C(_4718_),
    .Y(_4720_)
);

FILL FILL_2__8801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14446_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6947_),
    .B(_6951_),
    .C(_6833__bF$buf1),
    .Y(_6953_)
);

FILL FILL_0__14026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6595_),
    .B(_6611_),
    .Y(_6612_)
);

FILL FILL_2__7193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8380_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2769_),
    .B(_3324_),
    .C(_3339_),
    .Y(_2569_)
);

FILL FILL_0__10366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2961_)
);

OAI21X1 _7858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_814_)
);

NAND2X1 _7438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_426_),
    .Y(_427_)
);

FILL FILL_2__13165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9585_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4360_),
    .B(_4385_),
    .C(_4403_),
    .Y(_4424_)
);

FILL FILL_0__9165_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4024_),
    .C(_4064_),
    .Y(_4065_)
);

AOI22X1 _11016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .B(_3510__bF$buf1),
    .C(_3666_),
    .D(_3582_),
    .Y(_3359_)
);

FILL FILL_0__12932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14304_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .S(gnd),
    .Y(_192_)
);

FILL FILL_0__13717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf0),
    .B(_1297_),
    .C(_1290_),
    .Y(_1298_)
);

FILL FILL_1__10644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10224_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf53)
);

FILL FILL_0__7651_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf52)
);

FILL FILL_0__7231_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf48)
);

OR2X2 _12394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4933_),
    .B(\genblk1[5].u_ce.Ain12b [6]),
    .Y(_4935_)
);

FILL FILL_2__8610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8016_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10707_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2533_),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.Xcalc [6])
);

MUX2X1 _13599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5976_),
    .B(_5973_),
    .S(_5926__bF$buf1),
    .Y(_5977_)
);

OAI21X1 _13179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5555_),
    .C(_5601_),
    .Y(_5638_)
);

FILL FILL_0__14675_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14540_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6528_),
    .CLK(clk_bF$buf51),
    .Q(\u_ot.Yin12b [6])
);

FILL FILL_0__14255_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5930_),
    .B(_6466_),
    .C(_6467_),
    .Y(_5866_)
);

FILL FILL_1__7812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11182_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3535_),
    .C(_3536_),
    .Y(_3537_)
);

FILL FILL_0__10595_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_3176_),
    .Y(_3179_)
);

FILL FILL_0__10175_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2778_),
    .B(_2777_),
    .Y(_2779_)
);

FILL FILL_2__10922_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_640_),
    .Y(_646_)
);

INVX1 _7247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .Y(_245_)
);

FILL FILL_2__13394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9394_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11665_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3405_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Yin12b [6])
);

NAND2X1 _11245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(_3884_),
    .Y(_3886_)
);

FILL FILL_2__11707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7707_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9813_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1725_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Yin12b [10])
);

FILL FILL_1__8770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13946_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6162_),
    .B(_6166_),
    .C(_6178_),
    .Y(_6179_)
);

FILL FILL_0__13526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8665_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf2),
    .B(_3541_),
    .Y(_3590_)
);

FILL FILL_0__8245_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3210_),
    .B(_3218_),
    .C(_3217_),
    .Y(_3231_)
);

FILL FILL_2__9624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10311_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_803_),
    .C(_834_),
    .Y(_63_)
);

OAI21X1 _7476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_443_),
    .C(_463_),
    .Y(_464_)
);

FILL FILL_1__12196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4459_),
    .B(_4460_),
    .C(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4461_)
);

FILL FILL_0__11189_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4099_),
    .B(_4090_),
    .Y(_4101_)
);

NAND3X1 _11054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3702_),
    .C(_3701_),
    .Y(_3703_)
);

FILL FILL_2__11936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .B(\genblk1[2].u_ce.Ain12b [6]),
    .Y(_2421_)
);

AOI21X1 _9202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2022_),
    .B(_1996_),
    .C(_2021_),
    .Y(_2023_)
);

NAND2X1 _12679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5160_)
);

NAND2X1 _12259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [9]),
    .B(_4348__bF$buf2),
    .Y(_4809_)
);

FILL FILL256650x86550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13335_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Vld ),
    .B(_5995_),
    .C(_5996_),
    .Y(_5837_)
);

OAI21X1 _13200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5638_),
    .B(_5657_),
    .C(_5188__bF$buf2),
    .Y(_5658_)
);

FILL FILL_1__9364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10262_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7032_),
    .Y(_7040_)
);

OAI21X1 _14405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf3),
    .B(_6692_),
    .C(_6693_),
    .Y(_6508_)
);

FILL FILL_1__11887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8054_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10745_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2571_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Yin1 [0])
);

NAND2X1 _10325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3035_),
    .B(_3039_),
    .Y(_3051_)
);

FILL FILL_0__11821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert211 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert212 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert214 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert216 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert217 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert219 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14818_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf3),
    .B(_191_),
    .Y(_281_)
);

OAI21X1 _11283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3883_),
    .B(_3866_),
    .C(_3921_),
    .Y(_3922_)
);

FILL FILL_2__11745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7745_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(\genblk1[3].u_ce.Acalc [8]),
    .C(_2600_),
    .Y(_2601_)
);

FILL FILL_0__7325_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1812_),
    .B(_2236_),
    .C(_2239_),
    .Y(_2242_)
);

INVX2 _9011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_1840_)
);

INVX1 _12488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [0]),
    .Y(_5009_)
);

NAND2X1 _12068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4626_),
    .Y(_4627_)
);

FILL FILL_1__14571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14349_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6863_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(_6856_),
    .Y(_6770_)
);

DFFPOSX1 _14214_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.LoadCtl [5])
);

FILL FILL_2__7096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11276_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3457_),
    .B(_3510__bF$buf1),
    .C(_3626_),
    .D(_3582_),
    .Y(_3357_)
);

FILL FILL_0__8283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3258_),
    .B(_3263_),
    .Y(_3266_)
);

FILL FILL_0__10269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2862_),
    .B(_2868_),
    .C(_2865_),
    .Y(_2869_)
);

FILL FILL_2__9662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11210_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_1576_),
    .Y(_1587_)
);

FILL FILL_0__9488_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4329_),
    .C(_4330_),
    .Y(_4331_)
);

FILL FILL_0__9068_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .Y(_3975_)
);

FILL FILL_1__13842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x180150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12835_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_5180_)
);

FILL FILL_0__12415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2651_)
);

FILL FILL_1__8444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14627_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Acalc [1]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Acalc [3]),
    .Y(_101_)
);

FILL FILL257550x147750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_6267_),
    .C(_6268_),
    .Y(_6269_)
);

INVX1 _11092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3738_),
    .Y(_3739_)
);

FILL FILL_1__9649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11134_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1204_),
    .C(_1202_),
    .Y(_1205_)
);

FILL FILL_1__10967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7554_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [9]),
    .B(_1848__bF$buf1),
    .Y(_2456_)
);

FILL FILL_0__7134_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2059_),
    .B(_2058_),
    .C(_1906_),
    .Y(_2060_)
);

AOI21X1 _12297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4828_),
    .B(_4838_),
    .C(_4844_),
    .Y(_4845_)
);

FILL FILL_2__8933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14578_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6803_),
    .B(_6833__bF$buf2),
    .C(_7067_),
    .Y(_6795_)
);

FILL FILL_0__14158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6633_),
    .B(_6724_),
    .C(_6726_),
    .Y(_6513_)
);

NAND3X1 _14023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(_6378_),
    .C(_6381_),
    .Y(_6382_)
);

FILL FILL_1__7715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11085_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [9]),
    .Y(_3446_)
);

FILL FILL_0__8092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10078_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3041_),
    .B(_3044_),
    .Y(_3088_)
);

OAI21X1 _8931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1760_),
    .B(_1763_),
    .C(_1766_),
    .Y(_1767_)
);

OAI21X1 _8511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1352_),
    .C(_1407_),
    .Y(_1408_)
);

AOI21X1 _11988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4537_),
    .B(_4550_),
    .C(_4350_),
    .Y(_4551_)
);

FILL FILL_0__9297_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_4174_)
);

NAND2X1 _11148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3785_),
    .Y(_3793_)
);

FILL FILL_1__13651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12224_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [0]),
    .Y(_2495_)
);

FILL FILL_1__8673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13849_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .Y(_6086_)
);

FILL FILL_0__13009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10356_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[9]),
    .Y(Dout[9])
);

FILL FILL_0__7783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8568_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3495_),
    .C(_3496_),
    .Y(_3497_)
);

FILL FILL_0__8148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(_3139_),
    .C(_3140_),
    .Y(_3141_)
);

FILL FILL_1__12922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6894_),
    .B(_6888_),
    .C(_6889_),
    .Y(_6898_)
);

INVX1 _14252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin0 [0]),
    .Y(_6561_)
);

FILL FILL_1__7524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x223350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13707_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3300_),
    .Y(_3301_)
);

NAND2X1 _10172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2900_),
    .Y(_2905_)
);

FILL FILL_1__8729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8309_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_701_),
    .C(\genblk1[0].u_ce.Ain12b [8]),
    .Y(_768_)
);

NOR3X1 _7379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_350_),
    .C(_323_),
    .Y(_371_)
);

OAI22X1 _8740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_1621_),
    .D(_1620_),
    .Y(_872_)
);

INVX1 _8320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1224_),
    .Y(_1225_)
);

FILL FILL_1__12099_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4366_),
    .C(_4367_),
    .Y(_4368_)
);

NOR2X1 _11377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4010_),
    .B(_4009_),
    .Y(_4011_)
);

FILL FILL_1__13880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_2688_)
);

AOI21X1 _9525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2324_),
    .C(_2330_),
    .Y(_2331_)
);

AOI21X1 _9105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(_1924_),
    .C(_1925_),
    .Y(_1930_)
);

FILL FILL_1__8482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6285_),
    .B(_6300_),
    .C(_6298_),
    .Y(_6305_)
);

FILL FILL_0__13658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [7]),
    .B(_5891_),
    .Y(_5905_)
);

FILL FILL_0_BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5192_),
    .B(_5563_),
    .C(_5559_),
    .Y(_5566_)
);

FILL FILL_0_BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10165_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6949_),
    .B(_6948_),
    .Y(_6950_)
);

OAI21X1 _14308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6603_),
    .B(\u_ot.LoadCtl_6_bF$buf4 ),
    .C(_6609_),
    .Y(_6495_)
);

FILL FILL_0__7592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x133350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(_3321_),
    .Y(_3338_)
);

OAI21X1 _10228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2958_),
    .B(_2953_),
    .C(_2937_),
    .Y(_2527_)
);

FILL FILL_1__12731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11304_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6749_),
    .B(_6729_),
    .C(_6750_),
    .Y(_6527_)
);

NAND3X1 _14061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .B(_6416_),
    .C(_6417_),
    .Y(_6418_)
);

FILL FILL_1__7753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8118_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .S(gnd),
    .Y(_189_)
);

NAND2X1 _11186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf0),
    .B(_3785_),
    .Y(_3829_)
);

FILL FILL_2__7822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7648_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [1]),
    .B(_2486_),
    .Y(_1751_)
);

FILL FILL_0__7228_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2143_),
    .C(_2141_),
    .Y(_2149_)
);

FILL FILL_1__8291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13887_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6113_),
    .B(_6119_),
    .C(_6122_),
    .Y(_6123_)
);

FILL FILL_0__13047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _13332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5110_),
    .B(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .C(_5783_),
    .D(_5782_),
    .Y(_5057_)
);

FILL FILL_1__9496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10394_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14537_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6525_),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.Yin12b [11])
);

OAI21X1 _14117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6461_),
    .B(_6463_),
    .C(_6465_),
    .Y(_5865_)
);

FILL FILL_1__7809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12186_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .Y(_787_)
);

FILL FILL_1__11599_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_386_),
    .Y(_391_)
);

FILL FILL_1__11179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3532_),
    .C(_3533_),
    .Y(_3534_)
);

FILL FILL_0__8186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2649__bF$buf4),
    .C(_2668_),
    .Y(_3176_)
);

OAI21X1 _10037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf0),
    .B(_2774_),
    .C(_2775_),
    .Y(_2776_)
);

FILL FILL_1__12960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11113_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf4),
    .B(_6593_),
    .Y(_6594_)
);

NOR2X1 _8605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1495_),
    .Y(_1497_)
);

FILL FILL_1__7562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12738_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12603_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4257_),
    .CLK(clk_bF$buf47),
    .Q(\genblk1[5].u_ce.Ain12b [4])
);

FILL FILL_0__12318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8347_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [10]),
    .Y(_6176_)
);

FILL FILL_2__11877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7877_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .S(vdd),
    .Y(_2724_)
);

FILL FILL_0__7457_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2365_),
    .Y(_2366_)
);

AND2X2 _9143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1951_),
    .B(_1966_),
    .Y(_1967_)
);

FILL FILL_1__11811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6341_),
    .B(_6340_),
    .Y(_6342_)
);

FILL FILL_0__13696_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5939_),
    .B(_5936_),
    .S(_5926__bF$buf4),
    .Y(_5940_)
);

FILL FILL_0__13276_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5514_),
    .C(_5601_),
    .Y(_5602_)
);

FILL FILL_2__13603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9603_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6981_),
    .B(_6982_),
    .C(_6980_),
    .Y(_6985_)
);

NAND3X1 _14346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6643_),
    .C(_6640_),
    .Y(_6644_)
);

FILL FILL_1__7618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[3] [1]),
    .Y(_2593_)
);

NAND2X1 _10266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2993_),
    .B(_2994_),
    .Y(_2995_)
);

FILL FILL_0__11762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11342_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_915_)
);

NAND2X1 _8414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf2),
    .B(_1271_),
    .Y(_1315_)
);

FILL FILL_1__7791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12967_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5291_),
    .B(_5306_),
    .Y(_5307_)
);

FILL FILL_0__12127_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4942_),
    .B(_4950_),
    .C(_4348__bF$buf3),
    .Y(_4952_)
);

OAI21X1 _9619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2375_),
    .C(_1848__bF$buf3),
    .Y(_2418_)
);

FILL FILL_1__8996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949__bF$buf1),
    .B(_5994_),
    .C(_5950_),
    .Y(_5836_)
);

FILL FILL_2_BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9792_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1704_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Acalc [3])
);

FILL FILL_0__7266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2184_),
    .Y(_2186_)
);

FILL FILL_1__11200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14092_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6149_),
    .Y(_6159_)
);

FILL FILL_0__13085_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5811_)
);

FILL FILL_2__13832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9412_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6804_),
    .B(_6816_),
    .C(_6805_),
    .Y(_6817_)
);

NAND2X1 _14155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6486_)
);

FILL FILL_1__7847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert180 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert181 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert183 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert185 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert186 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert188 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3210_),
    .Y(_3211_)
);

NAND2X1 _10075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf2),
    .B(_2723_),
    .Y(_2812_)
);

FILL FILL_0__11991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11151_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .B(_1531_),
    .Y(_1532_)
);

INVX1 _8223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [6]),
    .Y(_1132_)
);

FILL FILL_1__7180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12776_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5125_),
    .B(_5124_),
    .Y(\genblk1[6].u_ce.Y_ [0])
);

FILL FILL_0__12356_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .B(_4751_),
    .Y(_4773_)
);

NOR2X1 _9848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [10]),
    .Y(_2598_)
);

OAI21X1 _9428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2237_),
    .C(_2238_),
    .Y(_2239_)
);

MUX2X1 _9008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(\genblk1[2].u_ce.Xin12b [6]),
    .S(gnd),
    .Y(_1837_)
);

FILL FILL_1__8385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14148_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6210_),
    .B(_6212_),
    .C(_6021_),
    .Y(_6213_)
);

NAND2X1 _13426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[6] [1]),
    .Y(_5101_)
);

OAI21X1 _13006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5292_),
    .C(_5472_),
    .Y(_5473_)
);

FILL FILL_1__10488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7075_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1915_),
    .C(_2002_),
    .Y(_2003_)
);

FILL FILL_0__10842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10002_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[0] [1]),
    .Y(_79_)
);

FILL FILL_1__12634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9641_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4476_),
    .B(_4473_),
    .C(_4466_),
    .Y(_4478_)
);

FILL FILL_0__9221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(\u_ot.Yin12b [6]),
    .C(_6674_),
    .Y(_6675_)
);

FILL FILL_1__7656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11380_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8872_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_870_),
    .CLK(clk_bF$buf46),
    .Q(\genblk1[1].u_ce.Acalc [7])
);

AOI22X1 _8452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(_996__bF$buf4),
    .C(_1351_),
    .D(_994_),
    .Y(_854_)
);

INVX1 _8032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [5]),
    .Y(_951_)
);

OAI21X1 _11089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3462_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3736_),
    .Y(_3362_)
);

FILL FILL_2__7725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13172_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5255_),
    .C(_5342_),
    .Y(_5343_)
);

FILL FILL_0__12165_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4982_),
    .B(_4978_),
    .C(_4981_),
    .Y(_4986_)
);

NAND3X1 _12030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4549_),
    .B(_4571_),
    .C(_4557_),
    .Y(_4591_)
);

FILL FILL_2__12912_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2453_),
    .C(_2439_),
    .Y(_1709_)
);

AND2X2 _9237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2056_),
    .Y(_2057_)
);

FILL FILL_1__8194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14377_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf2),
    .B(_6028_),
    .C(_6029_),
    .Y(_6030_)
);

NAND2X1 _13235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5690_),
    .B(_5689_),
    .Y(_5691_)
);

FILL FILL_0__14731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12089_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .Y(_697_)
);

NAND2X1 _7303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf3),
    .B(_209_),
    .Y(_298_)
);

FILL FILL_2__13870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11436_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(_4295_),
    .C(_4296_),
    .Y(_4297_)
);

FILL FILL_0__9030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11016_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3938_),
    .C(_3935_),
    .Y(_3939_)
);

DFFPOSX1 _14193_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5869_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Xin1 [1])
);

INVX2 _8928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_1764_)
);

NAND2X1 _8508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1404_),
    .B(_1403_),
    .Y(_1405_)
);

FILL FILL_1__7885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13228_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5393_),
    .B(_5396_),
    .Y(_5397_)
);

NAND2X1 _12506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.Y_ [0]),
    .Y(_5019_)
);

FILL FILL_2__10575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9611_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .Y(_1567_)
);

NAND2X1 _8261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(_1168_),
    .Y(_1169_)
);

BUFX2 BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .Y(_5926__bF$buf2)
);

FILL FILL_2__7534_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .Y(_5926__bF$buf1)
);

BUFX2 BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .Y(_5926__bF$buf0)
);

BUFX2 BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf4 )
);

BUFX2 BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf3 )
);

BUFX2 BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf2 )
);

BUFX2 BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf1 )
);

BUFX2 BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf0 )
);

BUFX2 BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .Y(_3510__bF$buf4)
);

BUFX2 BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .Y(_3510__bF$buf3)
);

FILL FILL_0__12394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12301_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [8]),
    .Y(_2632_)
);

AOI22X1 _9466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_1834__bF$buf4),
    .C(_2275_),
    .D(_2272_),
    .Y(_1696_)
);

NAND3X1 _9046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1847_),
    .B(_1864_),
    .C(_1872_),
    .Y(_1875_)
);

FILL FILL_1__11714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8301_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf1),
    .B(_6248_),
    .Y(_6249_)
);

FILL FILL_0__13599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13179_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13464_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5064_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin12b [7])
);

OAI21X1 _13044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174__bF$buf3),
    .B(_5509_),
    .C(_5488_),
    .Y(_5043_)
);

FILL FILL_2__13506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6895_),
    .B(_6892_),
    .Y(_6896_)
);

INVX1 _14249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [11]),
    .Y(_6559_)
);

FILL FILL_0__10880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10040_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7952_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[0].u_ce.Acalc [11])
);

NAND2X1 _7532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_516_),
    .Y(_517_)
);

AOI22X1 _7112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Ycalc [1]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_117_)
);

NAND2X1 _10589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [10]),
    .B(_2672__bF$buf3),
    .Y(_3298_)
);

AOI21X1 _10169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2885_),
    .B(_2889_),
    .C(_2901_),
    .Y(_2902_)
);

FILL FILL_1__12672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12252_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4514_)
);

NOR2X1 _11530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4149_),
    .B(_4150_),
    .Y(_4151_)
);

FILL FILL_0__11245_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3756_),
    .B(_3699_),
    .C(_3752_),
    .Y(_3757_)
);

NAND2X1 _8737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1617_),
    .Y(_1619_)
);

OAI21X1 _8317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_948_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1222_),
    .Y(_848_)
);

FILL FILL_1__7694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13037_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5187_),
    .B(_5204_),
    .C(_5212_),
    .Y(_5215_)
);

NOR2X1 _12315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .Y(_4861_)
);

FILL FILL_0__13811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9000_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1385_),
    .C(_1381_),
    .Y(_1388_)
);

OAI21X1 _8070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_984_),
    .C(_985_),
    .Y(_986_)
);

FILL FILL_2__7763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7589_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(_2483_),
    .Y(_2484_)
);

FILL FILL_0__7169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2092_),
    .Y(_2093_)
);

FILL FILL_1__11943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8548_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [9]),
    .Y(_3462_)
);

FILL FILL_0__8110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6063_),
    .B(_6045_),
    .C(_6062_),
    .Y(_6066_)
);

OAI21X1 _13273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5725_),
    .B(_5726_),
    .C(_5723_),
    .Y(_5727_)
);

FILL FILL_2__13315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9315_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14898_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6789_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.Atmp [2])
);

OAI21X1 _14478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6729_),
    .C(_6748_),
    .Y(_6526_)
);

OAI21X1 _14058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6395_),
    .C(_5963__bF$buf0),
    .Y(_6415_)
);

OAI22X1 _7761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_730_),
    .D(_732_),
    .Y(_30_)
);

NAND3X1 _7341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(_333_),
    .C(_334_),
    .Y(_335_)
);

FILL FILL256050x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3120_),
    .Y(_3121_)
);

FILL FILL_1__12481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [6]),
    .B(_1765_),
    .Y(_1798_)
);

INVX1 _8546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1441_)
);

AOI21X1 _8126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_1039_),
    .C(_998_),
    .Y(_1041_)
);

FILL FILL_1__7083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5431_),
    .B(_5432_),
    .Y(_5433_)
);

FILL FILL_0__12679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12259_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12544_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4198_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[5].u_ce.Ycalc [7])
);

AND2X2 _12124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4680_),
    .B(_4663_),
    .Y(_4681_)
);

FILL FILL_0__13620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6118_),
    .Y(_6120_)
);

NAND2X1 _13329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5780_),
    .B(_5779_),
    .Y(_5781_)
);

FILL FILL_0__14825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1846_),
    .B(_1871_),
    .C(_1889_),
    .Y(_1910_)
);

FILL FILL_1__11752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8777_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2838_),
    .B(_3313_),
    .C(_3315_),
    .Y(_2552_)
);

FILL FILL_0__10325_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5155_),
    .B(_5545_),
    .C(_5544_),
    .Y(_5546_)
);

NAND2X1 _7817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [10]),
    .B(_158__bF$buf2),
    .Y(_784_)
);

FILL FILL_2__13544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9544_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4360_),
    .C(_4385_),
    .Y(_4386_)
);

FILL FILL_0__9124_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [4]),
    .B(_6583_),
    .C(\u_ot.ISreg_bF$buf0 ),
    .Y(_6591_)
);

FILL FILL_1__7559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8500_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7990_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.LoadCtl [1])
);

OAI21X1 _7570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_553_),
    .C(_156_),
    .Y(_554_)
);

NAND2X1 _7150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_150_),
    .Y(_152_)
);

FILL FILL_1__12290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9705_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_1648_)
);

OAI21X1 _8355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1255_),
    .B(_1258_),
    .C(_1065_),
    .Y(_1259_)
);

FILL FILL_1__10603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13075_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5186_),
    .B(_5211_),
    .C(_5229_),
    .Y(_5250_)
);

FILL FILL_0__12488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12068_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4896_),
    .B(_4887_),
    .C(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4897_)
);

FILL FILL_1__8097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8815_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6334_),
    .B(_6338_),
    .C(_5967_),
    .Y(_6339_)
);

INVX1 _13558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .Y(_5937_)
);

NAND2X1 _13138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5575_),
    .B(_5577_),
    .Y(_5599_)
);

FILL FILL_0__14634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10134_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .Y(_607_)
);

OAI21X1 _7206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_204_),
    .C(_205_),
    .Y(_2_)
);

FILL FILL_2__13773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9353_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11624_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3364_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Ycalc [11])
);

FILL FILL_0__11339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3841_),
    .B(_3825_),
    .C(_3839_),
    .Y(_3846_)
);

AND2X2 _14096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6446_),
    .B(_6450_),
    .Y(_6451_)
);

FILL FILL_0__12700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14558_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5302_),
    .B(_5299_),
    .C(_5292_),
    .Y(_5304_)
);

NAND2X1 _12409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4943_),
    .B(_4946_),
    .Y(_4949_)
);

FILL FILL_1__14912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1395_),
    .C(_1423_),
    .Y(_1477_)
);

NAND2X1 _8164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf1),
    .B(_1027_),
    .Y(_1076_)
);

FILL FILL_1__10832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12297_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12582_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4236_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xin1 [1])
);

NAND3X1 _12162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(_4716_),
    .C(_4714_),
    .Y(_4717_)
);

FILL FILL_2__12624_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9789_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1701_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Acalc [0])
);

AOI21X1 _9369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2181_),
    .B(_2182_),
    .C(_1856_),
    .Y(_2183_)
);

FILL FILL_0__8624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14089_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6095_),
    .B(_6098_),
    .Y(_6156_)
);

OAI21X1 _13367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5192_),
    .B(_5807_),
    .C(_5809_),
    .Y(_5066_)
);

FILL FILL_0__14863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10363_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_810_),
    .C(_812_),
    .Y(_44_)
);

INVX1 _7435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_424_)
);

FILL FILL_2__13582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11568_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4409_),
    .B(_4397_),
    .C(_4410_),
    .Y(_4421_)
);

FILL FILL_0__9162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11148_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [4]),
    .Y(_4062_)
);

NAND2X1 _11013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .B(_3663_),
    .Y(_3664_)
);

FILL FILL_1__7597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5121_),
    .C(_5122_),
    .Y(_5123_)
);

OAI21X1 _12218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4745_),
    .B(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .C(_4770_),
    .Y(_4209_)
);

FILL FILL_1__14721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9323_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1114_),
    .C(_1294_),
    .Y(_1295_)
);

FILL FILL_1__10641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7246_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf78)
);

OAI21X1 _12391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4889_),
    .C(_4362__bF$buf4),
    .Y(_4932_)
);

FILL FILL_2__12853_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2104_),
    .B(_1917_),
    .C(_1848__bF$buf1),
    .Y(_2398_)
);

INVX1 _9178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_2000_)
);

FILL FILL_1__11846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8013_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10704_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2530_),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.Xcalc [3])
);

FILL FILL_0__10419_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .Y(_5974_)
);

NAND2X1 _13176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [9]),
    .B(_5174__bF$buf4),
    .Y(_5635_)
);

FILL FILL_0__14672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9638_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4472_),
    .Y(_4475_)
);

FILL FILL_0__9218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_642_),
    .Y(_643_)
);

AOI22X1 _7244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(_241_),
    .C(_240_),
    .D(_178_),
    .Y(_242_)
);

FILL FILL_2__13391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9391_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11662_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3402_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Yin12b [11])
);

FILL FILL_0__11377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3879_),
    .B(_3882_),
    .Y(_3883_)
);

DFFPOSX1 _8869_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_867_),
    .CLK(clk_bF$buf46),
    .Q(\genblk1[1].u_ce.Acalc [4])
);

OR2X2 _8449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1348_),
    .B(_1333_),
    .Y(_1349_)
);

INVX1 _8029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [9]),
    .Y(_948_)
);

FILL FILL_2__14596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7704_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9810_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1722_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin1 [1])
);

FILL FILL_1__13589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13169_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5340_)
);

OAI21X1 _12447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4982_),
    .B(_4978_),
    .C(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4984_)
);

NAND2X1 _12027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4583_),
    .B(_4587_),
    .Y(_4588_)
);

FILL FILL_1__14110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8662_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .Y(_3587_)
);

FILL FILL_0__8242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10648_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3227_),
    .B(_3224_),
    .Y(_3228_)
);

FILL FILL_0__10228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9447_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4292_),
    .C(_4293_),
    .Y(_4294_)
);

FILL FILL_0__9027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8403_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf3),
    .B(_799_),
    .C(_832_),
    .Y(_62_)
);

NAND3X1 _7473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf0),
    .B(_460_),
    .C(_438_),
    .Y(_461_)
);

FILL FILL_1__12193_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4445_),
    .B(_4457_),
    .C(_4455_),
    .Y(_4458_)
);

FILL FILL_0__11186_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4097_),
    .Y(_4098_)
);

INVX1 _11051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3700_)
);

FILL FILL_1__9608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1563_),
    .B(_1559_),
    .Y(_1564_)
);

NAND3X1 _8258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1165_),
    .C(_1161_),
    .Y(_1166_)
);

FILL FILL_1__10926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13398_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5155_),
    .C(_5156_),
    .Y(_5157_)
);

OR2X2 _12256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4804_),
    .Y(_4807_)
);

FILL FILL_0__13752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9361_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [18]),
    .B(FCW[18]),
    .Y(_7037_)
);

FILL FILL_0__14117_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .B(_6689_),
    .Y(_6691_)
);

FILL FILL_2__7284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10457_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10742_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2568_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin12b [7])
);

FILL FILL_0__10037_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .B(_2672__bF$buf2),
    .C(_3048_),
    .D(_2670_),
    .Y(_2531_)
);

FILL FILL_2__9850_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7949_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Acalc [8])
);

AOI21X1 _7529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_509_),
    .C(_507_),
    .Y(_514_)
);

NAND2X1 _7109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [7]),
    .B(_89_),
    .Y(_114_)
);

FILL FILL_0__14290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9676_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4510_),
    .B(_4494_),
    .C(_4506_),
    .Y(_4511_)
);

FILL FILL_0__9256_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510__bF$buf2),
    .B(_4148_),
    .C(_4147_),
    .Y(_3388_)
);

AOI21X1 _11107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3753_),
    .B(_3752_),
    .C(_3750_),
    .Y(_3754_)
);

FILL FILL_1__13610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14815_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_278_)
);

FILL FILL_0__13808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3918_),
    .B(_3917_),
    .Y(_3919_)
);

FILL FILL_1__9417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1379_),
    .B(_1384_),
    .Y(_1385_)
);

OAI21X1 _8067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_981_),
    .C(_982_),
    .Y(_983_)
);

FILL FILL_1__10315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7322_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4575_),
    .B(_4989_),
    .C(_5007_),
    .Y(_4239_)
);

NAND2X1 _12065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4624_)
);

FILL FILL_2__8701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6849_),
    .B(_6852_),
    .Y(_6861_)
);

DFFPOSX1 _14211_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.LoadCtl [2])
);

FILL FILL_2__7093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11273_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3623_),
    .B(_3620_),
    .Y(_3624_)
);

FILL FILL_2__8298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10686_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .B(_3263_),
    .Y(_3264_)
);

FILL FILL_0__10266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2837_),
    .Y(_2866_)
);

NOR2X1 _7758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_720_),
    .Y(_730_)
);

NAND3X1 _7338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_328_),
    .C(_331_),
    .Y(_332_)
);

FILL FILL_2__13065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9485_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4326_),
    .C(_4327_),
    .Y(_4328_)
);

FILL FILL_0__9065_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3969_),
    .B(_3954_),
    .Y(_3972_)
);

FILL FILL_0__12832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12412_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _9904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_2648_)
);

FILL FILL_1__8441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14624_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [7]),
    .B(_89_),
    .Y(_98_)
);

NAND2X1 _13902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6161_),
    .Y(_6266_)
);

FILL FILL_0__13617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11551_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1201_),
    .B(_1173_),
    .Y(_1202_)
);

FILL FILL_1__10964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7131_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4823_),
    .B(_4348__bF$buf2),
    .C(_4842_),
    .D(_4346_),
    .Y(_4213_)
);

FILL FILL_2__8510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3313_),
    .Y(_3314_)
);

DFFPOSX1 _13499_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.LoadCtl [4])
);

NAND3X1 _13079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(_5542_),
    .C(_5540_),
    .Y(_5543_)
);

FILL FILL_2__9715_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [15]),
    .B(_6833__bF$buf4),
    .C(En_bF$buf4),
    .Y(_7066_)
);

FILL FILL_0__14575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.X_ [0]),
    .B(_6724_),
    .Y(_6725_)
);

INVX1 _14020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6377_),
    .Y(_6379_)
);

FILL FILL_1__7712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3444_)
);

FILL FILL_0__10495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10075_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3064_),
    .B(_3084_),
    .Y(_3085_)
);

FILL FILL_2__10822_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7987_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_71_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Ain0 [0])
);

NAND2X1 _7567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_549_),
    .Y(_551_)
);

MUX2X1 _7147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_145_),
    .S(_135__bF$buf4),
    .Y(_149_)
);

FILL FILL_1__12287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .B(_4547_),
    .C(_4546_),
    .Y(_4548_)
);

FILL FILL_0__9294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_4172_)
);

AND2X2 _11145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_3789_),
    .Y(_3790_)
);

FILL FILL_0__12641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7607_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2475_),
    .C(_2493_),
    .Y(_1725_)
);

FILL FILL_1__8670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13846_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6083_),
    .B(_6082_),
    .C(_6021_),
    .Y(_6084_)
);

FILL FILL_0__13426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10353_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[6]),
    .Y(Dout[6])
);

FILL FILL_0__7780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8565_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3493_),
    .B(_3490_),
    .S(_3487__bF$buf3),
    .Y(_3494_)
);

FILL FILL_0__8145_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3120_),
    .B(_3118_),
    .C(_2686__bF$buf5),
    .Y(_3138_)
);

FILL FILL257550x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14909_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .Y(_765_)
);

INVX1 _7376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .Y(_368_)
);

FILL FILL_1__12096_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4363_),
    .C(_4364_),
    .Y(_4365_)
);

FILL FILL_0__11089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf1),
    .B(_3995_),
    .Y(_4008_)
);

FILL FILL_2__11836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7836_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2685_)
);

FILL FILL_0__7416_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_1834__bF$buf3),
    .C(_2328_),
    .D(_1832_),
    .Y(_1699_)
);

AOI21X1 _9102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1927_),
    .B(_1908_),
    .C(_1836_),
    .Y(_1928_)
);

OAI21X1 _12999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5187_),
    .C(_5465_),
    .Y(_5466_)
);

DFFPOSX1 _12579_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4233_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[5].u_ce.Xin12b [4])
);

OR2X2 _12159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4713_),
    .B(_4711_),
    .Y(_4714_)
);

FILL FILL_1__14662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert221 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert223 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6286_),
    .B(_6301_),
    .Y(_6303_)
);

FILL FILL_0__13655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert224 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13235_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Ycalc [11]),
    .C(_5889_),
    .Y(_5902_)
);

NAND2X1 _13100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .B(_5562_),
    .Y(_5563_)
);

FILL FILL_0_BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x244950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6946_),
    .B(_6942_),
    .Y(_6947_)
);

NAND2X1 _14305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Xin12b [6]),
    .Y(_6607_)
);

FILL FILL_1__11787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8374_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3335_),
    .B(_3317_),
    .C(_3336_),
    .Y(_2566_)
);

NAND2X1 _10225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2954_),
    .B(_2955_),
    .Y(_2956_)
);

FILL FILL_2__9753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14718_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_182_),
    .S(_135__bF$buf3),
    .Y(_186_)
);

NAND2X1 _11183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3795_),
    .B(_3812_),
    .Y(_3826_)
);

FILL FILL_2__11225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7645_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_2483_),
    .C(_1749_),
    .Y(_1742_)
);

FILL FILL_0__7225_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2146_),
    .B(_2145_),
    .C(_1836_),
    .Y(_2147_)
);

OAI21X1 _12388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4354_),
    .C(_4324__bF$buf0),
    .Y(_4929_)
);

FILL FILL_1__14471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14669_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14534_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6522_),
    .CLK(clk_bF$buf38),
    .Q(\u_ot.Xin0 [0])
);

FILL FILL_0__14249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(_6463_),
    .Y(_6464_)
);

FILL FILL_1__7806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11176_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3530_),
    .B(_3527_),
    .S(_3487__bF$buf3),
    .Y(_3531_)
);

FILL FILL_0__10589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10169_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3169_),
    .B(_3173_),
    .Y(_3174_)
);

NAND2X1 _10034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf3),
    .B(_2722_),
    .Y(_2773_)
);

FILL FILL_0__11950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11110_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf3),
    .B(_1481_),
    .Y(_1494_)
);

FILL FILL_0__9388_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11659_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3399_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xin0 [0])
);

OR2X2 _11239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3875_),
    .B(_3872_),
    .Y(_3880_)
);

FILL FILL256650x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12315_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12600_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4254_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ain12b [9])
);

DFFPOSX1 _9807_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1719_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin12b [4])
);

FILL FILL_1__8764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14107_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6172_),
    .B(_6160_),
    .C(_6018_),
    .Y(_6174_)
);

FILL FILL_1__9969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .B(_1106_),
    .Y(_1110_)
);

FILL FILL_1__10867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7874_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .B(_2713_),
    .C(_2711_),
    .Y(_2721_)
);

FILL FILL_0__7454_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .B(gnd),
    .S(_2361_),
    .Y(_2363_)
);

AOI21X1 _9140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1962_),
    .B(_1959_),
    .C(_1952_),
    .Y(_1964_)
);

NAND3X1 _12197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf1),
    .B(_4749_),
    .C(_4746_),
    .Y(_4750_)
);

FILL FILL_0__10801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6982_)
);

FILL FILL_0__14058_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .C(\u_ot.ISreg_bF$buf4 ),
    .Y(_6641_)
);

FILL FILL_1__7615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3349_),
    .B(_2597_),
    .C(_2591_),
    .Y(_2584_)
);

FILL FILL_0__10398_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf3),
    .B(_2990_),
    .C(_2991_),
    .Y(_2992_)
);

OAI21X1 _8831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1559_),
    .B(_1648_),
    .C(_913_),
    .Y(_906_)
);

NAND2X1 _8411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1298_),
    .Y(_1312_)
);

OR2X2 _11888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4454_),
    .B(_4453_),
    .Y(_4455_)
);

FILL FILL_0__9197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4094_),
    .B(_4093_),
    .Y(_4095_)
);

OAI21X1 _11048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3659_),
    .B(_3688_),
    .C(_3687_),
    .Y(_3697_)
);

FILL FILL_1__13971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12124_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1840_),
    .C(_1810__bF$buf1),
    .Y(_2415_)
);

FILL FILL_1__8993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13749_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .B(_5961_),
    .C(_5991_),
    .Y(_5992_)
);

FILL FILL_0__13329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7032_),
    .B(_7021_),
    .C(_7033_),
    .Y(_7034_)
);

FILL FILL_2_BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8048_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10739_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2565_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Yin12b [8])
);

OR2X2 _10319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3028_),
    .B(_3045_),
    .Y(_3046_)
);

FILL FILL_1__12822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14287_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [0]),
    .B(_6813_),
    .C(_6814_),
    .Y(\a[0] [0])
);

OAI21X1 _14152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6477_),
    .B(_5887_),
    .C(_6484_),
    .Y(_5881_)
);

FILL FILL_1__7844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x133350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert152 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert154 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert155 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert157 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert159 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _10492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3206_),
    .D(_3208_),
    .Y(_2541_)
);

INVX1 _10072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2809_)
);

FILL FILL_1__8629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8209_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_672_),
    .Y(_675_)
);

OAI21X1 _7279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_254_),
    .C(_271_),
    .Y(_275_)
);

INVX1 _8640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .Y(_1529_)
);

OAI21X1 _8220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1128_),
    .B(_1113_),
    .C(_1065_),
    .Y(_1130_)
);

INVX4 _11697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .Y(_4275_)
);

NAND2X1 _11277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3912_),
    .B(_3915_),
    .Y(_3916_)
);

FILL FILL_2__7913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7739_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _9845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2595_)
);

FILL FILL_0__7319_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf2),
    .B(_2235_),
    .C(_2232_),
    .Y(_2236_)
);

INVX8 _9005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .Y(_1834_)
);

FILL FILL_1__8382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13558_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6200_),
    .B(_6209_),
    .C(_6193_),
    .Y(_6210_)
);

FILL FILL_0__13138_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5832_),
    .B(_5104_),
    .C(_5099_),
    .Y(_5092_)
);

OAI21X1 _13003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5338_),
    .C(_5469_),
    .Y(_5470_)
);

FILL FILL_1__9587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10065_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6858_)
);

DFFPOSX1 _14208_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5884_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Ain12b [11])
);

FILL FILL_0__7492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12277_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_83_),
    .C(_77_),
    .Y(_70_)
);

FILL FILL_0__8697_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3615_),
    .B(_3616_),
    .Y(_3621_)
);

FILL FILL_0__8277_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3260_),
    .Y(_3261_)
);

OR2X2 _10128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2837_),
    .B(_2841_),
    .Y(_2863_)
);

FILL FILL_1__12631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6547_),
    .B(_6562__bF$buf3),
    .C(_6671_),
    .D(_6672_),
    .Y(_6505_)
);

FILL FILL_1__7653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8018_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [11]),
    .C(_86_),
    .Y(_95_)
);

AND2X2 _11086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3721_),
    .B(_3733_),
    .Y(_3734_)
);

FILL FILL_2__7722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7548_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2450_),
    .Y(_2451_)
);

FILL FILL_0__7128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_2051_),
    .C(_2048_),
    .Y(_2054_)
);

FILL FILL_1__8191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13787_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [10]),
    .Y(_6027_)
);

FILL FILL_0__13367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5687_),
    .B(_5685_),
    .Y(_5688_)
);

FILL FILL_1__9396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10294_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .B(_6833__bF$buf2),
    .C(_7064_),
    .Y(_6792_)
);

NAND2X1 _14437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [5]),
    .B(_6721_),
    .Y(_6722_)
);

INVX1 _14017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6375_),
    .Y(_6376_)
);

FILL FILL_1__7709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12086_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _7720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .C(_692_),
    .D(_694_),
    .Y(_27_)
);

FILL FILL_1__11499_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_295_)
);

FILL FILL_1__11079_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(\genblk1[4].u_ce.LoadCtl [3]),
    .Y(_3441_)
);

FILL FILL_0__8086_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3042_),
    .B(_3043_),
    .C(_2653_),
    .Y(_3082_)
);

FILL FILL_1__12860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11013_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14190_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5866_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin12b [4])
);

INVX4 _8925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .Y(_1761_)
);

NAND2X1 _8505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1401_),
    .Y(_1402_)
);

FILL FILL_1__7882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5391_),
    .C(_5388_),
    .Y(_5394_)
);

FILL FILL_0__12638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5009_),
    .B(_4273_),
    .C(_5017_),
    .Y(_4247_)
);

FILL FILL_1__8667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8247_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6078_),
    .B(_6080_),
    .Y(_6081_)
);

BUFX2 BUFX2_insert200 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .Y(_4348__bF$buf4)
);

BUFX2 BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .Y(_4348__bF$buf3)
);

BUFX2 BUFX2_insert202 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .Y(_4348__bF$buf2)
);

BUFX2 BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .Y(_4348__bF$buf1)
);

BUFX2 BUFX2_insert204 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .Y(_4348__bF$buf0)
);

BUFX2 BUFX2_insert205 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert207 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf0 )
);

FILL FILL_0__12391_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert209 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1811__bF$buf4)
);

FILL FILL_0__7777_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(_2629_),
    .C(_2606_),
    .Y(_2630_)
);

FILL FILL_0__7357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2248_),
    .Y(_2273_)
);

OAI21X1 _9043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1846_),
    .C(_1871_),
    .Y(_1872_)
);

FILL FILL_1__11711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8736_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6245_),
    .Y(_6246_)
);

FILL FILL_0__13596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13176_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13461_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5061_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Xin12b [8])
);

AND2X2 _13041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5506_),
    .B(_5489_),
    .Y(_5507_)
);

FILL FILL_2__13923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9503_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .Y(_6893_)
);

INVX1 _14246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [10]),
    .Y(_6557_)
);

FILL FILL_1__7518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14708_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf4 )
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf3 )
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf2 )
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf1 )
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf0 )
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf4 )
);

AND2X2 _10586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3292_),
    .B(_3295_),
    .Y(_3296_)
);

INVX1 _10166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .Y(_2899_)
);

FILL FILL_2__10208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1607_),
    .C(_1605_),
    .Y(_1616_)
);

AND2X2 _8314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1207_),
    .B(_1219_),
    .Y(_1220_)
);

FILL FILL_1__7691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12867_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5186_),
    .C(_5211_),
    .Y(_5212_)
);

FILL FILL_0__12447_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348__bF$buf1),
    .B(_4857_),
    .C(_4858_),
    .Y(_4215_)
);

FILL FILL_0__12027_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(vdd),
    .C(_2649__bF$buf2),
    .Y(_2682_)
);

AND2X2 _9519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2325_),
    .Y(_2326_)
);

FILL FILL_1__8476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert190 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert192 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert193 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5971_),
    .B(_6297_),
    .C(_6296_),
    .Y(_6300_)
);

FILL FILL_0_BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert195 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[7].u_ce.Ycalc [0]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Ycalc [2]),
    .Y(_5900_)
);

FILL FILL_0_BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert197 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert199 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7586_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Xin12b [9]),
    .Y(_2482_)
);

FILL FILL_0__7166_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .Y(_2090_)
);

FILL FILL_1__11940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10513_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6063_),
    .C(_5951_),
    .Y(_6064_)
);

NAND2X1 _13270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5719_),
    .B(_5722_),
    .Y(_5724_)
);

FILL FILL_2__13732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9312_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14895_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6786_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.acc_reg [19])
);

OAI21X1 _14475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6707_),
    .B(_6724_),
    .C(_6746_),
    .Y(_6525_)
);

NOR2X1 _14055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6411_),
    .Y(_6412_)
);

FILL FILL_1__7747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7327_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3073_),
    .B(_3102_),
    .C(_3075_),
    .Y(_3118_)
);

FILL FILL_0__11891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11051_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Xcalc [10]),
    .C(_1762_),
    .Y(_1795_)
);

OAI21X1 _8543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1433_),
    .C(_1429_),
    .Y(_1438_)
);

AND2X2 _8123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1037_),
    .Y(_1038_)
);

FILL FILL_1__7080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13263_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5430_)
);

FILL FILL_0__12676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12256_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12541_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4195_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[5].u_ce.Ycalc [4])
);

INVX1 _12121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4677_),
    .Y(_4678_)
);

NAND2X1 _9748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [6]),
    .B(_2483_),
    .Y(_2513_)
);

AND2X2 _9328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2143_),
    .Y(_2144_)
);

FILL FILL_1__8285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14048_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6116_),
    .Y(_6117_)
);

AOI21X1 _13326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5777_),
    .B(_5772_),
    .C(_5770_),
    .Y(_5778_)
);

FILL FILL_0__14822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7395_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1895_),
    .B(_1883_),
    .C(_1896_),
    .Y(_1907_)
);

FILL FILL_0__10322_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_781_),
    .Y(_782_)
);

FILL FILL_2__13961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11527_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(\genblk1[5].u_ce.Xin0 [1]),
    .S(vdd),
    .Y(_4383_)
);

FILL FILL_0__9121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11107_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [4]),
    .B(_6562__bF$buf0),
    .Y(_6589_)
);

FILL FILL_1__7556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1640_),
    .B(_1645_),
    .C(_1646_),
    .Y(_879_)
);

INVX1 _8352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1255_),
    .Y(_1256_)
);

FILL FILL_1__10600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13072_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5235_),
    .B(_5223_),
    .C(_5236_),
    .Y(_5247_)
);

FILL FILL_0__12485_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4888_),
    .B(_4892_),
    .Y(_4894_)
);

FILL FILL_0__12065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12812_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(\genblk1[2].u_ce.ISout ),
    .Y(_2719_)
);

OAI21X1 _9557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .B(_2352_),
    .C(_2357_),
    .Y(_2360_)
);

INVX1 _9137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1958_),
    .Y(_1961_)
);

FILL FILL_1__8094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .B(_6335_),
    .C(_6276_),
    .Y(_6336_)
);

INVX1 _13555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_5934_)
);

OAI21X1 _13135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5571_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5596_),
    .Y(_5047_)
);

FILL FILL_0__14631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10131_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_588_),
    .C(_561_),
    .Y(_604_)
);

OAI21X1 _7203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158__bF$buf2),
    .B(_203_),
    .C(_159_),
    .Y(_1_)
);

FILL FILL_2__13770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9350_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11621_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3361_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Ycalc [8])
);

FILL FILL_0__11336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3825_),
    .B(_3842_),
    .Y(_3844_)
);

NOR2X1 _14093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6204_),
    .B(_6447_),
    .Y(_6448_)
);

NAND2X1 _8828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [0]),
    .B(_1648_),
    .Y(_912_)
);

OAI21X1 _8408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996__bF$buf1),
    .B(_1309_),
    .C(_1283_),
    .Y(_852_)
);

FILL FILL_1__7785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13128_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5298_),
    .Y(_5301_)
);

NAND2X1 _12406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4944_),
    .B(_4945_),
    .Y(_4946_)
);

FILL FILL_0__13902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9511_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1452_),
    .Y(_1474_)
);

INVX1 _8161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .Y(_1073_)
);

FILL FILL_2__7434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12201_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9786_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1698_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [9])
);

OAI21X1 _9366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2159_),
    .B(_2150_),
    .C(_1848__bF$buf2),
    .Y(_2180_)
);

FILL FILL_0__8621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14086_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6135_),
    .B(_5949__bF$buf2),
    .C(_6153_),
    .D(_6133_),
    .Y(_5844_)
);

FILL FILL_0__13079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5807_),
    .Y(_5808_)
);

FILL FILL_0__14860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [1]),
    .B(_6811_),
    .Y(_6812_)
);

OAI21X1 _14149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6483_)
);

FILL FILL_0__10780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10360_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_810_),
    .Y(_811_)
);

OAI21X1 _7432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_421_),
    .C(_230_),
    .Y(_422_)
);

NOR2X1 _10489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3198_),
    .Y(_3206_)
);

OAI21X1 _10069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2806_),
    .B(_2805_),
    .C(_2744_),
    .Y(_2807_)
);

FILL FILL_1__12992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11565_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4418_),
    .B(_4416_),
    .C(_4396_),
    .Y(_4193_)
);

FILL FILL_0__11145_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4049_),
    .B(_4058_),
    .C(_4059_),
    .Y(_4060_)
);

AOI21X1 _11010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3617_),
    .B(_3619_),
    .C(_3607_),
    .Y(_3661_)
);

NAND2X1 _8637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain1 [0]),
    .B(_1525_),
    .Y(_1526_)
);

INVX1 _8217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1126_),
    .Y(_1127_)
);

FILL FILL_1__7594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13357_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5118_),
    .C(_5119_),
    .Y(_5120_)
);

NOR2X1 _12215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4763_),
    .B(_4767_),
    .Y(_4768_)
);

FILL FILL_0__13711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9320_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1160_),
    .C(_1291_),
    .Y(_1292_)
);

FILL FILL_0__14916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7489_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2395_),
    .B(_2394_),
    .C(_2385_),
    .Y(_1705_)
);

AOI21X1 _9175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_1980_),
    .C(_1992_),
    .Y(_1997_)
);

FILL FILL_1__11843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8010_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10701_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2527_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xcalc [0])
);

FILL FILL_0__10416_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_5971_)
);

OR2X2 _13173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5630_),
    .Y(_5633_)
);

OAI21X1 _7908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_76_)
);

FILL FILL_2__13215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9635_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf1),
    .B(_4470_),
    .C(_4471_),
    .Y(_4472_)
);

FILL FILL_0__9215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7014_),
    .B(_6887_),
    .Y(_7015_)
);

OAI21X1 _14378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6661_),
    .C(_6664_),
    .Y(_6670_)
);

INVX1 _7661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_639_),
    .Y(_640_)
);

OAI21X1 _7241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf0),
    .B(_237_),
    .C(_238_),
    .Y(_239_)
);

NAND2X1 _10298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3009_),
    .B(_3024_),
    .Y(_3026_)
);

FILL FILL_1__12381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11374_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8866_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_864_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Acalc [1])
);

INVX1 _8446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1345_),
    .Y(_1346_)
);

OAI21X1 _8026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_945_),
    .C(_930_),
    .Y(_946_)
);

FILL FILL_2__14593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12999_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5336_),
    .B(_5320_),
    .C(_5332_),
    .Y(_5337_)
);

FILL FILL_0__12159_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .B(_4362__bF$buf4),
    .Y(_4981_)
);

AND2X2 _12024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4579_),
    .B(_4362__bF$buf3),
    .Y(_4585_)
);

FILL FILL_0__13940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8188_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6024_)
);

NOR2X1 _13229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5684_),
    .Y(_5685_)
);

FILL FILL_0__14725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8677_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3583_),
    .Y(_3584_)
);

FILL FILL_2__8257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10645_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(gnd),
    .C(_2686__bF$buf1),
    .Y(_3225_)
);

FILL FILL_0__10225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_684_),
    .Y(_692_)
);

FILL FILL_2__13024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9444_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4291_),
    .B(_4290_),
    .Y(\a[6] [1])
);

FILL FILL_0__9024_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14187_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5863_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xin12b [9])
);

FILL FILL_1__7879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8400_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [0]),
    .B(_799_),
    .Y(_831_)
);

NAND2X1 _7470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf1),
    .B(_457_),
    .Y(_458_)
);

FILL FILL_1__12190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9605_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(_992_),
    .Y(_1561_)
);

NOR2X1 _8255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf3),
    .B(_1162_),
    .Y(_1163_)
);

FILL FILL_1__10923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10503_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .Y(_972__bF$buf0)
);

FILL FILL_0__7510_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert171 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 )
);

FILL FILL_1__13395_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert173 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert174 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert176 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .Y(_2649__bF$buf4)
);

BUFX2 BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .Y(_2649__bF$buf3)
);

BUFX2 BUFX2_insert178 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .Y(_2649__bF$buf2)
);

OAI21X1 _12673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5152_),
    .C(_5153_),
    .Y(_5154_)
);

FILL FILL_0__12388_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .Y(_2649__bF$buf1)
);

AOI21X1 _12253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4803_),
    .B(_4802_),
    .C(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4804_)
);

FILL FILL_1__11708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8715_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf2),
    .B(_6242_),
    .Y(_6243_)
);

DFFPOSX1 _13458_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5058_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Acalc [11])
);

INVX1 _13038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .Y(_5504_)
);

FILL FILL_0__14114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10034_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7946_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Acalc [5])
);

NAND2X1 _7526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(_510_),
    .Y(_512_)
);

OAI21X1 _7106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Ycalc [11]),
    .C(_86_),
    .Y(_111_)
);

FILL FILL_2__13253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9673_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4479_),
    .C(_4507_),
    .Y(_4508_)
);

FILL FILL_0__9253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11239_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4146_),
    .B(_4145_),
    .C(_4136_),
    .Y(_3387_)
);

AOI21X1 _11104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3726_),
    .B(_3728_),
    .C(_3722_),
    .Y(_3751_)
);

FILL FILL_1__7688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7268_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(\genblk1[6].u_ce.Xin0 [1]),
    .S(gnd),
    .Y(_5209_)
);

NAND2X1 _12309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4854_),
    .B(_4855_),
    .Y(_4856_)
);

FILL FILL_1__14812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1340_),
    .B(_1337_),
    .Y(_1382_)
);

MUX2X1 _8064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(_976_),
    .S(_973__bF$buf4),
    .Y(_980_)
);

FILL FILL_1__10312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.X_ [1]),
    .Y(_5006_)
);

NAND3X1 _12062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf2),
    .B(_4617_),
    .C(_4620_),
    .Y(_4621_)
);

OAI21X1 _9689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2480_)
);

INVX1 _9269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2087_)
);

FILL FILL_1__11937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8104_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6055_),
    .B(_6054_),
    .Y(_6061_)
);

OAI21X1 _13267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5445_),
    .C(_5720_),
    .Y(_5721_)
);

FILL FILL_0__14763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10263_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_725_),
    .Y(_727_)
);

INVX1 _7335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .Y(_329_)
);

FILL FILL_2__13062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11468_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _11753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_4325_)
);

FILL FILL_0__9062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11048_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3969_),
    .B(_3954_),
    .C(_3508_),
    .Y(_3970_)
);

FILL FILL_1__7497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2640_),
    .B(_2597_),
    .C(_2645_),
    .Y(\genblk1[3].u_ce.X_ [1])
);

INVX1 _12958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5427_)
);

DFFPOSX1 _12538_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4192_),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[5].u_ce.ISout )
);

AOI21X1 _12118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4621_),
    .B(_4627_),
    .C(_4653_),
    .Y(_4675_)
);

FILL FILL_1__14621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1198_),
    .C(_1199_),
    .Y(_1200_)
);

FILL FILL_1__10961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7146_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4828_),
    .B(_4839_),
    .Y(_4840_)
);

NAND2X1 _9498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .B(_2305_),
    .Y(_2306_)
);

OAI21X1 _9078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1904_),
    .B(_1902_),
    .C(_1882_),
    .Y(_1679_)
);

FILL FILL_1__11746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8333_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [5]),
    .B(_2599_),
    .Y(_3311_)
);

FILL FILL_0__10319_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13496_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.LoadCtl [1])
);

OR2X2 _13076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .B(_5537_),
    .Y(_5540_)
);

FILL FILL_2__13958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9538_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .S(vdd),
    .Y(_4380_)
);

FILL FILL_0__9118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10072_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7984_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_68_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.Ain12b [5])
);

AOI21X1 _7564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_547_),
    .C(_176_),
    .Y(_548_)
);

INVX1 _7144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .Y(_146_)
);

FILL FILL_2__13291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4538_),
    .B(_4544_),
    .C(_4541_),
    .Y(_4545_)
);

FILL FILL_0__11697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9291_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4151_),
    .Y(_4170_)
);

FILL FILL_0__11277_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3607_),
    .C(_3786_),
    .Y(_3787_)
);

FILL FILL_2__11604_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1641_),
    .C(_1644_),
    .Y(_878_)
);

NAND2X1 _8349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1252_),
    .B(_1228_),
    .Y(_1253_)
);

FILL FILL_0__7604_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.X_ [1]),
    .Y(_2492_)
);

FILL FILL_1__13069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5244_),
    .B(_5242_),
    .C(_5222_),
    .Y(_5031_)
);

OAI21X1 _12347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_4891_)
);

FILL FILL_1__14850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10350_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[3]),
    .Y(Dout[3])
);

FILL FILL_0__14628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8562_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .Y(_3491_)
);

FILL FILL_0__8142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3134_),
    .Y(_3135_)
);

FILL FILL_0__14381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9347_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11618_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3358_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[4].u_ce.Ycalc [5])
);

FILL FILL_1__13701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8303_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(_158__bF$buf4),
    .C(_761_),
    .D(_762_),
    .Y(_32_)
);

AND2X2 _7373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_307_),
    .Y(_365_)
);

FILL FILL_1__12093_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _11791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4362_)
);

FILL FILL_0__11086_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [11]),
    .B(_3510__bF$buf4),
    .Y(_4005_)
);

FILL FILL_1__9928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1826_),
    .Y(_1828_)
);

INVX1 _8578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [10]),
    .Y(_1471_)
);

INVX1 _8158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .Y(_1070_)
);

FILL FILL_1__10826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5463_)
);

DFFPOSX1 _12576_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4230_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Xin12b [9])
);

INVX1 _12156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4710_),
    .Y(_4711_)
);

FILL FILL_0__13652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14437_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [10]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf1),
    .Y(_6945_)
);

FILL FILL_0__14017_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6598_),
    .B(_6595_),
    .C(_6586_),
    .Y(_6604_)
);

FILL FILL_2__7184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3333_),
    .B(_3317_),
    .C(_3334_),
    .Y(_2565_)
);

FILL FILL_0__10357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .B(_2952_),
    .Y(_2953_)
);

NAND2X1 _7849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(_807_),
    .Y(_809_)
);

NOR3X1 _7429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_418_),
    .C(_402_),
    .Y(_419_)
);

FILL FILL_1__12989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9576_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4414_),
    .B(_4415_),
    .C(_4350_),
    .Y(_4416_)
);

FILL FILL_0__9156_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4056_),
    .Y(_4057_)
);

NAND2X1 _11007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3651_),
    .B(_3654_),
    .Y(_3658_)
);

FILL FILL_1__13930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14715_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .Y(_183_)
);

FILL FILL_0__13708_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510__bF$buf4),
    .B(_3823_),
    .C(_3797_),
    .Y(_3366_)
);

FILL FILL_1__9737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11222_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1288_),
    .B(_1286_),
    .S(_973__bF$buf4),
    .Y(_1289_)
);

FILL FILL_1__10635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7222_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4904_),
    .B(_4918_),
    .C(_4916_),
    .Y(_4926_)
);

FILL FILL_2__8601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14666_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14531_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6519_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin12b [5])
);

FILL FILL_0__14246_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Xin12b [9]),
    .Y(_6462_)
);

FILL FILL_1__7803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11173_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3528_)
);

FILL FILL_2__8198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10166_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2927_),
    .B(_3170_),
    .Y(_3171_)
);

INVX1 _10031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2770_)
);

NAND3X1 _7658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_629_),
    .C(_636_),
    .Y(_637_)
);

NAND2X1 _7238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_236_)
);

FILL FILL_1__12798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9385_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11656_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3396_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [5])
);

NOR2X1 _11236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3855_),
    .B(_3874_),
    .Y(_3877_)
);

FILL FILL_0__12732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12312_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9804_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1716_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin12b [9])
);

FILL FILL_1__8761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13937_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [9]),
    .B(_6170_),
    .C(_6169_),
    .Y(_6171_)
);

FILL FILL_0__13517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11451_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .B(_1102_),
    .Y(_1107_)
);

FILL FILL_1__10864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7451_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4706_),
    .C(_4728_),
    .Y(_4747_)
);

FILL FILL_2__8410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8656_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3581_)
);

FILL FILL_0__8236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3209_),
    .B(_3222_),
    .Y(_2542_)
);

OAI21X1 _13399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5149_),
    .C(_5826_),
    .Y(_5081_)
);

FILL FILL_2__9615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14475_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6963_),
    .B(_6978_),
    .C(_6971_),
    .Y(_6979_)
);

FILL FILL_0__14055_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6637_),
    .Y(_6638_)
);

FILL FILL_1__7612_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_2590_)
);

FILL FILL_0__10395_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2884_),
    .Y(_2989_)
);

FILL FILL_1__8817_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_133_),
    .C(_829_),
    .Y(_59_)
);

INVX1 _7467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .Y(_455_)
);

FILL FILL_1__12187_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf2),
    .B(_4450_),
    .C(_4451_),
    .Y(_4452_)
);

FILL FILL_0__9194_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4091_),
    .B(_4051_),
    .Y(_4092_)
);

OAI21X1 _11045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3692_),
    .B(_3690_),
    .C(_3694_),
    .Y(_3695_)
);

FILL FILL_2__11927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7507_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2404_),
    .C(_2402_),
    .Y(_2412_)
);

FILL FILL_1__8990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13746_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5988_),
    .Y(_5989_)
);

FILL FILL_0__13326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10253_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7029_),
    .B(_7030_),
    .C(_7031_),
    .Y(_6784_)
);

FILL FILL_2__7698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8045_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10736_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2562_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Xin0 [1])
);

OAI21X1 _10316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3039_),
    .C(_3034_),
    .Y(_3043_)
);

FILL FILL_0__11812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert121 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert123 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert124 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert126 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert128 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10951_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(gnd),
    .C(_671_),
    .Y(_672_)
);

FILL FILL_1__14809_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_272_),
    .C(_160_),
    .Y(_273_)
);

NOR2X1 _11694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4271_),
    .Y(_4272_)
);

NOR3X1 _11274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .B(_3893_),
    .C(_3897_),
    .Y(_3913_)
);

FILL FILL_2__11736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7736_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9842_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.LoadCtl [5])
);

FILL FILL_0__7316_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf1),
    .B(_2192_),
    .C(_2214_),
    .Y(_2233_)
);

INVX2 _9002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1831_),
    .Y(_1832_)
);

NAND3X1 _12899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5364_),
    .B(_5370_),
    .C(_5367_),
    .Y(_5371_)
);

OAI21X1 _12479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4995_),
    .B(_4273_),
    .C(_5004_),
    .Y(_4236_)
);

NOR2X1 _12059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_4618_)
);

FILL FILL_1__14562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13555_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6204_),
    .B(_6186_),
    .Y(_6207_)
);

FILL FILL_0__13135_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Ain1 [0]),
    .Y(_5098_)
);

MUX2X1 _13000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .B(_5464_),
    .S(_5151__bF$buf3),
    .Y(_5467_)
);

FILL FILL_1__9584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x154950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6854_),
    .B(_6855_),
    .C(_6834_),
    .Y(_6769_)
);

DFFPOSX1 _14205_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5881_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Yin1 [1])
);

FILL FILL_1__11267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8694_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3586_),
    .Y(_3618_)
);

FILL FILL_0__8274_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [6]),
    .B(_3257_),
    .Y(_3258_)
);

NOR2X1 _10125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2822_),
    .B(_2850_),
    .Y(_2860_)
);

FILL FILL_2__9653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14618_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Acalc [0]),
    .C(_91_),
    .D(_92_),
    .Y(_93_)
);

OAI21X1 _11083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3723_),
    .C(_3725_),
    .Y(_3731_)
);

FILL FILL_2__11965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7545_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2412_),
    .C(_2446_),
    .Y(_2448_)
);

FILL FILL_0__7125_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .Y(_2051_)
);

NOR2X1 _12288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4830_),
    .B(_4832_),
    .Y(_4837_)
);

FILL FILL_2__8924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14569_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [12]),
    .B(_6833__bF$buf3),
    .C(En_bF$buf4),
    .Y(_7063_)
);

FILL FILL_0__14149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [2]),
    .B(\u_ot.LoadCtl [0]),
    .Y(_6719_)
);

INVX1 _14014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .Y(_6373_)
);

FILL FILL_1__7706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.LoadCtl [3]),
    .Y(_3438_)
);

FILL FILL_0__8083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(_3078_),
    .Y(_3079_)
);

FILL FILL_0__11850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11010_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1757_),
    .Y(_1758_)
);

NOR3X1 _8502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1379_),
    .C(_1383_),
    .Y(_1399_)
);

NOR2X1 _11979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4517_),
    .B(_4513_),
    .Y(_4542_)
);

FILL FILL_0__9288_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3535_),
    .C(_4168_),
    .Y(_3400_)
);

NAND2X1 _11139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3784_)
);

FILL FILL_1__13642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12635_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5389_),
    .Y(_5391_)
);

FILL FILL_0__12215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_5000_),
    .Y(_5016_)
);

OAI21X1 _9707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .B(_1759_),
    .C(_2490_),
    .Y(_1722_)
);

FILL FILL_1__8664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x230550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14007_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6067_),
    .B(_6074_),
    .C(_6077_),
    .Y(_6078_)
);

FILL FILL_1__9869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11774_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_1014_)
);

FILL FILL_1__10347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7774_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [5]),
    .Y(_2627_)
);

FILL FILL_0__7354_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1849_),
    .B(_2268_),
    .C(_2269_),
    .Y(_2270_)
);

MUX2X1 _9040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(\genblk1[2].u_ce.Xin0 [1]),
    .S(gnd),
    .Y(_1869_)
);

AOI21X1 _12097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4651_),
    .B(_4654_),
    .C(_4373_),
    .Y(_4655_)
);

FILL FILL_2__12979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6890_)
);

INVX1 _14243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [9]),
    .Y(_6555_)
);

FILL FILL_1__7515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14705_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf1),
    .B(\genblk1[3].u_ce.Ain12b [9]),
    .Y(_3293_)
);

FILL FILL_0__10298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2895_),
    .B(_2883_),
    .C(_2741_),
    .Y(_2897_)
);

FILL FILL257250x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10625_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_1612_),
    .Y(_1614_)
);

OAI21X1 _8311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1209_),
    .C(_1211_),
    .Y(_1217_)
);

NAND3X1 _11788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf0),
    .B(_4358_),
    .C(_4357_),
    .Y(_4359_)
);

FILL FILL_0__9097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .B(_3990_),
    .Y(_4003_)
);

FILL FILL_1__13871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(_2678_),
    .Y(_2679_)
);

NOR2X1 _9516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2318_),
    .Y(_2323_)
);

FILL FILL_1__8473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert161 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert162 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13649_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6290_),
    .B(_6293_),
    .C(_6295_),
    .Y(_6297_)
);

FILL FILL_0_BUFX2_insert164 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [6]),
    .B(_5891_),
    .Y(_5897_)
);

FILL FILL_0_BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert166 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert168 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert169 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10156_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6941_),
    .B(_6938_),
    .Y(_6942_)
);

FILL FILL_0__7583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2925_),
    .B(_3313_),
    .C(_3332_),
    .Y(_2564_)
);

MUX2X1 _10219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2949_),
    .B(_2947_),
    .S(_2649__bF$buf0),
    .Y(_2950_)
);

FILL FILL_1__12722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11715_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14892_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6783_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.acc_reg [16])
);

NAND2X1 _14472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Y_ [0]),
    .B(_6724_),
    .Y(_6745_)
);

OAI22X1 _14052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5909_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6409_),
    .D(_6407_),
    .Y(_5856_)
);

FILL FILL_1__7744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13507_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3081_),
    .B(_3109_),
    .Y(_3115_)
);

FILL FILL_1__8949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10434_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [7]),
    .Y(_581_)
);

INVX1 _7179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_180_)
);

AOI22X1 _8960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Ycalc [1]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1793_)
);

INVX1 _8540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .Y(_1436_)
);

AOI21X1 _8120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .B(_1026_),
    .C(_1009_),
    .Y(_1035_)
);

OAI21X1 _11597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4185_),
    .B(_4159_),
    .C(_4189_),
    .Y(_3417_)
);

NAND2X1 _11177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3820_),
    .Y(_3821_)
);

FILL FILL_2__7813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7639_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [1]),
    .Y(_2511_)
);

FILL FILL_0__7219_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2137_),
    .B(_2140_),
    .C(_1859_),
    .Y(_2141_)
);

FILL FILL_1__8282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13878_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6076_),
    .B(_6092_),
    .C(_6075_),
    .Y(_6114_)
);

FILL FILL_0__13038_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5774_),
    .B(_5742_),
    .C(_5773_),
    .Y(_5775_)
);

FILL FILL_1__9487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10385_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14528_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6516_),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.Xin12b [6])
);

OAI21X1 _14108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6460_)
);

FILL FILL_0__7392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf3),
    .B(\genblk1[0].u_ce.Ain12b [9]),
    .Y(_779_)
);

FILL FILL_0__8597_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3525_)
);

FILL FILL_0__8177_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3159_),
    .Y(_3168_)
);

AOI22X1 _10028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2743_),
    .B(_2672__bF$buf0),
    .C(_2767_),
    .D(_2744_),
    .Y(_2518_)
);

FILL FILL_1__12951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11104_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6573_),
    .B(_6582_),
    .Y(_6586_)
);

FILL FILL_1__7553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7868_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2716_),
    .B(_2715_),
    .C(_2674_),
    .Y(_2717_)
);

FILL FILL_0__7448_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .B(_2357_),
    .Y(_2358_)
);

OAI21X1 _9134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf2),
    .B(_1956_),
    .C(_1957_),
    .Y(_1958_)
);

FILL FILL_1__8091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14274_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6332_),
    .Y(_6333_)
);

FILL FILL_0__13687_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [5]),
    .Y(_5931_)
);

FILL FILL_0__13267_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5589_),
    .B(_5593_),
    .Y(_5594_)
);

FILL FILL_1__9296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10194_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6974_),
    .B(_6975_),
    .C(_6976_),
    .Y(_6780_)
);

INVX1 _14337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .Y(_6635_)
);

FILL FILL_1__7609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8160_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_595_),
    .Y(_601_)
);

FILL FILL256950x165750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .B(_170_),
    .C(_200_),
    .Y(_201_)
);

OAI21X1 _10677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3224_),
    .B(_3324_),
    .C(_2588_),
    .Y(_2581_)
);

NAND2X1 _10257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [2]),
    .B(_2672__bF$buf4),
    .Y(_2986_)
);

FILL FILL_1__12760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11333_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6436_),
    .Y(_6445_)
);

OAI21X1 _8825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(_1645_),
    .C(_1675_),
    .Y(_903_)
);

NAND2X1 _8405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1284_),
    .B(_1306_),
    .Y(_1307_)
);

FILL FILL_1__7782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12958_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf4),
    .B(_5296_),
    .C(_5297_),
    .Y(_5298_)
);

FILL FILL_0__12118_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .Y(_4943_)
);

FILL FILL_1__8987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8147_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5985_),
    .B(_5982_),
    .S(_5925__bF$buf1),
    .Y(_5986_)
);

FILL FILL_2__7851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7677_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9783_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1695_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [6])
);

FILL FILL_0__7257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_1916_),
    .Y(_2177_)
);

FILL FILL_1__11611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14083_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6150_),
    .Y(_6151_)
);

FILL FILL_0__13076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(_5804_),
    .Y(_5806_)
);

FILL FILL_2__13823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9403_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(_6808_),
    .Y(_6809_)
);

OAI21X1 _14146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6046_),
    .B(_6466_),
    .C(_6481_),
    .Y(_5878_)
);

FILL FILL_1__7838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .B(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_3203_)
);

NAND2X1 _10066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2803_),
    .Y(_2804_)
);

FILL FILL_2__10948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11142_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_973__bF$buf3),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_1523_)
);

OAI21X1 _8214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1122_),
    .C(_1123_),
    .Y(_1124_)
);

FILL FILL_1__7591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12767_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5117_),
    .B(_5116_),
    .Y(\a[7] [1])
);

FILL FILL_0__12347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4740_),
    .B(_4764_),
    .C(_4739_),
    .Y(_4765_)
);

DFFPOSX1 _9839_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.LoadCtl [2])
);

OAI21X1 _9419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2230_),
    .Y(_1694_)
);

FILL FILL_1__8796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6201_),
    .B(_6203_),
    .Y(_6204_)
);

OAI21X1 _13417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5719_),
    .B(_5807_),
    .C(_5096_),
    .Y(_5089_)
);

FILL FILL_0__14913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7486_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .B(_2380_),
    .C(_2379_),
    .Y(_2393_)
);

NAND3X1 _9172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1963_),
    .B(_1965_),
    .C(_1993_),
    .Y(_1994_)
);

FILL FILL_1__11840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [6]),
    .Y(_5968_)
);

AOI21X1 _13170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5629_),
    .B(_5628_),
    .C(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5630_)
);

OAI21X1 _7905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_810_),
    .C(_74_),
    .Y(_67_)
);

FILL FILL_2__13632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9632_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4468_),
    .Y(_4469_)
);

FILL FILL_0__9212_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7011_),
    .B(_7010_),
    .Y(_7012_)
);

NAND3X1 _14375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6667_),
    .C(_6665_),
    .Y(_6668_)
);

FILL FILL_1__7647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .B(_3020_),
    .C(_3019_),
    .Y(_3023_)
);

FILL FILL_0__11791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11371_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8863_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_861_),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.Xcalc [10])
);

OR2X2 _8443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1341_),
    .Y(_1343_)
);

INVX1 _8023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [4]),
    .Y(_943_)
);

FILL FILL_1__13583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12996_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5303_),
    .B(_5305_),
    .C(_5333_),
    .Y(_5334_)
);

FILL FILL_0__12156_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4964_),
    .B(_4977_),
    .C(_4975_),
    .Y(_4978_)
);

OAI21X1 _12021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4578_),
    .B(_4580_),
    .C(_4581_),
    .Y(_4582_)
);

FILL FILL_2__12903_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .B(_2443_),
    .Y(_2445_)
);

INVX1 _9228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .Y(_2048_)
);

FILL FILL_1__8185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14368_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6019_),
    .Y(_6021_)
);

INVX1 _13226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5679_),
    .Y(_5682_)
);

FILL FILL_0__14722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10222_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_689_)
);

FILL FILL_2__13861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11427_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(_4287_),
    .C(_4288_),
    .Y(_4289_)
);

FILL FILL_0__9021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11007_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14184_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5860_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Xin12b [10])
);

DFFPOSX1 _8919_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.Vld )
);

FILL FILL_1__7876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13219_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5387_),
    .Y(_5388_)
);

FILL FILL_2__10986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9602_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1555_),
    .C(_1552_),
    .Y(_1558_)
);

INVX1 _8252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1160_)
);

FILL FILL_1__10920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10500_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert140 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf0)
);

BUFX2 BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf4 )
);

FILL FILL_2__7105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13392_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert142 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert143 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert145 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .Y(_135__bF$buf4)
);

BUFX2 BUFX2_insert147 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .Y(_135__bF$buf3)
);

BUFX2 BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .Y(_135__bF$buf2)
);

INVX8 _12670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_5151_)
);

FILL FILL_0__12385_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert149 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .Y(_135__bF$buf1)
);

AOI21X1 _12250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4800_),
    .B(_4798_),
    .C(_4793_),
    .Y(_4801_)
);

FILL FILL_2__12712_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [9]),
    .Y(_2624_)
);

NAND3X1 _9457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(_2263_),
    .C(_2266_),
    .Y(_2267_)
);

MUX2X1 _9037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .S(gnd),
    .Y(_1866_)
);

FILL FILL_1__11705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14597_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6240_)
);

DFFPOSX1 _13455_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5055_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[6].u_ce.Acalc [5])
);

AOI21X1 _13035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5447_),
    .B(_5453_),
    .C(_5479_),
    .Y(_5501_)
);

FILL FILL_0__14111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10031_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7943_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Acalc [2])
);

NAND3X1 _7523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_506_),
    .C(_505_),
    .Y(_509_)
);

AOI22X1 _7103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Ycalc [0]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Ycalc [2]),
    .Y(_109_)
);

FILL FILL_2__13670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9670_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [7]),
    .Y(_4505_)
);

FILL FILL_0__9250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4142_),
    .B(_4143_),
    .Y(_4144_)
);

NAND2X1 _11101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3746_),
    .B(_3747_),
    .Y(_3748_)
);

NAND3X1 _8728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1572_),
    .B(_1567_),
    .C(_1609_),
    .Y(_1611_)
);

OAI21X1 _8308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1209_),
    .C(_1213_),
    .Y(_1214_)
);

FILL FILL_1__7685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13028_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .S(gnd),
    .Y(_5206_)
);

OAI21X1 _12306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4619_),
    .B(_4852_),
    .C(\genblk1[5].u_ce.Ain0 [0]),
    .Y(_4853_)
);

FILL FILL_0__13802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9411_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf4),
    .B(_1377_),
    .C(_1378_),
    .Y(_1379_)
);

INVX1 _8061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .Y(_977_)
);

FILL FILL_2__7334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12101_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2000_),
    .B(_2475_),
    .C(_2477_),
    .Y(_1714_)
);

NAND2X1 _9266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [11]),
    .B(_1834__bF$buf3),
    .Y(_2084_)
);

FILL FILL_1__11934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10507_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6057_),
    .C(_6054_),
    .Y(_6058_)
);

FILL FILL_0__13399_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5705_),
    .B(_5718_),
    .Y(_5054_)
);

FILL FILL_2__9900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9306_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14889_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6780_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.acc_reg [13])
);

OAI21X1 _14469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6561_),
    .C(_6743_),
    .Y(_6522_)
);

INVX1 _14049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6406_),
    .Y(_6407_)
);

FILL FILL_0__10680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10260_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_172__bF$buf3),
    .Y(_724_)
);

INVX1 _7332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .Y(_326_)
);

AOI21X1 _10389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3111_),
    .B(_3112_),
    .C(_2669_),
    .Y(_3113_)
);

FILL FILL_1__12892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11465_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [0]),
    .Y(_4322_)
);

FILL FILL_0__11045_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3966_),
    .C(_3954_),
    .Y(_3967_)
);

NAND2X1 _8957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [7]),
    .B(_1765_),
    .Y(_1790_)
);

NAND2X1 _8537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1429_),
    .B(_1432_),
    .Y(_1433_)
);

MUX2X1 _8117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(_1030_),
    .S(_973__bF$buf4),
    .Y(_1032_)
);

FILL FILL_1__7494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [11]),
    .B(_5174__bF$buf2),
    .Y(_5424_)
);

OAI21X1 _12535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4873_),
    .C(_4269_),
    .Y(_4262_)
);

AOI21X1 _12115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4668_),
    .B(vdd),
    .C(_4671_),
    .Y(_4672_)
);

FILL FILL_0__13611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9220_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1193_),
    .B(_1196_),
    .Y(_1197_)
);

FILL FILL_1_CLKBUF1_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(_2301_),
    .C(_2302_),
    .Y(_2303_)
);

AOI21X1 _9075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .B(_1901_),
    .C(_1836_),
    .Y(_1902_)
);

FILL FILL_1__11743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [11]),
    .B(_2672__bF$buf3),
    .Y(_3309_)
);

FILL FILL_0__10316_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13493_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5093_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain0 [0])
);

INVX1 _13073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5536_),
    .Y(_5537_)
);

NAND2X1 _7808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_776_),
    .Y(_777_)
);

FILL FILL_2__13115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9535_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4376_),
    .B(_4369_),
    .S(_4324__bF$buf4),
    .Y(_4377_)
);

FILL FILL_0__9115_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [8]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf0),
    .Y(_6923_)
);

NAND2X1 _14278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6573_),
    .B(_6582_),
    .Y(_6583_)
);

DFFPOSX1 _7981_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_65_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.Ain12b [6])
);

NAND3X1 _7561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_544_),
    .C(_485_),
    .Y(_545_)
);

INVX1 _7141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_143_)
);

NAND2X1 _10198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2927_),
    .B(_2909_),
    .Y(_2930_)
);

FILL FILL_1__12281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11601_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1640_),
    .B(_1641_),
    .C(_1642_),
    .Y(_877_)
);

NAND2X1 _8346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .B(_1249_),
    .Y(_1250_)
);

FILL FILL_2__14073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12899_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5240_),
    .B(_5241_),
    .C(_5176_),
    .Y(_5242_)
);

FILL FILL_0__12479_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_4888_)
);

FILL FILL_0__12059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8806_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_6288_),
    .C(_6329_),
    .Y(_6330_)
);

NAND2X1 _13549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [7]),
    .Y(_5928_)
);

NAND3X1 _13129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5590_),
    .C(_5565_),
    .Y(_5591_)
);

FILL FILL_0__14625_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[10]),
    .Y(Dout[10])
);

FILL FILL_2__7372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8577_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_3488_)
);

FILL FILL_2__8157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10125_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _10410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2632_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3132_),
    .D(_3130_),
    .Y(_2535_)
);

AOI21X1 _7617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(_598_),
    .C(_155_),
    .Y(_599_)
);

FILL FILL_1__12757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9344_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11615_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3355_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Ycalc [2])
);

NOR2X1 _14087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6441_),
    .B(_6442_),
    .Y(_6443_)
);

FILL FILL_1__7779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8300_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_758_),
    .Y(_760_)
);

AOI22X1 _7370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_158__bF$buf1),
    .C(_362_),
    .D(_342_),
    .Y(_9_)
);

FILL FILL_1__12090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11410_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_1821_),
    .S(_1811__bF$buf2),
    .Y(_1825_)
);

AND2X2 _8575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1468_),
    .Y(_1469_)
);

INVX1 _8155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_1067_)
);

FILL FILL_1__10823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13295_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .B(_5455_),
    .C(_5439_),
    .Y(_5041_)
);

FILL FILL_0__12288_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12573_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4227_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xin12b [10])
);

OAI21X1 _12153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4666_),
    .C(_4707_),
    .Y(_4708_)
);

FILL FILL_1__11608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8615_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6143_),
    .C(_6141_),
    .Y(_6148_)
);

NAND2X1 _13358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5109_),
    .B(_5108_),
    .Y(_5804_)
);

FILL FILL_0__14854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10354_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_89_),
    .Y(_807_)
);

NAND2X1 _7426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_395_),
    .Y(_416_)
);

FILL FILL_2__13153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11559_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4397_),
    .B(_4412_),
    .Y(_4413_)
);

FILL FILL_0__9153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11139_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3516_),
    .B(_4053_),
    .C(_4052_),
    .Y(_4054_)
);

NAND2X1 _11004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3653_),
    .B(_3654_),
    .Y(_3655_)
);

FILL FILL_0__12920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7168_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5113_),
    .C(_5114_),
    .Y(_5115_)
);

NOR2X1 _12209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4757_),
    .B(_4761_),
    .Y(_4762_)
);

FILL FILL_1__14712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9314_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1071_),
    .C(_1285_),
    .Y(_1286_)
);

FILL FILL_1__10632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10212_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [6]),
    .B(_4348__bF$buf3),
    .Y(_4923_)
);

FILL FILL_0__12097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2389_),
    .B(_2386_),
    .Y(_2390_)
);

INVX1 _9169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [7]),
    .Y(_1991_)
);

FILL FILL_1__11837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_5965_)
);

AOI21X1 _13167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5626_),
    .B(_5624_),
    .C(_5619_),
    .Y(_5627_)
);

FILL FILL_0__14663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10910_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .Y(_634_)
);

INVX1 _7235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_233_)
);

FILL FILL_2__13382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11368_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11653_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3393_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xin12b [6])
);

NAND3X1 _11233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3834_),
    .B(_3795_),
    .C(_3812_),
    .Y(_3874_)
);

FILL FILL_1__7397_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9801_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1713_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin12b [10])
);

INVX1 _12858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [7]),
    .Y(_5331_)
);

OAI21X1 _12438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4971_),
    .B(_4956_),
    .C(_4970_),
    .Y(_4975_)
);

NAND3X1 _12018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4565_),
    .B(_4577_),
    .C(_4561_),
    .Y(_4579_)
);

FILL FILL_1__14101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9123_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1081_),
    .B(_1072_),
    .Y(_1104_)
);

FILL FILL_1__10861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4725_),
    .B(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .C(_4744_),
    .Y(_4208_)
);

AOI22X1 _9398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1797_),
    .B(_1834__bF$buf3),
    .C(_2210_),
    .D(_1832_),
    .Y(_1693_)
);

FILL FILL_1__11226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8653_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3512_),
    .Y(_3579_)
);

FILL FILL_0__8233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10639_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3217_),
    .B(_3219_),
    .Y(_3220_)
);

FILL FILL_0__10219_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5825_)
);

FILL FILL_2__9612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9438_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4284_),
    .C(_4285_),
    .Y(_4286_)
);

FILL FILL_0__9018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8814_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_828_)
);

NAND2X1 _7464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf4),
    .B(_451_),
    .Y(_452_)
);

FILL FILL_2__13191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11597_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf1),
    .B(_4398_),
    .Y(_4449_)
);

FILL FILL_0__9191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11177_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4088_),
    .Y(_4089_)
);

OAI21X1 _11042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .B(_3691_),
    .C(_3579_),
    .Y(_3692_)
);

FILL FILL_2__11924_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1554_),
    .Y(_1556_)
);

AOI21X1 _8249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1147_),
    .B(_1125_),
    .C(_1126_),
    .Y(_1157_)
);

FILL FILL_1__10917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [6]),
    .B(_1834__bF$buf1),
    .Y(_2409_)
);

FILL FILL_1__13389_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [0]),
    .Y(_5148_)
);

NAND3X1 _12247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf2),
    .B(_4797_),
    .C(_4794_),
    .Y(_4798_)
);

FILL FILL_1__14750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10250_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7025_),
    .B(_7028_),
    .Y(_7029_)
);

FILL FILL_0__14108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8042_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10733_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2559_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Xin1 [0])
);

FILL FILL_0__10448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10028_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3039_),
    .C(_3035_),
    .Y(_3040_)
);

FILL FILL_0__14281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9667_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4502_),
    .B(_4498_),
    .C(_4350_),
    .Y(_4503_)
);

FILL FILL_0__9247_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .Y(_4141_)
);

FILL FILL_1__13601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8203_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [1]),
    .B(_158__bF$buf4),
    .Y(_669_)
);

FILL FILL_1__14806_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_263_),
    .Y(_270_)
);

DFFPOSX1 _11691_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.Vld )
);

NAND2X1 _11271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3909_),
    .Y(_3910_)
);

FILL FILL_1__9408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8898_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_896_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Yin1 [1])
);

NOR2X1 _8478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf0),
    .B(_1249_),
    .Y(_1376_)
);

FILL FILL_0_CLKBUF1_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_974_)
);

FILL FILL_0_CLKBUF1_insert98 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert99 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5343_),
    .B(_5339_),
    .Y(_5368_)
);

OAI21X1 _12476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_5003_)
);

NAND2X1 _12056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4615_)
);

FILL FILL_2__12938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833__bF$buf4),
    .B(_6852_),
    .Y(_6853_)
);

DFFPOSX1 _14202_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5878_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[7].u_ce.Yin12b [4])
);

FILL FILL_2__7084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8691_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3614_),
    .Y(_3615_)
);

FILL FILL_0__8271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10677_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3254_),
    .Y(_3255_)
);

FILL FILL_0__10257_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2829_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_2857_),
    .Y(_2522_)
);

INVX1 _7749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [5]),
    .Y(_721_)
);

NAND3X1 _7329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_301_),
    .C(_284_),
    .Y(_323_)
);

FILL FILL257550x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9476_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4317_),
    .B(_4318_),
    .C(_4319_),
    .Y(_4320_)
);

FILL FILL_0__9056_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3958_),
    .C(_3956_),
    .Y(_3964_)
);

FILL FILL_1__13830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14615_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.Acalc [4]),
    .C(_89_),
    .D(\genblk1[0].u_ce.Acalc [6]),
    .Y(_90_)
);

FILL FILL_0__13608_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3723_),
    .C(_3727_),
    .Y(_3728_)
);

FILL FILL_1__9637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11122_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1191_),
    .C(_1187_),
    .Y(_1194_)
);

FILL FILL_1__10955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7122_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4832_),
    .B(_4830_),
    .Y(_4834_)
);

FILL FILL_2__8921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9390_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6811_),
    .B(_6833__bF$buf4),
    .C(_7061_),
    .Y(_6789_)
);

FILL FILL_0__14566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14146_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6716_),
    .C(_6713_),
    .Y(_6717_)
);

NAND2X1 _14011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Vld ),
    .B(_6370_),
    .Y(_6371_)
);

FILL FILL_1__7703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11073_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3434_),
    .Y(_3435_)
);

FILL FILL_2__8098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10066_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3073_),
    .Y(_3076_)
);

DFFPOSX1 _7978_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_62_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Ain12b [11])
);

INVX1 _7558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .Y(_542_)
);

NAND2X1 _7138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_140_)
);

FILL FILL_1__12698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12278_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4513_),
    .B(_4517_),
    .Y(_4539_)
);

FILL FILL_0__9285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.X_ [0]),
    .Y(_4167_)
);

NOR2X1 _11136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3516_),
    .Y(_3781_)
);

FILL FILL_0__12632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_2489_)
);

FILL FILL_1__8661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13837_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6034_),
    .B(_6053_),
    .C(_6025_),
    .Y(_6075_)
);

FILL FILL_0__13417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11351_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1011_)
);

FILL FILL_1__10344_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14907_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6798_),
    .CLK(clk_bF$buf72),
    .Q(\genblk1[0].u_ce.ISin )
);

FILL FILL_2__7789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7351_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4647_),
    .B(_4644_),
    .S(_4325__bF$buf2),
    .Y(_4652_)
);

FILL FILL_2__8310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8556_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .Y(_3485_)
);

FILL FILL_0__8136_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3129_),
    .Y(_3130_)
);

FILL FILL_1__12910_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5750_),
    .B(_5751_),
    .Y(_5752_)
);

FILL FILL_2__9935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14375_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6872_),
    .B(_6879_),
    .Y(_6887_)
);

INVX1 _14240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [8]),
    .Y(_6553_)
);

FILL FILL_1__7512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .B(_3290_),
    .Y(_3291_)
);

FILL FILL_0__10295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .B(_2893_),
    .C(_2892_),
    .Y(_2894_)
);

FILL FILL_1__8717_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_756_),
    .Y(_757_)
);

INVX1 _7367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .Y(_360_)
);

FILL FILL_1__12087_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4355_),
    .B(_4334_),
    .C(_4325__bF$buf3),
    .Y(_4356_)
);

FILL FILL_0__9094_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3999_),
    .B(_3998_),
    .C(_3608_),
    .Y(_4000_)
);

FILL FILL_0__12861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7827_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .B(\genblk1[3].u_ce.Xin12b [4]),
    .S(vdd),
    .Y(_2676_)
);

FILL FILL_0__7407_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2316_),
    .Y(_2320_)
);

FILL FILL_1__8470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert130 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert131 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert133 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6290_),
    .B(_6293_),
    .Y(_6294_)
);

FILL FILL_0_BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert135 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(\genblk1[7].u_ce.Ycalc [8]),
    .C(_5889_),
    .Y(_5894_)
);

FILL FILL_0_BUFX2_insert136 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert138 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10153_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6939_)
);

FILL FILL_2__7598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3313_),
    .Y(_3331_)
);

OAI21X1 _10216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2809_),
    .C(_2946_),
    .Y(_2947_)
);

FILL FILL_0__11712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8106_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_572_),
    .C(_227_),
    .Y(_579_)
);

FILL FILL_1__14709_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_177_)
);

OAI21X1 _11594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Ain12b [9]),
    .Y(_4188_)
);

INVX1 _11174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3817_),
    .Y(_3818_)
);

FILL FILL_2__7810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7636_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [0]),
    .Y(_2509_)
);

FILL FILL_0__7216_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_2130_),
    .S(_1811__bF$buf3),
    .Y(_2138_)
);

NAND2X1 _12799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf2),
    .B(_5224_),
    .Y(_5275_)
);

NAND2X1 _12379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4919_),
    .B(_4910_),
    .Y(_4921_)
);

FILL FILL_1__14462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13875_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6109_),
    .C(_6110_),
    .Y(_6111_)
);

FILL FILL_0__13035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5771_),
    .B(_5770_),
    .Y(_5772_)
);

FILL FILL_1__9484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10382_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14525_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6513_),
    .CLK(clk_bF$buf47),
    .Q(\u_ot.Xin12b [11])
);

OAI21X1 _14105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6115_),
    .B(_6455_),
    .C(_6457_),
    .Y(_5861_)
);

FILL FILL_2__12174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8594_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _10865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3518_),
    .B(_3521_),
    .C(_3486__bF$buf3),
    .D(_3515_),
    .Y(_3522_)
);

FILL FILL_0__8174_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3164_),
    .B(_3165_),
    .Y(_3166_)
);

NAND2X1 _10025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2762_),
    .B(_2764_),
    .Y(_2765_)
);

FILL FILL_0__11941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7865_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2713_),
    .Y(_2714_)
);

FILL FILL_0__7445_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2354_),
    .B(_2353_),
    .Y(_2355_)
);

INVX1 _9131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .Y(_1955_)
);

NOR2X1 _12188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4741_),
    .B(_4726_),
    .Y(_4742_)
);

FILL FILL_1__14691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14469_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6970_),
    .B(_6973_),
    .Y(_6974_)
);

FILL FILL_0__14049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [11]),
    .B(_6562__bF$buf3),
    .Y(_6632_)
);

FILL FILL_1__7606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .B(_3321_),
    .Y(_2587_)
);

FILL FILL_0__10389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2982_),
    .B(_2960_),
    .Y(_2984_)
);

FILL FILL_0__11750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Ain12b [9]),
    .Y(_1674_)
);

INVX1 _8402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1303_),
    .Y(_1304_)
);

INVX1 _11879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4446_)
);

FILL FILL_0__9188_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4068_),
    .Y(_4086_)
);

INVX1 _11039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .Y(_3689_)
);

FILL FILL_1__13962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12955_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5294_),
    .Y(_5295_)
);

FILL FILL_0__12535_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4938_),
    .B(_4940_),
    .C(_4923_),
    .Y(_4221_)
);

FILL FILL_0__12115_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2396_),
    .Y(_2407_)
);

FILL FILL_1__8984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .B(\genblk1[7].u_ce.Xin1 [1]),
    .S(vdd),
    .Y(_5983_)
);

FILL FILL_1__9349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7254_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9780_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1692_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [3])
);

MUX2X1 _9360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2130_),
    .S(vdd),
    .Y(_2174_)
);

FILL FILL_0__10601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14278_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6803_),
    .B(_6804_),
    .C(_6805_),
    .Y(_6806_)
);

NAND2X1 _14143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .B(_6463_),
    .Y(_6480_)
);

FILL FILL_1__7835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14605_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .C(gnd),
    .Y(_3200_)
);

FILL FILL_0__10198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2790_),
    .B(_2797_),
    .C(_2800_),
    .Y(_2801_)
);

FILL FILL_2__9591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10525_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1520_),
    .C(_1507_),
    .Y(_864_)
);

NAND3X1 _8211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf2),
    .B(_1120_),
    .C(_1115_),
    .Y(_1121_)
);

DFFPOSX1 _11688_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.LoadCtl [3])
);

INVX1 _11268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [6]),
    .Y(_3907_)
);

FILL FILL_1__13771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12344_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9836_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1748_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[2].u_ce.Ain0 [1])
);

NOR2X1 _9416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2212_),
    .Y(_2228_)
);

FILL FILL_1__8793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13549_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [11]),
    .B(_6115_),
    .Y(_6201_)
);

FILL FILL_0__13129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [7]),
    .B(_5804_),
    .Y(_5095_)
);

FILL FILL_0__14910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10056_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6850_)
);

FILL FILL_0__7483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12688_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .B(_807_),
    .Y(_73_)
);

FILL FILL_0__8688_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf2),
    .B(_3610_),
    .C(_3611_),
    .Y(_3612_)
);

FILL FILL_0__8268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3249_),
    .B(_3231_),
    .C(_3251_),
    .Y(_3252_)
);

OAI21X1 _10119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf0),
    .B(_2741_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_2855_)
);

FILL FILL_1__12622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12202_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4466_)
);

OAI21X1 _14792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6916_),
    .B(_7001_),
    .C(_7008_),
    .Y(_7009_)
);

FILL FILL_0__14087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6664_),
    .B(_6661_),
    .Y(_6665_)
);

FILL FILL_1__7644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13407_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3013_),
    .B(_3016_),
    .C(_3018_),
    .Y(_3020_)
);

FILL FILL_1__8429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10334_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_485_),
    .C(_482_),
    .Y(_486_)
);

OAI21X1 _7079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(\genblk1[0].u_ce.Acalc [8]),
    .C(_86_),
    .Y(_87_)
);

DFFPOSX1 _8860_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_858_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[1].u_ce.Xcalc [7])
);

NAND2X1 _8440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(_1339_),
    .Y(_1340_)
);

INVX1 _8020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [10]),
    .Y(_940_)
);

OAI21X1 _11497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4112_),
    .C(_4110_),
    .Y(_4122_)
);

OAI21X1 _11077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3632_),
    .C(_3678_),
    .Y(_3725_)
);

FILL FILL_2__7713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7539_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [8]),
    .B(_2377_),
    .C(_2441_),
    .Y(_2442_)
);

FILL FILL_0__7119_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2043_),
    .B(_2031_),
    .C(_2044_),
    .Y(_2045_)
);

FILL FILL_1__8182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13358_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6018_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_6019_)
);

OAI21X1 _13223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5445_),
    .B(_5678_),
    .C(\genblk1[6].u_ce.Ain0 [0]),
    .Y(_5679_)
);

FILL FILL_1__9387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10285_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [9]),
    .B(_6833__bF$buf4),
    .C(En_bF$buf4),
    .Y(_7060_)
);

OAI21X1 _14428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .C(\u_ot.ISreg_bF$buf3 ),
    .Y(_6714_)
);

OAI21X1 _14008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6305_),
    .B(_6366_),
    .C(_6367_),
    .Y(_6368_)
);

FILL FILL_0__7292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(gnd),
    .Y(_686_)
);

FILL FILL_0__8497_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [2]),
    .Y(_3432_)
);

FILL FILL_0__8077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2992_),
    .C(_3072_),
    .Y(_3073_)
);

FILL FILL_1__12851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11004_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14181_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5857_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [9])
);

DFFPOSX1 _8916_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.LoadCtl [3])
);

FILL FILL_1__7873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13216_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5383_),
    .B(_5371_),
    .C(_5384_),
    .Y(_5385_)
);

FILL FILL_0__12629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10563_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562_),
    .Y(_6562__bF$buf2)
);

FILL FILL_2__7522_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert111 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562_),
    .Y(_6562__bF$buf1)
);

BUFX2 BUFX2_insert112 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562_),
    .Y(_6562__bF$buf0)
);

BUFX2 BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert114 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert116 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf3)
);

BUFX2 BUFX2_insert118 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf2)
);

FILL FILL_0__12382_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert119 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf1)
);

FILL FILL_0__7768_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2618_),
    .B(_2621_),
    .C(_2606_),
    .Y(_2622_)
);

FILL FILL_0__7348_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .Y(_2264_)
);

MUX2X1 _9034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .B(_1855_),
    .S(_1810__bF$buf0),
    .Y(_1863_)
);

FILL FILL_1__11702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14594_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5937_),
    .B(_6234_),
    .Y(_6237_)
);

FILL FILL_0__13587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13167_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13452_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5052_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [11])
);

AOI21X1 _13032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .B(vdd),
    .C(_5497_),
    .Y(_5498_)
);

FILL FILL_1__9196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10094_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6868_),
    .Y(_6884_)
);

INVX1 _14237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [7]),
    .Y(_6551_)
);

FILL FILL_1__7509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8060_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7940_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [11])
);

OAI21X1 _7520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_502_),
    .C(_504_),
    .Y(_506_)
);

FILL FILL_1__11299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [6]),
    .B(_89_),
    .Y(_106_)
);

NAND3X1 _10997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3615_),
    .B(_3637_),
    .C(_3618_),
    .Y(_3648_)
);

OAI21X1 _10577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3287_),
    .B(_3231_),
    .C(_3286_),
    .Y(_3288_)
);

NAND3X1 _10157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_2890_),
    .C(_2888_),
    .Y(_2891_)
);

FILL FILL_1__12660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11233_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1598_),
    .C(_1596_),
    .Y(_1608_)
);

OAI21X1 _8305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1118_),
    .C(_1164_),
    .Y(_1211_)
);

FILL FILL_1__7682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12858_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5202_),
    .B(_5195_),
    .S(_5150__bF$buf0),
    .Y(_5203_)
);

FILL FILL_0__12438_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4849_),
    .B(_4845_),
    .C(_4346_),
    .Y(_4851_)
);

FILL FILL_0__12018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10372_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(_6239_),
    .Y(_6291_)
);

AND2X2 _13508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(\genblk1[7].u_ce.LoadCtl [3]),
    .Y(_5891_)
);

FILL FILL_2__7751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7157_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2475_),
    .Y(_2476_)
);

OAI21X1 _9263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2079_),
    .B(_2081_),
    .C(_1903_),
    .Y(_2082_)
);

FILL FILL_1__11931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10504_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6034_),
    .B(_6025_),
    .C(_5963__bF$buf4),
    .Y(_6055_)
);

FILL FILL_0__13396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5713_),
    .B(_5715_),
    .Y(_5716_)
);

FILL FILL_2__13723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9303_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14886_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6777_),
    .CLK(clk_bF$buf50),
    .Q(\u_pa.acc_reg [10])
);

OAI21X1 _14466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Xin1 [1]),
    .Y(_6742_)
);

NAND2X1 _14046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6398_),
    .B(_6400_),
    .Y(_6404_)
);

FILL FILL_1__7738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7318_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3096_),
    .B(_3086_),
    .C(_3109_),
    .Y(_3110_)
);

FILL FILL_2__10848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11042_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Ycalc [11]),
    .C(_1762_),
    .Y(_1787_)
);

NAND3X1 _8534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf1),
    .B(_1426_),
    .C(_1421_),
    .Y(_1430_)
);

MUX2X1 _8114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1028_),
    .B(_1027_),
    .S(_973__bF$buf1),
    .Y(_1029_)
);

FILL FILL_1__7491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13254_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5419_),
    .B(_5421_),
    .C(_5243_),
    .Y(_5422_)
);

FILL FILL_0__12667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12247_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[5] [0]),
    .Y(_4268_)
);

NAND2X1 _12112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4431_),
    .B(_4616_),
    .Y(_4669_)
);

OAI21X1 _9739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .B(_2475_),
    .C(_2507_),
    .Y(_1737_)
);

OAI21X1 _9319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf1),
    .B(_2131_),
    .C(_2134_),
    .Y(_2135_)
);

FILL FILL_1__8696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14039_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6059_),
    .B(_6062_),
    .Y(_6108_)
);

NAND3X1 _13317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [8]),
    .B(_5711_),
    .C(_5768_),
    .Y(_5769_)
);

FILL FILL_1_CLKBUF1_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7386_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2282_),
    .B(_2280_),
    .C(_1848__bF$buf0),
    .Y(_2300_)
);

NOR2X1 _9072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1883_),
    .B(_1898_),
    .Y(_1899_)
);

FILL FILL_1__11740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13490_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5090_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain12b [5])
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5492_),
    .C(_5533_),
    .Y(_5534_)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_717_),
    .C(_772_),
    .Y(_774_)
);

FILL FILL_2__13532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4374_)
);

FILL FILL_0__9112_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6916_),
    .B(_6919_),
    .Y(_6920_)
);

NAND2X1 _14275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [3]),
    .B(_6562__bF$buf4),
    .Y(_6581_)
);

FILL FILL_1__7547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7127_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2924_),
    .B(_2926_),
    .Y(_2927_)
);

FILL FILL_2__10237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11271_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [0]),
    .Y(_1640_)
);

INVX1 _8343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1235_),
    .Y(_1247_)
);

FILL FILL_2__14490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12896_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5223_),
    .B(_5238_),
    .Y(_5239_)
);

FILL FILL_0__12476_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [3]),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4885_)
);

FILL FILL_0__12056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12803_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2710_),
    .B(_2702_),
    .C(_2685_),
    .Y(_2711_)
);

OR2X2 _9548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2349_),
    .Y(_2352_)
);

INVX1 _9128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_1952_)
);

FILL FILL_1__8085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6305_),
    .C(_6318_),
    .Y(_6327_)
);

INVX4 _13546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_5925_)
);

NOR2X1 _13126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5583_),
    .B(_5587_),
    .Y(_5588_)
);

FILL FILL_0__14622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10122_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_572_),
    .C(_595_),
    .Y(_596_)
);

FILL FILL_2__13761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11327_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11612_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3352_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Ycalc [0])
);

NAND2X1 _14084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6439_),
    .B(_6436_),
    .Y(_6440_)
);

OAI21X1 _8819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Ain12b [8]),
    .Y(_1672_)
);

FILL FILL_1__7776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13119_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5292_)
);

FILL FILL_2__10886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9502_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .Y(_1822_)
);

NAND2X1 _8572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1463_),
    .B(_1464_),
    .Y(_1466_)
);

INVX2 _8152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .Y(_1065_)
);

FILL FILL_1__10820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13292_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .B(_5457_),
    .Y(_5458_)
);

DFFPOSX1 _12570_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4224_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [9])
);

FILL FILL_0__12285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4705_)
);

DFFPOSX1 _9777_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1689_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Xcalc [0])
);

INVX1 _9357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .Y(_2171_)
);

FILL FILL_1__11605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6143_),
    .C(_6144_),
    .Y(_6145_)
);

INVX1 _13355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [1]),
    .Y(_5802_)
);

FILL FILL_0__14851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10351_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_805_)
);

NAND2X1 _7423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_412_),
    .Y(_413_)
);

FILL FILL_2__13570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .B(_4405_),
    .C(_4408_),
    .Y(_4410_)
);

FILL FILL_0__9150_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3487__bF$buf4),
    .Y(_4051_)
);

FILL FILL_0__11136_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3651_),
    .C(_3648_),
    .Y(_3652_)
);

NOR2X1 _8628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1508_),
    .B(_1517_),
    .Y(_1518_)
);

AOI21X1 _8208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1075_),
    .B(_973__bF$buf0),
    .C(_1117_),
    .Y(_1118_)
);

FILL FILL_1__7585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13348_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5110_),
    .C(_5111_),
    .Y(_5112_)
);

NOR2X1 _12206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4758_),
    .B(_4738_),
    .Y(_4759_)
);

FILL FILL_0__13702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9311_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [1]),
    .B(_996__bF$buf1),
    .Y(_1283_)
);

FILL FILL_2__7234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12841_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(gnd),
    .C(_1848__bF$buf3),
    .Y(_2387_)
);

AOI21X1 _9166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(_1984_),
    .C(_1836_),
    .Y(_1989_)
);

FILL FILL_1__11834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10407_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin0 [1]),
    .Y(_5962_)
);

FILL FILL_0__13299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf2),
    .B(_5623_),
    .C(_5620_),
    .Y(_5624_)
);

FILL FILL_0__14660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9206_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6995_),
    .B(_6981_),
    .C(_6990_),
    .Y(_7006_)
);

NOR2X1 _14369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin1 [0]),
    .B(\u_ot.Yin1 [1]),
    .Y(_6662_)
);

FILL FILL_0__10580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10160_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf5)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf4)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf3)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf2)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf1)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .Y(_1010__bF$buf0)
);

OAI21X1 _7652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_621_),
    .C(_156_),
    .Y(_632_)
);

INVX2 _7232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .Y(_230_)
);

OR2X2 _10289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3013_),
    .B(_3016_),
    .Y(_3017_)
);

FILL FILL_1__12792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11785_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11650_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3390_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [11])
);

FILL FILL_0__11365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3870_),
    .Y(_3871_)
);

DFFPOSX1 _8857_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_855_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Xcalc [4])
);

NOR2X1 _8437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf0),
    .B(_1336_),
    .Y(_1337_)
);

OAI21X1 _8017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_937_),
    .C(_930_),
    .Y(_938_)
);

FILL FILL_1__7394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13157_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5328_),
    .B(_5324_),
    .C(_5176_),
    .Y(_5329_)
);

OAI21X1 _12435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4971_),
    .B(_4968_),
    .C(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4973_)
);

OAI21X1 _12015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4487_),
    .C(_4516_),
    .Y(_4576_)
);

FILL FILL_0__13931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9120_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _8190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .Y(_1101_)
);

FILL FILL_0__14716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7289_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2207_),
    .Y(_2208_)
);

FILL FILL_1__11223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8650_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3575_),
    .Y(_3576_)
);

FILL FILL_2__8248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10636_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3212_),
    .B(_3216_),
    .Y(_3217_)
);

FILL FILL_0__10216_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5292_),
    .B(_5807_),
    .C(_5823_),
    .Y(_5078_)
);

INVX1 _7708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_683_)
);

FILL FILL_2__13015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9435_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4270_),
    .B(_4273_),
    .C(_4283_),
    .Y(\a[6] [0])
);

FILL FILL_0__9015_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(_6834_),
    .Y(_6763_)
);

DFFPOSX1 _14178_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5854_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [6])
);

FILL FILL_1__8811_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_810_),
    .C(_826_),
    .Y(_56_)
);

NAND2X1 _7461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_449_)
);

OAI21X1 _10098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2832_),
    .C(_2833_),
    .Y(_2834_)
);

FILL FILL_1__12181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11501_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1548_),
    .B(_1551_),
    .Y(_1553_)
);

AOI21X1 _8246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1138_),
    .C(_1133_),
    .Y(_1154_)
);

FILL FILL_1__10914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12799_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5143_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5146_)
);

FILL FILL_0__12379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4708_),
    .Y(_4795_)
);

FILL FILL_0__13740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8706_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5937_),
    .B(_6234_),
    .C(_5947_),
    .Y(_6235_)
);

DFFPOSX1 _13449_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5049_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [8])
);

NAND2X1 _13029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5257_),
    .B(_5442_),
    .Y(_5495_)
);

AND2X2 _14810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_7026_)
);

FILL FILL_0__14105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8057_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10730_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2556_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xin12b [7])
);

FILL FILL_0__10445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10025_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3017_),
    .B(_3036_),
    .C(_2686__bF$buf3),
    .Y(_3037_)
);

DFFPOSX1 _7937_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [8])
);

OR2X2 _7517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_502_),
    .Y(_503_)
);

FILL FILL_1__12657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9664_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4499_),
    .B(_4478_),
    .Y(_4500_)
);

FILL FILL_0__9244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4131_),
    .B(_4132_),
    .C(_4121_),
    .Y(_4138_)
);

FILL FILL_1__7679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_666_),
    .Y(_667_)
);

FILL FILL_1__14803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_266_),
    .C(_263_),
    .Y(_267_)
);

FILL FILL_1__9405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8895_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_893_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[1].u_ce.Yin12b [4])
);

FILL FILL_0_CLKBUF1_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [5]),
    .Y(_1373_)
);

INVX1 _8055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .Y(_971_)
);

FILL FILL_0_CLKBUF1_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13195_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5339_),
    .B(_5343_),
    .Y(_5365_)
);

OAI21X1 _12473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4329_),
    .B(_5000_),
    .C(_5001_),
    .Y(_4233_)
);

FILL FILL_0__12188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4598_),
    .B(_4612_),
    .Y(_4202_)
);

FILL FILL_2__12515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8515_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf0),
    .B(_5954_),
    .Y(_6052_)
);

NOR2X1 _13258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5708_),
    .B(_5712_),
    .Y(_5713_)
);

FILL FILL_0__14754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10254_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_717_),
    .C(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .Y(_719_)
);

OAI21X1 _7326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_318_),
    .C(_319_),
    .Y(_320_)
);

FILL FILL_2__13053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Xcalc [11]),
    .Y(_4317_)
);

FILL FILL_0__9053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .B(_3935_),
    .C(_3524__bF$buf1),
    .Y(_3961_)
);

FILL FILL_0__12820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7488_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5413_),
    .B(_5409_),
    .Y(_5419_)
);

OAI21X1 _12529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5023_),
    .B(_4273_),
    .C(_4266_),
    .Y(_4259_)
);

OAI21X1 _12109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .C(_4665_),
    .Y(_4666_)
);

FILL FILL_1__14612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9214_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1188_),
    .Y(_1191_)
);

FILL FILL_1__10952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10112_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4794_),
    .B(_4796_),
    .Y(_4831_)
);

NOR2X1 _9489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2296_),
    .Y(_2297_)
);

NAND3X1 _9069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .B(_1891_),
    .C(_1894_),
    .Y(_1896_)
);

FILL FILL_1__11737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8324_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13487_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5087_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Ain12b [6])
);

NAND2X1 _13067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5531_)
);

FILL FILL_2__9703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10810_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7975_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_59_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin0 [0])
);

AOI21X1 _7555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf2),
    .B(_497_),
    .C(_538_),
    .Y(_539_)
);

NAND2X1 _7135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_137_)
);

FILL FILL_2__13282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12275_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4498_),
    .B(_4526_),
    .Y(_4536_)
);

FILL FILL_0__9282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4154_),
    .B(_3435_),
    .C(_4165_),
    .Y(_3397_)
);

FILL FILL_0__11268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3776_),
    .C(_3777_),
    .Y(_3778_)
);

FILL FILL_1__7297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14487_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_2486_),
    .C(_2487_),
    .Y(_1719_)
);

NAND3X1 _12758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .B(_5231_),
    .C(_5234_),
    .Y(_5236_)
);

NAND2X1 _12338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4881_),
    .B(_4874_),
    .Y(_4883_)
);

FILL FILL257250x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9023_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _8093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1004_),
    .B(_1007_),
    .C(_972__bF$buf1),
    .D(_1001_),
    .Y(_1008_)
);

FILL FILL_1__10341_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14904_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6795_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [8])
);

FILL FILL_0__14619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4645_),
    .C(_4648_),
    .Y(_4649_)
);

NOR2X1 _9298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .B(_2114_),
    .Y(_2115_)
);

FILL FILL_1__11966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8553_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.Xcalc [1]),
    .C(_3482_),
    .D(_3444_),
    .Y(_3483_)
);

FILL FILL_0__8133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3121_),
    .B(_3123_),
    .Y(_3127_)
);

NAND2X1 _13296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5748_),
    .B(_5747_),
    .Y(_5749_)
);

FILL FILL_0__11900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9338_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4016_),
    .C(_3430_),
    .Y(_3423_)
);

FILL FILL_0__10292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8714_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf5),
    .B(_671_),
    .Y(_754_)
);

OAI21X1 _7364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_352_),
    .C(_350_),
    .Y(_357_)
);

FILL FILL_2__13091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11497_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4352_),
    .B(_4351_),
    .S(_4325__bF$buf4),
    .Y(_4353_)
);

FILL FILL_0__9091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11077_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [10]),
    .B(_3995_),
    .C(_3996_),
    .Y(_3997_)
);

FILL FILL_1__9919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1819_)
);

NAND2X1 _8569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1461_),
    .B(_1462_),
    .Y(_1463_)
);

INVX1 _8149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1061_),
    .Y(_1062_)
);

FILL FILL_1__10817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7824_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [1]),
    .B(_2672__bF$buf4),
    .Y(_2673_)
);

FILL FILL_0__7404_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2280_),
    .B(_2282_),
    .Y(_2317_)
);

FILL FILL_1__13289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .B(_5454_),
    .Y(_5455_)
);

DFFPOSX1 _12567_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4221_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [6])
);

NAND2X1 _12147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4702_),
    .B(_4701_),
    .Y(_4703_)
);

FILL FILL_1__14650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14428_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6935_),
    .Y(_6936_)
);

FILL FILL_0__14008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8362_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2660_),
    .C(_3329_),
    .Y(_2561_)
);

FILL FILL_0__10348_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .B(_2942_),
    .C(_2943_),
    .D(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2944_)
);

FILL FILL_2__9741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9567_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4340_),
    .B(_4377_),
    .C(_4362__bF$buf5),
    .Y(_4407_)
);

FILL FILL_0__9147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4040_),
    .B(_4045_),
    .Y(_4048_)
);

FILL FILL_1__13921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8103_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .B(_550_),
    .C(_548_),
    .Y(_576_)
);

FILL FILL_1__14706_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_174_)
);

OAI21X1 _11591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Ain12b [8]),
    .Y(_4186_)
);

MUX2X1 _11171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3814_),
    .B(_3803_),
    .S(vdd),
    .Y(_3815_)
);

FILL FILL_1__9728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .B(_1645_),
    .Y(_1661_)
);

OAI21X1 _8378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf0),
    .B(_1280_),
    .C(_1269_),
    .Y(_1281_)
);

FILL FILL_1__10626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13098_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5272_)
);

NAND2X1 _12376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4917_),
    .B(_4916_),
    .Y(_4918_)
);

FILL FILL_2__12838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14657_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14522_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6510_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Ycalc [10])
);

FILL FILL_0__14237_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [0]),
    .B(_6455_),
    .Y(_6456_)
);

FILL FILL_1__11584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8591_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .B(_3516_),
    .C(_3487__bF$buf4),
    .Y(_3519_)
);

FILL FILL_0__8171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10157_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3162_),
    .B(_3159_),
    .Y(_3163_)
);

NAND3X1 _10022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2747_),
    .B(_2758_),
    .C(_2761_),
    .Y(_2762_)
);

FILL FILL_2__9550_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_628_),
    .Y(_629_)
);

OAI21X1 _7229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_227_),
    .C(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Y(_228_)
);

FILL FILL_2__13796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9376_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11647_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3387_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [10])
);

OAI21X1 _11227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3737_),
    .C(_3867_),
    .Y(_3868_)
);

FILL FILL_1__13730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11022_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf0),
    .B(_1096_),
    .C(_1097_),
    .Y(_1098_)
);

FILL FILL_1__10855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7442_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4738_),
    .Y(_4739_)
);

FILL FILL_0__13681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8647_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3572_),
    .Y(_3573_)
);

FILL FILL_0__8227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14466_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6971_)
);

FILL FILL_0__14046_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6628_),
    .B(_6629_),
    .Y(_6630_)
);

FILL FILL_1__7603_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert384 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert385 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert386 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert387 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert388 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert389 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

FILL FILL_1__11393_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3349_),
    .B(_3317_),
    .C(_3350_),
    .Y(_2578_)
);

FILL FILL_0__10386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2697_),
    .B(_2978_),
    .C(_2975_),
    .Y(_2981_)
);

FILL FILL_1__8808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_810_),
    .Y(_825_)
);

NOR2X1 _7458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_443_),
    .Y(_446_)
);

FILL FILL_1__12178_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4419_),
    .B(_4348__bF$buf4),
    .C(_4443_),
    .D(_4420_),
    .Y(_4194_)
);

FILL FILL_0__9185_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(_4083_),
    .Y(_4084_)
);

NAND2X1 _11036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .B(_3682_),
    .Y(_3686_)
);

FILL FILL_0__12952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x97350 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .B(_2402_),
    .Y(_2404_)
);

FILL FILL_1__8981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13737_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [8]),
    .B(\genblk1[7].u_ce.Xin12b [7]),
    .S(vdd),
    .Y(_5980_)
);

FILL FILL_0__13317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10244_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [16]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf2),
    .Y(_7024_)
);

FILL FILL_2__7689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8036_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10727_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2553_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xin12b [8])
);

OAI21X1 _10307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2950_),
    .C(_3033_),
    .Y(_3034_)
);

FILL FILL_1__12810_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5620_),
    .B(_5622_),
    .Y(_5657_)
);

FILL FILL_0__11803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14275_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [8]),
    .Y(_6803_)
);

OAI21X1 _14140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6477_),
    .B(_6459_),
    .C(_6478_),
    .Y(_5875_)
);

FILL FILL_1__7832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7412_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3197_)
);

FILL FILL_0__10195_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _10060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2776_),
    .C(_2748_),
    .Y(_2798_)
);

FILL FILL_1__8617_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain0 [0]),
    .Y(_664_)
);

OAI21X1 _7267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_234_),
    .C(_172__bF$buf2),
    .Y(_264_)
);

DFFPOSX1 _11685_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .CLK(clk_bF$buf38),
    .Q(\genblk1[4].u_ce.LoadCtl [0])
);

AND2X2 _11265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3888_),
    .B(_3903_),
    .Y(_3905_)
);

FILL FILL_2__7901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7727_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9833_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1745_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Ain1 [0])
);

FILL FILL_0__7307_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .Y(_2225_)
);

FILL FILL_1__8790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13546_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .B(_5949__bF$buf2),
    .C(_6198_),
    .D(_6021_),
    .Y(_5846_)
);

FILL FILL_0__13126_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5832_),
    .B(_5800_),
    .C(_5833_),
    .Y(_5086_)
);

FILL FILL_1__9995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10053_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6846_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(_6847_),
    .Y(_6768_)
);

FILL FILL_0__7480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8685_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3609_)
);

FILL FILL_0__8265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3243_),
    .B(_3248_),
    .Y(_3249_)
);

NOR2X1 _10116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2851_),
    .B(_2835_),
    .Y(_2852_)
);

FILL FILL_2__9224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14609_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .Y(_483_)
);

NOR2X1 _7076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [10]),
    .Y(_84_)
);

INVX1 _11494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4118_),
    .Y(_4119_)
);

INVX1 _11074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_3722_)
);

FILL FILL_2__7710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7536_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [8]),
    .B(_1834__bF$buf2),
    .Y(_2439_)
);

FILL FILL_0__7116_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_2011_),
    .C(_2041_),
    .Y(_2042_)
);

MUX2X1 _12699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5178_),
    .B(_5177_),
    .S(_5151__bF$buf0),
    .Y(_5179_)
);

OAI21X1 _12279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4792_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4828_)
);

FILL FILL_1__14782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13775_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6010_),
    .B(_6012_),
    .C(_5998_),
    .Y(_6016_)
);

FILL FILL_0__13355_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5675_),
    .B(_5671_),
    .C(_5172_),
    .Y(_5677_)
);

FILL FILL_1__9384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10282_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [8]),
    .B(_6833__bF$buf2),
    .C(En_bF$buf3),
    .Y(_7058_)
);

INVX1 _14425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6710_),
    .Y(_6711_)
);

AND2X2 _14005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6318_),
    .B(_6321_),
    .Y(_6365_)
);

FILL FILL_2__12494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8074_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10765_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.LoadCtl [4])
);

NAND3X1 _10345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3035_),
    .B(_3056_),
    .C(_3039_),
    .Y(_3070_)
);

FILL FILL_0__11841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13279_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8913_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[1].u_ce.LoadCtl [0])
);

FILL FILL_1__7870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5348_),
    .B(_5351_),
    .C(_5381_),
    .Y(_5382_)
);

FILL FILL_0__12626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7765_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [4]),
    .Y(_2619_)
);

FILL FILL_0__7345_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2260_),
    .Y(_2261_)
);

NAND2X1 _9031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1860_)
);

NAND2X1 _12088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4646_)
);

FILL FILL_1__14591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833__bF$buf1),
    .B(_6881_),
    .Y(_6882_)
);

INVX1 _14234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [6]),
    .Y(_6549_)
);

FILL FILL_1__7506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11296_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3465_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3645_),
    .Y(_3358_)
);

NOR2X1 _10574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3274_),
    .B(_3260_),
    .Y(_3285_)
);

FILL FILL_0__10289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2887_),
    .C(_2886_),
    .Y(_2888_)
);

FILL FILL_2__10616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11230_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .Y(_1605_)
);

INVX1 _8302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1208_)
);

NOR2X1 _11779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4344_),
    .Y(_4350_)
);

FILL FILL_0__9088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_3993_),
    .C(_3524__bF$buf1),
    .Y(_3994_)
);

FILL FILL_1__13862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12435_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5200_)
);

AOI21X1 _12300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4833_),
    .B(_4362__bF$buf2),
    .C(_4604_),
    .Y(_4848_)
);

FILL FILL_0__12015_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2665_),
    .B(_2667_),
    .C(_2670_),
    .Y(_2671_)
);

OAI21X1 _9507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .B(_2313_),
    .C(_2311_),
    .Y(_2314_)
);

FILL FILL_1__8464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14227_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6161_),
    .C(_6287_),
    .Y(_6288_)
);

INVX2 _13505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .Y(_5888_)
);

FILL FILL_1__9669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7574_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [5]),
    .B(_1761_),
    .Y(_2473_)
);

FILL FILL_0__7154_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2069_),
    .Y(_2079_)
);

FILL FILL_0__10921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14598_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14883_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6774_),
    .CLK(clk_bF$buf50),
    .Q(\u_pa.acc_reg [7])
);

NAND2X1 _14463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [1]),
    .B(_6736_),
    .Y(_6740_)
);

NAND2X1 _14043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6400_),
    .Y(_6401_)
);

FILL FILL_1__7735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3100_),
    .B(_3103_),
    .Y(_3107_)
);

FILL FILL_2__10425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9071_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Ycalc [0]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Ycalc [2]),
    .Y(_1785_)
);

OAI21X1 _8531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1400_),
    .B(_1394_),
    .C(_1010__bF$buf1),
    .Y(_1427_)
);

NAND3X1 _8111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf4),
    .B(_988_),
    .C(_1025_),
    .Y(_1026_)
);

NAND2X1 _11588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [1]),
    .B(_4151_),
    .Y(_4184_)
);

OAI21X1 _11168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf2),
    .B(_3811_),
    .C(_3804_),
    .Y(_3812_)
);

FILL FILL_1__13671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.Y_ [1]),
    .Y(_2506_)
);

NAND2X1 _9316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_2132_)
);

FILL FILL_1__8693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13869_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6085_),
    .B(_5949__bF$buf1),
    .C(_6105_),
    .D(_6021_),
    .Y(_5842_)
);

FILL FILL_0__13029_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5755_),
    .B(_5174__bF$buf0),
    .C(_5765_),
    .D(_5766_),
    .Y(_5056_)
);

FILL FILL_0__14810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10376_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14519_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6507_),
    .CLK(clk_bF$buf4),
    .Q(\u_ot.Ycalc [7])
);

FILL FILL_0__7383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10310_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_760_),
    .B(_746_),
    .Y(_771_)
);

FILL FILL_0__8588_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_3516_)
);

FILL FILL_0__8168_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3156_),
    .B(_3154_),
    .Y(_3160_)
);

INVX1 _10019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2748_),
    .Y(_2759_)
);

FILL FILL_1__12942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11515_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [4]),
    .Y(_4371_)
);

NAND2X1 _14692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6917_)
);

NAND2X1 _14272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin1 [1]),
    .B(_6577_),
    .Y(_6578_)
);

FILL FILL_1__7544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13307_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .B(_2838_),
    .Y(_2924_)
);

FILL FILL_1__8749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_389_),
    .Y(_390_)
);

OAI21X1 _8760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1094_),
    .B(_1637_),
    .C(_1638_),
    .Y(_875_)
);

OR2X2 _8340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1244_),
    .B(_1240_),
    .Y(_1245_)
);

OR2X2 _11397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4028_),
    .B(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4029_)
);

FILL FILL_2__7613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7859_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(_2706_),
    .S(_2649__bF$buf2),
    .Y(_2708_)
);

FILL FILL_0__7439_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2348_),
    .Y(_2349_)
);

OAI21X1 _9125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1950_)
);

FILL FILL_1__8082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6324_),
    .B(_6323_),
    .Y(_6325_)
);

FILL FILL_0__13678_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5917_),
    .B(_5887_),
    .C(_5922_),
    .Y(\genblk1[7].u_ce.X_ [1])
);

FILL FILL_0__13258_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5584_),
    .B(_5564_),
    .Y(_5585_)
);

FILL FILL_1__9287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10185_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6968_),
    .B(_6955_),
    .C(_6834_),
    .Y(_6779_)
);

NAND3X1 _14328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Xin12b [10]),
    .C(_6626_),
    .Y(_6627_)
);

FILL FILL_0__7192_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_589_),
    .Y(_593_)
);

FILL FILL_0__8397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3347_),
    .B(_3317_),
    .C(_3348_),
    .Y(_2577_)
);

OAI21X1 _10248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2957_),
    .C(_2977_),
    .Y(_2978_)
);

FILL FILL_1__12751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11324_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6433_),
    .B(_6431_),
    .Y(_6437_)
);

NAND2X1 _8816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [1]),
    .B(_1637_),
    .Y(_1670_)
);

FILL FILL_1__7773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12949_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5270_),
    .B(_5288_),
    .C(_5289_),
    .Y(_5290_)
);

FILL FILL_0__12529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7668_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9774_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1686_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Ycalc [9])
);

FILL FILL_0__7248_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2167_),
    .C(_1903_),
    .Y(_2169_)
);

FILL FILL_1__11602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14074_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf3),
    .B(_6141_),
    .C(_6140_),
    .Y(_6142_)
);

FILL FILL_0__13067_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5795_),
    .B(_5105_),
    .Y(_5800_)
);

FILL FILL_1__9096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12807_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [2]),
    .Y(_6800_)
);

OAI21X1 _14137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6475_),
    .B(_6459_),
    .C(_6476_),
    .Y(_5874_)
);

FILL FILL_1__7829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_85_),
    .Y(_803_)
);

NAND2X1 _7420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .B(_324_),
    .Y(_410_)
);

FILL FILL_1__11199_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3552_),
    .B(_3504_),
    .Y(_3554_)
);

NAND2X1 _10477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(_3193_),
    .Y(_3195_)
);

NAND2X1 _10057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf2),
    .B(_2705_),
    .Y(_2795_)
);

FILL FILL_1__12980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11133_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1514_),
    .B(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1515_)
);

NAND3X1 _8205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1084_),
    .B(_1101_),
    .C(_1083_),
    .Y(_1115_)
);

FILL FILL_1__7582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12758_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5109_)
);

FILL FILL_0__12338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4326_),
    .B(_4750_),
    .C(_4753_),
    .Y(_4756_)
);

FILL FILL257250x169350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10272_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6195_),
    .B(_6138_),
    .C(_6191_),
    .Y(_6196_)
);

OAI21X1 _13408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5830_),
    .B(_5800_),
    .C(_5831_),
    .Y(_5085_)
);

FILL FILL_2__7651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7477_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .B(_2384_),
    .Y(_1704_)
);

NOR2X1 _9163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .B(_1964_),
    .Y(_1986_)
);

FILL FILL_1__11831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .B(vdd),
    .C(_5926__bF$buf4),
    .Y(_5959_)
);

FILL FILL_0__13296_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5621_)
);

FILL FILL_2__13203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9203_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6983_),
    .B(_6996_),
    .Y(_7003_)
);

NAND3X1 _14366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6658_),
    .C(_6659_),
    .Y(_6660_)
);

FILL FILL_1__7638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2755_),
    .B(_2962_),
    .Y(_3014_)
);

FILL FILL_0__11782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11362_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8854_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_852_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Xcalc [1])
);

NAND2X1 _8434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [10]),
    .Y(_1334_)
);

INVX1 _8014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [5]),
    .Y(_935_)
);

FILL FILL_1__7391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12987_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_5304_),
    .Y(_5326_)
);

FILL FILL_0__12147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [9]),
    .B(_4362__bF$buf4),
    .Y(_4970_)
);

OAI21X1 _12012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4573_),
    .B(_4572_),
    .C(_4420_),
    .Y(_4574_)
);

OR2X2 _9639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2428_),
    .B(_2436_),
    .Y(_2437_)
);

NAND2X1 _9219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1992_),
    .B(_2008_),
    .Y(_2039_)
);

FILL FILL_1__8596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6012_),
    .B(_6010_),
    .Y(_6013_)
);

AOI21X1 _13217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5659_),
    .B(_5188__bF$buf1),
    .C(_5430_),
    .Y(_5674_)
);

FILL FILL_0__14713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256050x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2201_),
    .C(_2196_),
    .Y(_2205_)
);

FILL FILL_1__11220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256050x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5807_),
    .Y(_5822_)
);

NAND2X1 _7705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_679_),
    .Y(_681_)
);

FILL FILL_2__13012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4274_),
    .B(_4277_),
    .C(_4280_),
    .Y(_4281_)
);

FILL FILL_0__9012_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833__bF$buf0),
    .B(_6834_),
    .Y(_6760_)
);

DFFPOSX1 _14175_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5851_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Xcalc [3])
);

FILL FILL_1__7867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5332_),
    .B(_5348_),
    .Y(_5379_)
);

FILL FILL_1_BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2782_),
    .B(_2785_),
    .Y(_2831_)
);

FILL FILL_2__10977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11171_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1267_),
    .C(_1549_),
    .Y(_1550_)
);

OAI21X1 _8243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1150_),
    .C(_1151_),
    .Y(_1152_)
);

FILL FILL_1__10911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12796_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Xcalc [11]),
    .Y(_5143_)
);

FILL FILL_0__12376_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4791_),
    .B(_4767_),
    .C(_4790_),
    .Y(_4792_)
);

INVX1 _9868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [10]),
    .Y(_2616_)
);

INVX1 _9448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2241_),
    .Y(_2258_)
);

NAND2X1 _9028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [4]),
    .Y(_1857_)
);

FILL FILL_0__8703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14588_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6224_),
    .Y(_6232_)
);

DFFPOSX1 _13446_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5046_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [5])
);

OAI21X1 _13026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .C(_5491_),
    .Y(_5492_)
);

FILL FILL_2__13908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10022_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7934_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [5])
);

NAND2X1 _7514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_448_),
    .Y(_500_)
);

FILL FILL_2__13661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9661_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .B(_4495_),
    .C(_4496_),
    .Y(_4497_)
);

FILL FILL_0__9241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11227_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _11512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3446_),
    .B(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .C(_4135_),
    .D(_4134_),
    .Y(_3386_)
);

NOR2X1 _8719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_992_),
    .Y(_1602_)
);

FILL FILL_1__7676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [4]),
    .Y(_5197_)
);

FILL FILL_1__14800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8892_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_890_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Yin12b [9])
);

FILL FILL_0_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1352_),
    .Y(_1371_)
);

FILL FILL_0_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Xcalc [1]),
    .C(_968_),
    .D(_930_),
    .Y(_969_)
);

FILL FILL_0_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13192_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5324_),
    .B(_5352_),
    .Y(_5362_)
);

FILL FILL_0__12185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4995_),
    .B(_4997_),
    .C(_4999_),
    .Y(_4232_)
);

AOI21X1 _12050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4595_),
    .B(_4593_),
    .C(_4599_),
    .Y(_4610_)
);

FILL FILL256950x104550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [11]),
    .B(_1834__bF$buf1),
    .Y(_2471_)
);

AOI21X1 _9257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2044_),
    .B(_2053_),
    .C(_2075_),
    .Y(_2076_)
);

FILL FILL_1__11925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6047_),
    .C(_6048_),
    .Y(_6049_)
);

OAI21X1 _13255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf3),
    .B(_5709_),
    .C(_5188__bF$buf0),
    .Y(_5710_)
);

FILL FILL_0__14751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10251_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_714_),
    .Y(_716_)
);

AND2X2 _7323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_271_),
    .Y(_317_)
);

FILL FILL_2__13050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11456_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Xcalc [0]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Xcalc [2]),
    .Y(_4315_)
);

FILL FILL_0__9050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11036_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3957_),
    .C(_3937_),
    .Y(_3958_)
);

NAND2X1 _8948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [6]),
    .B(_1765_),
    .Y(_1782_)
);

OAI21X1 _8528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1336_),
    .C(_1423_),
    .Y(_1424_)
);

OAI21X1 _8108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1021_),
    .C(_1022_),
    .Y(_1023_)
);

FILL FILL_1__7485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13248_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5384_),
    .B(_5393_),
    .C(_5415_),
    .Y(_5416_)
);

NAND2X1 _12526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [1]),
    .B(_5000_),
    .Y(_4265_)
);

AOI21X1 _12106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4636_),
    .B(_4657_),
    .C(_4655_),
    .Y(_4663_)
);

FILL FILL_0__13602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9211_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1098_),
    .C(_1164_),
    .Y(_1188_)
);

FILL FILL_0__14807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12741_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _9486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1794_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2294_),
    .D(_2292_),
    .Y(_1697_)
);

OAI21X1 _9066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(_1863_),
    .C(_1848__bF$buf1),
    .Y(_1893_)
);

FILL FILL_1__11734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13199_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13484_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5084_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain12b [11])
);

NAND2X1 _13064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5528_),
    .B(_5527_),
    .Y(_5529_)
);

FILL FILL_0__14560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9106_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6913_),
    .Y(_6914_)
);

NAND2X1 _14269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [2]),
    .B(_6562__bF$buf4),
    .Y(_6576_)
);

FILL FILL_0__10480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10060_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7972_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_56_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Yin12b [5])
);

OAI21X1 _7552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_514_),
    .C(_527_),
    .Y(_536_)
);

INVX8 _7132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_134_)
);

AOI22X1 _10189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2616_),
    .B(_2672__bF$buf0),
    .C(_2921_),
    .D(_2744_),
    .Y(_2525_)
);

FILL FILL_1__12692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12272_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4505_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4533_),
    .Y(_4198_)
);

NAND2X1 _11550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4162_),
    .Y(_4164_)
);

FILL FILL_0__11265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [0]),
    .B(_3510__bF$buf3),
    .Y(_3775_)
);

NAND2X1 _8757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_924_),
    .B(_930_),
    .Y(_1636_)
);

NAND3X1 _8337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_1218_),
    .C(_1197_),
    .Y(_1242_)
);

FILL FILL_1__7294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13057_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5166_),
    .B(_5203_),
    .C(_5188__bF$buf0),
    .Y(_5233_)
);

NAND2X1 _12335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4878_),
    .B(_4879_),
    .Y(_4880_)
);

FILL FILL_0__13831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9020_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .B(_1002_),
    .C(_973__bF$buf3),
    .Y(_1005_)
);

FILL FILL_0__14616_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14901_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6792_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [5])
);

FILL FILL_2__11189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7189_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_2109_),
    .S(_1811__bF$buf3),
    .Y(_2112_)
);

FILL FILL_1__11963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8550_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(\genblk1[4].u_ce.Xcalc [9]),
    .C(_3438_),
    .Y(_3480_)
);

FILL FILL_2__8148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10116_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3120_),
    .B(_3123_),
    .Y(_3124_)
);

NOR2X1 _13293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5745_),
    .B(_5709_),
    .Y(_5746_)
);

NAND2X1 _7608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_589_),
    .Y(_590_)
);

FILL FILL_1__12748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9335_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_3429_)
);

NAND2X1 _14498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(\genblk1[7].u_ce.ISout ),
    .Y(_6759_)
);

NAND2X1 _14078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6431_),
    .B(_6433_),
    .Y(_6434_)
);

FILL FILL_1__8711_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [7]),
    .Y(_751_)
);

OAI21X1 _7361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_352_),
    .C(_353_),
    .Y(_354_)
);

FILL FILL_1__12081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11401_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1816_)
);

OAI21X1 _8566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1377_),
    .C(_1423_),
    .Y(_1460_)
);

INVX1 _8146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .Y(_1059_)
);

FILL FILL_1__10814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13286_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5451_),
    .B(_5449_),
    .S(_5151__bF$buf4),
    .Y(_5452_)
);

FILL FILL_0__12699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12279_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12564_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4218_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Acalc [3])
);

NAND2X1 _12144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4699_),
    .B(_4698_),
    .Y(_4700_)
);

FILL FILL_0__13640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8606_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6139_)
);

NAND2X1 _13349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5796_),
    .Y(_5798_)
);

FILL FILL_0__14845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14425_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6932_),
    .B(_6930_),
    .C(_6933_),
    .Y(_6776_)
);

FILL FILL_0__14005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8377_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_3328_)
);

FILL FILL_0__10345_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2940_),
    .Y(_2941_)
);

NAND2X1 _7837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_799_),
    .Y(_801_)
);

AOI22X1 _7417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_158__bF$buf1),
    .C(_407_),
    .D(_230_),
    .Y(_11_)
);

FILL FILL257250x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9564_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4385_),
    .B(_4360_),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4404_)
);

FILL FILL_0__9144_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .B(_4045_),
    .Y(_4046_)
);

FILL FILL256950x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8100_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_566_),
    .Y(_573_)
);

FILL FILL_1__14703_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_171_)
);

FILL FILL_1__9725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11210_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [1]),
    .Y(_1659_)
);

NAND2X1 _8375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf2),
    .B(_1273_),
    .Y(_1278_)
);

FILL FILL_1__10623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13095_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5245_),
    .B(_5174__bF$buf1),
    .C(_5269_),
    .D(_5246_),
    .Y(_5032_)
);

NAND2X1 _12373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4912_),
    .B(_4914_),
    .Y(_4915_)
);

FILL FILL_0__12088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6357_),
    .B(_6356_),
    .Y(_6358_)
);

NAND2X1 _13578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(_5955_),
    .Y(_5956_)
);

AOI21X1 _13158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5617_),
    .B(_5593_),
    .C(_5616_),
    .Y(_5618_)
);

FILL FILL_0__14654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10154_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_623_),
    .Y(_626_)
);

OAI21X1 _7226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_221_),
    .C(_207_),
    .Y(_225_)
);

FILL FILL_1__12786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11359_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11644_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3384_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[4].u_ce.Acalc [7])
);

AOI22X1 _11224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3478_),
    .B(_3510__bF$buf4),
    .C(_3865_),
    .D(_3508_),
    .Y(_3368_)
);

FILL FILL_0__12720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7388_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .B(_5321_),
    .C(_5322_),
    .Y(_5323_)
);

OAI21X1 _12429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4965_),
    .B(_4967_),
    .C(_4953_),
    .Y(_4223_)
);

AND2X2 _12009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4567_),
    .B(_4570_),
    .Y(_4571_)
);

FILL FILL_0__13925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1095_)
);

FILL FILL257550x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7877_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4710_),
    .B(_4735_),
    .C(_4362__bF$buf1),
    .Y(_4736_)
);

FILL FILL_2__12224_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2201_),
    .C(_2197_),
    .Y(_2202_)
);

FILL FILL_1__11217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8644_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3569_),
    .Y(_3570_)
);

FILL FILL_0__8224_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5816_),
    .B(_5804_),
    .C(_5820_),
    .Y(_5075_)
);

FILL FILL_2__9603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_807_),
    .C(_823_),
    .Y(_53_)
);

OAI21X1 _7455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_443_),
    .C(_156_),
    .Y(_444_)
);

FILL FILL_1__12175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11588_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4438_),
    .B(_4440_),
    .Y(_4441_)
);

FILL FILL_0__9182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11168_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4080_),
    .Y(_4081_)
);

NAND2X1 _11033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3681_),
    .B(_3682_),
    .Y(_3683_)
);

FILL FILL_2__11915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7915_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2400_),
    .Y(_2401_)
);

AOI22X1 _12658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Xcalc [0]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Xcalc [2]),
    .Y(_5141_)
);

AOI22X1 _12238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4771_),
    .B(_4348__bF$buf2),
    .C(_4789_),
    .D(_4786_),
    .Y(_4210_)
);

FILL FILL_1__14741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10241_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7017_),
    .B(_7018_),
    .C(_7020_),
    .Y(_7021_)
);

FILL FILL_2__12453_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1991_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2019_),
    .Y(_1684_)
);

FILL FILL_1__11866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8033_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10724_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2550_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Acalc [11])
);

FILL FILL_0__10439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3030_),
    .Y(_3031_)
);

OAI21X1 _13196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5618_),
    .B(_5653_),
    .C(_5651_),
    .Y(_5654_)
);

FILL FILL_0__11800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9658_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4485_),
    .B(_4490_),
    .C(_4493_),
    .Y(_4494_)
);

FILL FILL_0__9238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4132_),
    .B(_4131_),
    .Y(_4133_)
);

FILL FILL_0__10192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8614_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_661_),
    .B(_660_),
    .C(_653_),
    .Y(_24_)
);

NAND2X1 _7264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf1),
    .B(_163_),
    .Y(_261_)
);

DFFPOSX1 _11682_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3422_),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.Ain1 [1])
);

FILL FILL_0__11397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3899_),
    .C(_3895_),
    .Y(_3902_)
);

FILL FILL_2__11724_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8889_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_887_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[1].u_ce.Yin12b [10])
);

NAND3X1 _8469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .B(_1367_),
    .C(_1366_),
    .Y(_1368_)
);

OAI21X1 _8049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(\genblk1[1].u_ce.Xcalc [9]),
    .C(_924_),
    .Y(_966_)
);

FILL FILL_0__7724_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9830_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1742_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Ain12b [7])
);

FILL FILL_0__7304_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .B(_2221_),
    .C(_1848__bF$buf2),
    .Y(_2222_)
);

FILL FILL_1__13189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .C(_5359_),
    .Y(_5036_)
);

NAND2X1 _12467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(_4997_),
    .Y(_4998_)
);

NAND2X1 _12047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4605_),
    .B(_4606_),
    .Y(_4607_)
);

FILL FILL_1__14130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14328_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6844_),
    .Y(_6845_)
);

FILL FILL_1__11255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8682_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3583_),
    .B(_3600_),
    .C(_3601_),
    .Y(_3606_)
);

FILL FILL_0__8262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10668_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _10533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .B(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .C(_3244_),
    .D(_3246_),
    .Y(_2544_)
);

FILL FILL_0__10248_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(_2847_),
    .C(_2848_),
    .Y(_2849_)
);

FILL FILL_2__9641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9467_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [6]),
    .B(_4279_),
    .Y(_4312_)
);

FILL FILL_0__9047_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3955_)
);

FILL FILL_1__13821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14606_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_240_),
    .Y(_480_)
);

INVX2 _7073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_81_)
);

NOR2X1 _11491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3506_),
    .Y(_4116_)
);

OAI21X1 _11071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3664_),
    .B(_3718_),
    .C(_3716_),
    .Y(_3719_)
);

FILL FILL_1__9628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11113_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1581_),
    .B(\genblk1[1].u_ce.Ain12b [6]),
    .Y(_1583_)
);

AOI21X1 _8278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(_1158_),
    .C(_1183_),
    .Y(_1185_)
);

FILL FILL_1__10946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7113_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5170_),
    .Y(_5176_)
);

AOI21X1 _12276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4819_),
    .C(_4824_),
    .Y(_4825_)
);

FILL FILL_2__12738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14557_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7054_),
    .B(_7055_),
    .C(_6833__bF$buf0),
    .Y(_7056_)
);

FILL FILL_0__14137_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .B(_6707_),
    .Y(_6708_)
);

NAND2X1 _14002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6341_),
    .B(_6361_),
    .Y(_6362_)
);

FILL FILL_2__12491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10477_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10762_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.LoadCtl [1])
);

FILL FILL_0__10057_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3066_),
    .B(_3067_),
    .C(_2670_),
    .Y(_3068_)
);

FILL FILL_2__9450_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7969_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_53_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin12b [6])
);

NAND2X1 _7549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_532_),
    .Y(_534_)
);

OAI21X1 _7129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_83_),
    .C(_131_),
    .Y(\genblk1[0].u_ce.X_ [1])
);

FILL FILL_2__13696_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8910_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_908_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Ain1 [1])
);

FILL FILL_1__12689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9696_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf5),
    .B(_4417_),
    .C(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .Y(_4531_)
);

FILL FILL_0__9276_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3444_),
    .B(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_4162_)
);

OAI21X1 _11127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3769_),
    .B(_3772_),
    .C(_3579_),
    .Y(_3773_)
);

FILL FILL_1__13630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11762_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _8087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_1002_)
);

FILL FILL_1__10335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert101 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert103 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert106 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4643_)
);

FILL FILL_2__12967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8547_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3477_),
    .B(_3476_),
    .Y(\genblk1[4].u_ce.X_ [0])
);

FILL FILL_0__8127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6878_),
    .B(_6877_),
    .Y(_6879_)
);

INVX1 _14231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [5]),
    .Y(_6547_)
);

FILL FILL_1__7503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11293_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3627_),
    .B(_3642_),
    .Y(_3643_)
);

AOI21X1 _10571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3279_),
    .B(_3215_),
    .C(\genblk1[3].u_ce.Ain12b [8]),
    .Y(_3282_)
);

FILL FILL_0__10286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _10151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2864_),
    .C(_2837_),
    .Y(_2885_)
);

FILL FILL_1__8708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10613_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_738_),
    .Y(_749_)
);

NAND3X1 _7358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_350_),
    .C(_349_),
    .Y(_351_)
);

FILL FILL_1__12498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4322_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4347_),
    .Y(_4190_)
);

FILL FILL_0__9085_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3909_),
    .C(_3937_),
    .Y(_3991_)
);

FILL FILL_0__12852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7818_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf4),
    .B(_2649__bF$buf4),
    .Y(_2668_)
);

AOI21X1 _9504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2305_),
    .C(_2310_),
    .Y(_2311_)
);

FILL FILL_1__8461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13637_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6280_),
    .B(_6264_),
    .C(_6278_),
    .Y(_6285_)
);

FILL FILL_0__13217_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [1]),
    .Y(_5885_)
);

FILL FILL_1__9666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10144_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6929_),
    .B(_6924_),
    .Y(_6931_)
);

FILL FILL_0__7571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2690_),
    .B(_3324_),
    .C(_3326_),
    .Y(_2558_)
);

INVX1 _10207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2938_)
);

FILL FILL_1__12710_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5536_),
    .B(_5561_),
    .C(_5188__bF$buf3),
    .Y(_5562_)
);

FILL FILL_0__11703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9315_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14880_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6771_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [4])
);

FILL FILL_0__14595_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6727_),
    .B(_6737_),
    .C(_6738_),
    .Y(_6518_)
);

INVX1 _14040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .Y(_6398_)
);

FILL FILL_1__7732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3102_),
    .B(_3103_),
    .Y(_3104_)
);

FILL FILL_1__8937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8517_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_514_),
    .C(_569_),
    .Y(_570_)
);

NAND3X1 _7167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(gnd),
    .C(_135__bF$buf4),
    .Y(_168_)
);

OAI21X1 _11585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3523_),
    .C(_4182_),
    .Y(_3412_)
);

OAI21X1 _11165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3628_),
    .C(_3808_),
    .Y(_3809_)
);

FILL FILL_2__7801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7627_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_1759_),
    .C(_2504_),
    .Y(_1734_)
);

FILL FILL_0__7207_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2129_)
);

FILL FILL_1__8690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13866_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6078_),
    .B(_6102_),
    .Y(_6103_)
);

FILL FILL_0__13026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5763_),
    .B(_5762_),
    .Y(_5764_)
);

FILL FILL_1__9895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10373_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14516_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6504_),
    .CLK(clk_bF$buf4),
    .Q(\u_ot.Ycalc [4])
);

FILL FILL_2__7398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8585_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(\genblk1[4].u_ce.Xin12b [6]),
    .S(gnd),
    .Y(_3513_)
);

FILL FILL_0__8165_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3154_),
    .B(_3156_),
    .Y(_3157_)
);

AOI22X1 _10016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2696_),
    .B(_2755_),
    .C(_2754_),
    .D(_2692_),
    .Y(_2756_)
);

FILL FILL_2__9964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10651_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .Y(_387_)
);

OAI21X1 _11394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_4014_),
    .C(_3524__bF$buf4),
    .Y(_4026_)
);

FILL FILL_2__7610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7856_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_2703_),
    .S(_2649__bF$buf0),
    .Y(_2705_)
);

FILL FILL_0__7436_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2339_),
    .Y(_2346_)
);

OAI21X1 _9122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1945_),
    .B(_1946_),
    .C(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_1947_)
);

DFFPOSX1 _12599_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4253_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Ain12b [8])
);

NAND3X1 _12179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf1),
    .B(_4732_),
    .C(_4727_),
    .Y(_4733_)
);

FILL FILL_2__8815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14262_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6318_),
    .B(_6321_),
    .Y(_6322_)
);

FILL FILL_0__13675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13255_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .B(\genblk1[7].u_ce.Xcalc [5]),
    .C(_5891_),
    .D(\genblk1[7].u_ce.Xcalc [7]),
    .Y(_5920_)
);

NAND3X1 _13120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5152_),
    .B(_5576_),
    .C(_5579_),
    .Y(_5582_)
);

FILL FILL_1__9284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6965_),
    .B(_6962_),
    .Y(_6966_)
);

AND2X2 _14325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6595_),
    .B(_6611_),
    .Y(_6624_)
);

FILL FILL_2__12394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8394_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf0),
    .B(_3313_),
    .C(_3346_),
    .Y(_2576_)
);

NAND3X1 _10245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf3),
    .B(_2974_),
    .C(_2952_),
    .Y(_2975_)
);

FILL FILL_0__11741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1009_),
    .C(_1668_),
    .Y(_898_)
);

FILL FILL_1__7770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12946_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5285_),
    .B(_5286_),
    .C(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5287_)
);

FILL FILL_0__12526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7665_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9771_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1683_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Ycalc [6])
);

FILL FILL_0__7245_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2164_),
    .Y(_2166_)
);

FILL FILL_2__8624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14689_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14554_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [5]),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.LoadCtl [6])
);

FILL FILL_0__14269_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6202_),
    .B(_6455_),
    .C(_6474_),
    .Y(_5873_)
);

FILL FILL_1__7826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3523_),
    .B(_3540_),
    .C(_3548_),
    .Y(_3551_)
);

FILL FILL_0__10189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3187_),
    .B(_3189_),
    .C(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3192_)
);

NAND2X1 _10054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2792_)
);

FILL FILL_2__10936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11130_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1500_),
    .C(_1010__bF$buf4),
    .Y(_1512_)
);

AOI22X1 _8202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_943_),
    .B(_996__bF$buf4),
    .C(_1112_),
    .D(_1068_),
    .Y(_843_)
);

DFFPOSX1 _11679_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3419_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[4].u_ce.Ain12b [4])
);

NAND2X1 _11259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .B(_3898_),
    .Y(_3899_)
);

FILL FILL_1__13762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12755_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .B(\genblk1[6].u_ce.LoadCtl [3]),
    .Y(_5106_)
);

FILL FILL_0__12335_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4751_),
    .C(_4752_),
    .Y(_4753_)
);

DFFPOSX1 _9827_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1739_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Ain12b [8])
);

NAND3X1 _9407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf2),
    .B(_2218_),
    .C(_2213_),
    .Y(_2219_)
);

FILL FILL_1__8784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14127_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6192_),
    .B(_6191_),
    .C(_6189_),
    .Y(_6193_)
);

OAI21X1 _13405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf4),
    .B(_5796_),
    .C(_5829_),
    .Y(_5084_)
);

FILL FILL_1__9989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7474_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2381_),
    .Y(_2382_)
);

NAND3X1 _9160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .B(_1981_),
    .C(_1982_),
    .Y(_1983_)
);

FILL FILL_0__10821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14498_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6999_),
    .B(_6992_),
    .C(_6977_),
    .Y(_7000_)
);

FILL FILL_0__14078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6651_),
    .C(_6652_),
    .Y(_6657_)
);

FILL FILL_1__7635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13818_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2884_),
    .C(_3010_),
    .Y(_3011_)
);

FILL FILL_2__10325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9391_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8851_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_849_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Ycalc [10])
);

OAI21X1 _8431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996__bF$buf4),
    .B(_1331_),
    .C(_1310_),
    .Y(_853_)
);

INVX1 _8011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [9]),
    .Y(_932_)
);

AOI21X1 _11488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4104_),
    .B(_4112_),
    .C(_3510__bF$buf0),
    .Y(_4114_)
);

AND2X2 _11068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3715_),
    .B(_3687_),
    .Y(_3716_)
);

FILL FILL_1__13991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x100950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12144_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .Y(_2434_)
);

AOI21X1 _9216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2023_),
    .B(_2036_),
    .C(_1836_),
    .Y(_2037_)
);

FILL FILL_1__8593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13769_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6009_),
    .B(_6006_),
    .C(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6010_)
);

FILL FILL_0__13349_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5654_),
    .B(_5664_),
    .C(_5670_),
    .Y(_5671_)
);

FILL FILL_0__14710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .B(_7049_),
    .Y(_7053_)
);

OAI21X1 _14419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6557_),
    .B(\u_ot.LoadCtl_6_bF$buf0 ),
    .C(_6705_),
    .Y(_6510_)
);

FILL FILL_2_BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10210_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_675_),
    .C(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_678_)
);

FILL FILL_0__8488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8068_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10759_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2585_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[3].u_ce.Ain0 [0])
);

NAND2X1 _10339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3064_),
    .B(_3063_),
    .Y(_3065_)
);

FILL FILL_1__12842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11415_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_4278_)
);

OAI21X1 _14592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6826_),
    .B(_6831_),
    .C(_6832_),
    .Y(_6798_)
);

DFFPOSX1 _14172_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5848_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Xcalc [0])
);

DFFPOSX1 _8907_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_905_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Ain12b [4])
);

FILL FILL_1__7864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5363_),
    .B(_5376_),
    .C(_5176_),
    .Y(_5377_)
);

FILL FILL_1_BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2808_),
    .B(_2672__bF$buf0),
    .C(_2828_),
    .D(_2744_),
    .Y(_2521_)
);

FILL FILL_1__8649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10134_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [6]),
    .Y(_294_)
);

NAND2X1 _8660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [4]),
    .B(_996__bF$buf3),
    .Y(_1547_)
);

OAI21X1 _8240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1110_),
    .B(_1092_),
    .C(_1148_),
    .Y(_1149_)
);

NAND2X1 _11297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3911_),
    .B(_3913_),
    .Y(_3935_)
);

FILL FILL_2__7513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7759_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2613_),
    .C(_2606_),
    .Y(_2614_)
);

FILL FILL_0__7339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2255_),
    .Y(_2256_)
);

OAI21X1 _9025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1852_),
    .C(_1853_),
    .Y(_1854_)
);

FILL FILL_0__8700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13998_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6222_),
    .B(_6228_),
    .Y(_6229_)
);

FILL FILL_0__13578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13158_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13443_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5043_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Xcalc [2])
);

AOI21X1 _13023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .B(_5483_),
    .C(_5481_),
    .Y(_5489_)
);

FILL FILL_1__9187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10085_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6871_),
    .B(_6872_),
    .C(_6868_),
    .Y(_6876_)
);

INVX1 _14228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [4]),
    .Y(_6545_)
);

FILL FILL_0__7092_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7931_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xcalc [2])
);

OAI21X1 _7511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_370_),
    .C(_496_),
    .Y(_497_)
);

AOI21X1 _10988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3638_),
    .B(_3635_),
    .C(_3628_),
    .Y(_3640_)
);

FILL FILL_0__8297_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3278_),
    .Y(_3279_)
);

INVX1 _10148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2872_),
    .Y(_2882_)
);

FILL FILL_1__12651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11224_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(_1598_),
    .C(_996__bF$buf3),
    .Y(_1600_)
);

FILL FILL_1__7673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12849_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5192_),
    .C(_5193_),
    .Y(_5194_)
);

FILL FILL_0__12429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10363_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6264_),
    .B(_6281_),
    .Y(_6283_)
);

FILL FILL_2__7322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7568_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2464_),
    .B(_2468_),
    .Y(_2469_)
);

FILL FILL_0__7148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .B(_2067_),
    .C(_2072_),
    .Y(_2073_)
);

FILL FILL_1__11922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x169350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14394_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6046_)
);

FILL FILL_0__13387_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5706_),
    .Y(_5707_)
);

FILL FILL_1__12707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9714_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14877_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6768_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [1])
);

INVX1 _14457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .Y(_6736_)
);

NAND3X1 _14037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6350_),
    .B(_6379_),
    .C(_6352_),
    .Y(_6395_)
);

FILL FILL_1__7729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_672_),
    .C(_712_),
    .Y(_713_)
);

AOI22X1 _7320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_158__bF$buf1),
    .C(_314_),
    .D(_230_),
    .Y(_7_)
);

FILL FILL_1__11099_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3457_),
    .C(_3458_),
    .Y(_3459_)
);

NAND3X1 _10377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf3),
    .B(_3100_),
    .C(_3097_),
    .Y(_3101_)
);

FILL FILL_1__12880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11033_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(\genblk1[2].u_ce.Ycalc [8]),
    .C(_1762_),
    .Y(_1779_)
);

NAND2X1 _8525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .B(_1399_),
    .Y(_1421_)
);

OAI21X1 _8105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_)
);

FILL FILL_1__7482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13245_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .B(_5407_),
    .C(_5412_),
    .Y(_5413_)
);

FILL FILL_0__12658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12238_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5025_),
    .B(_4997_),
    .C(_4263_),
    .Y(_4256_)
);

AOI21X1 _12103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4660_),
    .B(_4659_),
    .C(_4350_),
    .Y(_4661_)
);

FILL FILL_1__8687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10172_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6056_),
    .B(_6058_),
    .C(_6046_),
    .Y(_6100_)
);

NOR2X1 _13308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5757_),
    .B(_5760_),
    .Y(_5761_)
);

FILL FILL_0__14804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7377_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .Y(_2292_)
);

AOI21X1 _9063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1871_),
    .B(_1846_),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1890_)
);

FILL FILL_1__11731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13196_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13481_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5081_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin0 [0])
);

NAND2X1 _13061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5525_),
    .B(_5524_),
    .Y(_5526_)
);

FILL FILL_2__13103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6878_),
    .Y(_6911_)
);

NOR2X1 _14266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .Y(_6573_)
);

FILL FILL_1__7538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2918_),
    .B(_2861_),
    .C(_2914_),
    .Y(_2919_)
);

FILL FILL_0__11262_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1626_),
    .C(_1629_),
    .Y(_1634_)
);

NAND3X1 _8334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1219_),
    .C(_1205_),
    .Y(_1239_)
);

FILL FILL_1__7291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12887_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5211_),
    .B(_5186_),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5230_)
);

FILL FILL_0__12467_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4876_),
    .B(vdd),
    .S(_4875_),
    .Y(_4877_)
);

FILL FILL_0__12047_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf0),
    .B(_2664_),
    .C(_2701_),
    .Y(_2702_)
);

NAND2X1 _9539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [0]),
    .B(_1834__bF$buf2),
    .Y(_2344_)
);

NAND3X1 _9119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1931_),
    .B(_1943_),
    .C(_1941_),
    .Y(_1944_)
);

FILL FILL_1__8496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6314_),
    .B(_6311_),
    .Y(_6319_)
);

INVX1 _13537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [3]),
    .Y(_5917_)
);

OAI21X1 _13117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5577_),
    .C(_5578_),
    .Y(_5579_)
);

FILL FILL_0__14613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1971_),
    .C(_2108_),
    .Y(_2109_)
);

FILL FILL_1__11960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10113_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5742_),
    .Y(_5743_)
);

NAND3X1 _7605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf4),
    .B(_586_),
    .C(_583_),
    .Y(_587_)
);

FILL FILL_2__13332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11318_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4073_),
    .B(_4162_),
    .C(_3427_),
    .Y(_3420_)
);

OAI21X1 _14495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6647_),
    .C(_6757_),
    .Y(_6534_)
);

INVX1 _14075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6430_),
    .Y(_6431_)
);

FILL FILL_1__7767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5271_),
    .B(_5283_),
    .C(_5281_),
    .Y(_5284_)
);

FILL FILL_2__10877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9913_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1813_)
);

NAND2X1 _8563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [9]),
    .B(_996__bF$buf1),
    .Y(_1457_)
);

NAND2X1 _8143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(_1055_),
    .Y(_1056_)
);

FILL FILL_1__10811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5311_),
    .C(_5448_),
    .Y(_5449_)
);

FILL FILL_0__12696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12276_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12561_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4215_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Acalc [0])
);

AOI21X1 _12141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4695_),
    .B(_4696_),
    .C(_4370_),
    .Y(_4697_)
);

DFFPOSX1 _9768_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1680_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Ycalc [3])
);

NAND3X1 _9348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(_2162_),
    .C(_2160_),
    .Y(_2163_)
);

FILL FILL_0__8603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x111750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6098_),
    .B(_6127_),
    .C(_6126_),
    .Y(_6136_)
);

NOR2X1 _13346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5794_),
    .B(_5795_),
    .Y(_5796_)
);

FILL FILL_2__13808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10342_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_797_),
    .B(_798_),
    .Y(_799_)
);

OAI21X1 _7414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_347_),
    .C(_400_),
    .Y(_405_)
);

FILL FILL_2__13141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11547_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4324__bF$buf4),
    .Y(_4401_)
);

FILL FILL_0__9141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11127_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .Y(_4043_)
);

NOR2X1 _8619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_1509_)
);

FILL FILL_1__7996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5102_),
    .Y(_5103_)
);

FILL FILL_1__14700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9302_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [0]),
    .Y(_1657_)
);

NAND2X1 _8372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1274_),
    .Y(_1275_)
);

FILL FILL_1__10620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13092_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5264_),
    .B(_5266_),
    .Y(_5267_)
);

OAI21X1 _12370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4618_),
    .B(_4431_),
    .C(_4362__bF$buf5),
    .Y(_4912_)
);

FILL FILL_0__12085_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .Y(_2738_)
);

NOR2X1 _9577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2374_),
    .B(_2378_),
    .Y(_2379_)
);

NAND3X1 _9157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1971_),
    .B(_1976_),
    .C(_1979_),
    .Y(_1980_)
);

FILL FILL_1__11825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6351_),
    .B(_6354_),
    .Y(_6355_)
);

MUX2X1 _13575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [5]),
    .B(\genblk1[7].u_ce.Xin12b [4]),
    .S(vdd),
    .Y(_5953_)
);

AOI22X1 _13155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5597_),
    .B(_5174__bF$buf4),
    .C(_5615_),
    .D(_5612_),
    .Y(_5048_)
);

FILL FILL_0__14651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10151_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .Y(_623_)
);

OR2X2 _7223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_219_),
    .Y(_222_)
);

FILL FILL_2__13370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11356_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11641_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3381_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [4])
);

OR2X2 _11221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3862_),
    .B(_3847_),
    .Y(_3863_)
);

DFFPOSX1 _8848_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_846_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Ycalc [7])
);

AND2X2 _8428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1328_),
    .B(_1311_),
    .Y(_1329_)
);

NOR2X1 _8008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_930_)
);

FILL FILL_1__7385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5311_),
    .B(_5316_),
    .C(_5319_),
    .Y(_5320_)
);

NOR2X1 _12426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4959_),
    .B(_4964_),
    .Y(_4965_)
);

NAND3X1 _12006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4565_),
    .C(_4562_),
    .Y(_4568_)
);

FILL FILL_0__13922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9111_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1092_)
);

FILL FILL_0__14707_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2179_),
    .B(_2198_),
    .C(_1848__bF$buf2),
    .Y(_2199_)
);

FILL FILL_1__11214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8641_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3565_),
    .B(_3566_),
    .Y(_3567_)
);

FILL FILL_0__8221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13099_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5819_)
);

FILL FILL_2__13846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9006_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(_6829_),
    .Y(_6830_)
);

DFFPOSX1 _14169_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5845_),
    .CLK(clk_bF$buf38),
    .Q(\genblk1[7].u_ce.Ycalc [9])
);

FILL FILL_0__10380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8802_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_822_)
);

NAND2X1 _7452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_433_),
    .Y(_441_)
);

NAND2X1 _10089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2825_),
    .Y(_2826_)
);

FILL FILL_1__12172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11585_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4423_),
    .B(_4434_),
    .C(_4437_),
    .Y(_4438_)
);

FILL FILL_0__11165_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4077_),
    .B(_4073_),
    .Y(_4078_)
);

NAND3X1 _11030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3679_),
    .C(_3675_),
    .Y(_3680_)
);

FILL FILL_2__11912_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1544_),
    .B(_1535_),
    .C(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_1545_)
);

NAND2X1 _8237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1145_),
    .Y(_1146_)
);

FILL FILL_1__7194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [6]),
    .B(_5108_),
    .Y(_5138_)
);

NOR2X1 _12235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4772_),
    .B(_4762_),
    .Y(_4787_)
);

FILL FILL_0__13731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9340_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6957_),
    .B(_7000_),
    .Y(_7018_)
);

FILL FILL_2__11089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7089_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_1903_),
    .C(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .Y(_2017_)
);

FILL FILL_1__11863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8450_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10721_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2547_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Acalc [8])
);

FILL FILL_0__8030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10016_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3008_),
    .B(_3023_),
    .C(_3021_),
    .Y(_3028_)
);

AOI21X1 _13193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5645_),
    .C(_5650_),
    .Y(_5651_)
);

DFFPOSX1 _7928_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ycalc [11])
);

OAI21X1 _7508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_473_),
    .C(_487_),
    .Y(_494_)
);

FILL FILL_1__12648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9655_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4489_),
    .Y(_4491_)
);

FILL FILL_0__9235_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4121_),
    .C(_4119_),
    .Y(_4130_)
);

NOR2X1 _14398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [6]),
    .B(\u_ot.Yin12b [7]),
    .Y(_6687_)
);

FILL FILL_1__8611_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

OAI21X1 _7261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_256_),
    .C(_257_),
    .Y(_258_)
);

FILL FILL_0__11394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11301_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8886_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_884_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Xin1 [1])
);

NAND3X1 _8466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(_1364_),
    .C(_1362_),
    .Y(_1365_)
);

NAND2X1 _8046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .B(_962_),
    .Y(\genblk1[1].u_ce.X_ [0])
);

FILL FILL_0__7721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5243_),
    .C(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .Y(_5357_)
);

FILL FILL_0__12179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Xin12b [9]),
    .Y(_4996_)
);

INVX1 _12044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4603_),
    .Y(_4604_)
);

FILL FILL_2__12926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8506_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6023_),
    .B(_6042_),
    .C(_6043_),
    .Y(_6044_)
);

NAND2X1 _13249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5703_),
    .B(_5696_),
    .Y(_5704_)
);

FILL FILL_0__14745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14325_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6841_),
    .B(_6840_),
    .C(_6838_),
    .Y(_6842_)
);

FILL FILL_2__7072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert384 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert385 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert386 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3603_),
    .B(_3584_),
    .C(_3512_),
    .Y(_3604_)
);

FILL FILL_2__8277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert387 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert388 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3243_),
    .B(_3234_),
    .Y(_3244_)
);

FILL FILL_0__10245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert389 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2836_),
    .B(_2842_),
    .C(_2845_),
    .Y(_2846_)
);

INVX1 _7737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [4]),
    .Y(_710_)
);

NAND2X1 _7317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_311_),
    .Y(_312_)
);

FILL FILL_1__12877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9464_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Xcalc [10]),
    .C(_4276_),
    .Y(_4309_)
);

FILL FILL_0__9044_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .B(_3947_),
    .C(_3943_),
    .Y(_3952_)
);

FILL FILL_0__12811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14603_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf2),
    .B(_433_),
    .Y(_477_)
);

FILL FILL_2__10589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11110_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1577_),
    .B(_1537_),
    .C(_1010__bF$buf5),
    .Y(_1580_)
);

INVX1 _8275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [8]),
    .Y(_1182_)
);

FILL FILL_1__10943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7548_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .Y(_6833__bF$buf3)
);

FILL FILL_0__7530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7110_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .Y(_6833__bF$buf2)
);

BUFX2 BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .Y(_6833__bF$buf1)
);

BUFX2 BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .Y(_6833__bF$buf0)
);

BUFX2 BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .Y(_973__bF$buf4)
);

BUFX2 BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .Y(_973__bF$buf3)
);

BUFX2 BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .Y(_973__bF$buf2)
);

BUFX2 BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .Y(_973__bF$buf1)
);

BUFX2 BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .Y(_973__bF$buf0)
);

OAI21X1 _12693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5148_),
    .B(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .C(_5173_),
    .Y(_5028_)
);

BUFX2 BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf4 )
);

OAI21X1 _12273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4822_),
    .B(_4821_),
    .C(_4809_),
    .Y(_4212_)
);

FILL FILL_2__12315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8315_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949__bF$buf3),
    .B(_6262_),
    .C(_6236_),
    .Y(_5849_)
);

DFFPOSX1 _13478_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5078_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [5])
);

AOI21X1 _13058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .B(_5522_),
    .C(_5196_),
    .Y(_5523_)
);

FILL FILL257250x226950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10054_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7966_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_50_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Yin12b [11])
);

NAND2X1 _7546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_530_),
    .Y(_531_)
);

AOI22X1 _7126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.Xcalc [5]),
    .C(_89_),
    .D(\genblk1[0].u_ce.Xcalc [7]),
    .Y(_129_)
);

FILL FILL_1__12686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9693_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4527_),
    .B(_4511_),
    .Y(_4528_)
);

FILL FILL_0__9273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4154_),
    .B(_4159_),
    .C(_4160_),
    .Y(_3393_)
);

INVX1 _11124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3769_),
    .Y(_3770_)
);

FILL FILL_0__12620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5150__bF$buf3),
    .Y(_5227_)
);

OAI21X1 _12329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4873_),
    .B(_4866_),
    .C(_4871_),
    .Y(_4874_)
);

FILL FILL_1__14832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9014_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(\genblk1[1].u_ce.Xin12b [6]),
    .S(vdd),
    .Y(_999_)
);

FILL FILL_1__10332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7777_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4361_),
    .C(_4639_),
    .Y(_4640_)
);

FILL FILL_2__12124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .B(_2104_),
    .C(_2105_),
    .D(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_2106_)
);

FILL FILL_1__11957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8544_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3473_),
    .C(_3474_),
    .Y(_3475_)
);

FILL FILL_0__8124_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5725_),
    .Y(_5740_)
);

FILL FILL_2__9503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8705_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_745_),
    .Y(_746_)
);

INVX1 _7355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_348_)
);

FILL FILL_1__12495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11488_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4344_),
    .C(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4345_)
);

FILL FILL_0__9082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11068_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3966_),
    .Y(_3988_)
);

FILL FILL_2__11815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7815_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .B(_2664_),
    .Y(_2665_)
);

OAI21X1 _9501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2308_),
    .B(_2307_),
    .C(_2295_),
    .Y(_1698_)
);

AOI22X1 _12978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .B(_5444_),
    .C(_5445_),
    .D(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5446_)
);

DFFPOSX1 _12558_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4212_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xcalc [9])
);

OAI21X1 _12138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4673_),
    .B(_4664_),
    .C(_4362__bF$buf1),
    .Y(_4694_)
);

FILL FILL_1__14641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6926_),
    .B(_6927_),
    .Y(_6928_)
);

FILL FILL_2__7586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12353_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1909_),
    .B(_1920_),
    .C(_1923_),
    .Y(_1924_)
);

FILL FILL_1__11766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8353_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3324_),
    .Y(_3325_)
);

FILL FILL_0__10339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2933_),
    .B(_2935_),
    .C(_2744_),
    .Y(_2936_)
);

NAND3X1 _13096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf3),
    .B(_5558_),
    .C(_5553_),
    .Y(_5559_)
);

FILL FILL_2__9732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9558_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(\genblk1[5].u_ce.Xin12b [8]),
    .S(vdd),
    .Y(_4398_)
);

FILL FILL_0__9138_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain1 [0]),
    .B(_4039_),
    .Y(_4040_)
);

FILL FILL_1__13912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8514_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_565_),
    .Y(_567_)
);

NAND2X1 _7164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(_164_),
    .Y(_165_)
);

FILL FILL_0__11297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.Y_ [0]),
    .Y(_4181_)
);

OAI21X1 _11162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3674_),
    .C(_3805_),
    .Y(_3806_)
);

FILL FILL_1__9719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1223_),
    .B(_1637_),
    .C(_1655_),
    .Y(_887_)
);

NAND2X1 _8369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1272_)
);

FILL FILL_1__10617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7204_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2503_)
);

OAI21X1 _9310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1847_),
    .C(_2125_),
    .Y(_2126_)
);

FILL FILL_1__13089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5249_),
    .B(_5260_),
    .C(_5263_),
    .Y(_5264_)
);

OAI21X1 _12367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4909_),
    .B(_4908_),
    .C(_4899_),
    .Y(_4219_)
);

FILL FILL_1__14450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14648_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14513_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6501_),
    .CLK(clk_bF$buf46),
    .Q(\u_ot.Ycalc [1])
);

FILL FILL_0__14228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8582_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _10853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_3510_)
);

FILL FILL_0__8162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10568_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .Y(_3154_)
);

FILL FILL_0__10148_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf3),
    .B(_2751_),
    .C(_2752_),
    .Y(_2753_)
);

FILL FILL_2__9541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9367_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11638_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3378_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [1])
);

INVX1 _11218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3859_),
    .Y(_3860_)
);

FILL FILL_1__13721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8323_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_384_),
    .Y(_10_)
);

FILL FILL_0__13919_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_4023_)
);

FILL FILL_1__9948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11853_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1471_),
    .B(_996__bF$buf2),
    .C(_1490_),
    .D(_994_),
    .Y(_861_)
);

AOI21X1 _8178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1070_),
    .C(_998_),
    .Y(_1090_)
);

FILL FILL_1__10846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7433_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12596_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4250_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin0 [1])
);

NAND2X1 _12176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf3),
    .B(_4649_),
    .Y(_4730_)
);

FILL FILL_2__12638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8638_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _10909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3563_),
    .B(_3514_),
    .C(_3562_),
    .D(_3506_),
    .Y(_3564_)
);

FILL FILL_0__8218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14457_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6963_)
);

FILL FILL_0__14037_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6620_),
    .B(_6619_),
    .C(_6562__bF$buf2),
    .Y(_6622_)
);

FILL FILL_2__12391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8391_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [0]),
    .B(_3313_),
    .Y(_3345_)
);

FILL FILL_0__10377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf1),
    .B(_2971_),
    .Y(_2972_)
);

FILL FILL_2__9350_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_820_)
);

AND2X2 _7449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_437_),
    .Y(_438_)
);

FILL FILL_2__13596_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.Y_ [0]),
    .Y(_1667_)
);

FILL FILL_1__12169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9596_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4424_),
    .Y(_4435_)
);

FILL FILL_0__9176_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(_3506_),
    .Y(_4075_)
);

NOR2X1 _11027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf4),
    .B(_3676_),
    .Y(_3677_)
);

FILL FILL_1__13950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8027_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10718_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2544_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Acalc [5])
);

FILL FILL_1__9090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14686_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14551_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [2]),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.LoadCtl [3])
);

FILL FILL_0__14266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [0]),
    .B(_6455_),
    .Y(_6473_)
);

FILL FILL_1__7823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11193_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3522_),
    .C(_3547_),
    .Y(_3548_)
);

FILL FILL_0__10186_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3188_),
    .B(_3186_),
    .Y(_3189_)
);

OAI21X1 _10051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .B(_2768_),
    .C(_2785_),
    .Y(_2789_)
);

FILL FILL_1__8608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10513_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf3),
    .B(_643_),
    .Y(_656_)
);

INVX1 _7258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_255_)
);

FILL FILL_1__12398_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11676_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3416_),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.Ain12b [9])
);

NOR2X1 _11256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3854_),
    .B(_3851_),
    .Y(_3896_)
);

FILL FILL_0__12752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7718_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9824_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1736_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Yin0 [1])
);

NAND2X1 _9404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf3),
    .B(_2135_),
    .Y(_2216_)
);

FILL FILL_1__8781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13957_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6165_),
    .B(_6167_),
    .C(_6161_),
    .Y(_6190_)
);

FILL FILL_0__13537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13117_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [0]),
    .B(_5796_),
    .Y(_5828_)
);

FILL FILL_1__9986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6839_)
);

FILL FILL_0__7891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8676_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3599_),
    .B(_3596_),
    .C(_3585_),
    .Y(_3601_)
);

FILL FILL_0__8256_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3235_),
    .B(_3239_),
    .Y(_3241_)
);

INVX1 _10107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .Y(_2843_)
);

FILL FILL_0__11603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14495_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [15]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf4),
    .Y(_6998_)
);

FILL FILL_0__14075_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6654_),
    .C(_6651_),
    .Y(_6655_)
);

FILL FILL_1__7632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12808_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3003_),
    .B(_2987_),
    .C(_3001_),
    .Y(_3008_)
);

FILL FILL_1__8837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_460_),
    .Y(_474_)
);

NAND2X1 _11485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4105_),
    .B(_4108_),
    .Y(_4111_)
);

OAI21X1 _11065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3699_),
    .B(_3712_),
    .C(_3713_),
    .Y(_3714_)
);

FILL FILL_2__7701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7527_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .B(_1848__bF$buf3),
    .Y(_2431_)
);

FILL FILL_0__7107_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .B(_2033_),
    .C(_2032_),
    .Y(_2034_)
);

FILL FILL_1__8590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13766_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6004_),
    .Y(_6007_)
);

FILL FILL_0__13346_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5649_),
    .B(_5174__bF$buf4),
    .C(_5668_),
    .D(_5172_),
    .Y(_5051_)
);

FILL FILL_1__9375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_7050_)
);

NAND2X1 _14416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(_6700_),
    .Y(_6703_)
);

FILL FILL_2_BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8065_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10756_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2582_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Ain12b [5])
);

AOI21X1 _10336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3057_),
    .B(_3061_),
    .C(_2690_),
    .Y(_3062_)
);

FILL FILL_2__9864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9024_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8904_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_902_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Ain12b [9])
);

FILL FILL_1__7861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .B(_5373_),
    .C(_5372_),
    .Y(_5374_)
);

FILL FILL_0__12617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_275_),
    .C(_227_),
    .Y(_292_)
);

OAI21X1 _11294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3907_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_3932_),
    .Y(_3371_)
);

FILL FILL_2__7510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7756_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [5]),
    .Y(_2611_)
);

FILL FILL_0__7336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2251_),
    .C(_2252_),
    .Y(_2253_)
);

OAI21X1 _9022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1849_),
    .C(_1850_),
    .Y(_1851_)
);

OAI21X1 _12499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4445_),
    .B(_5000_),
    .C(_5015_),
    .Y(_4245_)
);

NAND2X1 _12079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4637_)
);

FILL FILL_2__8715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13575_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6046_),
    .C(_6225_),
    .Y(_6226_)
);

FILL FILL_0__13155_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13440_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5040_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [11])
);

AOI21X1 _13020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .B(_5485_),
    .C(_5176_),
    .Y(_5487_)
);

FILL FILL_1__9184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6873_),
    .B(_6870_),
    .Y(_6874_)
);

INVX1 _14225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [3]),
    .Y(_6543_)
);

FILL FILL_2__12294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11287_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3634_),
    .Y(_3637_)
);

FILL FILL_0__8294_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3265_),
    .B(_2672__bF$buf1),
    .C(_3275_),
    .D(_3276_),
    .Y(_2546_)
);

AND2X2 _10145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2818_),
    .B(_2821_),
    .Y(_2879_)
);

FILL FILL_2__9253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .Y(_1597_)
);

FILL FILL_1__7670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12846_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5189_),
    .C(_5190_),
    .Y(_5191_)
);

FILL FILL_0__12426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12006_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2660_),
    .C(_2661_),
    .Y(_2662_)
);

FILL FILL_1__8455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14218_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6275_),
    .B(_6277_),
    .C(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_6280_)
);

FILL FILL_2__11565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7565_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2465_),
    .Y(_2466_)
);

FILL FILL_0__7145_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .Y(_2070_)
);

FILL FILL_0__10912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9729_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14874_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6765_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [5])
);

FILL FILL_0__14589_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6727_),
    .B(_6733_),
    .C(_6734_),
    .Y(_6516_)
);

NOR2X1 _14034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6358_),
    .B(_6386_),
    .Y(_6392_)
);

FILL FILL_1__7726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_3454_),
    .C(_3455_),
    .Y(_3456_)
);

FILL FILL_0__10089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf1),
    .B(_2925_),
    .Y(_3098_)
);

FILL FILL_2__10836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11030_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.Acalc [1]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Acalc [3]),
    .Y(_1777_)
);

OAI21X1 _8522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1393_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1418_),
    .Y(_857_)
);

MUX2X1 _8102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1016_),
    .B(_1013_),
    .S(_973__bF$buf4),
    .Y(_1017_)
);

NOR3X1 _11999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4517_),
    .B(_4540_),
    .C(_4513_),
    .Y(_4561_)
);

OAI21X1 _11579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4171_),
    .B(_3435_),
    .C(_4179_),
    .Y(_3409_)
);

MUX2X1 _11159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .B(_3800_),
    .S(_3487__bF$buf2),
    .Y(_3803_)
);

FILL FILL_1__13662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12655_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5404_),
    .Y(_5410_)
);

FILL FILL_0__12235_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [6]),
    .B(_4997_),
    .Y(_5027_)
);

AND2X2 _12100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4656_),
    .B(_4657_),
    .Y(_4658_)
);

OAI21X1 _9727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1931_),
    .B(_2486_),
    .C(_2501_),
    .Y(_1731_)
);

NAND2X1 _9307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_2123_)
);

FILL FILL_1__8684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14027_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6090_),
    .B(_6093_),
    .Y(_6097_)
);

NAND2X1 _13305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf4),
    .B(_5683_),
    .Y(_5758_)
);

FILL FILL_0__14801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x100950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2283_),
    .B(_2285_),
    .Y(_2289_)
);

NAND2X1 _9060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1810__bF$buf0),
    .Y(_1887_)
);

FILL FILL_2__8753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6907_),
    .B(_6906_),
    .Y(_6908_)
);

INVX1 _14263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin1 [0]),
    .Y(_6570_)
);

FILL FILL_1__7535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13718_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2915_),
    .B(_2914_),
    .C(_2912_),
    .Y(_2916_)
);

FILL FILL_2__10225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1626_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1632_)
);

NAND2X1 _8331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1231_),
    .B(_1235_),
    .Y(_1236_)
);

OAI21X1 _11388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510__bF$buf2),
    .B(_4019_),
    .C(_4020_),
    .Y(_3377_)
);

FILL FILL_1__13891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12044_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2697_),
    .C(_2698_),
    .Y(_2699_)
);

NOR2X1 _9536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(_2338_),
    .Y(_2341_)
);

OR2X2 _9116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1940_),
    .B(_1939_),
    .Y(_1941_)
);

FILL FILL_1__8493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6294_),
    .B(_6313_),
    .Y(_6316_)
);

FILL FILL_0__13669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13249_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5911_),
    .B(_5914_),
    .C(_5892_),
    .Y(_5915_)
);

NAND3X1 _13114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf3),
    .B(_5575_),
    .C(_5572_),
    .Y(_5576_)
);

FILL FILL_0_BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10176_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6959_),
    .B(_6939_),
    .C(_6948_),
    .Y(_6960_)
);

INVX1 _14319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [9]),
    .Y(_6619_)
);

FILL FILL_0__7183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10110_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf0),
    .B(_411_),
    .Y(_584_)
);

FILL FILL_0__8388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_2647_),
    .C(_3343_),
    .Y(_2573_)
);

INVX1 _10239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2968_),
    .Y(_2969_)
);

FILL FILL_1__12742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11315_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [0]),
    .B(_4162_),
    .Y(_3426_)
);

OAI21X1 _14492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Yin1 [1]),
    .Y(_6756_)
);

NAND3X1 _14072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6418_),
    .B(_6420_),
    .C(_6427_),
    .Y(_6428_)
);

OAI21X1 _8807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_921_),
    .C(_1665_),
    .Y(_895_)
);

FILL FILL_1__7764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13107_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5280_),
    .B(_5279_),
    .Y(_5281_)
);

FILL FILL_1__8969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9910_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_199_),
    .Y(_200_)
);

INVX8 _8980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_1810_)
);

OR2X2 _8560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1452_),
    .Y(_1455_)
);

NAND2X1 _8140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .B(_1052_),
    .Y(_1053_)
);

INVX1 _11197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3839_),
    .Y(_3840_)
);

FILL FILL_1__13280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7659_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9765_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1677_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Ycalc [1])
);

FILL FILL_0__7239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf2),
    .B(_2159_),
    .C(_2150_),
    .Y(_2160_)
);

FILL FILL_0__8600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13898_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6131_),
    .B(_6129_),
    .C(_6133_),
    .Y(_6134_)
);

FILL FILL_0__13058_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174__bF$buf0),
    .B(_5793_),
    .C(_5792_),
    .Y(_5058_)
);

FILL FILL257250x176550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9087_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14548_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.Vld ),
    .CLK(clk_bF$buf38),
    .Q(\u_ot.LoadCtl [0])
);

OAI21X1 _14128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5937_),
    .C(_6471_),
    .Y(_5870_)
);

FILL FILL_2__8791_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158__bF$buf2),
    .B(_796_),
    .C(_795_),
    .Y(_36_)
);

AOI21X1 _7411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_400_),
    .C(_398_),
    .Y(_402_)
);

MUX2X1 _10888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(\genblk1[4].u_ce.Xin0 [1]),
    .S(gnd),
    .Y(_3545_)
);

FILL FILL_0__8197_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(gnd),
    .C(_3185_),
    .Y(_3186_)
);

AOI21X1 _10048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2786_),
    .C(_2674_),
    .Y(_2787_)
);

FILL FILL_1__12971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11124_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996__bF$buf2),
    .B(_1505_),
    .C(_1506_),
    .Y(_863_)
);

FILL FILL_1__7573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12329_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12614_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.LoadCtl [5])
);

FILL FILL_1__8778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10263_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6185_),
    .B(_6186_),
    .Y(_6187_)
);

FILL FILL_2__7222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7888_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2734_),
    .Y(_2735_)
);

FILL FILL_0__7468_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf1),
    .B(_2375_),
    .C(_1848__bF$buf3),
    .Y(_2376_)
);

INVX1 _9154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .Y(_1977_)
);

FILL FILL_1__11822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14294_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6311_),
    .B(_6332_),
    .C(_6336_),
    .Y(_6352_)
);

NAND2X1 _13572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [1]),
    .B(_5949__bF$buf1),
    .Y(_5950_)
);

FILL FILL_0__13287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5598_),
    .B(_5588_),
    .Y(_5613_)
);

FILL FILL_0__9614_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6991_),
    .Y(_6995_)
);

OAI21X1 _14357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .C(\u_ot.ISreg_bF$buf2 ),
    .Y(_6652_)
);

FILL FILL_1__7629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_602_),
    .Y(_620_)
);

AOI21X1 _7220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_215_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_219_)
);

DFFPOSX1 _10697_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2523_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [8])
);

NOR2X1 _10277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2987_),
    .B(_3004_),
    .Y(_3006_)
);

FILL FILL_1__12780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11353_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8845_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_843_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Ycalc [4])
);

INVX1 _8425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1325_),
    .Y(_1326_)
);

AND2X2 _8005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(\genblk1[1].u_ce.LoadCtl [3]),
    .Y(_927_)
);

FILL FILL_1__7382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12978_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5317_)
);

FILL FILL_0__12138_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4961_),
    .B(_4926_),
    .C(_4960_),
    .Y(_4962_)
);

INVX1 _12003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4563_),
    .Y(_4565_)
);

FILL FILL_1__8587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6000_),
    .C(_6003_),
    .Y(_6004_)
);

AND2X2 _13208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5654_),
    .B(_5665_),
    .Y(_5666_)
);

FILL FILL_0__14704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2112_),
    .C(_2195_),
    .Y(_2196_)
);

FILL FILL_2_BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13096_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5817_)
);

FILL FILL_2__13003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9003_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [18]),
    .B(\u_pa.acc_reg [19]),
    .Y(_6827_)
);

DFFPOSX1 _14166_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5842_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[7].u_ce.Ycalc [6])
);

FILL FILL_1__7858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .B(_2781_),
    .C(_2769_),
    .Y(_2823_)
);

FILL FILL_0__11582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1540_),
    .Y(_1542_)
);

NAND3X1 _8234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf2),
    .B(_1139_),
    .C(_1134_),
    .Y(_1143_)
);

FILL FILL_1__7191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12787_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Xcalc [10]),
    .C(_5106_),
    .Y(_5135_)
);

FILL FILL_0__12367_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4363_),
    .B(_4782_),
    .C(_4783_),
    .Y(_4784_)
);

INVX1 _9859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [9]),
    .Y(_2608_)
);

AND2X2 _9439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2203_),
    .B(_2206_),
    .Y(_2250_)
);

INVX8 _9019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_1848_)
);

FILL FILL_1__8396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14579_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [7]),
    .Y(_6223_)
);

DFFPOSX1 _13437_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5037_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [8])
);

AND2X2 _13017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .B(_5483_),
    .Y(_5484_)
);

FILL FILL_2__7260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7086_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2013_),
    .B(_1997_),
    .Y(_2014_)
);

FILL FILL_1__11860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10013_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .B(_5647_),
    .C(_5635_),
    .Y(_5050_)
);

DFFPOSX1 _7925_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[0].u_ce.Ycalc [8])
);

NOR2X1 _7505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_490_),
    .Y(_492_)
);

FILL FILL256950x111750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9652_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf1),
    .B(_4399_),
    .Y(_4488_)
);

FILL FILL_0__9232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4121_),
    .B(_4126_),
    .Y(_4128_)
);

NAND3X1 _14395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6681_),
    .C(_6684_),
    .Y(_6685_)
);

FILL FILL_1__7667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14437_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _12708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_5188_)
);

FILL FILL_2__10777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11391_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8883_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_881_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[1].u_ce.Xin12b [4])
);

OR2X2 _8463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1359_),
    .Y(_1362_)
);

OAI21X1 _8043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(_959_),
    .C(_960_),
    .Y(_961_)
);

FILL FILL_1__13183_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5353_),
    .B(_5337_),
    .Y(_5354_)
);

FILL FILL_0__12176_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4994_)
);

INVX1 _12041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4601_)
);

FILL FILL_2__12503_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2463_)
);

NAND2X1 _9248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2062_),
    .Y(_2067_)
);

FILL FILL_1__11916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6041_)
);

OR2X2 _13246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5699_),
    .B(\genblk1[6].u_ce.Ain1 [0]),
    .Y(_5701_)
);

FILL FILL_2__13708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(_706_),
    .C(_707_),
    .Y(_708_)
);

AOI21X1 _7314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_267_),
    .C(_255_),
    .Y(_309_)
);

FILL FILL_2__13041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11447_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.Ycalc [1]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4307_)
);

FILL FILL_0__9041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11027_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947_),
    .Y(_3950_)
);

NAND2X1 _8939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [7]),
    .B(_1765_),
    .Y(_1774_)
);

NOR2X1 _8519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1411_),
    .B(_1415_),
    .Y(_1416_)
);

FILL FILL_1__7896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5402_),
    .Y(_5407_)
);

INVX1 _12517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [1]),
    .Y(_5025_)
);

FILL FILL_1__14600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9202_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1002_),
    .C(_972__bF$buf1),
    .Y(_1577_)
);

INVX1 _8272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .Y(_1180_)
);

FILL FILL_1__10940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10100_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .Y(_1810__bF$buf4)
);

BUFX2 BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .Y(_1810__bF$buf3)
);

BUFX2 BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .Y(_1810__bF$buf2)
);

BUFX2 BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .Y(_1810__bF$buf1)
);

BUFX2 BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .Y(_1810__bF$buf0)
);

BUFX2 BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf0 )
);

OAI21X1 _12690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5170_),
    .C(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .Y(_5171_)
);

BUFX2 BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925_),
    .Y(_5925__bF$buf3)
);

NAND2X1 _12270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4817_),
    .B(_4819_),
    .Y(_4820_)
);

FILL FILL_2_CLKBUF1_insert391 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(\genblk1[3].u_ce.Xcalc [9]),
    .C(_2600_),
    .Y(_2642_)
);

NAND2X1 _9477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2282_),
    .B(_2285_),
    .Y(_2286_)
);

MUX2X1 _9057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(\genblk1[2].u_ce.Xin12b [8]),
    .S(gnd),
    .Y(_1884_)
);

FILL FILL_1__11725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8312_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6237_),
    .B(_6259_),
    .Y(_6260_)
);

DFFPOSX1 _13475_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5075_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin12b [6])
);

OAI21X1 _13055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499_),
    .B(_5490_),
    .C(_5188__bF$buf3),
    .Y(_5520_)
);

FILL FILL_2__13937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x108150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10051_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7963_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_47_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin0 [0])
);

OR2X2 _7543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_520_),
    .Y(_528_)
);

INVX1 _7123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [3]),
    .Y(_126_)
);

FILL FILL_2__13270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9690_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(_4523_),
    .C(_4524_),
    .Y(_4525_)
);

FILL FILL_2__9288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11256_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4157_),
    .B(_4155_),
    .C(_4158_),
    .Y(_3392_)
);

NAND2X1 _11121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3766_),
    .B(_3742_),
    .Y(_3767_)
);

NAND2X1 _8748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .B(_1010__bF$buf5),
    .Y(_1629_)
);

AND2X2 _8328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1227_),
    .B(_1010__bF$buf3),
    .Y(_1233_)
);

FILL FILL_1__7285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13048_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(\genblk1[6].u_ce.Xin12b [8]),
    .S(gnd),
    .Y(_5224_)
);

NAND2X1 _12326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .B(_4871_),
    .Y(_4872_)
);

FILL FILL_0__13822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9011_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _8081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_996_)
);

FILL FILL_0__14607_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2102_),
    .Y(_2103_)
);

FILL FILL_1__11954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert384 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert385 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert386 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert387 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert388 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert389 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3470_),
    .C(_3471_),
    .Y(_3472_)
);

FILL FILL_0__8121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10107_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5736_),
    .B(_5727_),
    .Y(_5738_)
);

FILL FILL_2__9500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6749_),
    .B(_6737_),
    .C(_6754_),
    .Y(_6531_)
);

INVX1 _14069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6418_),
    .Y(_6425_)
);

FILL FILL_0__10280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8702_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_741_),
    .Y(_743_)
);

OAI21X1 _7352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_336_),
    .C(_335_),
    .Y(_345_)
);

FILL FILL_1__12492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11485_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4323_),
    .B(_4340_),
    .Y(_4342_)
);

FILL FILL_0__11065_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [10]),
    .Y(_3985_)
);

FILL FILL_1__9907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11812_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1759_),
    .C(_1807_),
    .Y(\genblk1[2].u_ce.X_ [1])
);

AOI21X1 _8557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1451_),
    .B(_1450_),
    .C(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1452_)
);

OAI22X1 _8137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1049_),
    .B(_1000_),
    .C(_1048_),
    .D(_992_),
    .Y(_1050_)
);

FILL FILL_1__7094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5442_),
    .Y(_5443_)
);

DFFPOSX1 _12555_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4209_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[5].u_ce.Xcalc [6])
);

NAND2X1 _12135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4647_),
    .B(_4430_),
    .Y(_4691_)
);

FILL FILL_0__13631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6925_)
);

INVX1 _9095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .Y(_1921_)
);

FILL FILL_1__11763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8350_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(_3321_),
    .Y(_3323_)
);

FILL FILL_0__10336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _10201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2923_),
    .B(_2932_),
    .C(_2916_),
    .Y(_2933_)
);

NAND2X1 _13093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf1),
    .B(_5475_),
    .Y(_5556_)
);

OAI21X1 _7828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_794_),
    .B(_793_),
    .C(_784_),
    .Y(_35_)
);

AOI21X1 _7408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_374_),
    .B(_376_),
    .C(_370_),
    .Y(_399_)
);

FILL FILL_2__13975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9555_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(_4394_),
    .C(_4395_),
    .Y(_4192_)
);

FILL FILL_0__9135_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3516_),
    .B(_3487__bF$buf4),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4037_)
);

FILL FILL256050x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6597_),
    .B(_6600_),
    .Y(_6601_)
);

FILL FILL_0__12902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8511_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_563_),
    .Y(_564_)
);

MUX2X1 _7161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .B(\genblk1[0].u_ce.Xin12b [4]),
    .S(gnd),
    .Y(_162_)
);

FILL FILL_0__11294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11201_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.X_ [1]),
    .Y(_1654_)
);

NAND3X1 _8366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf2),
    .B(_1265_),
    .C(_1268_),
    .Y(_1269_)
);

FILL FILL_1__10614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13086_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5250_),
    .Y(_5261_)
);

FILL FILL_0__12499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12079_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4886_),
    .B(_4894_),
    .C(_4893_),
    .Y(_4907_)
);

FILL FILL_2__12826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6348_),
    .Y(_6349_)
);

OAI21X1 _13569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5942_),
    .B(_5944_),
    .C(_5947_),
    .Y(_5948_)
);

NAND3X1 _13149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5189_),
    .B(_5608_),
    .C(_5609_),
    .Y(_5610_)
);

FILL FILL_0__14645_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14510_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6498_),
    .CLK(clk_bF$buf4),
    .Q(\u_ot.Xcalc [10])
);

FILL FILL_0__14225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10985_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3507_),
    .Y(_3508_)
);

FILL FILL_0__10565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10145_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3141_),
    .B(_3143_),
    .C(_3150_),
    .Y(_3151_)
);

NAND2X1 _10010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2750_)
);

OAI21X1 _7637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_602_),
    .C(_156_),
    .Y(_618_)
);

INVX1 _7217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .Y(_216_)
);

FILL FILL_2__13784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x226950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9364_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11635_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3375_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xcalc [10])
);

OR2X2 _11215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3856_),
    .B(_3855_),
    .Y(_3857_)
);

FILL FILL_0__12711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8320_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_381_),
    .Y(_382_)
);

FILL FILL_0__13916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11010_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_1487_),
    .Y(_1488_)
);

AOI21X1 _8175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_1082_),
    .C(_1071_),
    .Y(_1087_)
);

FILL FILL_1__10843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7448_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12593_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4247_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin1 [0])
);

NAND2X1 _12173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4711_),
    .B(_4715_),
    .Y(_4727_)
);

FILL FILL_2__12215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8635_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3560_),
    .B(_3513_),
    .S(gnd),
    .Y(_3561_)
);

FILL FILL_0__8215_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6162_),
    .C(_6166_),
    .Y(_6167_)
);

NAND2X1 _13378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5796_),
    .Y(_5815_)
);

FILL FILL_0__14454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10374_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_799_),
    .Y(_818_)
);

OAI21X1 _7446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_255_),
    .C(_434_),
    .Y(_435_)
);

FILL FILL_1__12166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11579_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4372_),
    .B(_4431_),
    .C(_4430_),
    .D(_4368_),
    .Y(_4432_)
);

FILL FILL_0__9173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11159_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4068_),
    .B(_4069_),
    .C(_4066_),
    .Y(_4072_)
);

INVX1 _11024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3674_)
);

FILL FILL_0__12940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7906_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Ycalc [1]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5133_)
);

NAND3X1 _12229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(_4777_),
    .C(_4780_),
    .Y(_4781_)
);

FILL FILL_1__14732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(_2009_),
    .C(_2010_),
    .Y(_2011_)
);

FILL FILL_1__11857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8024_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10715_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2541_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[3].u_ce.Acalc [2])
);

NAND2X1 _13187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5643_),
    .B(_5645_),
    .Y(_5646_)
);

FILL FILL_2__9403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8605_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [11]),
    .B(_158__bF$buf0),
    .Y(_653_)
);

OAI21X1 _7255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_251_),
    .C(_252_),
    .Y(_253_)
);

FILL FILL_1__12395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11388_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11673_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3413_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[4].u_ce.Ain12b [10])
);

OAI21X1 _11253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf2),
    .B(_3891_),
    .C(_3892_),
    .Y(_3893_)
);

FILL FILL_0__7715_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9821_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1733_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Yin1 [0])
);

NAND2X1 _9401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2201_),
    .Y(_2213_)
);

NAND3X1 _12878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(_5349_),
    .C(_5350_),
    .Y(_5351_)
);

OAI21X1 _12458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4514_),
    .B(_4989_),
    .C(_4991_),
    .Y(_4228_)
);

NAND2X1 _12038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [11]),
    .B(_4348__bF$buf4),
    .Y(_4598_)
);

FILL FILL257250x212550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6835_),
    .B(_6836_),
    .C(En_bF$buf0),
    .Y(_6837_)
);

FILL FILL_2__7486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8673_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .Y(_3598_)
);

FILL FILL_0__8253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10659_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3237_),
    .B(_2686__bF$buf0),
    .Y(_3238_)
);

FILL FILL_0__10239_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2839_),
    .Y(_2840_)
);

FILL FILL_0__11600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [7]),
    .B(_4279_),
    .Y(_4304_)
);

FILL FILL_0__9038_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3943_),
    .B(_3946_),
    .Y(_3947_)
);

FILL FILL_1__13812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8414_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158__bF$buf3),
    .B(_471_),
    .C(_445_),
    .Y(_14_)
);

FILL FILL_0__11197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_4107_),
    .Y(_4108_)
);

AND2X2 _11062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3707_),
    .B(_3710_),
    .Y(_3711_)
);

FILL FILL_1__9619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_1566_),
    .C(_1564_),
    .Y(_1574_)
);

OAI21X1 _8269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1150_),
    .C(_1145_),
    .Y(_1177_)
);

FILL FILL_1__10937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7524_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .B(_2425_),
    .Y(_2428_)
);

FILL FILL_0__7104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .B(_2030_),
    .C(_2027_),
    .Y(_2031_)
);

NAND2X1 _12687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5149_),
    .B(_5166_),
    .Y(_5168_)
);

NAND3X1 _12267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(_4815_),
    .C(_4816_),
    .Y(_4817_)
);

FILL FILL_1__14770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10270_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [19]),
    .B(En_bF$buf3),
    .Y(_7047_)
);

FILL FILL_0__14128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6699_),
    .B(_6666_),
    .C(_6698_),
    .Y(_6700_)
);

FILL FILL_2__12482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10468_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10753_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2579_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Ain12b [6])
);

FILL FILL_0__10048_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .B(_3058_),
    .C(_2999_),
    .Y(_3059_)
);

FILL FILL_2__9441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13267_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8901_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_899_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[1].u_ce.Ain12b [10])
);

FILL FILL_0__9687_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4512_),
    .B(_4518_),
    .C(_4521_),
    .Y(_4522_)
);

FILL FILL_0__9267_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4154_),
    .B(_4155_),
    .C(_4156_),
    .Y(_3391_)
);

NAND2X1 _11118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .B(_3763_),
    .Y(_3764_)
);

FILL FILL_1__13621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14406_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .Y(_289_)
);

FILL FILL_0__13819_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3925_),
    .B(_3929_),
    .Y(_3930_)
);

FILL FILL_1__9848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11753_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf0),
    .B(_1354_),
    .C(_1376_),
    .Y(_1395_)
);

INVX2 _8078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .Y(_994_)
);

FILL FILL_1__10326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7333_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(_4997_),
    .Y(_5014_)
);

OAI21X1 _12076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4634_),
    .B(_4629_),
    .C(_4613_),
    .Y(_4203_)
);

FILL FILL_0__13992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8538_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3469_),
    .B(_3468_),
    .Y(\genblk1[4].u_ce.Y_ [1])
);

FILL FILL_0__8118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6866_),
    .B(_6864_),
    .Y(_6871_)
);

INVX1 _14222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [2]),
    .Y(_6541_)
);

FILL FILL_1__7914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11284_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf4),
    .B(_3632_),
    .C(_3633_),
    .Y(_3634_)
);

FILL FILL_0__8291_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3273_),
    .B(_3272_),
    .Y(_3274_)
);

FILL FILL_0__10277_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2858_),
    .B(_2672__bF$buf0),
    .C(_2876_),
    .D(_2856_),
    .Y(_2523_)
);

FILL FILL_2__9670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9250_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_699_),
    .Y(_740_)
);

OAI21X1 _7349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_338_),
    .C(_342_),
    .Y(_343_)
);

NAND2X1 _8710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1593_),
    .Y(_1594_)
);

FILL FILL_1__12489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9496_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4338_),
    .B(_4335_),
    .S(_4325__bF$buf3),
    .Y(_4339_)
);

FILL FILL_0__9076_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3973_),
    .B(_3982_),
    .Y(_3983_)
);

FILL FILL_1__13850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2657_),
    .C(_2658_),
    .Y(_2659_)
);

FILL FILL_1__8452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14635_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_6276_),
    .C(_6273_),
    .Y(_6277_)
);

FILL FILL_0__13628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(_2603_),
    .Y(_3321_)
);

FILL FILL_1__12701_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14871_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6762_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [2])
);

FILL FILL_0__14586_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6731_),
    .B(_6729_),
    .C(_6732_),
    .Y(_6515_)
);

AOI21X1 _14031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6388_),
    .B(_6389_),
    .C(_5946_),
    .Y(_6390_)
);

FILL FILL_1__7723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11093_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3453_),
    .B(_3452_),
    .Y(\a[5] [1])
);

FILL FILL_0__10086_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [7]),
    .Y(_3095_)
);

FILL FILL_1__8928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_919_),
    .Y(_920_)
);

NOR3X1 _7578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_541_),
    .C(_545_),
    .Y(_561_)
);

NAND2X1 _7158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [1]),
    .B(_158__bF$buf2),
    .Y(_159_)
);

FILL FILL_1__12298_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4548_),
    .Y(_4558_)
);

NAND2X1 _11576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4162_),
    .Y(_4178_)
);

OAI21X1 _11156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3585_),
    .C(_3799_),
    .Y(_3800_)
);

FILL FILL_0__12652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x90150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(_2483_),
    .Y(_2500_)
);

OAI21X1 _9304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2120_),
    .B(_2115_),
    .C(_2099_),
    .Y(_1689_)
);

FILL FILL_1__8681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13857_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6092_),
    .B(_6093_),
    .Y(_6094_)
);

FILL FILL_0__13017_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [7]),
    .Y(_5755_)
);

FILL FILL_1__9886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10364_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14507_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6495_),
    .CLK(clk_bF$buf9),
    .Q(\u_ot.Xcalc [7])
);

FILL FILL_0__7791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8576_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3504_),
    .Y(_3505_)
);

FILL FILL_0__8156_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3141_),
    .Y(_3148_)
);

INVX1 _10007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2747_)
);

FILL FILL_1__12930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14395_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6872_),
    .B(_6879_),
    .Y(_6905_)
);

NAND2X1 _14260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6564_),
    .B(_6567_),
    .Y(_6568_)
);

FILL FILL_1__7532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12708_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2888_),
    .B(_2890_),
    .C(_2884_),
    .Y(_2913_)
);

FILL FILL_1__8737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10222_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_371_),
    .C(_373_),
    .Y(_379_)
);

NAND2X1 _11385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4016_),
    .B(_4017_),
    .Y(_4018_)
);

FILL FILL_2__7601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7847_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2694_),
    .C(_2695_),
    .Y(_2696_)
);

FILL FILL_0__7427_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1811__bF$buf0),
    .C(_1830_),
    .Y(_2338_)
);

OAI21X1 _9113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf4),
    .B(_1936_),
    .C(_1937_),
    .Y(_1938_)
);

FILL FILL_1__8490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13666_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .B(_6234_),
    .C(_6251_),
    .Y(_6313_)
);

FILL FILL_0_BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13246_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [4]),
    .Y(_5912_)
);

FILL FILL_0_BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5532_),
    .C(_5554_),
    .Y(_5573_)
);

FILL FILL_0_BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10173_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6941_),
    .B(_6950_),
    .C(_6956_),
    .Y(_6957_)
);

NAND2X1 _14316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [8]),
    .B(_6562__bF$buf0),
    .Y(_6617_)
);

FILL FILL_2_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8385_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_3342_)
);

NAND2X1 _10236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf0),
    .B(_2965_),
    .Y(_2966_)
);

FILL FILL_0__11732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11312_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1648_),
    .Y(_1664_)
);

FILL FILL_1__7761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12937_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf2),
    .B(_5276_),
    .C(_5277_),
    .Y(_5278_)
);

FILL FILL_0__12517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14309_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_188_),
    .C(_171_),
    .Y(_197_)
);

AOI21X1 _11194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_3789_),
    .C(_3815_),
    .Y(_3837_)
);

FILL FILL_2__7830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7656_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[2] [1]),
    .Y(_1755_)
);

FILL FILL_0__7236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2155_),
    .B(_2156_),
    .Y(_2157_)
);

NAND2X1 _12399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(_4939_),
    .Y(_4940_)
);

FILL FILL_2__8615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13895_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6127_),
    .B(_6130_),
    .C(_6018_),
    .Y(_6131_)
);

FILL FILL_0__13055_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5789_),
    .B(_5790_),
    .Y(_5791_)
);

FILL FILL_1__9084_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14545_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6533_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Yin1 [1])
);

OAI21X1 _14125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_6470_)
);

FILL FILL_1__7817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11187_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .S(gnd),
    .Y(_3542_)
);

FILL FILL_0__8194_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [1]),
    .B(_2672__bF$buf1),
    .Y(_3183_)
);

AND2X2 _10045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2778_),
    .B(_2777_),
    .Y(_2784_)
);

FILL FILL_2__10927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11121_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1502_),
    .B(_1503_),
    .Y(_1504_)
);

FILL FILL_1__7570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12326_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12611_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.LoadCtl [2])
);

DFFPOSX1 _9818_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1730_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Yin12b [7])
);

FILL FILL_1__8775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14118_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6176_),
    .B(_6183_),
    .Y(_6184_)
);

FILL FILL_2__11465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7885_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2730_),
    .B(_2731_),
    .Y(_2732_)
);

FILL FILL_0__7465_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .Y(_2373_)
);

NAND2X1 _9151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf4),
    .B(_1885_),
    .Y(_1974_)
);

FILL FILL_0__10812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14489_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6991_),
    .B(_6990_),
    .Y(_6992_)
);

FILL FILL_0__14069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6646_),
    .C(_6649_),
    .Y(_6650_)
);

FILL FILL_1__7626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13809_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10694_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2520_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [5])
);

AOI21X1 _10274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2998_),
    .B(_3000_),
    .C(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_3003_)
);

FILL FILL_0__11770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11350_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8842_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_840_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[1].u_ce.ISout )
);

AOI21X1 _8422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(_1275_),
    .C(_1301_),
    .Y(_1323_)
);

NOR2X1 _8002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.LoadCtl [3]),
    .Y(_924_)
);

OAI21X1 _11899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4462_),
    .B(_4444_),
    .C(_4461_),
    .Y(_4465_)
);

INVX1 _11479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .Y(_4105_)
);

NAND3X1 _11059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3705_),
    .C(_3701_),
    .Y(_3708_)
);

FILL FILL_1__13982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12975_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf2),
    .B(_5225_),
    .Y(_5314_)
);

NOR2X1 _12420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4958_),
    .B(_4957_),
    .Y(_4959_)
);

FILL FILL_0__12135_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4561_),
    .Y(_4562_)
);

NAND2X1 _9627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_2425_),
    .Y(_2426_)
);

NOR2X1 _9207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_1999_),
    .Y(_2028_)
);

FILL FILL_1__8584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14347_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [1]),
    .B(\genblk1[7].u_ce.Xin1 [0]),
    .S(vdd),
    .Y(_6001_)
);

NOR2X1 _13205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5656_),
    .B(_5658_),
    .Y(_5663_)
);

FILL FILL_0__14701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7274_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2192_),
    .Y(_2193_)
);

FILL FILL_2_BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [0]),
    .B(\u_pa.Atmp [1]),
    .Y(_6825_)
);

DFFPOSX1 _14163_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5839_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[7].u_ce.Ycalc [3])
);

FILL FILL_1__7855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .B(_2816_),
    .Y(_2820_)
);

FILL FILL_2__10965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9191_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1539_)
);

OAI21X1 _8231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1120_),
    .B(_1115_),
    .C(_1010__bF$buf2),
    .Y(_1140_)
);

NAND3X1 _11288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .B(_3926_),
    .C(_3901_),
    .Y(_3927_)
);

FILL FILL_1__13791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12364_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2606_)
);

NAND2X1 _9436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2246_),
    .Y(_2247_)
);

NAND3X1 _9016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf1),
    .B(_1844_),
    .C(_1843_),
    .Y(_1845_)
);

FILL FILL_1__8393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13989_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5955_),
    .Y(_6220_)
);

FILL FILL_0__13569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13149_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13434_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5034_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [5])
);

AOI21X1 _13014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5477_),
    .B(_5480_),
    .C(_5199_),
    .Y(_5481_)
);

FILL FILL_1__9598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10076_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6868_)
);

INVX1 _14219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [1]),
    .Y(_6539_)
);

FILL FILL_0__7083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10010_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7922_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ycalc [5])
);

AOI21X1 _7502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_486_),
    .C(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_489_)
);

INVX1 _10979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3630_),
    .Y(_3631_)
);

FILL FILL_0__8288_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .B(_3270_),
    .Y(_3271_)
);

INVX1 _10139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2873_),
    .Y(_2874_)
);

FILL FILL_1__12642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x176550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9667_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4485_)
);

FILL FILL_0__11215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4086_),
    .B(_4081_),
    .C(_4123_),
    .Y(_4125_)
);

INVX1 _14392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [7]),
    .Y(_6682_)
);

INVX1 _8707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .Y(_1591_)
);

FILL FILL_1__7664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13007_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf0),
    .B(_5184_),
    .C(_5183_),
    .Y(_5185_)
);

FILL FILL_1__8449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10774_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [4]),
    .Y(_105_)
);

DFFPOSX1 _8880_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_878_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Xin12b [9])
);

INVX1 _8460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .Y(_1359_)
);

AOI21X1 _8040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_956_),
    .C(_957_),
    .Y(_958_)
);

OAI21X1 _11097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3742_),
    .C(_3743_),
    .Y(_3744_)
);

FILL FILL_1__13180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7559_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [10]),
    .B(_1834__bF$buf2),
    .Y(_2460_)
);

FILL FILL_0__7139_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2051_),
    .C(_2063_),
    .Y(_2064_)
);

FILL FILL_1__11913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13798_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6036_),
    .C(_6037_),
    .Y(_6038_)
);

FILL FILL_0__13378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(vdd),
    .Y(_5698_)
);

FILL FILL_0__9705_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7069_),
    .B(_7070_),
    .Y(_6797_)
);

OAI21X1 _14448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6727_),
    .B(_6729_),
    .C(_6730_),
    .Y(_6514_)
);

OAI21X1 _14028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6373_),
    .B(_6363_),
    .C(_6386_),
    .Y(_6387_)
);

FILL FILL_2__8691_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .Y(_705_)
);

NAND2X1 _7311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_302_),
    .Y(_306_)
);

OAI21X1 _10788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3449_),
    .C(_3450_),
    .Y(_3451_)
);

FILL FILL_0__8097_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3092_),
    .B(_3086_),
    .C(_2741_),
    .Y(_3093_)
);

FILL FILL_1__12871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11024_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [11]),
    .C(_1762_),
    .Y(_1771_)
);

NAND3X1 _8516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1412_),
    .C(_1387_),
    .Y(_1413_)
);

FILL FILL_1__7893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13236_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5387_),
    .B(_5391_),
    .C(_5403_),
    .Y(_5404_)
);

FILL FILL_0__12649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12229_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [0]),
    .Y(_5023_)
);

FILL FILL_1__8678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10163_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf1),
    .B(_6090_),
    .C(_6087_),
    .Y(_6091_)
);

BUFX2 BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2648__bF$buf3)
);

BUFX2 BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2648__bF$buf2)
);

FILL FILL_2__7122_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2648__bF$buf1)
);

BUFX2 BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2648__bF$buf0)
);

BUFX2 BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf5)
);

BUFX2 BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf4)
);

BUFX2 BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf3)
);

FILL FILL_2__11788_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf2)
);

FILL FILL_2__11368_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf1)
);

BUFX2 BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .Y(_2686__bF$buf0)
);

FILL FILL256950x252150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7788_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2638_),
    .Y(\genblk1[3].u_ce.X_ [0])
);

FILL FILL_0__7368_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2282_),
    .Y(_2283_)
);

OAI21X1 _9054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_1880_),
    .C(_1881_),
    .Y(_1678_)
);

FILL FILL_1__11722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8327_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6256_),
    .Y(_6257_)
);

FILL FILL_0__13187_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13472_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5072_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [11])
);

NAND2X1 _13052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5473_),
    .B(_5256_),
    .Y(_5517_)
);

FILL FILL256950x219750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9514_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6898_),
    .B(_6901_),
    .C(_6833__bF$buf1),
    .Y(_6903_)
);

INVX4 _14257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf4 ),
    .Y(_6565_)
);

FILL FILL_1__7529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7109_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7960_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_44_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Xin12b [5])
);

NOR2X1 _7540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_522_),
    .Y(_525_)
);

OAI21X1 _7120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_123_),
    .C(_92_),
    .Y(_124_)
);

NAND2X1 _10597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3304_),
    .B(_3305_),
    .Y(_3306_)
);

NAND2X1 _10177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2908_),
    .B(_2909_),
    .Y(_2910_)
);

FILL FILL_1__12680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11253_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1625_),
    .C(_1623_),
    .Y(_1626_)
);

OAI21X1 _8325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1228_),
    .C(_1229_),
    .Y(_1230_)
);

FILL FILL_1__7282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12878_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .B(_5220_),
    .C(_5221_),
    .Y(_5030_)
);

FILL FILL_0__12458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4868_),
    .B(_4867_),
    .Y(_4869_)
);

FILL FILL_0__12038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10392_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6309_),
    .Y(_6310_)
);

INVX1 _13528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [8]),
    .Y(_5909_)
);

OAI21X1 _13108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5551_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5570_),
    .Y(_5046_)
);

FILL FILL257250x129750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7177_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2100_)
);

FILL FILL_1__11951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5734_),
    .B(_5733_),
    .Y(_5735_)
);

FILL FILL_1__12736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [4]),
    .B(_6737_),
    .Y(_6753_)
);

OAI21X1 _14066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6421_),
    .B(_6412_),
    .C(_5947_),
    .Y(_6423_)
);

FILL FILL_1__7758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9904_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.Xcalc [5]),
    .C(_1765_),
    .D(\genblk1[2].u_ce.Xcalc [7]),
    .Y(_1805_)
);

AOI21X1 _8554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1446_),
    .C(_1441_),
    .Y(_1449_)
);

MUX2X1 _8134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .B(_999_),
    .S(gnd),
    .Y(_1047_)
);

FILL FILL_1__7091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13274_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5440_)
);

FILL FILL_0__12687_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12552_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4206_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xcalc [3])
);

FILL FILL_0__12267_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .B(_4644_),
    .S(gnd),
    .Y(_4688_)
);

OAI21X1 _9759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_1759_),
    .C(_1753_),
    .Y(_1746_)
);

OAI21X1 _9339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf3),
    .B(_2152_),
    .C(_2153_),
    .Y(_2154_)
);

FILL FILL_1__8296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14059_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6127_),
    .Y(_6128_)
);

INVX1 _13337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [10]),
    .Y(_5788_)
);

FILL FILL_0__14833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10399_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(_1917_),
    .C(_1916_),
    .D(_1854_),
    .Y(_1918_)
);

FILL FILL_1__11760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10333_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5537_),
    .B(_5541_),
    .Y(_5553_)
);

NAND2X1 _7825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_791_),
    .Y(_792_)
);

NAND2X1 _7405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_395_),
    .Y(_396_)
);

FILL FILL_1__12965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11538_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348__bF$buf1),
    .B(_4393_),
    .C(_4349_),
    .Y(_4191_)
);

FILL FILL_0__9132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11118_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4032_),
    .B(_4034_),
    .C(_4021_),
    .Y(_3378_)
);

INVX1 _14295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [6]),
    .Y(_6598_)
);

FILL FILL_1__7567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14337_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12608_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4262_),
    .CLK(clk_bF$buf51),
    .Q(\genblk1[5].u_ce.Ain0 [1])
);

FILL FILL_0__11291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9713_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_921_),
    .C(_1652_),
    .Y(_884_)
);

NOR2X1 _8363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_1266_)
);

FILL FILL_1__10611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13083_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5198_),
    .B(_5257_),
    .C(_5256_),
    .D(_5194_),
    .Y(_5258_)
);

FILL FILL_0__12496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12076_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4903_),
    .B(_4900_),
    .Y(_4904_)
);

FILL FILL_2__12403_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .B(_2728_),
    .Y(_2729_)
);

OAI22X1 _9568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1756_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_2368_),
    .D(_2370_),
    .Y(_1703_)
);

INVX1 _9148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_1971_)
);

FILL FILL_1__11816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [6]),
    .Y(_6346_)
);

NAND2X1 _13566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_5926__bF$buf2),
    .Y(_5945_)
);

NAND3X1 _13146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(_5603_),
    .C(_5606_),
    .Y(_5607_)
);

FILL FILL_2__13608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10142_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_614_),
    .C(_602_),
    .Y(_615_)
);

AOI21X1 _7214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_209_),
    .C(_212_),
    .Y(_213_)
);

FILL FILL_1__12774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11347_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11632_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3372_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [7])
);

NAND2X1 _11212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3852_),
    .B(_3853_),
    .Y(_3854_)
);

OAI21X1 _8839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_1521_),
    .C(_917_),
    .Y(_910_)
);

AOI21X1 _8419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(gnd),
    .C(_1319_),
    .Y(_1320_)
);

FILL FILL_1__7796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x108150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13139_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5311_)
);

NAND3X1 _12417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [8]),
    .B(_4891_),
    .C(_4955_),
    .Y(_4956_)
);

FILL FILL_1__14920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9102_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(_1480_),
    .Y(_1485_)
);

INVX1 _8172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1081_),
    .Y(_1084_)
);

FILL FILL_1__10840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7865_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12590_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4244_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Yin12b [7])
);

AOI22X1 _12170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4311_),
    .B(_4348__bF$buf2),
    .C(_4724_),
    .D(_4346_),
    .Y(_4207_)
);

DFFPOSX1 _9797_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1709_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Acalc [8])
);

AOI21X1 _9377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .B(_2185_),
    .C(_2183_),
    .Y(_2190_)
);

FILL FILL_1__11205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8632_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [2]),
    .B(_3510__bF$buf0),
    .Y(_3558_)
);

FILL FILL_0__8212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14097_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6071_),
    .C(_6117_),
    .Y(_6164_)
);

OAI21X1 _13375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5199_),
    .C(_5813_),
    .Y(_5070_)
);

FILL FILL_2__13837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10371_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_183_),
    .C(_816_),
    .Y(_48_)
);

NAND2X1 _7443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_432_)
);

FILL FILL_2__13170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11576_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf1),
    .B(_4427_),
    .C(_4428_),
    .Y(_4429_)
);

FILL FILL_0__9170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11156_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4069_),
    .B(_4068_),
    .Y(_4070_)
);

AOI21X1 _11021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3661_),
    .B(_3639_),
    .C(_3640_),
    .Y(_3671_)
);

FILL FILL_2__11903_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_1536_)
);

OAI21X1 _8228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf3),
    .B(_1135_),
    .C(_1136_),
    .Y(_1137_)
);

FILL FILL_1__7185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [7]),
    .B(_5108_),
    .Y(_5130_)
);

INVX1 _12226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4776_),
    .Y(_4778_)
);

FILL FILL_0__13722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12441_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1998_),
    .B(_2004_),
    .C(_2007_),
    .Y(_2008_)
);

FILL FILL_1__11854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8021_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10712_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2538_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xcalc [11])
);

FILL FILL_0__10427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10007_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(_5641_),
    .C(_5642_),
    .Y(_5643_)
);

FILL FILL_2__9400_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7919_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ycalc [2])
);

FILL FILL_2__13646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9646_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4482_),
    .B(_4481_),
    .C(_4420_),
    .Y(_4483_)
);

FILL FILL_0__9226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6549_),
    .B(\u_ot.LoadCtl_6_bF$buf1 ),
    .C(_6679_),
    .Y(_6506_)
);

FILL FILL_0__10180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8602_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_638_),
    .Y(_651_)
);

INVX1 _7252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .Y(_250_)
);

FILL FILL_1__12392_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11670_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3410_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Yin1 [1])
);

FILL FILL_0__11385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf1),
    .B(_3763_),
    .Y(_3890_)
);

FILL FILL_2__11712_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8877_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_875_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[1].u_ce.Xin12b [10])
);

OAI21X1 _8457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1314_),
    .C(_1355_),
    .Y(_1356_)
);

NAND2X1 _8037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_954_),
    .Y(\genblk1[1].u_ce.Y_ [1])
);

FILL FILL_0__7712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13177_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5338_),
    .B(_5344_),
    .C(_5347_),
    .Y(_5348_)
);

NAND2X1 _12455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_4989_),
    .Y(_4990_)
);

OAI21X1 _12035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4593_),
    .B(_4595_),
    .C(_4417_),
    .Y(_4596_)
);

FILL FILL_2__12917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6826_),
    .B(_6834_),
    .Y(_6766_)
);

FILL FILL_1__11243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8670_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf1),
    .B(_3591_),
    .C(_3594_),
    .Y(_3595_)
);

FILL FILL_0__8250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10656_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [5]),
    .Y(_3235_)
);

FILL FILL_0__10236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .B(_2815_),
    .C(_2798_),
    .Y(_2837_)
);

OAI21X1 _7728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_701_),
    .C(_700_),
    .Y(_702_)
);

NAND2X1 _7308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_301_),
    .B(_302_),
    .Y(_303_)
);

FILL FILL_2__13875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9455_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Ycalc [11]),
    .C(_4276_),
    .Y(_4301_)
);

FILL FILL_0__9035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3940_),
    .C(_3935_),
    .Y(_3944_)
);

DFFPOSX1 _14198_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5874_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Yin12b [8])
);

FILL FILL_0__12802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8411_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_468_),
    .Y(_469_)
);

FILL FILL_0__11194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11101_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [6]),
    .B(_996__bF$buf3),
    .Y(_1571_)
);

NAND2X1 _8266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1170_),
    .B(_1173_),
    .Y(_1174_)
);

FILL FILL_1__10934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10514_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150_),
    .Y(_5150__bF$buf4)
);

FILL FILL_0__7521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7539_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150_),
    .Y(_5150__bF$buf3)
);

FILL FILL_2__7119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7101_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150_),
    .Y(_5150__bF$buf2)
);

BUFX2 BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150_),
    .Y(_5150__bF$buf1)
);

BUFX2 BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150_),
    .Y(_5150__bF$buf0)
);

BUFX2 BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .Y(_4324__bF$buf4)
);

BUFX2 BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .Y(_4324__bF$buf3)
);

BUFX2 BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .Y(_4324__bF$buf2)
);

BUFX2 BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .Y(_4324__bF$buf1)
);

MUX2X1 _12684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5164_),
    .B(_5161_),
    .S(_5151__bF$buf0),
    .Y(_5165_)
);

FILL FILL_0__12399_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .Y(_4324__bF$buf0)
);

OAI21X1 _12264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4796_),
    .B(_4794_),
    .C(_4362__bF$buf2),
    .Y(_4814_)
);

FILL FILL_2__12726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8306_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6253_),
    .B(_6242_),
    .S(vdd),
    .Y(_6254_)
);

DFFPOSX1 _13469_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5069_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin0 [0])
);

MUX2X1 _13049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5513_),
    .B(_5470_),
    .S(vdd),
    .Y(_5514_)
);

OAI21X1 _14830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [18]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(En_bF$buf2),
    .Y(_7045_)
);

FILL FILL_0__14125_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6555_),
    .B(_6562__bF$buf0),
    .C(_6696_),
    .D(_6697_),
    .Y(_6509_)
);

FILL FILL_1__11892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10465_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10750_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2576_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Ain12b [11])
);

FILL FILL_0__10045_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3055_),
    .Y(_3056_)
);

DFFPOSX1 _7957_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_41_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin12b [6])
);

NAND3X1 _7537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_443_),
    .C(_460_),
    .Y(_522_)
);

INVX1 _7117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [4]),
    .Y(_121_)
);

FILL FILL_2__13684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9684_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4517_),
    .Y(_4519_)
);

FILL FILL_0__9264_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [0]),
    .Y(_4154_)
);

INVX1 _11115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3749_),
    .Y(_3761_)
);

FILL FILL_1__7699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14403_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_284_),
    .C(_285_),
    .Y(_286_)
);

FILL FILL_0__13816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11750_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1373_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1392_),
    .Y(_856_)
);

INVX1 _8075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_990_),
    .Y(_991_)
);

FILL FILL_1__10323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5011_),
    .B(_4993_),
    .C(_5012_),
    .Y(_4242_)
);

NAND2X1 _12073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4630_),
    .B(_4631_),
    .Y(_4632_)
);

FILL FILL_2__12955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8535_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3465_),
    .C(_3466_),
    .Y(_3467_)
);

FILL FILL_0__8115_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6028_),
    .B(_5926__bF$buf2),
    .C(_6070_),
    .Y(_6071_)
);

NAND2X1 _13278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5729_),
    .B(_5731_),
    .Y(_5732_)
);

FILL FILL_2__9914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10601_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .Y(_737_)
);

OAI21X1 _7346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_339_),
    .C(_227_),
    .Y(_340_)
);

FILL FILL_1__12486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11479_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .Y(_4336_)
);

FILL FILL_0__9073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .B(_3978_),
    .Y(_3980_)
);

FILL FILL_0__12840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7806_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2652_),
    .S(_2649__bF$buf2),
    .Y(_2656_)
);

OAI21X1 _12969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_5437_),
    .C(_5246_),
    .Y(_5438_)
);

DFFPOSX1 _12549_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4203_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [0])
);

INVX1 _12129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4684_),
    .Y(_4685_)
);

FILL FILL_1__14632_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .Y(_6274_)
);

FILL FILL_0__13625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf4),
    .B(_1913_),
    .C(_1914_),
    .Y(_1915_)
);

FILL FILL_1__11757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x212550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8344_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [1]),
    .Y(_3319_)
);

AOI22X1 _13087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5137_),
    .B(_5174__bF$buf4),
    .C(_5550_),
    .D(_5172_),
    .Y(_5045_)
);

FILL FILL_2__9303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8505_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7995_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Vld )
);

NAND2X1 _7575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_557_),
    .Y(_558_)
);

OAI21X1 _7155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_153_),
    .C(_156_),
    .Y(_157_)
);

FILL FILL_1__12295_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4494_),
    .B(_4497_),
    .Y(_4555_)
);

FILL FILL_0__11288_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(_4159_),
    .C(_4176_),
    .Y(_3406_)
);

NAND2X1 _11153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [1]),
    .B(_3510__bF$buf4),
    .Y(_3797_)
);

FILL FILL_1__10608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7615_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_2479_),
    .C(_2498_),
    .Y(_1728_)
);

NAND2X1 _9301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_2117_),
    .Y(_2118_)
);

OAI21X1 _12778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf2),
    .B(_5253_),
    .C(_5254_),
    .Y(_5255_)
);

AOI21X1 _12358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4619_),
    .B(vdd),
    .C(_4362__bF$buf4),
    .Y(_4901_)
);

FILL FILL_1__14861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14219_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14504_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6492_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Xcalc [4])
);

FILL FILL_2__7386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8573_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3501_),
    .B(_3494_),
    .S(_3486__bF$buf3),
    .Y(_3502_)
);

FILL FILL_0__8153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10139_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3144_),
    .B(_3135_),
    .C(_2670_),
    .Y(_3146_)
);

INVX2 _10004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2742_),
    .Y(_2744_)
);

FILL FILL_2__9952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9358_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11629_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3369_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [4])
);

NOR2X1 _11209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf2),
    .B(_3850_),
    .Y(_3851_)
);

FILL FILL_1__13712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14917_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_371_),
    .C(_375_),
    .Y(_376_)
);

FILL FILL_0__11097_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_4014_),
    .C(\genblk1[4].u_ce.Ain0 [0]),
    .Y(_4015_)
);

FILL FILL_1__9939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9519_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(_1478_),
    .Y(_1482_)
);

OAI21X1 _8169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf4),
    .B(_1077_),
    .C(_1080_),
    .Y(_1081_)
);

FILL FILL_1__10837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7844_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2689_),
    .S(_2649__bF$buf2),
    .Y(_2693_)
);

FILL FILL_0__7424_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2331_),
    .B(_2335_),
    .Y(_2336_)
);

NAND2X1 _9110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf4),
    .B(_1884_),
    .Y(_1935_)
);

DFFPOSX1 _12587_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4241_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin12b [8])
);

OR2X2 _12167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4704_),
    .B(_4721_),
    .Y(_4722_)
);

FILL FILL_2__8803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14448_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6952_),
    .B(_6953_),
    .C(_6954_),
    .Y(_6778_)
);

FILL FILL_0__14028_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6613_),
    .B(_6610_),
    .Y(_6614_)
);

FILL FILL_2__12382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8382_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2790_),
    .B(_3324_),
    .C(_3340_),
    .Y(_2570_)
);

FILL FILL_0__10368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2963_)
);

FILL FILL_2__9341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13167_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1645_),
    .C(_1662_),
    .Y(_892_)
);

FILL FILL_0__9587_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4426_)
);

FILL FILL_0__9167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4062_),
    .B(_4065_),
    .Y(_4067_)
);

AOI21X1 _11018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3655_),
    .B(_3652_),
    .C(_3647_),
    .Y(_3668_)
);

FILL FILL_1__13941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14306_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .B(_192_),
    .S(_135__bF$buf3),
    .Y(_194_)
);

FILL FILL_0__13719_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3830_),
    .B(vdd),
    .C(_3833_),
    .Y(_3834_)
);

FILL FILL_1__9748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9328_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1292_),
    .S(_973__bF$buf1),
    .Y(_1300_)
);

FILL FILL_1__10646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10226_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf33)
);

FILL FILL_0__7653_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf32)
);

FILL FILL_0__7233_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf28)
);

INVX1 _12396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4936_),
    .Y(_4937_)
);

FILL FILL_0__13892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8018_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10709_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2535_),
    .CLK(clk_bF$buf34),
    .Q(\genblk1[3].u_ce.Xcalc [8])
);

FILL FILL_1__9081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14677_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14542_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6530_),
    .CLK(clk_bF$buf51),
    .Q(\u_ot.Yin12b [4])
);

FILL FILL_0__14257_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5967_),
    .B(_6466_),
    .C(_6468_),
    .Y(_5867_)
);

FILL FILL_1__7814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11184_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3538_),
    .B(_3531_),
    .S(_3486__bF$buf1),
    .Y(_3539_)
);

FILL FILL_0__8191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10597_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3177_),
    .B(_3180_),
    .Y(_3181_)
);

FILL FILL_0__10177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2780_),
    .C(_2777_),
    .Y(_2781_)
);

FILL FILL_2__10924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9150_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .B(_646_),
    .C(_256_),
    .Y(_648_)
);

OAI21X1 _7249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_245_),
    .C(_246_),
    .Y(_247_)
);

FILL FILL_2__13396_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1500_),
    .C(\genblk1[1].u_ce.Ain0 [0]),
    .Y(_1501_)
);

FILL FILL_1__12389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9396_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11667_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3407_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Yin12b [4])
);

INVX1 _11247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [5]),
    .Y(_3887_)
);

FILL FILL_1__13750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7709_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9815_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1727_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Yin12b [8])
);

FILL FILL_1__8772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13948_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf3),
    .B(_6180_),
    .Y(_6181_)
);

FILL FILL_0__13528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8667_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3487__bF$buf1),
    .Y(_3592_)
);

FILL FILL_0__8247_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3231_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_3233_)
);

FILL FILL_0__14486_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6989_)
);

FILL FILL_0__14066_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [0]),
    .Y(_6647_)
);

FILL FILL_1__7623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13806_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10691_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2517_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [2])
);

OAI21X1 _10271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2999_),
    .C(_2996_),
    .Y(_3000_)
);

FILL FILL_1__8828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10313_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Ain12b [9]),
    .Y(_836_)
);

INVX1 _7478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .Y(_466_)
);

FILL FILL_1__12198_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4444_),
    .B(_4462_),
    .C(_4350_),
    .Y(_4463_)
);

OAI21X1 _11476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4100_),
    .B(_4102_),
    .C(_4085_),
    .Y(_3383_)
);

INVX1 _11056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3702_),
    .Y(_3705_)
);

FILL FILL_2__11938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7518_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2422_),
    .Y(_2423_)
);

OR2X2 _9204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1999_),
    .B(_2003_),
    .Y(_2025_)
);

FILL FILL_1__8581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13757_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5943_),
    .B(_5990_),
    .C(_5988_),
    .Y(_5998_)
);

FILL FILL_0__13337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5658_),
    .B(_5656_),
    .Y(_5660_)
);

FILL FILL_1__9366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7009_),
    .B(_7040_),
    .C(_7041_),
    .Y(_7042_)
);

OAI21X1 _14407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6686_),
    .C(_6689_),
    .Y(_6695_)
);

FILL FILL_2_BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8056_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10747_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2573_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Yin0 [0])
);

AOI21X1 _10327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf1),
    .B(_3011_),
    .C(_3052_),
    .Y(_3053_)
);

FILL FILL_1__12830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14295_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [3]),
    .Y(_6822_)
);

DFFPOSX1 _14160_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5836_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[7].u_ce.Ycalc [1])
);

FILL FILL_1__7852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2815_),
    .B(_2816_),
    .Y(_2817_)
);

FILL FILL_1__8637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10122_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf2),
    .B(_282_),
    .C(_277_),
    .Y(_283_)
);

NOR2X1 _11285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3919_),
    .B(_3923_),
    .Y(_3924_)
);

FILL FILL_2__7501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7747_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(\genblk1[3].u_ce.LoadCtl [3]),
    .Y(_2603_)
);

FILL FILL_0__7327_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2204_),
    .B(_2205_),
    .C(_1815_),
    .Y(_2244_)
);

AOI21X1 _9013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1820_),
    .C(_1811__bF$buf0),
    .Y(_1842_)
);

FILL FILL_1__8390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13986_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6215_),
    .C(_6216_),
    .Y(_6217_)
);

FILL FILL_0__13566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13146_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13431_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5031_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Ycalc [2])
);

MUX2X1 _13011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5473_),
    .B(_5470_),
    .S(_5151__bF$buf3),
    .Y(_5478_)
);

FILL FILL_1__9595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10073_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6858_),
    .Y(_6865_)
);

INVX1 _14216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [0]),
    .Y(_6537_)
);

FILL FILL_0__7080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11278_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3628_)
);

FILL FILL_0__8285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf1),
    .B(_3185_),
    .Y(_3268_)
);

OAI21X1 _10136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2866_),
    .C(_2864_),
    .Y(_2871_)
);

FILL FILL_0__11212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1586_),
    .B(_1588_),
    .C(_1571_),
    .Y(_869_)
);

FILL FILL_1__7661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12837_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5181_),
    .B(_5160_),
    .C(_5151__bF$buf1),
    .Y(_5182_)
);

FILL FILL_0__12417_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .Y(_2653_)
);

FILL FILL_1__8446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14629_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [10]),
    .Y(_102_)
);

NAND2X1 _13907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6226_),
    .B(_6031_),
    .Y(_6271_)
);

NAND3X1 _11094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3727_),
    .B(_3739_),
    .C(_3723_),
    .Y(_3741_)
);

FILL FILL_2__7310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7556_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2454_),
    .B(_2457_),
    .Y(_2458_)
);

FILL FILL_0__7136_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .Y(_2061_)
);

FILL FILL_1__11910_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4603_),
    .B(_4846_),
    .Y(_4847_)
);

FILL FILL_0__10903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13795_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf4),
    .B(_6034_),
    .C(_6025_),
    .Y(_6035_)
);

FILL FILL_0__13375_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5695_)
);

FILL FILL_0__9702_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6816_),
    .B(_6833__bF$buf0),
    .C(_7068_),
    .Y(_6796_)
);

NOR2X1 _14445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [3]),
    .B(_6721_),
    .Y(_6728_)
);

NAND2X1 _14025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6377_),
    .B(_6380_),
    .Y(_6384_)
);

FILL FILL_1__7717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11087_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3446_),
    .C(_3447_),
    .Y(_3448_)
);

FILL FILL_0__8094_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3082_),
    .B(_3064_),
    .C(_3062_),
    .Y(_3090_)
);

FILL FILL_2__10827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11021_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.Acalc [0]),
    .C(_1767_),
    .D(_1768_),
    .Y(_1769_)
);

NOR2X1 _8513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1409_),
    .Y(_1410_)
);

FILL FILL_1__7890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12646_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .Y(_5401_)
);

FILL FILL_0__12226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4979_),
    .B(_4989_),
    .C(_5021_),
    .Y(_4251_)
);

OAI21X1 _9718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .B(_2479_),
    .C(_2496_),
    .Y(_1727_)
);

FILL FILL_1__8675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14018_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6049_),
    .B(_5926__bF$buf2),
    .C(_6070_),
    .Y(_6088_)
);

FILL FILL_2__11365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7785_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2635_),
    .C(_2636_),
    .Y(_2637_)
);

FILL FILL_0__7365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2264_),
    .C(_2237_),
    .Y(_2280_)
);

OAI21X1 _9051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834__bF$buf0),
    .B(_1879_),
    .C(_1835_),
    .Y(_1677_)
);

FILL FILL_2__8744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6900_)
);

NAND2X1 _14254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [0]),
    .B(_6562__bF$buf4),
    .Y(_6563_)
);

FILL FILL_1__7526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13709_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .Y(_3303_)
);

NAND2X1 _10174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2899_),
    .B(_2906_),
    .Y(_2907_)
);

FILL FILL_0__11250_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1619_),
    .B(_1604_),
    .C(_1618_),
    .Y(_1623_)
);

NAND3X1 _8322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_1225_),
    .C(_1209_),
    .Y(_1227_)
);

INVX1 _11799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4370_)
);

OAI21X1 _11379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4011_),
    .B(_4007_),
    .C(_3508_),
    .Y(_4013_)
);

FILL FILL_1__13882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12875_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174__bF$buf1),
    .B(_5219_),
    .C(_5175_),
    .Y(_5029_)
);

FILL FILL_0__12455_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4865_),
    .B(_4863_),
    .Y(_4866_)
);

FILL FILL_0__12035_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2690_)
);

NOR2X1 _9527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2332_),
    .Y(_2333_)
);

INVX1 _9107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_1932_)
);

FILL FILL_1__8484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6176_),
    .C(_6306_),
    .Y(_6307_)
);

FILL FILL_0_BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5903_),
    .B(_5906_),
    .C(_5892_),
    .Y(_5907_)
);

FILL FILL_0_BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(_5552_),
    .Y(_5568_)
);

FILL FILL_0_BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7174_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2095_),
    .B(_2097_),
    .C(_1906_),
    .Y(_2098_)
);

FILL FILL_0__10941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11306_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6733_),
    .C(_6751_),
    .Y(_6528_)
);

NAND2X1 _14063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6026_),
    .B(_6419_),
    .Y(_6420_)
);

FILL FILL257250x183750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9901_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [3]),
    .Y(_1802_)
);

NAND3X1 _8551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf3),
    .B(_1445_),
    .C(_1442_),
    .Y(_1446_)
);

NAND2X1 _8131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [2]),
    .B(_996__bF$buf0),
    .Y(_1044_)
);

NAND2X1 _11188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3593_),
    .B(_3778_),
    .Y(_3831_)
);

FILL FILL_1__13691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12264_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_1752_)
);

NAND2X1 _9336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2046_),
    .Y(_2151_)
);

FILL FILL_1__8293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13889_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6118_),
    .B(_6121_),
    .Y(_6125_)
);

FILL FILL_0__13049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5779_),
    .B(_5780_),
    .C(_5772_),
    .Y(_5785_)
);

FILL FILL_0__14830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10396_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14539_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6527_),
    .CLK(clk_bF$buf47),
    .Q(\u_ot.Yin12b [9])
);

NAND2X1 _14119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [0]),
    .B(_6466_),
    .Y(_6467_)
);

FILL FILL_2__8782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10330_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .Y(_789_)
);

NAND2X1 _7402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_392_),
    .Y(_393_)
);

NAND2X1 _10879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3536_)
);

FILL FILL_0__8188_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain0 [0]),
    .Y(_3178_)
);

OAI21X1 _10039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2748_),
    .C(_2686__bF$buf2),
    .Y(_2778_)
);

FILL FILL_1__12962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11535_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .B(_4360_),
    .C(_4390_),
    .Y(_4391_)
);

FILL FILL_0__11115_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4022_),
    .B(_4031_),
    .Y(_4032_)
);

NOR2X1 _14292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [4]),
    .B(\u_ot.Xin12b [5]),
    .Y(_6595_)
);

OAI21X1 _8607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .B(_1493_),
    .C(_994_),
    .Y(_1499_)
);

FILL FILL_1__7564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13327_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12605_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4259_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Ain1 [0])
);

FILL FILL_1__8769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9710_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1651_)
);

NAND2X1 _8360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1263_)
);

FILL FILL_1__13080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7879_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _9985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .B(_2676_),
    .C(_2724_),
    .D(_2668_),
    .Y(_2726_)
);

FILL FILL_0__7459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2367_),
    .B(_2360_),
    .Y(_2368_)
);

OAI21X1 _9145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1968_),
    .B(_1967_),
    .C(_1906_),
    .Y(_1969_)
);

FILL FILL_1__11813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14285_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6327_),
    .B(_6342_),
    .Y(_6344_)
);

FILL FILL_0__13698_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5924_),
    .B(_5941_),
    .Y(_5942_)
);

FILL FILL_0__13278_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5602_),
    .Y(_5604_)
);

FILL FILL_0__9605_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [14]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf4),
    .Y(_6987_)
);

NAND2X1 _14348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.LoadCtl_6_bF$buf4 ),
    .Y(_6645_)
);

FILL FILL_2__8591_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf0),
    .B(_606_),
    .C(_604_),
    .Y(_612_)
);

MUX2X1 _7211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .S(gnd),
    .Y(_210_)
);

DFFPOSX1 _10688_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2514_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Ycalc [0])
);

INVX1 _10268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .Y(_2997_)
);

FILL FILL_1__12771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11344_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[1] [0]),
    .Y(_916_)
);

NAND2X1 _8416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1079_),
    .B(_1264_),
    .Y(_1317_)
);

FILL FILL_1__7793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12969_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5308_),
    .B(_5307_),
    .C(_5246_),
    .Y(_5309_)
);

FILL FILL_0__12129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [8]),
    .B(_4348__bF$buf1),
    .Y(_4953_)
);

FILL FILL_0__13910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10063_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Vld ),
    .B(\genblk1[6].u_ce.ISout ),
    .Y(_5996_)
);

FILL FILL_2_BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7688_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9794_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1706_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[2].u_ce.Acalc [5])
);

FILL FILL_2_BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7268_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2186_),
    .Y(_2188_)
);

FILL FILL_2_BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11202_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.ISout ),
    .Y(_3556_)
);

FILL FILL_0__10615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14094_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [9]),
    .Y(_6161_)
);

FILL FILL_0__13087_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.X_ [0]),
    .Y(_5812_)
);

FILL FILL_1__12827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x129750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9414_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6818_),
    .B(\u_pa.RdyCtl [3]),
    .C(\u_pa.RdyCtl [2]),
    .Y(_6819_)
);

NAND2X1 _14157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[7] [1]),
    .B(_6455_),
    .Y(_6487_)
);

FILL FILL_1__7849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7429_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(gnd),
    .Y(_815_)
);

NOR2X1 _7440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_164_),
    .Y(_429_)
);

NOR2X1 _10497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2649__bF$buf4),
    .Y(_3213_)
);

NAND3X1 _10077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf2),
    .B(_2813_),
    .C(_2810_),
    .Y(_2814_)
);

FILL FILL_1__12160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11900_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [3]),
    .B(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_1533_)
);

NAND3X1 _8225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .B(_1123_),
    .C(_1104_),
    .Y(_1134_)
);

FILL FILL_1__7182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12778_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Ycalc [11]),
    .C(_5106_),
    .Y(_5127_)
);

FILL FILL_0__12358_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4774_),
    .Y(_4775_)
);

FILL FILL_1__8387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [0]),
    .B(_5949__bF$buf2),
    .Y(_6214_)
);

DFFPOSX1 _13428_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5028_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Ycalc [0])
);

OAI21X1 _13008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf3),
    .B(_5471_),
    .C(_5474_),
    .Y(_5475_)
);

FILL FILL_2__11077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7077_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .Y(_2005_)
);

FILL FILL_1__11851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10004_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5622_),
    .B(_5620_),
    .C(_5188__bF$buf2),
    .Y(_5640_)
);

DFFPOSX1 _7916_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Ycalc [0])
);

FILL FILL_1__12636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9643_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4479_),
    .Y(_4480_)
);

FILL FILL_0__9223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(_6674_),
    .Y(_6677_)
);

FILL FILL_1__7658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11382_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8874_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_872_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[1].u_ce.Acalc [9])
);

NAND2X1 _8454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1353_)
);

OAI21X1 _8034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(_951_),
    .C(_952_),
    .Y(_953_)
);

FILL FILL256950x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13174_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5343_),
    .Y(_5345_)
);

FILL FILL_0__12167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [5]),
    .B(_4275_),
    .Y(_4987_)
);

AND2X2 _12032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4587_),
    .B(_4583_),
    .Y(_4593_)
);

OR2X2 _9659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf1),
    .B(\genblk1[2].u_ce.Ain12b [9]),
    .Y(_2455_)
);

OAI21X1 _9239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2057_),
    .B(_2045_),
    .C(_1903_),
    .Y(_2059_)
);

FILL FILL_1__8196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .Y(_6032_)
);

NAND2X1 _13237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5682_),
    .B(_5691_),
    .Y(_5693_)
);

FILL FILL_0__14733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10233_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_135__bF$buf4),
    .Y(_699_)
);

NAND3X1 _7305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf2),
    .B(_299_),
    .C(_296_),
    .Y(_300_)
);

FILL FILL_1__12865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11438_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.Ycalc [0]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Ycalc [2]),
    .Y(_4299_)
);

FILL FILL_0__9032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11018_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3914_),
    .B(_3908_),
    .C(_3524__bF$buf5),
    .Y(_3941_)
);

DFFPOSX1 _14195_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5871_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin0 [1])
);

FILL FILL_1__7887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14237_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5397_),
    .B(_5385_),
    .C(_5243_),
    .Y(_5399_)
);

NAND2X1 _12508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.Y_ [1]),
    .Y(_5020_)
);

FILL FILL257250x115350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9613_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1558_),
    .Y(_1569_)
);

NAND3X1 _8263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1167_),
    .C(_1161_),
    .Y(_1171_)
);

FILL FILL_1__10931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10511_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .Y(_3486__bF$buf2)
);

FILL FILL_2__7536_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .Y(_3486__bF$buf1)
);

BUFX2 BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .Y(_3486__bF$buf0)
);

BUFX2 BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf5)
);

BUFX2 BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188_),
    .Y(_5188__bF$buf4)
);

INVX1 _12681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .Y(_5162_)
);

FILL FILL_0__12396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4810_),
    .Y(_4811_)
);

FILL FILL_2__12303_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2632_),
    .C(_2633_),
    .Y(_2634_)
);

NOR2X1 _9468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .B(_2271_),
    .Y(_2277_)
);

OAI21X1 _9048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .B(_1846_),
    .C(_1876_),
    .Y(_1877_)
);

FILL FILL_1__11716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8303_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf2),
    .B(_6250_),
    .C(_6243_),
    .Y(_6251_)
);

DFFPOSX1 _13466_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5066_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin12b [5])
);

INVX1 _13046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5511_)
);

FILL FILL_2__13508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10042_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7954_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Xin12b [11])
);

NAND2X1 _7534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_518_),
    .Y(_519_)
);

INVX1 _7114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [8]),
    .Y(_118_)
);

FILL FILL_1__12674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9681_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4515_),
    .Y(_4516_)
);

FILL FILL_0__9261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3608_),
    .B(_4151_),
    .C(_4152_),
    .Y(_3389_)
);

FILL FILL_0__11247_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3758_),
    .B(_3754_),
    .Y(_3759_)
);

OAI21X1 _8739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1619_),
    .B(_1616_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1621_)
);

OAI21X1 _8319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1135_),
    .C(_1164_),
    .Y(_1224_)
);

FILL FILL_1__7696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .B(_5186_),
    .C(_5216_),
    .Y(_5217_)
);

NOR2X1 _12317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4862_),
    .Y(_4863_)
);

FILL FILL_1__14820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9002_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .B(_1374_),
    .Y(_1390_)
);

MUX2X1 _8072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_987_),
    .B(_980_),
    .S(_972__bF$buf2),
    .Y(_988_)
);

FILL FILL_1__10320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7765_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5009_),
    .B(_4993_),
    .C(_5010_),
    .Y(_4241_)
);

NOR2X1 _12070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .B(_4628_),
    .Y(_4629_)
);

FILL FILL_2__12532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12112_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(_2483_),
    .Y(_2485_)
);

NOR3X1 _9277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2094_),
    .C(_2078_),
    .Y(_2095_)
);

FILL FILL_1__11945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8532_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3462_),
    .C(_3463_),
    .Y(_3464_)
);

FILL FILL_0__8112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6037_),
    .B(_6054_),
    .C(_6036_),
    .Y(_6068_)
);

OAI21X1 _13275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .B(_5257_),
    .C(_5188__bF$buf0),
    .Y(_5729_)
);

FILL FILL_2__13737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10271_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .Y(_734_)
);

INVX1 _7343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .Y(_337_)
);

FILL FILL_1__12483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11476_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4333_)
);

FILL FILL_0__9070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11056_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3975_),
    .B(_3976_),
    .Y(_3977_)
);

FILL FILL_2__11803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1796_),
    .B(_1799_),
    .C(_1768_),
    .Y(_1800_)
);

INVX1 _8548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .Y(_1443_)
);

INVX1 _8128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.ISout ),
    .Y(_1042_)
);

FILL FILL_1__7085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13268_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5425_),
    .B(_5434_),
    .C(_5418_),
    .Y(_5435_)
);

DFFPOSX1 _12546_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4200_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[5].u_ce.Ycalc [9])
);

OAI21X1 _12126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4682_),
    .B(_4681_),
    .C(_4417_),
    .Y(_4683_)
);

FILL FILL_0__13622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12341_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_1912_)
);

FILL FILL_1__11754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8341_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3312_),
    .B(_2599_),
    .Y(_3317_)
);

FILL FILL_0__10327_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .B(_5547_),
    .Y(_5548_)
);

FILL FILL_2__9720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9300_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_780_),
    .C(_769_),
    .Y(_786_)
);

FILL FILL_2__13966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9546_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4387_),
    .Y(_4388_)
);

FILL FILL_0__9126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13900_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [5]),
    .B(_6591_),
    .Y(_6593_)
);

FILL FILL_0__10080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8502_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7992_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[0].u_ce.LoadCtl [3])
);

INVX1 _7572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [6]),
    .Y(_555_)
);

NAND2X1 _7152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf1),
    .B(_135__bF$buf3),
    .Y(_154_)
);

FILL FILL_1__12292_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4534_),
    .B(_4348__bF$buf4),
    .C(_4552_),
    .D(_4532_),
    .Y(_4199_)
);

NAND2X1 _11570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .B(_4159_),
    .Y(_4175_)
);

FILL FILL_0__11285_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf1),
    .B(_3794_),
    .C(_3783_),
    .Y(_3795_)
);

FILL FILL_1__9707_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .B(_1648_),
    .C(_1649_),
    .Y(_881_)
);

NAND2X1 _8357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1246_),
    .B(_1260_),
    .Y(_850_)
);

FILL FILL_1__10605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13077_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5252_)
);

NOR2X1 _12355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4885_),
    .B(_4898_),
    .Y(_4218_)
);

FILL FILL_2__12817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14636_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14501_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6489_),
    .CLK(clk_bF$buf46),
    .Q(\u_ot.Xcalc [1])
);

FILL FILL_0__14216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8570_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(gnd),
    .Y(_3499_)
);

FILL FILL_0__8150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10136_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2749_),
    .B(_3142_),
    .Y(_3143_)
);

OAI21X1 _10001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2741_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_2742_)
);

OAI21X1 _7628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_583_),
    .C(_172__bF$buf4),
    .Y(_609_)
);

AOI21X1 _7208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_199_),
    .C(_197_),
    .Y(_207_)
);

FILL FILL_2__13775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9355_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11626_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3366_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[4].u_ce.Xcalc [1])
);

NAND2X1 _11206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [10]),
    .Y(_3848_)
);

OAI21X1 _14098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6452_),
    .B(_6451_),
    .C(_6444_),
    .Y(_5859_)
);

FILL FILL_0__12702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_280_),
    .C(_326_),
    .Y(_373_)
);

FILL FILL_0__13907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11001_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(_1444_),
    .Y(_1479_)
);

NOR2X1 _8166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_973__bF$buf2),
    .Y(_1078_)
);

FILL FILL_1__10834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7421_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12584_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4238_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xin0 [1])
);

FILL FILL_0__12299_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4715_),
    .C(_4710_),
    .Y(_4719_)
);

FILL FILL_2__12626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8206_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6103_),
    .B(_6157_),
    .C(_6155_),
    .Y(_6158_)
);

OAI21X1 _13369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5799_),
    .B(_5104_),
    .C(_5810_),
    .Y(_5067_)
);

FILL FILL_0__14865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14445_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6947_),
    .B(_6951_),
    .Y(_6952_)
);

FILL FILL_0__14025_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [6]),
    .B(\u_ot.Xin12b [7]),
    .Y(_6611_)
);

FILL FILL_1__11792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10785_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3324_),
    .Y(_3339_)
);

FILL FILL_0__10365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .B(_2957_),
    .Y(_2960_)
);

OAI21X1 _7857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_83_),
    .C(_813_),
    .Y(_45_)
);

OAI21X1 _7437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_424_),
    .C(_425_),
    .Y(_426_)
);

FILL FILL_2__13584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9584_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4423_)
);

FILL FILL_0__9164_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3781_),
    .C(_4063_),
    .Y(_4064_)
);

OAI21X1 _11015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3660_),
    .B(_3664_),
    .C(_3665_),
    .Y(_3666_)
);

FILL FILL_0__12931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14303_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_189_),
    .S(_135__bF$buf0),
    .Y(_191_)
);

FILL FILL_0__13716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9325_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf2),
    .B(_1293_),
    .C(_1296_),
    .Y(_1297_)
);

FILL FILL256650x126150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10223_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf63)
);

FILL FILL_0__7650_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf62)
);

FILL FILL_0__7230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7248_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf60)
);

CLKBUF1 CLKBUF1_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf58)
);

NAND2X1 _12393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [6]),
    .B(_4933_),
    .Y(_4934_)
);

FILL FILL_2__12855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8015_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10706_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2532_),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.Xcalc [5])
);

OAI21X1 _13598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5974_),
    .C(_5975_),
    .Y(_5976_)
);

NOR2X1 _13178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5636_),
    .Y(_5637_)
);

FILL FILL_0__14674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10501_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [10]),
    .B(_643_),
    .C(_644_),
    .Y(_645_)
);

NAND3X1 _7246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_243_),
    .C(_234_),
    .Y(_244_)
);

FILL FILL_1__12386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9393_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11664_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3404_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Yin12b [9])
);

FILL FILL_0__11379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3883_),
    .B(_3866_),
    .Y(_3885_)
);

FILL FILL_0__12740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7706_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9812_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1724_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin0 [1])
);

INVX1 _12869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5341_),
    .Y(_5342_)
);

NAND2X1 _12449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [11]),
    .B(_4348__bF$buf0),
    .Y(_4985_)
);

AOI21X1 _12029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4558_),
    .B(_4567_),
    .C(_4589_),
    .Y(_4590_)
);

FILL FILL_1__14112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13945_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6177_),
    .Y(_6178_)
);

FILL FILL_0__13525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8664_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3587_),
    .C(_3588_),
    .Y(_3589_)
);

FILL FILL_0__8244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3229_),
    .B(_3228_),
    .Y(_3230_)
);

FILL FILL_2__9203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8405_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Ain12b [8]),
    .Y(_834_)
);

MUX2X1 _7475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_451_),
    .S(gnd),
    .Y(_463_)
);

FILL FILL_1__12195_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4454_),
    .B(_4453_),
    .Y(_4460_)
);

FILL FILL_0__11188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4099_),
    .B(_4090_),
    .Y(_4100_)
);

OAI21X1 _11053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3612_),
    .C(_3678_),
    .Y(_3702_)
);

FILL FILL_2__11515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7515_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [6]),
    .B(_2419_),
    .Y(_2420_)
);

NOR2X1 _9201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .B(_2012_),
    .Y(_2022_)
);

INVX1 _12678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5159_)
);

OAI22X1 _12258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4308_),
    .B(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .C(_4808_),
    .D(_4806_),
    .Y(_4211_)
);

FILL FILL_1__14761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10261_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7038_),
    .B(_7034_),
    .Y(_7039_)
);

FILL FILL_0__14119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Ycalc [8]),
    .B(_6562__bF$buf1),
    .Y(_6693_)
);

FILL FILL_2__7286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10459_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10744_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2570_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin12b [5])
);

FILL FILL_0__10039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3045_),
    .B(_3028_),
    .C(_3041_),
    .Y(_3050_)
);

FILL FILL_2__9852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9678_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4475_),
    .B(_4491_),
    .C(_4474_),
    .Y(_4513_)
);

FILL FILL_0__9258_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3438_),
    .B(_3444_),
    .Y(_4150_)
);

NAND3X1 _11109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3729_),
    .B(_3732_),
    .C(_3711_),
    .Y(_3756_)
);

FILL FILL_1__13612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert200 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert202 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert204 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert205 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert207 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert209 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14817_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_135__bF$buf0),
    .C(_279_),
    .Y(_280_)
);

NOR2X1 _11282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3920_),
    .B(_3900_),
    .Y(_3921_)
);

FILL FILL_1__9419_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1386_),
    .Y(_1387_)
);

NAND2X1 _8069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(vdd),
    .Y(_985_)
);

FILL FILL_1__10317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7744_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.LoadCtl [3]),
    .Y(_2600_)
);

FILL FILL_0__7324_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(_2240_),
    .Y(_2241_)
);

MUX2X1 _9010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1838_),
    .B(_1837_),
    .S(_1811__bF$buf4),
    .Y(_1839_)
);

OAI21X1 _12487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4601_),
    .B(_4989_),
    .C(_5008_),
    .Y(_4240_)
);

MUX2X1 _12067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4625_),
    .B(_4623_),
    .S(_4325__bF$buf2),
    .Y(_4626_)
);

FILL FILL_2__8703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6860_),
    .B(_6862_),
    .Y(_6863_)
);

DFFPOSX1 _14213_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.LoadCtl [4])
);

FILL FILL_1__7905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11275_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(_3624_),
    .C(_3625_),
    .Y(_3626_)
);

FILL FILL_0__8282_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [7]),
    .Y(_3265_)
);

FILL FILL_0__10268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2866_),
    .C(_2867_),
    .Y(_2868_)
);

FILL FILL_2__9241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13067_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_1576_),
    .Y(_1586_)
);

FILL FILL_0__9487_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4330_)
);

FILL FILL_0__9067_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3891_),
    .C(_3937_),
    .Y(_3974_)
);

FILL FILL_1__13841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12414_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_2650_)
);

FILL FILL_1__8443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14626_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_99_),
    .C(_92_),
    .Y(_100_)
);

NAND2X1 _13904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf0),
    .B(_6224_),
    .Y(_6268_)
);

FILL FILL_0__13619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3649_),
    .C(_3678_),
    .Y(_3738_)
);

FILL FILL_1__9648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11553_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1170_),
    .B(_1173_),
    .C(_1203_),
    .Y(_1204_)
);

FILL FILL_1__10966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7133_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4835_),
    .Y(_4844_)
);

FILL FILL_0__10900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3313_),
    .Y(_3315_)
);

FILL FILL_2__9717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14577_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [16]),
    .B(_6833__bF$buf2),
    .C(En_bF$buf2),
    .Y(_7067_)
);

FILL FILL_0__14157_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.X_ [1]),
    .B(_6724_),
    .Y(_6726_)
);

NAND2X1 _14022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6379_),
    .B(_6380_),
    .Y(_6381_)
);

FILL FILL_1__7714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11084_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3432_),
    .B(_3435_),
    .C(_3445_),
    .Y(\a[5] [0])
);

FILL FILL_0__8091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10077_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3079_),
    .B(_3080_),
    .Y(_3087_)
);

FILL FILL_2__10824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9050_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7989_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[0].u_ce.LoadCtl [0])
);

AND2X2 _7569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_551_),
    .Y(_553_)
);

NOR2X1 _7149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_150_),
    .Y(_151_)
);

FILL FILL_2__13296_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.Acalc [4]),
    .C(_1765_),
    .D(\genblk1[2].u_ce.Acalc [6]),
    .Y(_1766_)
);

NOR2X1 _8510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1406_),
    .B(_1386_),
    .Y(_1407_)
);

FILL FILL_1__12289_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4549_),
    .Y(_4550_)
);

FILL FILL_0__9296_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [1]),
    .Y(_4173_)
);

NAND2X1 _11147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf0),
    .B(_3787_),
    .Y(_3792_)
);

FILL FILL_1__13650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7609_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2087_),
    .B(_2475_),
    .C(_2494_),
    .Y(_1726_)
);

FILL FILL_1__8672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13848_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [6]),
    .Y(_6085_)
);

FILL FILL_0__13008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10355_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[8]),
    .Y(Dout[8])
);

FILL FILL_0__7782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3496_)
);

FILL FILL_0__8147_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3138_),
    .B(_3137_),
    .Y(_3140_)
);

FILL FILL_1__12921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14386_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6896_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(_6897_),
    .Y(_6773_)
);

OAI21X1 _14251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_6559_),
    .C(_6560_),
    .Y(_7071_[11])
);

FILL FILL_1__7523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13706_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3293_),
    .B(_3294_),
    .C(_3283_),
    .Y(_3300_)
);

NAND2X1 _10171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2903_),
    .Y(_2904_)
);

FILL FILL_1__8728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10213_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .Y(_767_)
);

INVX1 _7378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_370_)
);

FILL FILL_1__12098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_4367_)
);

AOI21X1 _11376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .B(_3524__bF$buf2),
    .C(_3766_),
    .Y(_4010_)
);

FILL FILL_2__11838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7418_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2687_)
);

INVX1 _9524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2321_),
    .Y(_2330_)
);

AOI22X1 _9104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .B(_1834__bF$buf0),
    .C(_1929_),
    .D(_1906_),
    .Y(_1680_)
);

FILL FILL_1__8481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13657_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5917_),
    .B(_5949__bF$buf3),
    .C(_6304_),
    .D(_5947_),
    .Y(_5851_)
);

FILL FILL_0_BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13237_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [5]),
    .Y(_5904_)
);

FILL FILL_0_BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5564_),
    .Y(_5565_)
);

FILL FILL_0_BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10164_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6949_)
);

NAND3X1 _14307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6605_),
    .C(_6608_),
    .Y(_6609_)
);

FILL FILL_0__7591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3333_),
    .B(_3321_),
    .C(_3337_),
    .Y(_2567_)
);

OAI21X1 _10227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .B(_2957_),
    .C(_2670_),
    .Y(_2958_)
);

FILL FILL_1__12730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11303_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [9]),
    .B(_6729_),
    .Y(_6750_)
);

OR2X2 _14060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6415_),
    .B(_6414_),
    .Y(_6417_)
);

FILL FILL_1__7752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10022_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf5),
    .B(_150_),
    .C(_187_),
    .Y(_188_)
);

OAI21X1 _11185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .C(_3827_),
    .Y(_3828_)
);

FILL FILL_2__7401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7647_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2486_),
    .C(_1750_),
    .Y(_1743_)
);

FILL FILL_0__7227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [2]),
    .B(_1834__bF$buf4),
    .Y(_2148_)
);

FILL FILL_1__8290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13886_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6120_),
    .B(_6121_),
    .Y(_6122_)
);

FILL FILL_0__13046_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5781_),
    .B(_5778_),
    .C(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .Y(_5783_)
);

FILL FILL_1__9495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10393_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14536_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6524_),
    .CLK(clk_bF$buf47),
    .Q(\u_ot.Yin12b [10])
);

NAND2X1 _14116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(_6463_),
    .Y(_6465_)
);

FILL FILL_1__7808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [4]),
    .Y(_3533_)
);

FILL FILL_0__8185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3175_),
    .B(_3174_),
    .C(_3167_),
    .Y(_2538_)
);

NAND2X1 _10036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf0),
    .B(_2677_),
    .Y(_2775_)
);

FILL FILL_0__11952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11112_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1010__bF$buf3),
    .C(_1252_),
    .Y(_1496_)
);

FILL FILL_1__7561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12317_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12602_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4256_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Ain12b [7])
);

DFFPOSX1 _9809_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1721_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin1 [0])
);

FILL FILL_1__8766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14109_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5901_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6175_),
    .Y(_5845_)
);

FILL FILL_2__7210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7876_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2675_),
    .S(vdd),
    .Y(_2723_)
);

FILL FILL_0__7456_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .B(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_2365_)
);

NAND2X1 _9142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1963_),
    .B(_1965_),
    .Y(_1966_)
);

FILL FILL_1__11810_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .Y(_4752_)
);

FILL FILL_0__10803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14282_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5967_),
    .B(_6338_),
    .C(_6334_),
    .Y(_6341_)
);

FILL FILL_0__13695_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5937_),
    .C(_5938_),
    .Y(_5939_)
);

FILL FILL_0__13275_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5600_),
    .Y(_5601_)
);

FILL FILL_0__9602_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6980_),
    .B(_6983_),
    .Y(_6984_)
);

NAND2X1 _14345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6637_),
    .B(_6642_),
    .Y(_6643_)
);

FILL FILL256650x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7617_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3178_),
    .C(_2592_),
    .Y(_2585_)
);

NAND2X1 _10265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2949_),
    .B(_2754_),
    .Y(_2994_)
);

FILL FILL_0__11761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11341_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(_921_),
    .C(_914_),
    .Y(_907_)
);

OAI21X1 _8413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .C(_1313_),
    .Y(_1314_)
);

FILL FILL_1__7790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12966_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5303_),
    .B(_5305_),
    .Y(_5306_)
);

FILL FILL_0__12126_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4942_),
    .B(_4950_),
    .Y(_4951_)
);

NAND2X1 _9618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2416_),
    .Y(_2417_)
);

FILL FILL_1__8995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14338_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .B(_5992_),
    .C(_5951_),
    .Y(_5994_)
);

FILL FILL_2__11265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7685_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9791_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1703_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[2].u_ce.Acalc [2])
);

FILL FILL_0__7265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1856_),
    .B(_2182_),
    .C(_2181_),
    .Y(_2185_)
);

FILL FILL_2__8644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14289_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [9]),
    .Y(_6816_)
);

OAI21X1 _14154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5924_),
    .C(_6485_),
    .Y(_5882_)
);

FILL FILL_1__7846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert171 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert173 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert174 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert176 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert178 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3202_),
    .B(_3207_),
    .Y(_3210_)
);

AOI21X1 _10074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2772_),
    .B(_2649__bF$buf3),
    .C(_2793_),
    .Y(_2811_)
);

FILL FILL_0__11990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11150_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_1522_),
    .Y(_1531_)
);

OAI21X1 _8222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1131_),
    .Y(_844_)
);

OAI21X1 _11699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(\genblk1[5].u_ce.Acalc [8]),
    .C(_4276_),
    .Y(_4277_)
);

NAND3X1 _11279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3488_),
    .B(_3912_),
    .C(_3915_),
    .Y(_3918_)
);

FILL FILL_2__7915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x183750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12775_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Ycalc [0]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Ycalc [2]),
    .Y(_5125_)
);

FILL FILL_0__12355_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4755_),
    .Y(_4772_)
);

INVX2 _9847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .Y(_2597_)
);

INVX1 _9427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .Y(_2238_)
);

NOR2X1 _9007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1830_),
    .Y(_1836_)
);

FILL FILL_1__8384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14147_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6208_),
    .B(_6211_),
    .C(_6018_),
    .Y(_6212_)
);

OAI21X1 _13425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5680_),
    .C(_5100_),
    .Y(_5093_)
);

NAND2X1 _13005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5472_)
);

FILL FILL_1__9589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7074_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2001_),
    .Y(_2002_)
);

FILL FILL_0__10841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_664_),
    .C(_78_),
    .Y(_71_)
);

FILL FILL_2__13220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9658_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4466_),
    .B(_4473_),
    .C(_4476_),
    .Y(_4477_)
);

FILL FILL_0__9220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6673_),
    .B(_6666_),
    .Y(_6674_)
);

FILL FILL_1__7655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13418_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8871_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_869_),
    .CLK(clk_bF$buf46),
    .Q(\genblk1[1].u_ce.Acalc [6])
);

NAND2X1 _8451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1349_),
    .Y(_1351_)
);

AOI21X1 _8031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_948_),
    .C(_949_),
    .Y(_950_)
);

OAI21X1 _11088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3735_),
    .B(_3734_),
    .C(_3582_),
    .Y(_3736_)
);

FILL FILL_1__13591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12164_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .B(_2452_),
    .Y(_2453_)
);

NAND3X1 _9236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .B(_2055_),
    .C(_2054_),
    .Y(_2056_)
);

FILL FILL_1__8193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13789_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf2),
    .B(_5980_),
    .Y(_6029_)
);

FILL FILL_0__13369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(_5687_),
    .C(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5690_)
);

FILL FILL_0__14730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10296_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6801_),
    .B(_6833__bF$buf4),
    .C(_7065_),
    .Y(_6793_)
);

AND2X2 _14439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6723_),
    .B(_6720_),
    .Y(_6724_)
);

NAND3X1 _14019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf5),
    .B(_6377_),
    .C(_6374_),
    .Y(_6378_)
);

FILL FILL_2__8682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10230_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(_693_),
    .Y(_696_)
);

AOI21X1 _7302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_135__bF$buf0),
    .C(_279_),
    .Y(_297_)
);

OAI21X1 _10779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3436_),
    .B(_3439_),
    .C(_3442_),
    .Y(_3443_)
);

FILL FILL_0__8088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3045_),
    .B(_3028_),
    .C(_3083_),
    .Y(_3084_)
);

FILL FILL_1__12862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11435_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [6]),
    .B(_4279_),
    .Y(_4296_)
);

FILL FILL_0__11015_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3850_),
    .C(_3937_),
    .Y(_3938_)
);

DFFPOSX1 _14192_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5868_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin1 [0])
);

OAI21X1 _8927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(\genblk1[2].u_ce.Acalc [8]),
    .C(_1762_),
    .Y(_1763_)
);

NAND3X1 _8507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_1398_),
    .C(_1401_),
    .Y(_1404_)
);

FILL FILL_1__7884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .B(_5395_),
    .C(_5394_),
    .Y(_5396_)
);

OAI21X1 _12505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5011_),
    .B(_4273_),
    .C(_5018_),
    .Y(_4248_)
);

FILL FILL_1__8669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9610_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1565_),
    .B(_1564_),
    .Y(_1566_)
);

OAI21X1 _8260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1134_),
    .C(_1010__bF$buf0),
    .Y(_1168_)
);

BUFX2 BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .Y(_2672__bF$buf3)
);

BUFX2 BUFX2_insert221 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .Y(_2672__bF$buf2)
);

BUFX2 BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .Y(_2672__bF$buf1)
);

BUFX2 BUFX2_insert223 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .Y(_2672__bF$buf0)
);

BUFX2 BUFX2_insert224 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf0 )
);

FILL FILL_2__11779_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .Y(_5926__bF$buf4)
);

BUFX2 BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .Y(_5926__bF$buf3)
);

FILL FILL_0__12393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7779_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_2630_),
    .Y(\genblk1[3].u_ce.Y_ [1])
);

FILL FILL_0__7359_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2273_),
    .B(_2274_),
    .C(_1831_),
    .Y(_2275_)
);

INVX1 _9045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1873_),
    .Y(_1874_)
);

FILL FILL_1__11713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6067_),
    .C(_6247_),
    .Y(_6248_)
);

FILL FILL_0__13178_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13463_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5063_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin12b [6])
);

OAI21X1 _13043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5508_),
    .B(_5507_),
    .C(_5243_),
    .Y(_5509_)
);

FILL FILL_2__13925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9505_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6893_),
    .B(_6894_),
    .C(_6888_),
    .Y(_6895_)
);

OAI21X1 _14248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_6557_),
    .C(_6558_),
    .Y(_7071_[10])
);

FILL FILL257250x136950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8491_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7951_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Acalc [10])
);

OAI21X1 _7531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_385_),
    .C(_515_),
    .Y(_516_)
);

OAI21X1 _7111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_115_),
    .C(_92_),
    .Y(_116_)
);

OAI22X1 _10588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2608_),
    .B(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .C(_3297_),
    .D(_3296_),
    .Y(_2548_)
);

INVX1 _10168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2900_),
    .Y(_2901_)
);

FILL FILL_1__12671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [9]),
    .B(_1010__bF$buf5),
    .Y(_1618_)
);

OAI21X1 _8316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .B(_1220_),
    .C(_1068_),
    .Y(_1222_)
);

FILL FILL_1__7693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12869_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5213_),
    .Y(_5214_)
);

FILL FILL_0__12449_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4853_),
    .Y(_4860_)
);

FILL FILL_0__12029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8058_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6301_),
    .B(_6286_),
    .Y(_6302_)
);

INVX1 _13519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [9]),
    .Y(_5901_)
);

FILL FILL_0__7588_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(_1765_),
    .Y(_2483_)
);

FILL FILL_0__7168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2071_),
    .Y(_2092_)
);

FILL FILL_1__11942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10935_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3461_),
    .B(_3460_),
    .Y(\genblk1[4].u_ce.Y_ [0])
);

FILL FILL_0__10515_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5896_),
    .B(_5949__bF$buf1),
    .C(_6065_),
    .D(_6021_),
    .Y(_5840_)
);

AOI21X1 _13272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5706_),
    .B(_5714_),
    .C(_5713_),
    .Y(_5726_)
);

FILL FILL_2__13734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9314_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14897_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6788_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.Atmp [1])
);

NAND2X1 _14477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [8]),
    .B(_6729_),
    .Y(_6748_)
);

INVX1 _14057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6413_),
    .Y(_6414_)
);

FILL FILL_1__7749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_731_),
    .Y(_732_)
);

NAND2X1 _7340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_330_),
    .Y(_334_)
);

OAI21X1 _10397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3119_),
    .C(_3099_),
    .Y(_3120_)
);

FILL FILL_1__12480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11800_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [4]),
    .Y(_1797_)
);

AOI21X1 _8545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .B(_1415_),
    .C(_1438_),
    .Y(_1440_)
);

OR2X2 _8125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1038_),
    .B(_990_),
    .Y(_1040_)
);

FILL FILL_1__7082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .B(_5411_),
    .Y(_5432_)
);

FILL FILL_0__12678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12258_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12543_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4197_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[5].u_ce.Ycalc [6])
);

NOR2X1 _12123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4679_),
    .B(_4678_),
    .Y(_4680_)
);

FILL FILL_1__8287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf1),
    .B(_6118_),
    .C(_6114_),
    .Y(_6119_)
);

NAND2X1 _13328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [9]),
    .B(_5188__bF$buf4),
    .Y(_5780_)
);

FILL FILL_0__14824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7397_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_1909_)
);

FILL FILL_1__11751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10324_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5541_),
    .C(_5536_),
    .Y(_5545_)
);

OAI22X1 _7816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_783_),
    .D(_782_),
    .Y(_34_)
);

FILL FILL_2__13963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11529_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4384_),
    .B(_4381_),
    .S(_4324__bF$buf4),
    .Y(_4385_)
);

FILL FILL_0__9123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11109_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [5]),
    .Y(_6590_)
);

FILL FILL_1__7558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9704_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1645_),
    .C(_1647_),
    .Y(_880_)
);

AOI21X1 _8354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(_1241_),
    .C(_1247_),
    .Y(_1258_)
);

FILL FILL_1__10602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13074_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5249_)
);

FILL FILL_0__12487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12067_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4893_),
    .B(_4895_),
    .Y(_4896_)
);

FILL FILL_2__12814_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [2]),
    .B(_2672__bF$buf0),
    .Y(_2720_)
);

OAI21X1 _9559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(gnd),
    .Y(_2362_)
);

NAND3X1 _9139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1952_),
    .B(_1959_),
    .C(_1962_),
    .Y(_1963_)
);

FILL FILL_1__8096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x115350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6332_),
    .B(_6337_),
    .Y(_6338_)
);

OAI21X1 _13557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5934_),
    .C(_5935_),
    .Y(_5936_)
);

INVX1 _13137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .Y(_5598_)
);

FILL FILL_0__14633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10133_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_605_),
    .C(_585_),
    .Y(_606_)
);

NAND2X1 _7205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .B(\genblk1[0].u_ce.ISin ),
    .Y(_205_)
);

FILL FILL_1__12765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11338_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11623_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3363_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[4].u_ce.Ycalc [10])
);

OAI21X1 _11203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510__bF$buf3),
    .B(_3845_),
    .C(_3824_),
    .Y(_3367_)
);

NOR2X1 _14095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6449_),
    .B(_6448_),
    .Y(_6450_)
);

FILL FILL_1__7787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14137_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5292_),
    .B(_5299_),
    .C(_5302_),
    .Y(_5303_)
);

INVX1 _12408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4947_),
    .Y(_4948_)
);

FILL FILL_1__14911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1475_),
    .C(_1473_),
    .Y(_1476_)
);

OAI21X1 _8163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1073_),
    .C(_1074_),
    .Y(_1075_)
);

FILL FILL_1__10831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12296_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12581_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4235_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xin1 [0])
);

OAI21X1 _12161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4715_),
    .C(_4711_),
    .Y(_4716_)
);

FILL FILL_2__12203_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9788_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1700_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [11])
);

OAI21X1 _9368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2175_),
    .B(_2178_),
    .C(_2180_),
    .Y(_2182_)
);

FILL FILL_0__8623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14088_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6154_),
    .B(_6126_),
    .Y(_6155_)
);

NAND2X1 _13366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5807_),
    .Y(_5809_)
);

FILL FILL_2__13408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10362_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_810_),
    .Y(_812_)
);

NAND2X1 _7434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [0]),
    .B(_158__bF$buf3),
    .Y(_423_)
);

FILL FILL_1__12994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11567_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4418_),
    .Y(_4420_)
);

FILL FILL_0__9161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [4]),
    .B(_3510__bF$buf0),
    .Y(_4061_)
);

OAI21X1 _11012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3624_),
    .B(_3606_),
    .C(_3662_),
    .Y(_3663_)
);

NAND2X1 _8639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1526_),
    .B(_1527_),
    .Y(_1528_)
);

AND2X2 _8219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1113_),
    .B(_1128_),
    .Y(_1129_)
);

FILL FILL_1__7596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [6]),
    .B(_5108_),
    .Y(_5122_)
);

NAND2X1 _12217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .B(_4769_),
    .Y(_4770_)
);

FILL FILL_1__14720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1294_)
);

FILL FILL_1__10640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7665_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4930_),
    .Y(_4931_)
);

FILL FILL_2__12432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12012_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [5]),
    .Y(_2397_)
);

NAND3X1 _9177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1961_),
    .B(_1977_),
    .C(_1960_),
    .Y(_1999_)
);

FILL FILL_1__11845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8012_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10703_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2529_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xcalc [2])
);

OAI21X1 _13595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5971_),
    .C(_5972_),
    .Y(_5973_)
);

OAI22X1 _13175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5134_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5634_),
    .D(_5632_),
    .Y(_5049_)
);

FILL FILL_2__13637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9637_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _11908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .B(_4452_),
    .C(_4424_),
    .Y(_4474_)
);

FILL FILL_0__9217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10171_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_641_),
    .C(_172__bF$buf0),
    .Y(_642_)
);

NOR2X1 _7243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_241_)
);

FILL FILL_1__12383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9390_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11661_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3401_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Yin12b [10])
);

FILL FILL_0__11376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_3881_),
    .C(_3880_),
    .Y(_3882_)
);

FILL FILL_2__11703_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8868_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_866_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Acalc [3])
);

NAND2X1 _8448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1347_),
    .B(_1346_),
    .Y(_1348_)
);

NAND2X1 _8028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_947_),
    .B(_946_),
    .Y(\genblk1[1].u_ce.Y_ [0])
);

FILL FILL_0__7703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5301_),
    .B(_5317_),
    .C(_5300_),
    .Y(_5339_)
);

AND2X2 _12446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4978_),
    .B(_4982_),
    .Y(_4983_)
);

NAND3X1 _12026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .B(_4581_),
    .C(_4586_),
    .Y(_4587_)
);

FILL FILL_0__13942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8661_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3522_),
    .B(_3547_),
    .C(_3565_),
    .Y(_3586_)
);

FILL FILL_0__8241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10647_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3186_),
    .C(_3226_),
    .Y(_3227_)
);

FILL FILL_0__10227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_693_),
    .Y(_694_)
);

FILL FILL_2__13866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9446_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(\genblk1[5].u_ce.Ycalc [8]),
    .C(_4276_),
    .Y(_4293_)
);

FILL FILL_0__9026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13800_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14189_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5865_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Xin12b [7])
);

FILL FILL_1__8822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8402_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [1]),
    .B(_799_),
    .Y(_832_)
);

OAI21X1 _7472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf0),
    .B(_459_),
    .C(_452_),
    .Y(_460_)
);

FILL FILL_1__12192_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4456_),
    .C(_4453_),
    .Y(_4457_)
);

FILL FILL_0__11185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4095_),
    .B(\genblk1[4].u_ce.Ain12b [6]),
    .Y(_4097_)
);

AOI21X1 _11050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3698_),
    .B(_3672_),
    .C(_3697_),
    .Y(_3699_)
);

FILL FILL_1__9607_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .B(_1562_),
    .Y(_1563_)
);

OAI21X1 _8257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1077_),
    .C(_1164_),
    .Y(_1165_)
);

FILL FILL_1__10925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10505_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert190 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_158__bF$buf0)
);

FILL FILL_0__7512_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .Y(_5174__bF$buf4)
);

BUFX2 BUFX2_insert192 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .Y(_5174__bF$buf3)
);

FILL FILL_1__13397_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert193 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .Y(_5174__bF$buf2)
);

BUFX2 BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .Y(_5174__bF$buf1)
);

BUFX2 BUFX2_insert195 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .Y(_5174__bF$buf0)
);

BUFX2 BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert197 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf1 )
);

NAND2X1 _12675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5156_)
);

BUFX2 BUFX2_insert199 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf0 )
);

INVX1 _12255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4805_),
    .Y(_4806_)
);

FILL FILL_2__12717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9360_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(_7035_),
    .Y(_7036_)
);

FILL FILL_0__14116_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6689_),
    .B(_6686_),
    .Y(_6690_)
);

FILL FILL_2__12470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8050_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10741_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2567_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Yin12b [6])
);

FILL FILL_0__10456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10036_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3047_),
    .B(_3046_),
    .Y(_3048_)
);

DFFPOSX1 _7948_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Acalc [7])
);

AOI22X1 _7528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_158__bF$buf0),
    .C(_513_),
    .D(_156_),
    .Y(_16_)
);

INVX1 _7108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [5]),
    .Y(_113_)
);

FILL FILL_2__13675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9675_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4444_),
    .B(_4508_),
    .C(_4509_),
    .Y(_4510_)
);

FILL FILL_0__9255_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4144_),
    .B(_4140_),
    .C(_4143_),
    .Y(_4148_)
);

NAND3X1 _11106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3711_),
    .B(_3733_),
    .C(_3719_),
    .Y(_3753_)
);

FILL FILL_1__8631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14814_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_263_),
    .C(_245_),
    .Y(_277_)
);

FILL FILL_0__13807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11741_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1383_),
    .C(_1010__bF$buf2),
    .Y(_1384_)
);

NAND2X1 _8066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_982_)
);

FILL FILL_1__10314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_4989_),
    .Y(_5007_)
);

OAI21X1 _12064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4485_),
    .C(_4622_),
    .Y(_4623_)
);

FILL FILL_2__12946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8106_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6062_),
    .B(_6059_),
    .Y(_6063_)
);

OR2X2 _13269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5722_),
    .B(_5719_),
    .Y(_5723_)
);

FILL FILL_2__9905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14345_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6849_),
    .B(_6852_),
    .C(_6859_),
    .Y(_6860_)
);

DFFPOSX1 _14210_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.LoadCtl [1])
);

FILL FILL_1__7902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x126150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11272_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3621_),
    .B(_3622_),
    .C(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3623_)
);

FILL FILL_0__10685_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .B(_3252_),
    .Y(_3263_)
);

FILL FILL_0__10265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2864_),
    .C(_2863_),
    .Y(_2865_)
);

INVX1 _7757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .Y(_729_)
);

NAND2X1 _7337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_330_),
    .Y(_331_)
);

FILL FILL_1__12897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9484_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4327_)
);

FILL FILL_0__9064_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [9]),
    .B(_3510__bF$buf4),
    .Y(_3971_)
);

FILL FILL_0__12831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14689_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .Y(_2647_)
);

FILL FILL_1__8440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14623_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [5]),
    .Y(_97_)
);

NAND2X1 _13901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6234_),
    .B(_6251_),
    .Y(_6265_)
);

FILL FILL_0__13616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1170_),
    .Y(_1201_)
);

FILL FILL_1__10963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4840_),
    .B(_4841_),
    .Y(_4842_)
);

FILL FILL_2__12755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8335_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3311_),
    .B(_3312_),
    .Y(_3313_)
);

DFFPOSX1 _13498_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.LoadCtl [3])
);

OAI21X1 _13078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5541_),
    .C(_5537_),
    .Y(_5542_)
);

FILL FILL_0__14574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10401_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7986_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_70_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Ain1 [1])
);

NAND3X1 _7566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_547_),
    .C(_543_),
    .Y(_550_)
);

OAI21X1 _7146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_146_),
    .C(_147_),
    .Y(_148_)
);

FILL FILL_2__13293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11699_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4542_),
    .C(_4540_),
    .Y(_4547_)
);

FILL FILL_0__9293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11279_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [0]),
    .Y(_4171_)
);

NAND2X1 _11144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3788_),
    .Y(_3789_)
);

FILL FILL_2__11606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7606_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2475_),
    .Y(_2493_)
);

INVX2 _12769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5244_),
    .Y(_5246_)
);

NOR2X1 _12349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4888_),
    .B(_4892_),
    .Y(_4893_)
);

FILL FILL_1__14852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13845_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6081_),
    .B(_6066_),
    .C(_6018_),
    .Y(_6083_)
);

FILL FILL_0__13425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10352_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[5]),
    .Y(Dout[5])
);

FILL FILL_2__7377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8564_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3491_),
    .C(_3492_),
    .Y(_3493_)
);

FILL FILL_0__8144_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3136_),
    .Y(_3137_)
);

FILL FILL_2__9943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14908_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_154_),
    .Y(_764_)
);

OAI21X1 _7375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_366_),
    .C(_364_),
    .Y(_367_)
);

FILL FILL_1__12095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4364_)
);

FILL FILL_0__11088_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3990_),
    .B(_4000_),
    .C(_4006_),
    .Y(_4007_)
);

FILL FILL_2__11415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7835_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _9941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .B(_2683_),
    .C(_2648__bF$buf3),
    .D(_2677_),
    .Y(_2684_)
);

FILL FILL_0__7415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2326_),
    .B(_2327_),
    .Y(_2328_)
);

NAND2X1 _9101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1924_),
    .B(_1926_),
    .Y(_1927_)
);

NAND2X1 _12998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5465_)
);

DFFPOSX1 _12578_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4232_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xin12b [7])
);

OAI21X1 _12158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4693_),
    .B(_4712_),
    .C(_4362__bF$buf1),
    .Y(_4713_)
);

FILL FILL_1__14661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert211 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert212 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert214 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert216 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert217 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert219 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14439_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6946_)
);

FILL FILL_0__14019_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [7]),
    .Y(_6606_)
);

FILL FILL_2__7186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8373_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_3336_)
);

FILL FILL_0__10359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2947_),
    .Y(_2955_)
);

FILL FILL_0__11720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9578_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4417_),
    .C(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .Y(_4418_)
);

FILL FILL_0__9158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4058_),
    .B(_4049_),
    .C(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_4059_)
);

NAND2X1 _11009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3656_),
    .B(_3659_),
    .Y(_3660_)
);

FILL FILL_1__13932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14717_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_183_),
    .C(_184_),
    .Y(_185_)
);

AOI21X1 _11182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3819_),
    .C(_3817_),
    .Y(_3825_)
);

FILL FILL_1__9739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9319_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1291_)
);

FILL FILL_1__10637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7644_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .B(_2483_),
    .Y(_1749_)
);

FILL FILL_0__7224_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .B(_2122_),
    .Y(_2146_)
);

OAI21X1 _12387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4925_),
    .B(_4907_),
    .C(_4927_),
    .Y(_4928_)
);

FILL FILL_2__8603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14668_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14533_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6521_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin1 [1])
);

FILL FILL_0__14248_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .B(_5891_),
    .Y(_6463_)
);

FILL FILL_1__7805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11175_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3528_),
    .C(_3529_),
    .Y(_3530_)
);

FILL FILL_0__8182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(_3171_),
    .Y(_3173_)
);

OAI21X1 _10033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2770_),
    .C(_2771_),
    .Y(_2772_)
);

FILL FILL_2__10915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9141_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_1486_),
    .C(_1492_),
    .Y(_1493_)
);

FILL FILL_0__9387_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11658_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3398_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Xin1 [1])
);

NAND3X1 _11238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(_3878_),
    .C(_3876_),
    .Y(_3879_)
);

FILL FILL_1__13741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12314_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9806_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1718_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin12b [7])
);

FILL FILL_1__8763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13939_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6160_),
    .B(_6172_),
    .Y(_6173_)
);

FILL FILL_0__13519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11453_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1107_),
    .B(_1108_),
    .C(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1109_)
);

FILL FILL_1__10866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7453_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4668_),
    .C(_4748_),
    .Y(_4749_)
);

FILL FILL_2__8832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8658_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3571_),
    .B(_3559_),
    .C(_3572_),
    .Y(_3583_)
);

FILL FILL_0__8238_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [4]),
    .Y(_3224_)
);

FILL FILL_2__9617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14477_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6981_)
);

FILL FILL_0__14057_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6638_),
    .B(_6639_),
    .C(_6629_),
    .Y(_6640_)
);

FILL FILL_1__7614_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_2591_)
);

FILL FILL_0__10397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf3),
    .B(_2947_),
    .Y(_2991_)
);

FILL FILL_1__8819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_171_),
    .C(_830_),
    .Y(_60_)
);

OAI21X1 _7469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_276_),
    .C(_456_),
    .Y(_457_)
);

FILL FILL_2__13196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [1]),
    .B(_1648_),
    .Y(_913_)
);

AOI21X1 _8410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1284_),
    .B(_1305_),
    .C(_1303_),
    .Y(_1311_)
);

FILL FILL_1__12189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .B(_4424_),
    .C(_4362__bF$buf0),
    .Y(_4454_)
);

FILL FILL_0__9196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4091_),
    .B(_4051_),
    .C(_3524__bF$buf2),
    .Y(_4094_)
);

INVX1 _11047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [8]),
    .Y(_3696_)
);

FILL FILL_1__13970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2411_),
    .B(_2393_),
    .C(_2413_),
    .Y(_2414_)
);

FILL FILL_1__8992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13748_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5989_),
    .B(_5990_),
    .Y(_5991_)
);

FILL FILL_0__13328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7028_),
    .B(_7010_),
    .C(_7026_),
    .Y(_7033_)
);

FILL FILL_2_BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8047_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10738_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2564_),
    .CLK(clk_bF$buf50),
    .Q(\genblk1[3].u_ce.Yin12b [11])
);

NAND2X1 _10318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3041_),
    .B(_3044_),
    .Y(_3045_)
);

FILL FILL_1__12821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [0]),
    .B(\u_pa.RdyCtl [0]),
    .Y(_6814_)
);

OAI21X1 _14151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6484_)
);

FILL FILL_1__7843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert140 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert142 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert143 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert145 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert147 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert149 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .B(_3207_),
    .Y(_3208_)
);

INVX1 _10071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [6]),
    .Y(_2808_)
);

FILL FILL_1__8628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10113_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_662_),
    .C(_172__bF$buf5),
    .Y(_674_)
);

AOI22X1 _7278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_158__bF$buf1),
    .C(_274_),
    .D(_230_),
    .Y(_5_)
);

NOR2X1 _11696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Acalc [10]),
    .Y(_4274_)
);

OAI21X1 _11276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3913_),
    .C(_3914_),
    .Y(_3915_)
);

FILL FILL_2__11738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7738_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [2]),
    .Y(_2594_)
);

FILL FILL_0__7318_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2154_),
    .C(_2234_),
    .Y(_2235_)
);

OAI21X1 _9004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1808_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_1833_),
    .Y(_1676_)
);

FILL FILL_1__8381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13557_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6208_),
    .Y(_6209_)
);

FILL FILL_0__13137_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Ain1 [1]),
    .Y(_5099_)
);

NAND2X1 _13002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5469_)
);

FILL FILL_1__9586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10064_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6857_)
);

DFFPOSX1 _14207_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5883_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[7].u_ce.Yin0 [1])
);

FILL FILL_0__7491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8450_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_77_)
);

FILL FILL_1__11269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8696_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3607_),
    .B(_3619_),
    .C(_3617_),
    .Y(_3620_)
);

FILL FILL_0__8276_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3258_),
    .B(_3259_),
    .Y(_3260_)
);

INVX1 _10127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_2862_)
);

FILL FILL_1__12630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14095_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6670_),
    .B(_6669_),
    .C(_6562__bF$buf3),
    .Y(_6672_)
);

FILL FILL_1__7652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8017_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [9]),
    .Y(_94_)
);

AND2X2 _11085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3729_),
    .B(_3732_),
    .Y(_3733_)
);

FILL FILL_2__11967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7547_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .B(_2393_),
    .C(_2448_),
    .Y(_2450_)
);

FILL FILL_0__7127_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_2052_),
    .C(_2050_),
    .Y(_2053_)
);

FILL FILL_1__8190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13366_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .Y(_6026_)
);

AND2X2 _13231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5686_),
    .B(_5684_),
    .Y(_5687_)
);

FILL FILL_1__9395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10293_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [13]),
    .B(_6833__bF$buf2),
    .C(En_bF$buf2),
    .Y(_7064_)
);

INVX1 _14436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [4]),
    .Y(_6721_)
);

NOR2X1 _14016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_6202_),
    .Y(_6375_)
);

FILL FILL_1__7708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11078_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_3440_)
);

FILL FILL_0__8085_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3080_),
    .B(_3079_),
    .Y(_3081_)
);

FILL FILL_0__11852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11012_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [10]),
    .Y(_1760_)
);

OAI21X1 _8504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1399_),
    .C(_1400_),
    .Y(_1401_)
);

FILL FILL_1__7881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13224_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5386_),
    .B(_5392_),
    .C(_5390_),
    .Y(_5393_)
);

FILL FILL_0__12637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12217_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_5017_)
);

OAI21X1 _9709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1822_),
    .C(_2491_),
    .Y(_1723_)
);

FILL FILL_1__8666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14009_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6079_),
    .Y(_6080_)
);

FILL FILL_2__7110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7776_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2627_),
    .C(_2628_),
    .Y(_2629_)
);

FILL FILL_0__7356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2248_),
    .C(_2271_),
    .Y(_2272_)
);

MUX2X1 _9042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .B(_1867_),
    .S(_1810__bF$buf0),
    .Y(_1871_)
);

FILL FILL_1__11710_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4373_),
    .B(_4654_),
    .C(_4651_),
    .Y(_4657_)
);

FILL FILL_2__8315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13595_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6113_),
    .C(_6244_),
    .Y(_6245_)
);

FILL FILL_0__13175_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13460_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5060_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Xin12b [11])
);

NOR2X1 _13040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .B(_5504_),
    .Y(_5506_)
);

FILL FILL_1__12915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9502_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6888_),
    .B(_6891_),
    .Y(_6892_)
);

OAI21X1 _14245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_6555_),
    .C(_6556_),
    .Y(_7071_[9])
);

FILL FILL_1__7517_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3294_),
    .B(_3293_),
    .Y(_3295_)
);

OAI21X1 _10165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2624_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_2898_),
    .Y(_2524_)
);

FILL FILL_2__9693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11241_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1613_),
    .B(_1615_),
    .C(_1601_),
    .Y(_871_)
);

AND2X2 _8313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_1218_),
    .Y(_1219_)
);

FILL FILL_1__7690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12866_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5210_),
    .B(_5207_),
    .S(_5150__bF$buf0),
    .Y(_5211_)
);

FILL FILL_0__12446_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [0]),
    .B(_4348__bF$buf1),
    .Y(_4858_)
);

FILL FILL_0__12026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x190950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .B(_2678_),
    .C(_2649__bF$buf4),
    .Y(_2681_)
);

NAND2X1 _9518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .B(_2321_),
    .Y(_2325_)
);

FILL FILL_1__8475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert180 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert181 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert183 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6298_),
    .Y(_6299_)
);

FILL FILL_0_BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5895_),
    .B(_5898_),
    .C(_5892_),
    .Y(_5899_)
);

FILL FILL_0_BUFX2_insert185 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert186 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert188 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7585_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [1]),
    .Y(_2481_)
);

FILL FILL_0__7165_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2086_),
    .B(_2088_),
    .Y(_2089_)
);

FILL FILL_2__8964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9311_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14894_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6785_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.acc_reg [18])
);

NAND2X1 _14474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Y_ [1]),
    .B(_6724_),
    .Y(_6746_)
);

NOR2X1 _14054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6408_),
    .B(_6393_),
    .Y(_6411_)
);

FILL FILL_1__7746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13509_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3117_)
);

FILL FILL_0__11890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11050_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [8]),
    .Y(_1794_)
);

AOI22X1 _8542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(_996__bF$buf0),
    .C(_1437_),
    .D(_1434_),
    .Y(_858_)
);

NAND3X1 _8122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1009_),
    .B(_1026_),
    .C(_1034_),
    .Y(_1037_)
);

OAI21X1 _11599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4187_),
    .B(_4159_),
    .C(_3425_),
    .Y(_3418_)
);

AOI21X1 _11179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3822_),
    .B(_3821_),
    .C(_3512_),
    .Y(_3823_)
);

FILL FILL256650x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13262_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5426_),
    .B(_5428_),
    .Y(_5429_)
);

FILL FILL_0__12675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12255_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12540_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4194_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ycalc [3])
);

NAND3X1 _12120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(_4676_),
    .C(_4674_),
    .Y(_4677_)
);

OAI21X1 _9747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_2479_),
    .C(_2512_),
    .Y(_1740_)
);

NAND3X1 _9327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1859_),
    .B(_2140_),
    .C(_2137_),
    .Y(_2143_)
);

FILL FILL_1__8284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14047_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_6115_),
    .Y(_6116_)
);

OAI21X1 _13325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5776_),
    .B(_5726_),
    .C(_5775_),
    .Y(_5777_)
);

FILL FILL_0__14821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7394_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _9080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1904_),
    .Y(_1906_)
);

FILL FILL_2__8353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12179_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_779_),
    .Y(_781_)
);

FILL FILL_0__8599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11526_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .S(vdd),
    .Y(_4382_)
);

FILL FILL_0__9120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11106_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6584_),
    .B(_6587_),
    .Y(_6588_)
);

FILL FILL_1__7555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9701_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(_1645_),
    .Y(_1646_)
);

NAND2X1 _8351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .B(_1254_),
    .Y(_1255_)
);

FILL FILL_1__13071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12064_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.ISout ),
    .Y(_2718_)
);

INVX1 _9556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2359_)
);

NOR3X1 _9136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1938_),
    .C(_1910_),
    .Y(_1960_)
);

FILL FILL_1__8093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14276_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6293_),
    .B(_6290_),
    .Y(_6335_)
);

FILL FILL_0__13689_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5932_),
    .B(_5929_),
    .S(_5926__bF$buf0),
    .Y(_5933_)
);

FILL FILL_0__13269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .B(_5595_),
    .Y(_5596_)
);

FILL FILL_0__14630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert98 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6978_)
);

NAND2X1 _14339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6634_),
    .B(_6636_),
    .Y(_6637_)
);

FILL FILL_0__10970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10130_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_603_)
);

AOI21X1 _7202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_201_),
    .C(_160_),
    .Y(_203_)
);

OAI21X1 _10679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3235_),
    .B(_3324_),
    .C(_2589_),
    .Y(_2582_)
);

NAND2X1 _10259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2957_),
    .B(_2974_),
    .Y(_2988_)
);

FILL FILL_1__12762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9367_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11620_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3360_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[4].u_ce.Ycalc [7])
);

FILL FILL_0__11335_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3842_),
    .B(_3825_),
    .Y(_3843_)
);

NAND2X1 _14092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf0),
    .B(_6434_),
    .Y(_6447_)
);

OAI21X1 _8827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1645_),
    .C(_911_),
    .Y(_904_)
);

AOI21X1 _8407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1308_),
    .B(_1307_),
    .C(_998_),
    .Y(_1309_)
);

FILL FILL_1__7784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x136950 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5259_),
    .B(_5278_),
    .C(_5250_),
    .Y(_5300_)
);

OR2X2 _12405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4861_),
    .B(_4362__bF$buf4),
    .Y(_4945_)
);

FILL FILL_0__13901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9510_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1467_),
    .C(_1472_),
    .Y(_1473_)
);

NAND3X1 _8160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1033_),
    .C(_1051_),
    .Y(_1072_)
);

FILL FILL_2__7853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7259_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9785_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1697_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [8])
);

OR2X2 _9365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2175_),
    .B(_2178_),
    .Y(_2179_)
);

FILL FILL_0__8620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14085_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6138_),
    .B(_6151_),
    .C(_6152_),
    .Y(_6153_)
);

FILL FILL_0__13078_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5109_),
    .B(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5807_)
);

FILL FILL_2__13825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9405_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [2]),
    .Y(_6811_)
);

OAI21X1 _14148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6067_),
    .B(_6466_),
    .C(_6482_),
    .Y(_5879_)
);

FILL FILL_2__8391_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_810_)
);

OAI21X1 _7431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_420_),
    .C(_227_),
    .Y(_421_)
);

INVX1 _10488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3204_),
    .Y(_3205_)
);

OAI21X1 _10068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2804_),
    .B(_2789_),
    .C(_2741_),
    .Y(_2806_)
);

FILL FILL_1__12991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11144_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1524_),
    .B(gnd),
    .S(_1523_),
    .Y(_1525_)
);

AOI21X1 _8216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1121_),
    .C(_1114_),
    .Y(_1126_)
);

FILL FILL_1__7593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12769_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(\genblk1[6].u_ce.Ycalc [8]),
    .C(_5106_),
    .Y(_5119_)
);

FILL FILL_0__12349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4704_),
    .B(_4765_),
    .C(_4766_),
    .Y(_4767_)
);

FILL FILL_0__13710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6205_),
    .B(_6181_),
    .Y(_6206_)
);

OAI21X1 _13419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5728_),
    .B(_5807_),
    .C(_5097_),
    .Y(_5090_)
);

FILL FILL_0__14915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7488_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2393_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2395_)
);

OAI21X1 _9174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1994_),
    .C(_1995_),
    .Y(_1996_)
);

FILL FILL_1__11842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10835_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10700_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2526_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Ycalc [11])
);

FILL FILL_0__10415_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5969_),
    .B(_5966_),
    .S(_5926__bF$buf0),
    .Y(_5970_)
);

INVX1 _13172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5631_),
    .Y(_5632_)
);

OAI21X1 _7907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_810_),
    .C(_75_),
    .Y(_68_)
);

FILL FILL_2__13634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9634_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf1),
    .B(_4381_),
    .Y(_4471_)
);

FILL FILL_0__9214_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6901_),
    .B(_6891_),
    .Y(_7014_)
);

INVX1 _14377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [5]),
    .Y(_6669_)
);

FILL FILL_1__7649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14839_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_557_),
    .C(_585_),
    .Y(_639_)
);

NAND2X1 _7240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf0),
    .B(_189_),
    .Y(_238_)
);

OR2X2 _10297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3024_),
    .B(_3009_),
    .Y(_3025_)
);

FILL FILL_1__12380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11700_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8865_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_863_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Acalc [0])
);

AOI21X1 _8445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1343_),
    .B(_1344_),
    .C(_1018_),
    .Y(_1345_)
);

OAI21X1 _8025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(_943_),
    .C(_944_),
    .Y(_945_)
);

FILL FILL_2__7718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12998_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5270_),
    .B(_5334_),
    .C(_5335_),
    .Y(_5336_)
);

FILL FILL_0__12158_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4979_),
    .Y(_4980_)
);

INVX1 _12023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4578_),
    .Y(_4584_)
);

FILL FILL_2__12905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8187_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6022_),
    .Y(_6023_)
);

AOI21X1 _13228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5445_),
    .B(vdd),
    .C(_5683_),
    .Y(_5684_)
);

FILL FILL257250x122550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10224_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .Y(_691_)
);

FILL FILL_2__13863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11429_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Acalc [1]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Acalc [3]),
    .Y(_4291_)
);

FILL FILL_0__9023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11009_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14186_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5862_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Xin12b [8])
);

FILL FILL_1__7878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14228_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5389_),
    .C(_5388_),
    .Y(_5390_)
);

FILL FILL_2__10568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9604_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1079_),
    .C(_1010__bF$buf4),
    .Y(_1560_)
);

INVX1 _8254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1162_)
);

FILL FILL_1__10922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10502_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .Y(_4325__bF$buf0)
);

FILL FILL_2__7527_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert161 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 )
);

FILL FILL_2__7107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13394_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert162 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert164 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert166 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .Y(_972__bF$buf4)
);

BUFX2 BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .Y(_972__bF$buf3)
);

BUFX2 BUFX2_insert168 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .Y(_972__bF$buf2)
);

NAND2X1 _12672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5153_)
);

FILL FILL_0__12387_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert169 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .Y(_972__bF$buf1)
);

NAND2X1 _12252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4797_),
    .B(_4799_),
    .Y(_4803_)
);

FILL FILL_2__12714_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2624_),
    .C(_2625_),
    .Y(_2626_)
);

NAND2X1 _9459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2265_),
    .Y(_2269_)
);

MUX2X1 _9039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .S(gnd),
    .Y(_1868_)
);

FILL FILL_1__11707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14599_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6241_),
    .B(_6239_),
    .S(_5926__bF$buf1),
    .Y(_6242_)
);

DFFPOSX1 _13457_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5057_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Acalc [9])
);

NAND3X1 _13037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(_5502_),
    .C(_5500_),
    .Y(_5503_)
);

FILL FILL_0__14113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10033_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7945_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .CLK(clk_bF$buf9),
    .Q(\genblk1[0].u_ce.Acalc [4])
);

OR2X2 _7525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_495_),
    .Y(_511_)
);

INVX1 _7105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [9]),
    .Y(_110_)
);

FILL FILL_2__13672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9672_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4458_),
    .B(_4461_),
    .Y(_4507_)
);

FILL FILL_0__9252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11238_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4144_),
    .B(_4140_),
    .C(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Y(_4146_)
);

NAND2X1 _11103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3745_),
    .B(_3749_),
    .Y(_3750_)
);

FILL FILL_1__7687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14037_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .S(gnd),
    .Y(_5208_)
);

NOR2X1 _12308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4619_),
    .B(_4852_),
    .Y(_4855_)
);

FILL FILL_1__14811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf1),
    .B(_1380_),
    .C(_1375_),
    .Y(_1381_)
);

OAI21X1 _8063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_977_),
    .C(_978_),
    .Y(_979_)
);

FILL FILL_1__10311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4336_),
    .C(_5005_),
    .Y(_4237_)
);

AOI22X1 _12061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .B(_4618_),
    .C(_4619_),
    .D(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4620_)
);

FILL FILL_2__12943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12103_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_1761_),
    .Y(_2479_)
);

NAND2X1 _9268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .B(_2000_),
    .Y(_2086_)
);

FILL FILL_1__11936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6054_),
    .B(_6055_),
    .Y(_6060_)
);

AOI21X1 _13266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5445_),
    .B(vdd),
    .C(_5188__bF$buf4),
    .Y(_5720_)
);

FILL FILL_2__9902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10262_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_721_),
    .Y(_726_)
);

NAND3X1 _7334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf2),
    .B(_327_),
    .C(_323_),
    .Y(_328_)
);

FILL FILL_1__12894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11467_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _11752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_4324_)
);

FILL FILL_2__9079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3966_),
    .Y(_3969_)
);

OAI21X1 _8959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1788_),
    .B(_1791_),
    .C(_1768_),
    .Y(_1792_)
);

NOR2X1 _8539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1410_),
    .Y(_1435_)
);

OAI21X1 _8119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1008_),
    .C(_1033_),
    .Y(_1034_)
);

FILL FILL_1__7496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14266_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Xcalc [1]),
    .C(_2644_),
    .D(_2606_),
    .Y(_2645_)
);

FILL FILL_1__13679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .B(_5340_),
    .Y(_5426_)
);

DFFPOSX1 _12537_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4191_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ycalc [1])
);

NAND3X1 _12117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf1),
    .B(_4673_),
    .C(_4664_),
    .Y(_4674_)
);

FILL FILL_1__14620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x147750 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1198_),
    .C(_998_),
    .Y(_1199_)
);

FILL FILL_1__10960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7565_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4838_),
    .B(_4835_),
    .Y(_4839_)
);

FILL FILL_2__12752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1911_),
    .B(_2304_),
    .Y(_2305_)
);

OAI21X1 _9077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1903_),
    .C(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .Y(_1904_)
);

FILL FILL_1__11745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8332_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672__bF$buf3),
    .B(_3310_),
    .C(_3309_),
    .Y(_2550_)
);

FILL FILL_0__10318_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13495_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.LoadCtl [0])
);

OAI21X1 _13075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5519_),
    .B(_5538_),
    .C(_5188__bF$buf3),
    .Y(_5539_)
);

FILL FILL_2__13537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9537_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .S(vdd),
    .Y(_4379_)
);

FILL FILL_0__9117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10071_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7983_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_67_),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.Ain12b [4])
);

NAND2X1 _7563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_546_),
    .Y(_547_)
);

OAI21X1 _7143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_143_),
    .C(_144_),
    .Y(_145_)
);

FILL FILL_1__12283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11696_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4542_),
    .C(_4543_),
    .Y(_4544_)
);

FILL FILL_0__9290_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3737_),
    .B(_4151_),
    .C(_4169_),
    .Y(_3401_)
);

FILL FILL_0__11276_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3786_)
);

OAI21X1 _8768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Xin12b [9]),
    .Y(_1644_)
);

INVX1 _8348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .Y(_1252_)
);

FILL FILL_2__14075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13068_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5243_),
    .C(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .Y(_5244_)
);

OAI21X1 _12346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf0),
    .B(_4889_),
    .C(_4362__bF$buf5),
    .Y(_4890_)
);

FILL FILL_0__13842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9031_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[2]),
    .Y(Dout[2])
);

FILL FILL_0__14627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8561_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3488_),
    .C(_3489_),
    .Y(_3490_)
);

FILL FILL_0__8141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10127_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3131_),
    .B(_3116_),
    .Y(_3134_)
);

FILL FILL_2__9940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9100_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_595_),
    .C(_591_),
    .Y(_600_)
);

FILL FILL_2__13346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9346_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11617_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3357_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Ycalc [4])
);

FILL FILL_1__13700_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [11]),
    .B(_5949__bF$buf0),
    .Y(_6444_)
);

FILL FILL_1__8722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8302_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_760_),
    .C(_158__bF$buf4),
    .Y(_762_)
);

AND2X2 _7372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_335_),
    .Y(_364_)
);

FILL FILL_1__12092_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4361_)
);

FILL FILL_0__11085_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3985_),
    .B(_3510__bF$buf3),
    .C(_4004_),
    .D(_3508_),
    .Y(_3375_)
);

FILL FILL_1__9927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9507_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1826_),
    .Y(_1827_)
);

OAI21X1 _8577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(_1469_),
    .C(_1457_),
    .Y(_860_)
);

OAI21X1 _8157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1057_),
    .B(_1045_),
    .C(_1058_),
    .Y(_1069_)
);

FILL FILL_1__10825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5162_),
    .B(_5459_),
    .Y(_5462_)
);

DFFPOSX1 _12575_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4229_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Xin12b [8])
);

OAI21X1 _12155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4626_),
    .C(_4709_),
    .Y(_4710_)
);

FILL FILL_2__12617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14436_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6942_),
    .B(_6943_),
    .Y(_6944_)
);

FILL FILL_0__14016_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [7]),
    .Y(_6603_)
);

FILL FILL_2__12370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8370_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_3334_)
);

FILL FILL_0__10356_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2945_),
    .B(_2951_),
    .Y(_2952_)
);

OAI21X1 _7848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_807_),
    .C(_808_),
    .Y(_41_)
);

INVX1 _7428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .Y(_418_)
);

FILL FILL_2__13575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9575_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4409_),
    .B(_4411_),
    .C(_4397_),
    .Y(_4415_)
);

FILL FILL_0__9155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4050_),
    .B(_4054_),
    .Y(_4056_)
);

NAND3X1 _11006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3653_),
    .C(_3648_),
    .Y(_3657_)
);

FILL FILL_0__12922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14714_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_180_),
    .C(_181_),
    .Y(_182_)
);

FILL FILL_0__13707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9316_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1009_),
    .C(_1287_),
    .Y(_1288_)
);

FILL FILL_1__10634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4919_),
    .B(_4924_),
    .Y(_4925_)
);

FILL FILL_0__12099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8006_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [5]),
    .Y(_5967_)
);

NAND2X1 _13169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5623_),
    .B(_5625_),
    .Y(_5629_)
);

FILL FILL_0__14665_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14530_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6518_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin12b [4])
);

FILL FILL_0__14245_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [1]),
    .Y(_6461_)
);

FILL FILL_1__7802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11172_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3525_),
    .C(_3526_),
    .Y(_3527_)
);

FILL FILL_0__10585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10165_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf5),
    .B(_3157_),
    .Y(_3170_)
);

INVX1 _10030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2769_)
);

FILL FILL_2__10912_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_614_),
    .Y(_636_)
);

INVX1 _7237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .Y(_235_)
);

FILL FILL_2__13384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9384_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11655_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3395_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [4])
);

OR2X2 _11235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3875_),
    .B(_3873_),
    .Y(_3876_)
);

FILL FILL_0__12731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14589_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9803_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1715_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin12b [8])
);

FILL FILL_1__8760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13936_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6162_),
    .C(_6164_),
    .Y(_6170_)
);

FILL FILL_0__13516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1093_),
    .B(_1105_),
    .C(_1103_),
    .Y(_1106_)
);

FILL FILL_1__10863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7450_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4711_),
    .B(_4732_),
    .C(_4715_),
    .Y(_4746_)
);

FILL FILL_2__12655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8655_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3580_),
    .B(_3578_),
    .C(_3558_),
    .Y(_3355_)
);

FILL FILL_0__8235_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3211_),
    .B(_3220_),
    .C(_3221_),
    .Y(_3222_)
);

NAND2X1 _13398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5826_)
);

FILL FILL_0__14474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10301_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(gnd),
    .Y(_829_)
);

OAI21X1 _7466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_322_),
    .C(_453_),
    .Y(_454_)
);

FILL FILL_2__13193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11599_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf2),
    .B(_4353_),
    .Y(_4451_)
);

FILL FILL_0__9193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3516_),
    .C(_3486__bF$buf3),
    .Y(_4091_)
);

INVX1 _11044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3693_),
    .Y(_3694_)
);

FILL FILL_0__12960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2410_),
    .Y(_2411_)
);

INVX8 _12669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_5150_)
);

NAND2X1 _12249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

FILL FILL_1__14752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13745_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5987_),
    .B(_5979_),
    .C(_5962_),
    .Y(_5988_)
);

FILL FILL_0__13325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10252_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [17]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf2),
    .Y(_7031_)
);

FILL FILL_2__7277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8044_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10735_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2561_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Xin0 [0])
);

OR2X2 _10315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .B(_3034_),
    .Y(_3042_)
);

FILL FILL_0__11811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert111 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert112 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert114 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert116 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert118 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert119 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10110_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_671_)
);

FILL FILL_1__14808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_268_),
    .Y(_272_)
);

INVX2 _11693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4271_)
);

NAND3X1 _11273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3911_),
    .C(_3908_),
    .Y(_3912_)
);

FILL FILL_2__11315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7735_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9841_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[2].u_ce.LoadCtl [4])
);

FILL FILL_0__7315_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2218_),
    .C(_2201_),
    .Y(_2232_)
);

OAI21X1 _9001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1830_),
    .C(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .Y(_1831_)
);

OAI21X1 _12898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5368_),
    .C(_5369_),
    .Y(_5370_)
);

OAI21X1 _12478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_5004_)
);

NAND2X1 _12058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4616_),
    .Y(_4617_)
);

FILL FILL_1__14561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [2]),
    .B(_6833__bF$buf4),
    .Y(_6855_)
);

DFFPOSX1 _14204_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5880_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Yin1 [0])
);

FILL FILL_2__7086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8693_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3616_),
    .B(_3615_),
    .Y(_3617_)
);

FILL FILL_0__8273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10679_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3256_),
    .B(_3255_),
    .Y(_3257_)
);

FILL FILL_0__10259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2821_),
    .B(_2850_),
    .C(_2849_),
    .Y(_2859_)
);

FILL FILL_0__11200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9478_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4273_),
    .C(_4321_),
    .Y(\genblk1[5].u_ce.X_ [1])
);

FILL FILL_0__9058_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3965_),
    .B(_3964_),
    .C(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3966_)
);

FILL FILL_1__13832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14617_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_92_)
);

NAND3X1 _11082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf3),
    .B(_3727_),
    .C(_3724_),
    .Y(_3730_)
);

FILL FILL_1__9639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11544_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .B(_1195_),
    .C(_1194_),
    .Y(_1196_)
);

FILL FILL_1__10957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7544_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2422_),
    .Y(_2447_)
);

FILL FILL_0__7124_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_2049_),
    .C(_2048_),
    .Y(_2050_)
);

AND2X2 _12287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4832_),
    .B(_4830_),
    .Y(_4836_)
);

FILL FILL_2__8503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14568_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6822_),
    .B(_6833__bF$buf3),
    .C(_7062_),
    .Y(_6790_)
);

FILL FILL_0__14148_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [1]),
    .Y(_6718_)
);

INVX1 _14013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [7]),
    .Y(_6372_)
);

FILL FILL_1__7705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x248550 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _10773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .Y(_3437_)
);

FILL FILL_0__8082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10068_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3074_),
    .B(_3077_),
    .Y(_3078_)
);

FILL FILL_2__10815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9881_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _8921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1757_)
);

NAND3X1 _8501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf1),
    .B(_1397_),
    .C(_1394_),
    .Y(_1398_)
);

NAND3X1 _11978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4540_),
    .C(_4539_),
    .Y(_4541_)
);

FILL FILL_0__9287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.X_ [1]),
    .Y(_4168_)
);

NAND3X1 _11138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf1),
    .B(_3779_),
    .C(_3782_),
    .Y(_3783_)
);

FILL FILL_1__13641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12214_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_2490_)
);

FILL FILL_1__8663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13839_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6075_),
    .C(_6076_),
    .Y(_6077_)
);

FILL FILL_0__13419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11353_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1011_),
    .C(_1012_),
    .Y(_1013_)
);

FILL FILL_1__10346_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[1]),
    .Y(Dout[1])
);

FILL FILL_0__7773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7353_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4633_),
    .C(_4653_),
    .Y(_4654_)
);

FILL FILL_2__8732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8558_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _10829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_3487_)
);

FILL FILL_0__8138_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3131_),
    .B(_3116_),
    .C(_2670_),
    .Y(_3132_)
);

FILL FILL_1__12912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6889_)
);

OAI21X1 _14242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_6553_),
    .C(_6554_),
    .Y(_7071_[8])
);

FILL FILL_1__7514_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3288_),
    .B(_3283_),
    .C(_3281_),
    .Y(_3292_)
);

FILL FILL_0__10297_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2883_),
    .B(_2895_),
    .Y(_2896_)
);

FILL FILL_1__8719_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_756_),
    .Y(_759_)
);

OAI21X1 _7369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_360_),
    .C(_361_),
    .Y(_362_)
);

FILL FILL_2__13096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_1612_),
    .Y(_1613_)
);

NAND3X1 _8310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf0),
    .B(_1213_),
    .C(_1210_),
    .Y(_1216_)
);

FILL FILL_1__12089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(vdd),
    .C(_4325__bF$buf3),
    .Y(_4358_)
);

FILL FILL_0__9096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3990_),
    .B(_4001_),
    .Y(_4002_)
);

FILL FILL_1__13870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7829_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _9935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_2678_)
);

FILL FILL_0__7409_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2316_),
    .Y(_2322_)
);

FILL FILL_1__8472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert152 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13648_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6295_),
    .B(_6294_),
    .Y(_6296_)
);

FILL FILL_0_BUFX2_insert154 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert155 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [4]),
    .Y(_5896_)
);

FILL FILL_0__13228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert157 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert159 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6940_),
    .B(_6939_),
    .Y(_6941_)
);

FILL FILL_0__7582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8367_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3313_),
    .Y(_3332_)
);

OAI21X1 _10218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2769_),
    .C(_2948_),
    .Y(_2949_)
);

FILL FILL_1__12721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9326_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14891_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6782_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [15])
);

OAI21X1 _14471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6566_),
    .C(_6744_),
    .Y(_6523_)
);

OAI21X1 _14051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6408_),
    .B(_6393_),
    .C(_5947_),
    .Y(_6409_)
);

FILL FILL_1__7743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12919_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3079_),
    .B(_3109_),
    .C(_3105_),
    .Y(_3114_)
);

FILL FILL_1__8948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10013_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_580_),
    .Y(_19_)
);

MUX2X1 _7178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_175_),
    .S(_135__bF$buf3),
    .Y(_179_)
);

NAND2X1 _11596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [6]),
    .B(_4159_),
    .Y(_4189_)
);

AND2X2 _11176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3818_),
    .B(_3819_),
    .Y(_3820_)
);

FILL FILL_0__12672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7638_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_2479_),
    .C(_2510_),
    .Y(_1739_)
);

FILL FILL_0__7218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2119_),
    .C(_2139_),
    .Y(_2140_)
);

FILL FILL_1__8281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13877_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .Y(_6113_)
);

NOR2X1 _13322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5764_),
    .B(_5752_),
    .Y(_5774_)
);

FILL FILL_0__13037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10384_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14527_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6515_),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.Xin12b [9])
);

OR2X2 _14107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6454_),
    .B(_5888_),
    .Y(_6459_)
);

FILL FILL_0__7391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8350_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_769_),
    .C(_767_),
    .Y(_778_)
);

FILL FILL_1__11589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8596_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _10867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_3524_)
);

FILL FILL_0__8176_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [11]),
    .B(_2672__bF$buf2),
    .Y(_3167_)
);

OAI21X1 _10027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2746_),
    .B(_2765_),
    .C(_2766_),
    .Y(_2767_)
);

FILL FILL_1__12950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11103_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [4]),
    .Y(_6585_)
);

FILL FILL_1__7552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7867_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_2666_),
    .Y(_2716_)
);

FILL FILL_0__7447_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .B(_2355_),
    .Y(_2357_)
);

NAND2X1 _9133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf4),
    .B(_1867_),
    .Y(_1957_)
);

FILL FILL_1__8090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14273_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_6330_),
    .C(_6331_),
    .Y(_6332_)
);

FILL FILL_0__13686_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .Y(_5930_)
);

FILL FILL_0__13266_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .B(_5591_),
    .C(_5592_),
    .Y(_5593_)
);

FILL FILL_1__9295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10193_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [13]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf2),
    .Y(_6976_)
);

NAND2X1 _14336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .B(_6633_),
    .Y(_6634_)
);

FILL FILL_1__7608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [0]),
    .B(_3324_),
    .Y(_2588_)
);

OAI21X1 _10256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672__bF$buf4),
    .B(_2985_),
    .C(_2959_),
    .Y(_2528_)
);

FILL FILL_0__11752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [6]),
    .B(_1645_),
    .Y(_1675_)
);

AND2X2 _8404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1304_),
    .B(_1305_),
    .Y(_1306_)
);

FILL FILL_1__7781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12957_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf0),
    .B(_5207_),
    .Y(_5297_)
);

FILL FILL_0__12117_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4934_),
    .B(_4939_),
    .Y(_4942_)
);

OAI22X1 _9609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1773_),
    .B(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .C(_2406_),
    .D(_2408_),
    .Y(_1706_)
);

FILL FILL_1__8986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14329_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5984_),
    .B(_5983_),
    .S(_5926__bF$buf0),
    .Y(_5985_)
);

FILL FILL_2__11256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7256_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9782_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1694_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [5])
);

NAND2X1 _9362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_2124_),
    .Y(_2176_)
);

FILL FILL_1__11610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x190950 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6146_),
    .B(_6149_),
    .Y(_6150_)
);

FILL FILL_0__13075_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5799_),
    .B(_5804_),
    .C(_5805_),
    .Y(_5063_)
);

FILL FILL_1__12815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9402_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6801_),
    .B(_6802_),
    .C(_6807_),
    .Y(_6808_)
);

NAND2X1 _14145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [0]),
    .B(_6466_),
    .Y(_6481_)
);

FILL FILL_1__7837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain1 [0]),
    .B(_3201_),
    .Y(_3202_)
);

INVX1 _10065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2802_),
    .Y(_2803_)
);

FILL FILL_0__11981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11141_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1521_),
    .B(_1514_),
    .C(_1519_),
    .Y(_1522_)
);

INVX1 _8213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1120_),
    .Y(_1123_)
);

FILL FILL_1__7590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12766_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Acalc [1]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Acalc [3]),
    .Y(_5117_)
);

FILL FILL_0__12346_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4717_),
    .B(_4720_),
    .Y(_4764_)
);

DFFPOSX1 _9838_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.LoadCtl [1])
);

OAI21X1 _9418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2228_),
    .B(_2229_),
    .C(_1832_),
    .Y(_2230_)
);

FILL FILL_1__8795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14138_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [11]),
    .B(_6202_),
    .Y(_6203_)
);

NAND2X1 _13416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [0]),
    .B(_5807_),
    .Y(_5096_)
);

FILL FILL_0__14912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7485_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2390_),
    .Y(_2392_)
);

AND2X2 _9171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1944_),
    .B(_1947_),
    .Y(_1993_)
);

FILL FILL_0__10832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10412_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [0]),
    .B(_810_),
    .Y(_74_)
);

FILL FILL_1__12624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9631_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4468_)
);

FILL FILL_2__9229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9211_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_7011_)
);

FILL FILL_0__14089_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6666_),
    .C(_6661_),
    .Y(_6667_)
);

FILL FILL_1__7646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13409_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3021_),
    .Y(_3022_)
);

FILL FILL_0__11790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11370_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8862_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_860_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Xcalc [9])
);

OAI21X1 _8442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .B(_1312_),
    .C(_1010__bF$buf2),
    .Y(_1342_)
);

AOI21X1 _8022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_940_),
    .C(_941_),
    .Y(_942_)
);

AOI21X1 _11499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4123_),
    .B(_4088_),
    .C(_4122_),
    .Y(_4124_)
);

INVX1 _11079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3725_),
    .Y(_3727_)
);

FILL FILL_2__7715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12995_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5284_),
    .B(_5287_),
    .Y(_5333_)
);

INVX1 _12440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4976_),
    .Y(_4977_)
);

FILL FILL_0__12155_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4576_),
    .Y(_4581_)
);

AOI21X1 _9647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2441_),
    .B(_2377_),
    .C(\genblk1[2].u_ce.Ain12b [8]),
    .Y(_2444_)
);

NOR3X1 _9227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_2026_),
    .C(_1999_),
    .Y(_2047_)
);

FILL FILL_1__8184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14367_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [3]),
    .Y(_6020_)
);

NAND2X1 _13225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [1]),
    .B(_5174__bF$buf0),
    .Y(_5681_)
);

FILL FILL_0__14721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain1 [0]),
    .B(_687_),
    .Y(_688_)
);

FILL FILL_0__8499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11426_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [7]),
    .B(_4279_),
    .Y(_4288_)
);

FILL FILL_2__9038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11006_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14183_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5859_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [11])
);

DFFPOSX1 _8918_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.LoadCtl [5])
);

FILL FILL_1__7875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5343_),
    .B(_5366_),
    .C(_5339_),
    .Y(_5387_)
);

FILL FILL_1__9601_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1556_),
    .C(_1547_),
    .Y(_867_)
);

AOI21X1 _8251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1142_),
    .C(_1154_),
    .Y(_1159_)
);

BUFX2 BUFX2_insert130 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 )
);

FILL FILL_2__7524_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert131 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .Y(_3487__bF$buf4)
);

BUFX2 BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .Y(_3487__bF$buf3)
);

FILL FILL_1__13391_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert133 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .Y(_3487__bF$buf2)
);

BUFX2 BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .Y(_3487__bF$buf1)
);

BUFX2 BUFX2_insert135 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .Y(_3487__bF$buf0)
);

BUFX2 BUFX2_insert136 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf4)
);

BUFX2 BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf3)
);

BUFX2 BUFX2_insert138 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf2)
);

FILL FILL_0__12384_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf1)
);

NAND2X1 _9876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2622_),
    .Y(\genblk1[3].u_ce.Y_ [0])
);

NAND2X1 _9456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2264_),
    .B(_2265_),
    .Y(_2266_)
);

MUX2X1 _9036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .S(gnd),
    .Y(_1865_)
);

FILL FILL_1__11704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14596_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6024_),
    .C(_6238_),
    .Y(_6239_)
);

FILL FILL_0__13589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13169_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13454_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5054_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Acalc [3])
);

NAND3X1 _13034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf3),
    .B(_5499_),
    .C(_5490_),
    .Y(_5500_)
);

FILL FILL_2__13916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10096_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6878_),
    .B(_6884_),
    .C(_6885_),
    .Y(_6886_)
);

OAI21X1 _14239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_6551_),
    .C(_6552_),
    .Y(_7071_[7])
);

FILL FILL_0__10870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10030_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7942_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[0].u_ce.Acalc [1])
);

INVX1 _7522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .Y(_508_)
);

OAI21X1 _7102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_107_),
    .C(_92_),
    .Y(_108_)
);

NAND2X1 _10999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf0),
    .B(_3561_),
    .Y(_3650_)
);

NAND2X1 _10579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3283_),
    .B(_3288_),
    .Y(_3290_)
);

OAI21X1 _10159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2885_),
    .C(_2887_),
    .Y(_2893_)
);

FILL FILL_1__12662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4484_),
    .B(_4348__bF$buf4),
    .C(_4504_),
    .D(_4420_),
    .Y(_4197_)
);

FILL FILL_2__9267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11235_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .B(_3524__bF$buf4),
    .Y(_4143_)
);

AND2X2 _11100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3741_),
    .B(_3524__bF$buf3),
    .Y(_3747_)
);

AOI21X1 _8727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1609_),
    .B(_1574_),
    .C(_1608_),
    .Y(_1610_)
);

INVX1 _8307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1211_),
    .Y(_1213_)
);

FILL FILL_1__7684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13027_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .S(gnd),
    .Y(_5205_)
);

OAI21X1 _12305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4325__bF$buf3),
    .C(_4344_),
    .Y(_4852_)
);

FILL FILL_0__13801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9410_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf4),
    .B(_1297_),
    .Y(_1378_)
);

OAI21X1 _8060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_974_),
    .C(_975_),
    .Y(_976_)
);

FILL FILL_2__7753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7579_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2475_),
    .Y(_2477_)
);

FILL FILL_0__7159_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1778_),
    .B(_1834__bF$buf4),
    .C(_2083_),
    .D(_1906_),
    .Y(_1687_)
);

FILL FILL_1__11933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6034_),
    .B(_6025_),
    .Y(_6057_)
);

FILL FILL_0__13398_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5707_),
    .B(_5716_),
    .C(_5717_),
    .Y(_5718_)
);

FILL FILL_2__13725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9305_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14888_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6779_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.acc_reg [12])
);

NAND2X1 _14468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.X_ [0]),
    .Y(_6743_)
);

OAI21X1 _14048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6405_),
    .C(_6393_),
    .Y(_6406_)
);

FILL FILL_2__8291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(_154_),
    .Y(_723_)
);

NOR2X1 _7331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf4),
    .B(_324_),
    .Y(_325_)
);

INVX1 _10388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3109_),
    .Y(_3112_)
);

FILL FILL_1__12891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11044_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [5]),
    .Y(_1789_)
);

NAND3X1 _8536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(_1430_),
    .C(_1431_),
    .Y(_1432_)
);

MUX2X1 _8116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(\genblk1[1].u_ce.Xin0 [1]),
    .S(vdd),
    .Y(_1031_)
);

FILL FILL_1__7493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13256_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5118_),
    .B(_5174__bF$buf2),
    .C(_5423_),
    .D(_5246_),
    .Y(_5039_)
);

FILL FILL_0__12669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[5] [1]),
    .Y(_4269_)
);

NAND2X1 _12114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4669_),
    .B(_4670_),
    .Y(_4671_)
);

FILL FILL_0__13610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8278_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6100_),
    .B(_6078_),
    .C(_6079_),
    .Y(_6110_)
);

AOI21X1 _13319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5768_),
    .B(_5711_),
    .C(\genblk1[6].u_ce.Ain12b [8]),
    .Y(_5771_)
);

FILL FILL_1_CLKBUF1_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2299_),
    .Y(_2302_)
);

OAI21X1 _9074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1895_),
    .B(_1897_),
    .C(_1883_),
    .Y(_1901_)
);

FILL FILL_1__11742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8767_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3308_),
    .B(_3307_),
    .C(_3298_),
    .Y(_2549_)
);

FILL FILL_0__10315_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13492_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5092_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain1 [1])
);

OAI21X1 _13072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5452_),
    .C(_5535_),
    .Y(_5536_)
);

NAND2X1 _7807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_774_),
    .Y(_776_)
);

FILL FILL_2__13954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x122550 (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4375_),
    .B(_4372_),
    .S(_4325__bF$buf4),
    .Y(_4376_)
);

FILL FILL_0__9114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6921_),
    .B(_6920_),
    .Y(_6922_)
);

NOR2X1 _14277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin1 [0]),
    .B(\u_ot.Xin1 [1]),
    .Y(_6582_)
);

FILL FILL_1__7549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14739_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7980_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_64_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Ain12b [9])
);

NOR2X1 _7560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_499_),
    .Y(_544_)
);

MUX2X1 _7140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_138_),
    .S(_135__bF$buf3),
    .Y(_142_)
);

NAND2X1 _10197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2928_),
    .B(_2904_),
    .Y(_2929_)
);

FILL FILL_1__12280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11273_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1642_)
);

INVX1 _8345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1249_)
);

FILL FILL_2__14492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12898_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5235_),
    .B(_5237_),
    .C(_5223_),
    .Y(_5241_)
);

FILL FILL_0__12478_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4886_),
    .Y(_4887_)
);

FILL FILL_0__12058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8805_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_6202_),
    .Y(_6329_)
);

INVX1 _13548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .Y(_5927_)
);

AND2X2 _13128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5543_),
    .B(_5546_),
    .Y(_5590_)
);

FILL FILL_0__14624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10124_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_598_)
);

FILL FILL_2__13763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11329_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11614_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3354_),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[4].u_ce.ISout )
);

NOR2X1 _14086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6440_),
    .B(_6429_),
    .Y(_6442_)
);

FILL FILL_1__7778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5294_)
);

FILL FILL_2__10468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9504_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1822_),
    .C(_1823_),
    .Y(_1824_)
);

NAND2X1 _8574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1465_),
    .B(_1467_),
    .Y(_1468_)
);

OAI21X1 _8154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(_1064_),
    .C(_1044_),
    .Y(_841_)
);

FILL FILL_1__10822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5162_),
    .B(_5459_),
    .C(_5172_),
    .Y(_5460_)
);

DFFPOSX1 _12572_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4226_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [11])
);

FILL FILL_0__12287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4706_),
    .Y(_4707_)
);

DFFPOSX1 _9779_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1691_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Xcalc [2])
);

OAI21X1 _9359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2046_),
    .C(_2172_),
    .Y(_2173_)
);

FILL FILL_1__11607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf3),
    .B(_6144_),
    .C(_6140_),
    .Y(_6147_)
);

OAI21X1 _13357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5802_),
    .B(_5800_),
    .C(_5803_),
    .Y(_5062_)
);

FILL FILL_0__14853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x198150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10353_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_803_),
    .C(_806_),
    .Y(_40_)
);

NAND2X1 _7425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_390_),
    .Y(_415_)
);

FILL FILL_2__13992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11558_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4411_),
    .B(_4409_),
    .Y(_4412_)
);

FILL FILL_0__9152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11138_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4053_)
);

OAI21X1 _11003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3634_),
    .B(_3629_),
    .C(_3524__bF$buf3),
    .Y(_3654_)
);

FILL FILL_1__7587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14777_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Acalc [7]),
    .B(_5108_),
    .Y(_5114_)
);

NAND2X1 _12208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4740_),
    .B(_4760_),
    .Y(_4761_)
);

FILL FILL_1__14711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9313_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1285_)
);

FILL FILL_1__10631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7236_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _12381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4287_),
    .B(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .C(_4920_),
    .D(_4922_),
    .Y(_4220_)
);

FILL FILL_0__12096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12003_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2348_),
    .C(_2388_),
    .Y(_2389_)
);

AOI22X1 _9168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .B(_1834__bF$buf3),
    .C(_1990_),
    .D(_1906_),
    .Y(_1683_)
);

FILL FILL_1__11836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10409_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .Y(_5964_)
);

NAND2X1 _13166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5622_),
    .B(_5625_),
    .Y(_5626_)
);

FILL FILL_2__13208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10162_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [10]),
    .Y(_633_)
);

INVX1 _7234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .Y(_232_)
);

FILL FILL_1__12794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9381_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11652_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3392_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [9])
);

FILL FILL_0__11367_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .Y(_3873_)
);

DFFPOSX1 _8859_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_857_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Xcalc [6])
);

NAND2X1 _8439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1078_),
    .Y(_1339_)
);

NAND2X1 _8019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_939_),
    .B(_938_),
    .Y(\a[2] [1])
);

FILL FILL_1__7396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13999_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9800_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1712_),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[2].u_ce.Acalc [11])
);

FILL FILL_1__13579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13159_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5310_),
    .B(_5174__bF$buf2),
    .C(_5330_),
    .D(_5246_),
    .Y(_5035_)
);

NAND2X1 _12437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [10]),
    .B(_4348__bF$buf3),
    .Y(_4974_)
);

AOI21X1 _12017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4561_),
    .B(_4565_),
    .C(_4577_),
    .Y(_4578_)
);

FILL FILL_1__14100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9122_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1101_),
    .Y(_1103_)
);

FILL FILL_1__10860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7465_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4742_),
    .B(_4743_),
    .C(_4346_),
    .Y(_4744_)
);

FILL FILL_2__12652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12232_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2208_),
    .Y(_2210_)
);

FILL FILL_1__11225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8652_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3576_),
    .B(_3577_),
    .C(_3512_),
    .Y(_3578_)
);

FILL FILL_0__8232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10638_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3218_),
    .Y(_3219_)
);

FILL FILL_0__10218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5816_),
    .B(_5104_),
    .C(_5824_),
    .Y(_5079_)
);

FILL FILL_2__13017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9437_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Acalc [11]),
    .C(_4276_),
    .Y(_4285_)
);

FILL FILL_0__9017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8813_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_83_),
    .C(_827_),
    .Y(_57_)
);

MUX2X1 _7463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(_448_),
    .S(_135__bF$buf1),
    .Y(_451_)
);

FILL FILL_1__12183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11596_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4446_),
    .C(_4447_),
    .Y(_4448_)
);

FILL FILL_0__9190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11176_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4066_),
    .B(_4080_),
    .C(_4078_),
    .Y(_4088_)
);

OAI21X1 _11041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3660_),
    .B(_3664_),
    .C(_3659_),
    .Y(_3691_)
);

FILL FILL_2__11503_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .B(_1542_),
    .C(_1541_),
    .Y(_1555_)
);

NAND3X1 _8248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1127_),
    .C(_1155_),
    .Y(_1156_)
);

FILL FILL_1__10916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5142_),
    .B(_5104_),
    .C(_5147_),
    .Y(\genblk1[6].u_ce.X_ [1])
);

INVX1 _12246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4796_),
    .Y(_4797_)
);

FILL FILL_0__13742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9351_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7027_),
    .B(_7026_),
    .Y(_7028_)
);

FILL FILL_0__14107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8041_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10732_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2558_),
    .CLK(clk_bF$buf50),
    .Q(\genblk1[3].u_ce.Xin12b [5])
);

FILL FILL_0__10447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10027_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3017_),
    .B(_3036_),
    .Y(_3039_)
);

DFFPOSX1 _7939_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [10])
);

FILL FILL_2__9000_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_503_),
    .Y(_505_)
);

FILL FILL_2__13246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9666_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4501_),
    .Y(_4502_)
);

FILL FILL_0__9246_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4139_),
    .C(_4137_),
    .Y(_4140_)
);

FILL FILL_1__13600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8202_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158__bF$buf4),
    .B(_667_),
    .C(_668_),
    .Y(_25_)
);

FILL FILL_1__14805_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_264_),
    .Y(_269_)
);

DFFPOSX1 _11690_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.LoadCtl [5])
);

AOI21X1 _11270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf1),
    .B(_3868_),
    .C(_3890_),
    .Y(_3909_)
);

FILL FILL_1__9407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8897_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_895_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Yin1 [0])
);

NAND2X1 _8477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1363_),
    .Y(_1375_)
);

FILL FILL_0_CLKBUF1_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _8057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_973_)
);

FILL FILL_0_CLKBUF1_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5366_),
    .C(_5365_),
    .Y(_5367_)
);

OAI21X1 _12475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4366_),
    .B(_5000_),
    .C(_5002_),
    .Y(_4234_)
);

INVX1 _12055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4614_)
);

FILL FILL_0__13971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14336_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6851_),
    .B(_6848_),
    .Y(_6852_)
);

DFFPOSX1 _14201_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5877_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Yin12b [7])
);

FILL FILL_2__12270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8690_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf4),
    .B(_3612_),
    .C(_3613_),
    .Y(_3614_)
);

FILL FILL_0__8270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10676_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .B(_3213_),
    .Y(_3254_)
);

FILL FILL_0__10256_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2854_),
    .B(_2852_),
    .C(_2856_),
    .Y(_2857_)
);

OAI21X1 _7748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_717_),
    .C(_714_),
    .Y(_720_)
);

INVX1 _7328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_322_)
);

FILL FILL_2__13055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9475_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.Xcalc [5]),
    .C(_4279_),
    .D(\genblk1[5].u_ce.Xcalc [7]),
    .Y(_4319_)
);

FILL FILL_0__9055_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3962_),
    .B(_3960_),
    .C(_3955_),
    .Y(_3963_)
);

FILL FILL_0__12822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14614_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(\genblk1[0].u_ce.LoadCtl [3]),
    .Y(_89_)
);

FILL FILL_0__13607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9216_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1186_),
    .B(_1192_),
    .C(_1189_),
    .Y(_1193_)
);

FILL FILL_1__10954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7121_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4830_),
    .B(_4832_),
    .Y(_4833_)
);

FILL FILL_0__13780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8326_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13489_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5089_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain12b [4])
);

NAND2X1 _13069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5532_),
    .Y(_5533_)
);

FILL FILL_2__9705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14565_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [10]),
    .B(_6833__bF$buf1),
    .C(En_bF$buf0),
    .Y(_7061_)
);

FILL FILL_0__14145_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6710_),
    .B(_6715_),
    .Y(_6716_)
);

OAI21X1 _14010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6369_),
    .B(_6363_),
    .C(_6018_),
    .Y(_6370_)
);

FILL FILL_1__7702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11072_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3433_),
    .Y(_3434_)
);

FILL FILL_0__10485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10065_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _10350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .B(_3055_),
    .C(_3059_),
    .Y(_3075_)
);

FILL FILL_2__10812_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7977_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_61_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ain12b [10])
);

OAI21X1 _7557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf0),
    .B(_539_),
    .C(_540_),
    .Y(_541_)
);

INVX1 _7137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .Y(_139_)
);

FILL FILL_2__13284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12277_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4538_)
);

FILL FILL_0__9284_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4157_),
    .B(_3435_),
    .C(_4166_),
    .Y(_3398_)
);

NOR2X1 _11135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_3780_)
);

FILL FILL_0__12631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7299_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_2486_),
    .C(_2488_),
    .Y(_1720_)
);

FILL FILL_1__8660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13836_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf4),
    .B(_6073_),
    .C(_6068_),
    .Y(_6074_)
);

FILL FILL_0__13416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9025_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _8095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_1010_)
);

FILL FILL_1__10343_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14906_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6797_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.Atmp [11])
);

FILL FILL_0__7770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7350_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf2),
    .B(_4650_),
    .C(_4628_),
    .Y(_4651_)
);

FILL FILL_1__11968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8555_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [0]),
    .Y(_3484_)
);

FILL FILL_0__8135_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3128_),
    .C(_3116_),
    .Y(_3129_)
);

OR2X2 _13298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5749_),
    .B(\genblk1[6].u_ce.Ain12b [6]),
    .Y(_5751_)
);

FILL FILL_0__11902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10201_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_755_),
    .Y(_756_)
);

AND2X2 _7366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_358_),
    .Y(_359_)
);

FILL FILL_2__13093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11499_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(_4354_),
    .Y(_4355_)
);

FILL FILL_0__9093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3992_),
    .B(_3994_),
    .Y(_3999_)
);

FILL FILL_2__11826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7826_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(\genblk1[3].u_ce.Xin12b [6]),
    .S(vdd),
    .Y(_2675_)
);

FILL FILL_0__7406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2318_),
    .Y(_2319_)
);

NAND2X1 _12989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5449_),
    .Y(_5457_)
);

DFFPOSX1 _12569_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4223_),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.Acalc [8])
);

AOI21X1 _12149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4684_),
    .B(_4699_),
    .C(_4697_),
    .Y(_4704_)
);

FILL FILL_1__14652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert121 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert123 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6291_),
    .B(_6292_),
    .Y(_6293_)
);

FILL FILL_0__13645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert124 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13225_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [10]),
    .Y(_5893_)
);

FILL FILL_0_BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert126 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert128 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10152_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6937_),
    .B(_6916_),
    .C(_6936_),
    .Y(_6938_)
);

FILL FILL_2__7177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8364_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2697_),
    .C(_3330_),
    .Y(_2562_)
);

NAND2X1 _10215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2946_)
);

FILL FILL_2__9743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10010_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_573_),
    .B(_577_),
    .Y(_578_)
);

FILL FILL_1__14708_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_176_)
);

INVX1 _11593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [1]),
    .Y(_4187_)
);

AOI21X1 _11173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3813_),
    .B(_3816_),
    .C(_3535_),
    .Y(_3817_)
);

FILL FILL_2__11215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7635_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf3),
    .B(_2475_),
    .C(_2508_),
    .Y(_1738_)
);

FILL FILL_0__7215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf1),
    .B(_2136_),
    .C(_2114_),
    .Y(_2137_)
);

OAI21X1 _12798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5272_),
    .C(_5273_),
    .Y(_5274_)
);

NOR2X1 _12378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4919_),
    .B(_4910_),
    .Y(_4920_)
);

FILL FILL_1__14461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14659_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14524_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6512_),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.Xin12b [10])
);

FILL FILL_0__14239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [1]),
    .B(_6455_),
    .Y(_6457_)
);

FILL FILL_1__11586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8593_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf0),
    .B(_3520_),
    .C(_3519_),
    .Y(_3521_)
);

FILL FILL_0__8173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10159_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3163_),
    .B(_3152_),
    .Y(_3165_)
);

INVX1 _10024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2763_),
    .Y(_2764_)
);

FILL FILL_0__11940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9378_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11649_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3389_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [10])
);

OAI21X1 _11229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3828_),
    .C(_3869_),
    .Y(_3870_)
);

FILL FILL_1__13732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x248550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11024_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf4),
    .B(_1098_),
    .C(_1099_),
    .Y(_1100_)
);

FILL FILL_1__10857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7864_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2685_),
    .B(_2702_),
    .C(_2710_),
    .Y(_2713_)
);

FILL FILL_0__7444_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2351_),
    .C(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2354_)
);

NAND2X1 _9130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_1954_)
);

NAND2X1 _12187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4740_),
    .B(_4739_),
    .Y(_4741_)
);

FILL FILL_2__8403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14468_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6971_),
    .B(_6972_),
    .Y(_6973_)
);

FILL FILL_0__14048_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6623_),
    .B(\u_ot.LoadCtl_6_bF$buf1 ),
    .C(_6631_),
    .Y(_6498_)
);

FILL FILL_1__7605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11395_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3347_),
    .B(_3321_),
    .C(_3351_),
    .Y(_2579_)
);

FILL FILL_0__10388_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2960_),
    .B(_2982_),
    .Y(_2983_)
);

INVX1 _8821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [1]),
    .Y(_1673_)
);

AOI21X1 _8401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(_1302_),
    .C(_1021_),
    .Y(_1303_)
);

INVX1 _11878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4445_)
);

FILL FILL_0__9187_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [6]),
    .B(_3510__bF$buf0),
    .Y(_4085_)
);

NAND2X1 _11038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3684_),
    .B(_3687_),
    .Y(_3688_)
);

FILL FILL_1__13961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2396_),
    .Y(_2406_)
);

FILL FILL_1__8983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13739_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5981_),
    .B(_5980_),
    .S(_5926__bF$buf0),
    .Y(_5982_)
);

FILL FILL_0__13319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10246_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7009_),
    .B(_7012_),
    .C(_7010_),
    .Y(_7025_)
);

FILL FILL_0__7673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8038_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10729_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2555_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xin12b [6])
);

NAND3X1 _10309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .B(_2957_),
    .C(_2974_),
    .Y(_3036_)
);

FILL FILL_1__12812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [11]),
    .B(_6804_),
    .Y(_6805_)
);

OAI21X1 _14142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6475_),
    .B(_6463_),
    .C(_6479_),
    .Y(_5876_)
);

FILL FILL_1__7834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10197_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2678_),
    .B(_2649__bF$buf4),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_3199_)
);

OAI21X1 _10062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2798_),
    .C(_2799_),
    .Y(_2800_)
);

FILL FILL_1__8619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_665_),
    .Y(_666_)
);

NOR2X1 _7269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_234_),
    .Y(_266_)
);

NAND2X1 _8630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1519_),
    .Y(_1520_)
);

OAI21X1 _8210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf3),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_)
);

DFFPOSX1 _11687_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[4].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.LoadCtl [2])
);

OAI21X1 _11267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3887_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_3906_),
    .Y(_3370_)
);

FILL FILL_2__7903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7729_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9835_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1747_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[2].u_ce.Ain0 [0])
);

FILL FILL_0__7309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2225_),
    .Y(_2227_)
);

FILL FILL_1__8792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13548_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6188_),
    .Y(_6200_)
);

FILL FILL_0__13128_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5830_),
    .B(_5804_),
    .C(_5834_),
    .Y(_5087_)
);

FILL FILL_1__9997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10055_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6849_)
);

FILL FILL_0__7482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x234150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12267_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_807_),
    .C(_837_),
    .Y(_65_)
);

FILL FILL_0__8687_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf2),
    .B(_3560_),
    .Y(_3611_)
);

FILL FILL_0__8267_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3251_)
);

OAI21X1 _10118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2850_),
    .B(_2853_),
    .C(_2741_),
    .Y(_2854_)
);

FILL FILL_1__12621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9226_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7004_),
    .B(_7002_),
    .C(_7007_),
    .Y(_7008_)
);

FILL FILL_0__14086_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(_6663_),
    .Y(_6664_)
);

FILL FILL_1__7643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3018_),
    .B(_3017_),
    .Y(_3019_)
);

FILL FILL_1__8428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8008_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_437_),
    .C(_463_),
    .Y(_485_)
);

NOR2X1 _7078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.LoadCtl [3]),
    .Y(_86_)
);

NOR2X1 _11496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4120_),
    .B(_4119_),
    .Y(_4121_)
);

INVX1 _11076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3723_),
    .Y(_3724_)
);

FILL FILL_2__11958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7538_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .Y(_2441_)
);

FILL FILL_0__7118_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2034_),
    .Y(_2044_)
);

FILL FILL_1__8181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13777_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5951_),
    .Y(_6018_)
);

FILL FILL_0__13357_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5151__bF$buf1),
    .C(_5170_),
    .Y(_5678_)
);

FILL FILL_1__9386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [1]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .Y(_7059_)
);

NAND3X1 _14427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6711_),
    .B(_6712_),
    .C(_6703_),
    .Y(_6713_)
);

AOI21X1 _14007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6359_),
    .B(_6341_),
    .C(_6339_),
    .Y(_6367_)
);

FILL FILL_0__7291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12496_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_135__bF$buf4),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_685_)
);

FILL FILL_1__11489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8076_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10767_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Vld )
);

NAND2X1 _10347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3071_),
    .Y(_3072_)
);

FILL FILL_1__12850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11003_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14180_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5856_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [8])
);

DFFPOSX1 _8915_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[1].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.LoadCtl [2])
);

FILL FILL_1__7872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13215_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5374_),
    .Y(_5384_)
);

FILL FILL_0__12628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11767_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562_),
    .Y(_6562__bF$buf4)
);

FILL FILL_0__12381_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562_),
    .Y(_6562__bF$buf3)
);

FILL FILL_0__7767_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2619_),
    .C(_2620_),
    .Y(_2621_)
);

FILL FILL_0__7347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf0),
    .B(_2262_),
    .C(_2259_),
    .Y(_2263_)
);

MUX2X1 _9033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1861_),
    .B(_1858_),
    .S(_1811__bF$buf2),
    .Y(_1862_)
);

FILL FILL_1__11701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13586_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [1]),
    .B(_5949__bF$buf3),
    .Y(_6236_)
);

DFFPOSX1 _13451_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5051_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [10])
);

FILL FILL_0__13166_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .B(_5496_),
    .Y(_5497_)
);

FILL FILL_2__13913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10093_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6882_),
    .B(_6880_),
    .C(_6883_),
    .Y(_6772_)
);

OAI21X1 _14236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_6549_),
    .C(_6550_),
    .Y(_7071_[6])
);

FILL FILL_1__7508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11298_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3647_)
);

NAND3X1 _10576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3248_),
    .B(_3243_),
    .C(_3285_),
    .Y(_3287_)
);

OAI21X1 _10156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2885_),
    .C(_2889_),
    .Y(_2890_)
);

FILL FILL_2__10618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11232_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(_1605_),
    .Y(_1607_)
);

INVX1 _8304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1209_),
    .Y(_1210_)
);

FILL FILL_1__7681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12857_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5201_),
    .B(_5198_),
    .S(_5151__bF$buf3),
    .Y(_5202_)
);

FILL FILL_0__12437_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4845_),
    .B(_4849_),
    .Y(_4850_)
);

FILL FILL_0__12017_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _9929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .Y(_2672_)
);

INVX1 _9509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2315_),
    .Y(_2316_)
);

FILL FILL_1__8466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_6289_),
    .Y(_6290_)
);

INVX1 _13507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .Y(_5890_)
);

FILL FILL_2__11996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7576_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2473_),
    .B(_2474_),
    .Y(_2475_)
);

FILL FILL_0__7156_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_2023_),
    .C(_2076_),
    .Y(_2081_)
);

FILL FILL_1__11930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10503_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6053_),
    .Y(_6054_)
);

FILL FILL_0__13395_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5714_),
    .Y(_5715_)
);

FILL FILL_1__12715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9302_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14885_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6776_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [9])
);

OAI21X1 _14465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6727_),
    .B(_6740_),
    .C(_6741_),
    .Y(_6520_)
);

NAND3X1 _14045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf0),
    .B(_6397_),
    .C(_6395_),
    .Y(_6403_)
);

FILL FILL_1__7737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3105_),
    .B(_3108_),
    .Y(_3109_)
);

FILL FILL_0__11881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11041_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [9]),
    .Y(_1786_)
);

NAND3X1 _8533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(_1425_),
    .C(_1428_),
    .Y(_1429_)
);

MUX2X1 _8113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .S(vdd),
    .Y(_1028_)
);

FILL FILL_1__7490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13253_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420_),
    .B(_5363_),
    .C(_5416_),
    .Y(_5421_)
);

FILL FILL_0__12666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12246_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5025_),
    .B(_4273_),
    .C(_4267_),
    .Y(_4260_)
);

OAI21X1 _12111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4666_),
    .C(_4667_),
    .Y(_4668_)
);

NAND2X1 _9738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [0]),
    .B(_2475_),
    .Y(_2507_)
);

NAND2X1 _9318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf3),
    .B(_2133_),
    .Y(_2134_)
);

FILL FILL_1__8695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14038_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6094_),
    .B(_6091_),
    .C(_6086_),
    .Y(_6107_)
);

INVX1 _13316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5767_),
    .Y(_5768_)
);

FILL FILL_1_CLKBUF1_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7385_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2298_),
    .Y(_2299_)
);

OR2X2 _9071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1897_),
    .B(_1895_),
    .Y(_1898_)
);

FILL FILL_0__10312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x79350 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_729_),
    .C(_771_),
    .Y(_773_)
);

FILL FILL_2__13951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11517_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .Y(_4373_)
);

FILL FILL_2__9129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9111_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6917_),
    .B(_6918_),
    .Y(_6919_)
);

NAND2X1 _14274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6578_),
    .B(_6579_),
    .Y(_6580_)
);

FILL FILL_1__7546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .B(_2925_),
    .Y(_2926_)
);

FILL FILL_2__10656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11270_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1162_),
    .B(_1637_),
    .C(_1639_),
    .Y(_876_)
);

NAND2X1 _8342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [11]),
    .B(_996__bF$buf1),
    .Y(_1246_)
);

NAND2X1 _11399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4030_),
    .B(_4029_),
    .Y(_4031_)
);

FILL FILL_2__7615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12895_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5237_),
    .B(_5235_),
    .Y(_5238_)
);

FILL FILL_0__12475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12055_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _12340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4270_),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .C(_4882_),
    .D(_4884_),
    .Y(_4217_)
);

OAI21X1 _9967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2684_),
    .C(_2709_),
    .Y(_2710_)
);

AND2X2 _9547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2350_),
    .B(_2348_),
    .Y(_2351_)
);

OAI21X1 _9127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_1930_),
    .C(_1947_),
    .Y(_1951_)
);

FILL FILL_1__8084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14267_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [5]),
    .Y(_6326_)
);

INVX1 _13545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .Y(_5924_)
);

NAND2X1 _13125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5586_),
    .Y(_5587_)
);

FILL FILL_0__14621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10121_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_594_),
    .Y(_595_)
);

FILL FILL_0__8399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4035_),
    .C(_3431_),
    .Y(_3424_)
);

OAI21X1 _14083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6438_),
    .B(_6437_),
    .C(_6047_),
    .Y(_6439_)
);

INVX1 _8818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[1] [0]),
    .Y(_1671_)
);

FILL FILL_1__7775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13118_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5288_),
    .B(_5270_),
    .C(_5287_),
    .Y(_5291_)
);

FILL FILL_2__10465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9501_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1819_),
    .C(_1820_),
    .Y(_1821_)
);

NAND3X1 _8571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(_1463_),
    .C(_1464_),
    .Y(_1465_)
);

AOI21X1 _8151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1062_),
    .B(_1063_),
    .C(_998_),
    .Y(_1064_)
);

FILL FILL_2__7844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12284_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9776_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1688_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Ycalc [11])
);

OAI21X1 _9356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2149_),
    .C(_2163_),
    .Y(_2170_)
);

FILL FILL_1__11604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14076_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6144_)
);

FILL FILL_0__13069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5799_),
    .B(_5800_),
    .C(_5801_),
    .Y(_5061_)
);

FILL FILL_0__14850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12809_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [3]),
    .Y(_6802_)
);

OAI21X1 _14139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Yin12b [9]),
    .Y(_6478_)
);

FILL FILL_0__10770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10350_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_803_),
    .C(_804_),
    .Y(_39_)
);

NAND2X1 _7422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .B(_411_),
    .Y(_412_)
);

OAI21X1 _10899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510__bF$buf3),
    .B(_3555_),
    .C(_3511_),
    .Y(_3353_)
);

OAI21X1 _10479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3194_),
    .B(_3196_),
    .C(_3183_),
    .Y(_2540_)
);

NAND3X1 _10059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf2),
    .B(_2796_),
    .C(_2791_),
    .Y(_2797_)
);

FILL FILL_1__12982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11555_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4408_),
    .B(_4405_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4409_)
);

FILL FILL_2__9167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11135_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_4050_)
);

OAI21X1 _11000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf4),
    .B(_3649_),
    .C(_3650_),
    .Y(_3651_)
);

NAND2X1 _8627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1516_),
    .B(_1515_),
    .Y(_1517_)
);

INVX1 _8207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .Y(_1117_)
);

FILL FILL_1__7584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13347_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Acalc [11]),
    .C(_5106_),
    .Y(_5111_)
);

AOI21X1 _12205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4718_),
    .B(_4719_),
    .C(_4329_),
    .Y(_4758_)
);

FILL FILL_0__13701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9310_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1282_),
    .B(_1277_),
    .C(_1261_),
    .Y(_851_)
);

FILL FILL_2__7653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7479_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [4]),
    .Y(_2386_)
);

NAND2X1 _9165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1963_),
    .B(_1987_),
    .Y(_1988_)
);

FILL FILL_1__11833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10406_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _13583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5957_),
    .B(_5960_),
    .C(_5925__bF$buf1),
    .D(_5954_),
    .Y(_5961_)
);

FILL FILL_0__13298_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5622_),
    .Y(_5623_)
);

FILL FILL_2__13625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9205_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6979_),
    .B(_6999_),
    .C(_6992_),
    .Y(_7005_)
);

INVX1 _14368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [4]),
    .Y(_6661_)
);

FILL FILL_2__8191_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_996__bF$buf4)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_996__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_996__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_996__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_996__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf3 )
);

AND2X2 _7651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_621_),
    .B(_630_),
    .Y(_631_)
);

INVX1 _7231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_229_)
);

NAND2X1 _10288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3014_),
    .B(_3015_),
    .Y(_3016_)
);

FILL FILL_1__12791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11364_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8856_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_854_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Xcalc [3])
);

MUX2X1 _8436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1292_),
    .S(gnd),
    .Y(_1336_)
);

OAI21X1 _8016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(_935_),
    .C(_936_),
    .Y(_937_)
);

FILL FILL_1__7393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12989_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5303_),
    .B(_5327_),
    .Y(_5328_)
);

FILL FILL_0__12149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4968_),
    .B(_4971_),
    .Y(_4972_)
);

INVX1 _12014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .Y(_4575_)
);

FILL FILL_0__13930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8178_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6014_),
    .Y(_6015_)
);

AND2X2 _13219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5671_),
    .B(_5675_),
    .Y(_5676_)
);

FILL FILL_0__14715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7288_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2203_),
    .B(_2206_),
    .Y(_2207_)
);

FILL FILL_1__11222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8667_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3559_),
    .B(_3574_),
    .Y(_3575_)
);

FILL FILL_0__10635_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2678_),
    .B(_3215_),
    .C(_3214_),
    .Y(_3216_)
);

FILL FILL_0__10215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5807_),
    .Y(_5823_)
);

OAI21X1 _7707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .B(_682_),
    .C(_669_),
    .Y(_26_)
);

FILL FILL_2__13854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9434_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Acalc [0]),
    .C(_4281_),
    .D(_4282_),
    .Y(_4283_)
);

FILL FILL_0__9014_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [1]),
    .B(En_bF$buf3),
    .Y(_6762_)
);

DFFPOSX1 _14177_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5853_),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.Xcalc [5])
);

FILL FILL_1__7869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8810_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_810_),
    .Y(_826_)
);

OAI21X1 _7460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_233_),
    .C(_447_),
    .Y(_448_)
);

AOI21X1 _10097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2823_),
    .B(_2801_),
    .C(_2802_),
    .Y(_2833_)
);

FILL FILL_1__12180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11173_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1551_),
    .B(_1548_),
    .Y(_1552_)
);

INVX1 _8245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [7]),
    .Y(_1153_)
);

FILL FILL_1__10913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12798_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .B(\genblk1[6].u_ce.Xcalc [5]),
    .C(_5108_),
    .D(\genblk1[6].u_ce.Xcalc [7]),
    .Y(_5145_)
);

FILL FILL_0__12378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .B(_4778_),
    .C(_4751_),
    .Y(_4794_)
);

FILL FILL_2__12705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8705_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf2),
    .B(_6233_),
    .C(_6222_),
    .Y(_6234_)
);

DFFPOSX1 _13448_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5048_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [7])
);

OAI21X1 _13028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5492_),
    .C(_5493_),
    .Y(_5494_)
);

FILL FILL_0__14104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10024_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7936_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [7])
);

NAND2X1 _7516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .B(_501_),
    .Y(_502_)
);

FILL FILL_2__13663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9663_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4455_),
    .B(_4457_),
    .C(_4445_),
    .Y(_4499_)
);

FILL FILL_0__9243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11229_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4133_),
    .B(_4118_),
    .C(_4132_),
    .Y(_4137_)
);

FILL FILL_1__7678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14028_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .Y(_5199_)
);

FILL FILL_1__14802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x198150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8894_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_892_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Yin12b [7])
);

AOI22X1 _8474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_959_),
    .B(_996__bF$buf0),
    .C(_1372_),
    .D(_994_),
    .Y(_855_)
);

FILL FILL_0_CLKBUF1_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [0]),
    .Y(_970_)
);

FILL FILL_0_CLKBUF1_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13194_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5364_)
);

NAND2X1 _12472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_5000_),
    .Y(_5001_)
);

FILL FILL_0__12187_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4609_),
    .B(_4611_),
    .C(_4420_),
    .Y(_4612_)
);

FILL FILL_2__12934_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834__bF$buf1),
    .B(_2472_),
    .C(_2471_),
    .Y(_1712_)
);

AOI21X1 _9259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2076_),
    .C(_2074_),
    .Y(_2078_)
);

FILL FILL_1__11927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_6049_),
    .C(_6050_),
    .Y(_6051_)
);

OAI21X1 _13257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5180_),
    .B(_5711_),
    .C(_5710_),
    .Y(_5712_)
);

FILL FILL_0__14753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10253_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_717_),
    .B(_716_),
    .Y(_718_)
);

AOI21X1 _7325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_287_),
    .C(_288_),
    .Y(_319_)
);

FILL FILL_2__13892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9472_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [3]),
    .Y(_4316_)
);

FILL FILL_0__11458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11038_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3959_),
    .C(_3956_),
    .Y(_3960_)
);

FILL FILL_1__7487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14677_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5417_),
    .B(_5416_),
    .C(_5414_),
    .Y(_5418_)
);

OAI21X1 _12528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_4266_)
);

NAND2X1 _12108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4560_),
    .Y(_4665_)
);

FILL FILL_1__14611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(_1161_),
    .Y(_1190_)
);

FILL FILL_1__10951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7136_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4829_),
    .Y(_4830_)
);

FILL FILL_2__12743_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2278_),
    .Y(_2296_)
);

AOI21X1 _9068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1894_),
    .B(_1891_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_1895_)
);

FILL FILL_1__11736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10309_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13486_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5086_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Ain12b [9])
);

AOI21X1 _13066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5530_)
);

FILL FILL_2__13108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10062_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7974_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_58_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin1 [1])
);

NOR2X1 _7554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf2),
    .B(_411_),
    .Y(_538_)
);

INVX1 _7134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_136_)
);

FILL FILL_1__12694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12274_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4497_),
    .B(_4526_),
    .C(_4525_),
    .Y(_4535_)
);

FILL FILL_0__9281_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_4165_)
);

FILL FILL_0__11267_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3777_)
);

NAND2X1 _8759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1637_),
    .Y(_1638_)
);

OAI21X1 _8339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1243_),
    .C(_1065_),
    .Y(_1244_)
);

FILL FILL_1__7296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13899_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2486_),
    .Y(_2487_)
);

FILL FILL_1__13059_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5234_),
    .B(_5231_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5235_)
);

NOR2X1 _12337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4881_),
    .B(_4874_),
    .Y(_4882_)
);

FILL FILL_1__14840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9022_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf1),
    .B(_1006_),
    .C(_1005_),
    .Y(_1007_)
);

FILL FILL_1__10340_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14903_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6794_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [7])
);

FILL FILL_0__14618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf2),
    .B(_4647_),
    .Y(_4648_)
);

FILL FILL_2__12972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12132_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2113_),
    .Y(_2114_)
);

FILL FILL_1__11965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8552_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3479_),
    .B(_3480_),
    .C(_3481_),
    .Y(_3482_)
);

FILL FILL_0__8132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10118_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf5),
    .B(_3120_),
    .C(_3118_),
    .Y(_3126_)
);

OAI21X1 _13295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5745_),
    .B(_5709_),
    .C(_5188__bF$buf0),
    .Y(_5748_)
);

FILL FILL_2__9931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[4] [0]),
    .Y(_3430_)
);

FILL FILL_0__10291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8713_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .Y(_753_)
);

NAND3X1 _7363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_353_),
    .C(_349_),
    .Y(_356_)
);

FILL FILL_1__12083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11496_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .B(\genblk1[5].u_ce.Xin12b [4]),
    .S(vdd),
    .Y(_4352_)
);

FILL FILL_0__9090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11076_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3994_),
    .B(_3992_),
    .Y(_3996_)
);

FILL FILL_1__9918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11403_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .B(_1814_),
    .S(_1811__bF$buf2),
    .Y(_1818_)
);

OAI21X1 _8568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1444_),
    .B(_1442_),
    .C(_1010__bF$buf3),
    .Y(_1462_)
);

NOR2X1 _8148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1060_),
    .Y(_1061_)
);

FILL FILL_1__10816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13288_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5447_),
    .B(_5453_),
    .Y(_5454_)
);

DFFPOSX1 _12566_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4220_),
    .CLK(clk_bF$buf47),
    .Q(\genblk1[5].u_ce.Acalc [5])
);

NAND2X1 _12146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4685_),
    .B(_4700_),
    .Y(_4702_)
);

FILL FILL_0__13642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14427_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6917_),
    .B(_6934_),
    .C(_6925_),
    .Y(_6935_)
);

FILL FILL_0__14007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[2].u_ce.X_ [0]),
    .Y(_3329_)
);

FILL FILL_0__10347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2678_),
    .Y(_2943_)
);

INVX1 _7839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_802_)
);

INVX1 _7419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .Y(_409_)
);

FILL FILL_2__13146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9566_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4403_),
    .Y(_4406_)
);

FILL FILL_0__9146_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [3]),
    .B(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_4047_)
);

FILL FILL_1__13920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8102_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_574_),
    .C(_549_),
    .Y(_575_)
);

FILL FILL_1__14705_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_173_)
);

INVX1 _11590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [0]),
    .Y(_4185_)
);

MUX2X1 _11170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .B(_3806_),
    .S(_3487__bF$buf1),
    .Y(_3814_)
);

FILL FILL_1__9727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9307_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1641_),
    .C(_1660_),
    .Y(_890_)
);

NAND2X1 _8377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1278_),
    .B(_1279_),
    .Y(_1280_)
);

FILL FILL_1__10625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13097_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5271_)
);

NAND2X1 _12375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4911_),
    .B(_4915_),
    .Y(_4917_)
);

FILL FILL_0__13871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14656_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14521_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6509_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Ycalc [9])
);

FILL FILL_0__14236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6453_),
    .B(_6454_),
    .Y(_6455_)
);

FILL FILL_2__12170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8590_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3517_),
    .B(_3496_),
    .C(_3487__bF$buf4),
    .Y(_3518_)
);

FILL FILL_0__8170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10156_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3161_),
    .B(_3160_),
    .C(_2770_),
    .Y(_3162_)
);

OAI21X1 _10021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2759_),
    .C(_2760_),
    .Y(_2761_)
);

FILL FILL_2__10903_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(_626_),
    .Y(_628_)
);

INVX2 _7228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .Y(_227_)
);

FILL FILL_1__12788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9375_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11646_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3386_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [9])
);

NAND2X1 _11226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_3867_)
);

FILL FILL_0__12722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11441_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf1),
    .B(_1046_),
    .Y(_1097_)
);

FILL FILL_1__10854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7441_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4733_),
    .B(_4737_),
    .C(_4366_),
    .Y(_4738_)
);

FILL FILL_2__8820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8646_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .B(_3567_),
    .C(_3570_),
    .Y(_3572_)
);

FILL FILL_0__8226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5804_),
    .C(_5821_),
    .Y(_5076_)
);

FILL FILL_2__9605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14465_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6965_),
    .B(_6969_),
    .C(_6963_),
    .Y(_6970_)
);

FILL FILL_0__14045_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(_6626_),
    .Y(_6629_)
);

FILL FILL_1__7602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11392_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Ain12b [9]),
    .Y(_3350_)
);

FILL FILL_0__10385_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2979_),
    .Y(_2980_)
);

FILL FILL_1__8807_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_807_),
    .C(_824_),
    .Y(_54_)
);

NAND2X1 _7457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [1]),
    .B(_158__bF$buf3),
    .Y(_445_)
);

FILL FILL_2__13184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4422_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4443_)
);

FILL FILL_0__9184_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4072_),
    .Y(_4083_)
);

NAND3X1 _11035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf0),
    .B(_3681_),
    .C(_3675_),
    .Y(_3685_)
);

FILL FILL_2__11917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2401_),
    .Y(_2403_)
);

FILL FILL_1__8980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13736_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf4),
    .B(_5941_),
    .C(_5978_),
    .Y(_5979_)
);

FILL FILL_0__13316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10243_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7022_),
    .B(_7013_),
    .Y(_7023_)
);

FILL FILL_0__7670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8455_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10726_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2552_),
    .CLK(clk_bF$buf50),
    .Q(\genblk1[3].u_ce.Xin12b [11])
);

FILL FILL_0__8035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3032_),
    .Y(_3033_)
);

INVX1 _13198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5655_),
    .Y(_5656_)
);

FILL FILL_0__11802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10101_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_662_),
    .C(\genblk1[0].u_ce.Ain0 [0]),
    .Y(_663_)
);

INVX2 _7266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .Y(_263_)
);

FILL FILL_0__11399_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11684_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3424_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Ain0 [1])
);

NOR2X1 _11264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3903_),
    .B(_3888_),
    .Y(_3904_)
);

FILL FILL_2__11726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7726_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9832_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1744_),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[2].u_ce.Ain12b [5])
);

FILL FILL_0__7306_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2219_),
    .B(_2223_),
    .C(_1852_),
    .Y(_2224_)
);

OAI21X1 _12889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5323_),
    .B(_5352_),
    .C(_5351_),
    .Y(_5361_)
);

NAND2X1 _12469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(_4997_),
    .Y(_4999_)
);

NOR3X1 _12049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4599_),
    .B(_4608_),
    .C(_4592_),
    .Y(_4609_)
);

FILL FILL_1__14132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13545_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6197_),
    .B(_6193_),
    .Y(_6198_)
);

FILL FILL_0__13125_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Ain12b [9]),
    .Y(_5833_)
);

FILL FILL_1__9994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10052_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [1]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf0),
    .Y(_6847_)
);

FILL FILL_1__11257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8684_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3608_)
);

FILL FILL_0__8264_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .Y(_3248_)
);

INVX1 _10115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2850_),
    .Y(_2851_)
);

FILL FILL_2__9643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14608_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(gnd),
    .C(_481_),
    .Y(_482_)
);

INVX2 _7075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .Y(_83_)
);

NAND3X1 _11493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [8]),
    .B(_4053_),
    .C(_4117_),
    .Y(_4118_)
);

AOI21X1 _11073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3719_),
    .B(_3707_),
    .C(_3720_),
    .Y(_3721_)
);

FILL FILL_2__11955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7535_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2427_),
    .B(_1834__bF$buf1),
    .C(_2437_),
    .D(_2438_),
    .Y(_1708_)
);

FILL FILL_0__7115_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1980_),
    .B(_1983_),
    .Y(_2041_)
);

MUX2X1 _12698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .B(\genblk1[6].u_ce.Xin12b [4]),
    .S(gnd),
    .Y(_5178_)
);

NAND3X1 _12278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4817_),
    .B(_4819_),
    .C(_4826_),
    .Y(_4827_)
);

FILL FILL_1__14781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14559_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [0]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .Y(_7057_)
);

FILL FILL_0__14139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6708_),
    .B(_6709_),
    .Y(_6710_)
);

AND2X2 _14004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .B(_6357_),
    .Y(_6364_)
);

FILL FILL_1__11486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10479_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10764_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[3].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.LoadCtl [3])
);

FILL FILL_0__10059_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [6]),
    .Y(_3069_)
);

FILL FILL_0__11840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11000_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8912_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_910_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Ain0 [1])
);

FILL FILL_0__9698_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4530_),
    .B(_4528_),
    .C(_4532_),
    .Y(_4533_)
);

FILL FILL_0__9278_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_4162_),
    .C(_4163_),
    .Y(_3395_)
);

NAND2X1 _11129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3760_),
    .B(_3774_),
    .Y(_3364_)
);

FILL FILL_1__13632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13212_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5320_),
    .B(_5323_),
    .Y(_5381_)
);

FILL FILL_0__12625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x90150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11344_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1003_),
    .B(_982_),
    .C(_973__bF$buf3),
    .Y(_1004_)
);

FILL FILL_1__10337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7764_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_2616_),
    .C(_2617_),
    .Y(_2618_)
);

FILL FILL_0__7344_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf3),
    .B(_2087_),
    .Y(_2260_)
);

INVX1 _9030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .Y(_1859_)
);

INVX1 _12087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4644_),
    .Y(_4645_)
);

FILL FILL_2__8303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6879_),
    .B(_6876_),
    .Y(_6881_)
);

OAI21X1 _14233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_6547_),
    .C(_6548_),
    .Y(_7071_[5])
);

FILL FILL_1__7505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11295_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3644_),
    .B(_3643_),
    .C(_3582_),
    .Y(_3645_)
);

OAI21X1 _10573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3258_),
    .B(_3274_),
    .C(_3272_),
    .Y(_3284_)
);

FILL FILL_0__10288_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2794_),
    .C(_2840_),
    .Y(_2887_)
);

NAND3X1 _8721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [8]),
    .B(_1539_),
    .C(_1603_),
    .Y(_1604_)
);

AOI21X1 _8301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1193_),
    .C(_1206_),
    .Y(_1207_)
);

NAND2X1 _11778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [1]),
    .B(_4348__bF$buf1),
    .Y(_4349_)
);

FILL FILL_0__9087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3956_),
    .B(_3958_),
    .Y(_3993_)
);

FILL FILL_1__13861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12014_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _9926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .Y(_2670_)
);

NAND3X1 _9506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .B(_2305_),
    .C(_2312_),
    .Y(_2313_)
);

FILL FILL_1__8463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13639_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [10]),
    .Y(_6287_)
);

FILL FILL_0__13219_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5886_),
    .Y(_5887_)
);

FILL FILL_1__9668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10146_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [9]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf0),
    .Y(_6933_)
);

FILL FILL_0__7573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8358_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3316_),
    .B(_2597_),
    .C(_3327_),
    .Y(_2559_)
);

OAI21X1 _10209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2938_),
    .C(_2939_),
    .Y(_2940_)
);

FILL FILL_1__12712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14597_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14882_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6773_),
    .CLK(clk_bF$buf50),
    .Q(\u_pa.acc_reg [6])
);

OAI21X1 _14462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6731_),
    .B(_6737_),
    .C(_6739_),
    .Y(_6519_)
);

OAI21X1 _14042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6377_),
    .B(_6374_),
    .C(_5963__bF$buf5),
    .Y(_6400_)
);

FILL FILL_1__7734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x234150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf3),
    .B(_3102_),
    .C(_3097_),
    .Y(_3106_)
);

FILL FILL_1__8939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_571_),
    .Y(_572_)
);

OAI22X1 _7169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_169_),
    .C(_134__bF$buf2),
    .D(_163_),
    .Y(_170_)
);

OAI21X1 _8950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1780_),
    .B(_1783_),
    .C(_1768_),
    .Y(_1784_)
);

INVX1 _8530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1424_),
    .Y(_1426_)
);

MUX2X1 _8110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1017_),
    .S(_972__bF$buf2),
    .Y(_1025_)
);

OAI21X1 _11587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4141_),
    .B(_4151_),
    .C(_4183_),
    .Y(_3413_)
);

OAI21X1 _11167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf0),
    .B(_3807_),
    .C(_3810_),
    .Y(_3811_)
);

FILL FILL_2__7803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7629_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1809_),
    .C(_2505_),
    .Y(_1735_)
);

FILL FILL_0__7209_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2130_),
    .Y(_2131_)
);

FILL FILL_1__8692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13868_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6099_),
    .B(_6103_),
    .C(_6104_),
    .Y(_6105_)
);

FILL FILL_0__13028_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5756_),
    .B(_5764_),
    .C(_5174__bF$buf0),
    .Y(_5766_)
);

FILL FILL_1__9897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10375_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14518_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6506_),
    .CLK(clk_bF$buf4),
    .Q(\u_ot.Ycalc [6])
);

FILL FILL_0__7382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12167_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_760_),
    .C(_758_),
    .Y(_770_)
);

FILL FILL_0__8587_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3514_),
    .B(_3513_),
    .S(_3487__bF$buf4),
    .Y(_3515_)
);

FILL FILL_0__8167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [10]),
    .B(_3157_),
    .C(_3158_),
    .Y(_3159_)
);

NAND3X1 _10018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf2),
    .B(_2757_),
    .C(_2748_),
    .Y(_2758_)
);

FILL FILL_1__12941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9126_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6910_),
    .B(_6871_),
    .C(_6915_),
    .Y(_6916_)
);

OAI21X1 _14271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6570_),
    .C(_6571_),
    .Y(_6577_)
);

FILL FILL_1__7543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12719_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2911_),
    .Y(_2923_)
);

FILL FILL_1__8748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_387_),
    .C(_371_),
    .Y(_389_)
);

OR2X2 _11396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_4025_),
    .Y(_4028_)
);

FILL FILL_0__12892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7858_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(\genblk1[3].u_ce.Xin0 [1]),
    .S(vdd),
    .Y(_2707_)
);

FILL FILL_0__7438_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(gnd),
    .C(_2347_),
    .Y(_2348_)
);

AOI21X1 _9124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1948_),
    .C(_1836_),
    .Y(_1949_)
);

FILL FILL_1__8081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14264_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6305_),
    .Y(_6324_)
);

FILL FILL_0__13677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13257_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _13542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[7].u_ce.Xcalc [1]),
    .C(_5921_),
    .D(_5892_),
    .Y(_5922_)
);

AOI21X1 _13122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .B(_5545_),
    .C(_5155_),
    .Y(_5584_)
);

FILL FILL_1__9286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10184_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6966_),
    .B(_6967_),
    .C(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .Y(_6968_)
);

NAND3X1 _14327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6625_),
    .B(_6586_),
    .C(_6624_),
    .Y(_6626_)
);

FILL FILL_0__7191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf4),
    .B(_588_),
    .C(_583_),
    .Y(_592_)
);

FILL FILL_1__11389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8396_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Ain12b [8]),
    .Y(_3348_)
);

MUX2X1 _10247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2976_),
    .B(_2965_),
    .S(gnd),
    .Y(_2977_)
);

FILL FILL_1__12750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11323_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [10]),
    .B(_6434_),
    .C(_6435_),
    .Y(_6436_)
);

OAI21X1 _8815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1637_),
    .C(_1669_),
    .Y(_899_)
);

FILL FILL_1__7772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12948_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5270_),
    .B(_5288_),
    .C(_5176_),
    .Y(_5289_)
);

FILL FILL_0__12528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7667_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9773_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1685_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Ycalc [8])
);

FILL FILL_0__7247_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2149_),
    .B(_2166_),
    .Y(_2168_)
);

FILL FILL_1__11601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14073_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6051_),
    .C(_6117_),
    .Y(_6141_)
);

FILL FILL_0__13066_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.X_ [0]),
    .Y(_5799_)
);

FILL FILL_2__13813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12806_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [4]),
    .Y(_6799_)
);

OAI21X1 _14136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6476_)
);

FILL FILL_1__7828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11198_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .B(_3522_),
    .C(_3552_),
    .Y(_3553_)
);

NOR2X1 _10476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(_3193_),
    .Y(_3194_)
);

AOI21X1 _10056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2751_),
    .B(_2649__bF$buf3),
    .C(_2793_),
    .Y(_2794_)
);

FILL FILL257550x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11132_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1511_),
    .Y(_1514_)
);

INVX1 _8204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1114_)
);

FILL FILL_1__7581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12757_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(\genblk1[6].u_ce.LoadCtl [3]),
    .Y(_5108_)
);

FILL FILL_0__12337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(_4754_),
    .Y(_4755_)
);

DFFPOSX1 _9829_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1741_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[2].u_ce.Ain12b [6])
);

NAND3X1 _9409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .B(_2220_),
    .C(_2161_),
    .Y(_2221_)
);

FILL FILL_1__8786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6168_),
    .B(_6171_),
    .C(_6150_),
    .Y(_6195_)
);

OAI21X1 _13407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Ain12b [8]),
    .Y(_5831_)
);

FILL FILL_2__11896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7476_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2382_),
    .C(_2383_),
    .Y(_2384_)
);

AOI21X1 _9162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1941_),
    .B(_1943_),
    .C(_1931_),
    .Y(_1985_)
);

FILL FILL_1__11830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10403_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .B(_5955_),
    .C(_5926__bF$buf4),
    .Y(_5958_)
);

FILL FILL_0__13295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5575_),
    .B(_5604_),
    .C(_5577_),
    .Y(_5620_)
);

FILL FILL_2__13622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9202_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6960_),
    .B(_6958_),
    .Y(_7002_)
);

OR2X2 _14365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6657_),
    .B(\u_ot.Yin1 [1]),
    .Y(_6659_)
);

FILL FILL_1__7637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14827_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf1),
    .B(_3012_),
    .Y(_3013_)
);

FILL FILL_0__11781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11361_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8853_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_851_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Xcalc [0])
);

INVX1 _8433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1332_),
    .Y(_1333_)
);

AOI21X1 _8013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_932_),
    .C(_933_),
    .Y(_934_)
);

FILL FILL_1__7390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12986_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5281_),
    .B(_5283_),
    .C(_5271_),
    .Y(_5325_)
);

FILL FILL_0__12146_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf4),
    .B(\genblk1[5].u_ce.Ain12b [9]),
    .Y(_4969_)
);

OAI21X1 _12011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4571_),
    .B(_4559_),
    .C(_4417_),
    .Y(_4573_)
);

NAND2X1 _9638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2434_),
    .Y(_2436_)
);

AOI22X1 _9218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2020_),
    .B(_1834__bF$buf4),
    .C(_2038_),
    .D(_2018_),
    .Y(_1685_)
);

FILL FILL_1__8595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14358_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6011_),
    .Y(_6012_)
);

NOR2X1 _13216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .B(_5672_),
    .Y(_5673_)
);

FILL FILL_0__14712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .B(_2196_),
    .Y(_2204_)
);

FILL FILL_0__10632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10212_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_679_),
    .Y(_680_)
);

FILL FILL_2__13851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11417_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.Acalc [4]),
    .C(_4279_),
    .D(\genblk1[5].u_ce.Acalc [6]),
    .Y(_4280_)
);

FILL FILL_0__9011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9029_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(En_bF$buf3),
    .Y(_6834_)
);

DFFPOSX1 _14174_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5850_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Xcalc [2])
);

DFFPOSX1 _8909_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_907_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Ain1 [0])
);

FILL FILL_1__7866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5360_),
    .B(_5174__bF$buf2),
    .C(_5378_),
    .D(_5358_),
    .Y(_5037_)
);

FILL FILL_1_BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2817_),
    .B(_2814_),
    .C(_2809_),
    .Y(_2830_)
);

FILL FILL_2__10556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11170_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(gnd),
    .C(_1010__bF$buf4),
    .Y(_1549_)
);

AOI21X1 _8242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1146_),
    .C(_998_),
    .Y(_1151_)
);

FILL FILL_1__10910_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3937_)
);

FILL FILL_2__7515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12795_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [3]),
    .Y(_5142_)
);

FILL FILL_0__12375_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4757_),
    .B(_4785_),
    .Y(_4791_)
);

FILL FILL_2__12702_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2615_),
    .B(_2614_),
    .Y(\a[4] [1])
);

INVX1 _9447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [7]),
    .Y(_2257_)
);

INVX1 _9027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1856_)
);

FILL FILL_0__8702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14587_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf1),
    .B(_6226_),
    .Y(_6231_)
);

DFFPOSX1 _13445_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5045_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Xcalc [4])
);

NAND2X1 _13025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5386_),
    .Y(_5491_)
);

FILL FILL_0__14101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10021_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7933_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf35),
    .Q(\genblk1[0].u_ce.Xcalc [4])
);

NOR2X1 _7513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf0),
    .B(_498_),
    .Y(_499_)
);

FILL FILL_0__8299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9660_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4489_),
    .B(_4492_),
    .Y(_4496_)
);

FILL FILL_0__9240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4133_),
    .B(_4130_),
    .C(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_4135_)
);

NAND2X1 _8718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [8]),
    .B(_996__bF$buf3),
    .Y(_1601_)
);

FILL FILL_1__7675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13018_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5196_)
);

FILL FILL_2__10365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9401_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8891_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_889_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Yin12b [8])
);

OR2X2 _8471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1369_),
    .Y(_1370_)
);

OAI21X1 _8051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_966_),
    .C(_967_),
    .Y(_968_)
);

FILL FILL_0_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12931_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .B(_2469_),
    .C(_2460_),
    .Y(_1711_)
);

AOI21X1 _9256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2050_),
    .B(_2052_),
    .C(_2046_),
    .Y(_2075_)
);

FILL FILL_1__11924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6048_)
);

FILL FILL_0__13389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5151__bF$buf1),
    .Y(_5709_)
);

FILL FILL_0__14750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9716_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14879_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6770_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [3])
);

NAND2X1 _14459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [4]),
    .B(_6737_),
    .Y(_6738_)
);

OAI21X1 _14039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6396_),
    .C(_6376_),
    .Y(_6397_)
);

FILL FILL_0__10670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10250_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_713_),
    .Y(_715_)
);

AOI21X1 _7322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_300_),
    .C(_295_),
    .Y(_316_)
);

AOI22X1 _10799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Ycalc [0]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Ycalc [2]),
    .Y(_3461_)
);

OAI21X1 _10379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3076_),
    .B(_3070_),
    .C(_2686__bF$buf3),
    .Y(_3103_)
);

FILL FILL_1__12882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11875_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4310_),
    .B(_4313_),
    .C(_4282_),
    .Y(_4314_)
);

FILL FILL_0__11455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11035_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3870_),
    .Y(_3957_)
);

INVX1 _8947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [4]),
    .Y(_1781_)
);

INVX1 _8527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1422_),
    .Y(_1423_)
);

NAND2X1 _8107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1022_)
);

FILL FILL_1__7484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13247_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5390_),
    .B(_5392_),
    .C(_5386_),
    .Y(_5415_)
);

OAI21X1 _12525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4900_),
    .B(_5000_),
    .C(_4264_),
    .Y(_4257_)
);

NAND2X1 _12105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [2]),
    .B(_4348__bF$buf0),
    .Y(_4662_)
);

FILL FILL_0__13601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9210_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1161_),
    .B(_1165_),
    .Y(_1187_)
);

FILL FILL_0__14806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2278_),
    .C(_1832_),
    .Y(_2294_)
);

INVX1 _9065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1889_),
    .Y(_1892_)
);

FILL FILL_1__11733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13198_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13483_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5083_),
    .CLK(clk_bF$buf57),
    .Q(\genblk1[6].u_ce.Ain12b [10])
);

NAND2X1 _13063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5511_),
    .B(_5526_),
    .Y(_5528_)
);

FILL FILL_2__13525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9105_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .B(_6907_),
    .C(_6899_),
    .Y(_6913_)
);

NAND2X1 _14268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6574_),
    .B(_6572_),
    .Y(_6575_)
);

FILL FILL_2__8091_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7971_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_55_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Yin12b [4])
);

INVX1 _7551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [5]),
    .Y(_535_)
);

INVX1 _7131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .Y(_133_)
);

OR2X2 _10188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2920_),
    .B(_2916_),
    .Y(_2921_)
);

FILL FILL_1__12691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11264_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [5]),
    .B(_923_),
    .Y(_1635_)
);

AND2X2 _8336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1235_),
    .B(_1231_),
    .Y(_1241_)
);

FILL FILL_1__7293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12889_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5229_),
    .Y(_5232_)
);

FILL FILL_0__12469_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4877_),
    .B(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_4879_)
);

FILL FILL_0__12049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8078_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5930_),
    .B(_6320_),
    .C(_6319_),
    .Y(_6321_)
);

OAI21X1 _13539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(\genblk1[7].u_ce.Xcalc [9]),
    .C(_5889_),
    .Y(_5919_)
);

NAND2X1 _13119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(_5580_),
    .Y(_5581_)
);

DFFPOSX1 _14900_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6791_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [4])
);

FILL FILL_0__14615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7188_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1931_),
    .C(_2110_),
    .Y(_2111_)
);

FILL FILL_1__11962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Xcalc [11]),
    .Y(_3479_)
);

FILL FILL_0__10535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10115_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3100_),
    .B(_3097_),
    .C(_2686__bF$buf5),
    .Y(_3123_)
);

OAI21X1 _13292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5180_),
    .C(_5150__bF$buf3),
    .Y(_5745_)
);

OAI21X1 _7607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_556_),
    .C(_172__bF$buf4),
    .Y(_589_)
);

FILL FILL_2__13754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9334_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4185_),
    .B(_3435_),
    .C(_3428_),
    .Y(_3421_)
);

OAI21X1 _14497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(_6648_),
    .C(_6758_),
    .Y(_6535_)
);

OAI21X1 _14077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6413_),
    .B(_6432_),
    .C(_5963__bF$buf0),
    .Y(_6433_)
);

FILL FILL_1__7769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8710_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_750_),
    .C(_733_),
    .Y(_31_)
);

INVX1 _7360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .Y(_353_)
);

FILL FILL_1__12080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9915_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .Y(_1815_)
);

NOR2X1 _8565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1458_),
    .Y(_1459_)
);

NAND3X1 _8145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .B(_1053_),
    .C(_1056_),
    .Y(_1058_)
);

FILL FILL_1__10813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13285_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5271_),
    .C(_5450_),
    .Y(_5451_)
);

FILL FILL_0__12698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12278_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12563_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4217_),
    .CLK(clk_bF$buf51),
    .Q(\genblk1[5].u_ce.Acalc [2])
);

NAND3X1 _12143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4370_),
    .B(_4696_),
    .C(_4695_),
    .Y(_4699_)
);

FILL FILL_0__8605_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6137_),
    .B(_6111_),
    .C(_6136_),
    .Y(_6138_)
);

OAI21X1 _13348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5272_),
    .B(_5796_),
    .C(_5797_),
    .Y(_5059_)
);

FILL FILL_0__14844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_799_),
    .C(_800_),
    .Y(_37_)
);

OR2X2 _7416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_402_),
    .Y(_407_)
);

FILL FILL_2__13563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11549_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4399_),
    .C(_4402_),
    .Y(_4403_)
);

FILL FILL_0__9143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4043_),
    .B(_4036_),
    .Y(_4045_)
);

FILL FILL_0__12910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7158_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _12619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .Y(_5105_)
);

FILL FILL_1__14702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9304_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1641_),
    .C(_1658_),
    .Y(_889_)
);

NOR2X1 _8374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .B(_1276_),
    .Y(_1277_)
);

FILL FILL_1__10622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13094_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5248_),
    .B(_5267_),
    .C(_5268_),
    .Y(_5269_)
);

FILL FILL_0__12087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4913_),
    .B(_4362__bF$buf5),
    .Y(_4914_)
);

FILL FILL_2__12834_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2738_),
    .B(_2739_),
    .C(_2674_),
    .Y(_2740_)
);

INVX1 _9579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .Y(_2381_)
);

NAND2X1 _9159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .B(_1978_),
    .Y(_1982_)
);

FILL FILL_1__11827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .B(_6351_),
    .C(_6354_),
    .Y(_6357_)
);

INVX1 _13577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_5955_)
);

NOR2X1 _13157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5583_),
    .B(_5611_),
    .Y(_5617_)
);

FILL FILL_0__14653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10900_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_624_),
    .Y(_625_)
);

INVX1 _7225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .Y(_224_)
);

FILL FILL_2__13792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x248550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11358_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11643_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3383_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[4].u_ce.Acalc [6])
);

NAND2X1 _11223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3864_),
    .B(_3863_),
    .Y(_3865_)
);

FILL FILL_1__7387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14577_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .B(_5318_),
    .Y(_5322_)
);

NAND2X1 _12428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .B(_4966_),
    .Y(_4967_)
);

NAND3X1 _12008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .B(_4569_),
    .C(_4568_),
    .Y(_4570_)
);

FILL FILL_0__13924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9113_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1094_)
);

FILL FILL_1__10851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14709_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .B(_4734_),
    .C(_4675_),
    .Y(_4735_)
);

FILL FILL_2__12643_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2179_),
    .B(_2198_),
    .Y(_2201_)
);

FILL FILL_1__11216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8643_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3502_),
    .B(_3539_),
    .C(_3524__bF$buf2),
    .Y(_3569_)
);

FILL FILL_0__8223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .B(_5804_),
    .Y(_5820_)
);

FILL FILL_0__14462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .B(_807_),
    .Y(_823_)
);

OAI21X1 _7454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf4),
    .B(_442_),
    .C(_431_),
    .Y(_443_)
);

FILL FILL_2__13181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11587_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4439_),
    .Y(_4440_)
);

FILL FILL_0__9181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4079_),
    .B(_4078_),
    .Y(_4080_)
);

OAI21X1 _11032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3651_),
    .B(_3648_),
    .C(_3524__bF$buf0),
    .Y(_3682_)
);

NOR2X1 _8659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .B(_1546_),
    .Y(_866_)
);

NOR2X1 _8239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1147_),
    .B(_1126_),
    .Y(_1148_)
);

FILL FILL_1__7196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13799_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2399_),
    .B(_1848__bF$buf3),
    .Y(_2400_)
);

FILL FILL_1__13379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5136_),
    .B(_5139_),
    .C(_5109_),
    .Y(_5140_)
);

AOI21X1 _12237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4787_),
    .B(_4788_),
    .C(_4345_),
    .Y(_4789_)
);

FILL FILL_1__14740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10240_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7000_),
    .B(_6961_),
    .C(_7019_),
    .Y(_7020_)
);

FILL FILL_2__7265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12872_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(_2014_),
    .C(_2018_),
    .Y(_2019_)
);

FILL FILL_1__11865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8032_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10723_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2549_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Acalc [10])
);

FILL FILL_0__10438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10018_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2899_),
    .C(_3029_),
    .Y(_3030_)
);

NAND3X1 _13195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5643_),
    .B(_5645_),
    .C(_5652_),
    .Y(_5653_)
);

FILL FILL_0__14691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9657_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4491_),
    .B(_4492_),
    .Y(_4493_)
);

FILL FILL_0__9237_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [9]),
    .B(_3524__bF$buf4),
    .Y(_4132_)
);

FILL FILL_0__10191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8613_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_655_),
    .C(_156_),
    .Y(_661_)
);

OAI21X1 _7263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf0),
    .B(_258_),
    .C(_259_),
    .Y(_260_)
);

DFFPOSX1 _11681_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3421_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Ain1 [0])
);

FILL FILL_0__11396_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3900_),
    .Y(_3901_)
);

FILL FILL_2__11303_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8888_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_886_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Xin0 [1])
);

OAI21X1 _8468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1363_),
    .C(_1358_),
    .Y(_1367_)
);

NOR2X1 _8048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Xcalc [11]),
    .Y(_965_)
);

FILL FILL_0__7723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13188_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5356_),
    .B(_5354_),
    .C(_5358_),
    .Y(_5359_)
);

NAND2X1 _12466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4282_),
    .B(_4279_),
    .Y(_4997_)
);

NAND2X1 _12046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4603_),
    .B(_4585_),
    .Y(_4606_)
);

FILL FILL_0__13962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14327_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6838_),
    .B(_6843_),
    .Y(_6844_)
);

FILL FILL_2__7494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8681_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3581_),
    .B(_3510__bF$buf1),
    .C(_3605_),
    .D(_3582_),
    .Y(_3356_)
);

FILL FILL_0__8261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10667_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_3245_),
    .Y(_3246_)
);

FILL FILL_0__10247_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2844_),
    .Y(_2848_)
);

OAI21X1 _7739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_429_),
    .C(_711_),
    .Y(_712_)
);

OAI21X1 _7319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_312_),
    .C(_313_),
    .Y(_314_)
);

FILL FILL_2__13046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9466_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [4]),
    .Y(_4311_)
);

FILL FILL_0__9046_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3953_),
    .B(_3929_),
    .C(_3952_),
    .Y(_3954_)
);

FILL FILL_1__13820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14605_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_426_),
    .Y(_479_)
);

INVX1 _7072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [2]),
    .Y(_80_)
);

NAND2X1 _11490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [8]),
    .B(_3510__bF$buf0),
    .Y(_4115_)
);

NAND3X1 _11070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3684_),
    .B(_3687_),
    .C(_3717_),
    .Y(_3718_)
);

FILL FILL_1__9627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11532_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [6]),
    .B(_1581_),
    .Y(_1582_)
);

NOR2X1 _8277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1174_),
    .Y(_1184_)
);

FILL FILL_1__10945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7112_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [1]),
    .B(_5174__bF$buf1),
    .Y(_5175_)
);

INVX1 _12275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4817_),
    .Y(_4824_)
);

FILL FILL_0__13771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14556_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .Y(_7055_)
);

FILL FILL_0__14136_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [11]),
    .Y(_6707_)
);

OAI21X1 _14001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6305_),
    .C(_6360_),
    .Y(_6361_)
);

FILL FILL_2__12070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10476_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10761_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .CLK(clk_bF$buf9),
    .Q(\genblk1[3].u_ce.LoadCtl [0])
);

FILL FILL_0__10056_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3050_),
    .B(_3065_),
    .Y(_3067_)
);

FILL FILL_2__10803_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7968_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_52_),
    .CLK(clk_bF$buf18),
    .Q(\genblk1[0].u_ce.Yin12b [9])
);

NAND2X1 _7548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_514_),
    .Y(_533_)
);

AOI22X1 _7128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.Xcalc [1]),
    .C(_130_),
    .D(_92_),
    .Y(_131_)
);

FILL FILL_1__12688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9695_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4526_),
    .B(_4529_),
    .C(_4417_),
    .Y(_4530_)
);

FILL FILL_0__9275_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4157_),
    .B(_4159_),
    .C(_4161_),
    .Y(_3394_)
);

AOI21X1 _11126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3757_),
    .B(_3755_),
    .C(_3761_),
    .Y(_3772_)
);

FILL FILL_0__12622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11341_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1000_),
    .B(_999_),
    .S(_973__bF$buf4),
    .Y(_1001_)
);

FILL FILL_1__10334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7341_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf2),
    .B(_4641_),
    .Y(_4642_)
);

FILL FILL_2__8720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8546_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.Xcalc [0]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Xcalc [2]),
    .Y(_3477_)
);

FILL FILL_0__8126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12900_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5723_),
    .B(_5735_),
    .C(_5733_),
    .Y(_5742_)
);

FILL FILL_2__9505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14785_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6878_)
);

FILL FILL_0__14365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_6545_),
    .C(_6546_),
    .Y(_7071_[4])
);

FILL FILL_1__7502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11292_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .B(_3641_),
    .Y(_3642_)
);

INVX1 _10570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3280_),
    .Y(_3281_)
);

FILL FILL_0__10285_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_2884_)
);

FILL FILL_1__8707_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_738_),
    .Y(_748_)
);

OAI21X1 _7357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_260_),
    .C(_326_),
    .Y(_350_)
);

FILL FILL_2__13084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4343_),
    .C(_4346_),
    .Y(_4347_)
);

FILL FILL_0__9084_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .B(_3989_),
    .C(_3987_),
    .Y(_3990_)
);

FILL FILL_2__11817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7817_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .Y(_2667_)
);

INVX1 _9503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .Y(_2310_)
);

FILL FILL_1__8460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13636_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949__bF$buf3),
    .B(_6284_),
    .C(_6263_),
    .Y(_5850_)
);

FILL FILL_0__13216_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13501_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[6].u_ce.Vld )
);

FILL FILL_1__9665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10143_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6929_),
    .B(_6924_),
    .Y(_6930_)
);

FILL FILL_0__7570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3324_),
    .Y(_3326_)
);

NAND2X1 _10206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [0]),
    .B(_2672__bF$buf4),
    .Y(_2937_)
);

NAND3X1 _13098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .B(_5560_),
    .C(_5501_),
    .Y(_5561_)
);

FILL FILL_2__9734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10001_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .B(_548_),
    .Y(_569_)
);

NAND3X1 _7166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .B(_164_),
    .C(_135__bF$buf4),
    .Y(_167_)
);

FILL FILL_0__11299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Y_ [1]),
    .Y(_4182_)
);

NAND2X1 _11164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3808_)
);

FILL FILL_2__11206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7206_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2504_)
);

NAND2X1 _9312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf2),
    .B(_2127_),
    .Y(_2128_)
);

INVX1 _12789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5265_),
    .Y(_5266_)
);

INVX1 _12369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [5]),
    .Y(_4911_)
);

FILL FILL_1__14452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13865_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6063_),
    .B(_6045_),
    .C(_6101_),
    .Y(_6102_)
);

FILL FILL_0__13025_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5757_),
    .B(_5760_),
    .Y(_5763_)
);

FILL FILL_1__9894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10372_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14515_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6503_),
    .CLK(clk_bF$buf58),
    .Q(\u_ot.Ycalc [3])
);

FILL FILL_1__11997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8584_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3506_),
    .Y(_3512_)
);

FILL FILL_0__8164_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3136_),
    .B(_3155_),
    .C(_2686__bF$buf5),
    .Y(_3156_)
);

NOR2X1 _10015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_2755_)
);

FILL FILL_0__11931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8325_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_297_),
    .C(_326_),
    .Y(_386_)
);

NOR2X1 _11393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4024_),
    .Y(_4025_)
);

FILL FILL_2__11855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7855_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .S(vdd),
    .Y(_2704_)
);

FILL FILL_0__7435_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [1]),
    .B(_1834__bF$buf2),
    .Y(_2345_)
);

AND2X2 _9121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1940_),
    .B(_1939_),
    .Y(_1946_)
);

DFFPOSX1 _12598_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4252_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ain12b [11])
);

INVX1 _12178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4731_),
    .Y(_4732_)
);

FILL FILL_1__14681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6963_),
    .B(_6964_),
    .Y(_6965_)
);

FILL FILL_0__14039_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [10]),
    .Y(_6623_)
);

FILL FILL_1__11386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8393_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [1]),
    .B(_3313_),
    .Y(_3346_)
);

FILL FILL_0__10379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf1),
    .B(_2973_),
    .C(_2966_),
    .Y(_2974_)
);

FILL FILL_0__11740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11320_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.Y_ [1]),
    .Y(_1668_)
);

FILL FILL_0__9598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4435_),
    .C(_4436_),
    .Y(_4437_)
);

FILL FILL_0__9178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4074_),
    .B(_4076_),
    .Y(_4077_)
);

OAI21X1 _11029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3591_),
    .C(_3678_),
    .Y(_3679_)
);

FILL FILL_1__13952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12945_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5280_),
    .B(_5279_),
    .Y(_5286_)
);

FILL FILL_0__12525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7664_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9770_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1682_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[2].u_ce.Ycalc [5])
);

FILL FILL_0__7244_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2162_),
    .C(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_2165_)
);

FILL FILL_2__8203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14688_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14553_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [4]),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.LoadCtl [5])
);

FILL FILL_0__14268_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [1]),
    .B(_6455_),
    .Y(_6474_)
);

FILL FILL_1__7825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11195_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3549_),
    .Y(_3550_)
);

FILL FILL257250x241350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10188_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3191_)
);

NAND3X1 _10053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2760_),
    .B(_2777_),
    .C(_2759_),
    .Y(_2791_)
);

FILL FILL_2__10515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9581_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1510_),
    .Y(_1511_)
);

OAI21X1 _8201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(_1110_),
    .C(_1111_),
    .Y(_1112_)
);

DFFPOSX1 _11678_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3418_),
    .CLK(clk_bF$buf26),
    .Q(\genblk1[4].u_ce.Ain12b [7])
);

OAI21X1 _11258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .B(_3897_),
    .C(_3524__bF$buf1),
    .Y(_3898_)
);

FILL FILL257250x208950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12334_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9826_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1738_),
    .CLK(clk_bF$buf76),
    .Q(\genblk1[2].u_ce.Ain12b [11])
);

INVX1 _9406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .Y(_2218_)
);

FILL FILL_1__8783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13959_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6150_),
    .B(_6172_),
    .C(_6158_),
    .Y(_6192_)
);

FILL FILL_0__13539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [1]),
    .B(_5796_),
    .Y(_5829_)
);

FILL FILL_1__9988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10046_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6841_)
);

FILL FILL_0__7893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8678_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3600_),
    .B(_3602_),
    .Y(_3603_)
);

FILL FILL_0__8258_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3242_),
    .Y(_3243_)
);

NAND2X1 _10109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2843_),
    .B(_2844_),
    .Y(_2845_)
);

FILL FILL_0__11605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14497_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6982_),
    .B(_6981_),
    .Y(_6999_)
);

FILL FILL_0__14077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6541_),
    .B(\u_ot.LoadCtl_6_bF$buf4 ),
    .C(_6656_),
    .Y(_6502_)
);

FILL FILL_1__7634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13817_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [10]),
    .Y(_3010_)
);

FILL FILL_1__8839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .C(_475_),
    .Y(_476_)
);

DFFPOSX1 _8850_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_848_),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.Ycalc [9])
);

OAI21X1 _8430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .B(_1329_),
    .C(_1065_),
    .Y(_1331_)
);

OAI21X1 _8010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(_921_),
    .C(_931_),
    .Y(\a[2] [0])
);

OR2X2 _11487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4104_),
    .B(_4112_),
    .Y(_4113_)
);

NAND2X1 _11067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3668_),
    .B(_3684_),
    .Y(_3715_)
);

FILL FILL_2__7703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7529_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2429_),
    .B(_2432_),
    .Y(_2433_)
);

FILL FILL_0__7109_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2035_),
    .Y(_2036_)
);

FILL FILL_1__8592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13768_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6007_),
    .B(_6008_),
    .Y(_6009_)
);

FILL FILL_0__13348_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5661_),
    .Y(_5670_)
);

FILL FILL_1__9377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7050_),
    .B(_7051_),
    .Y(_7052_)
);

NAND3X1 _14418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6701_),
    .C(_6704_),
    .Y(_6705_)
);

FILL FILL_2_BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12067_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_677_)
);

FILL FILL_0__8487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8067_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10758_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2584_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Ain1 [1])
);

NAND3X1 _10338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2690_),
    .B(_3061_),
    .C(_3057_),
    .Y(_3064_)
);

FILL FILL_1__12841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.ISin ),
    .B(_6826_),
    .Y(_6832_)
);

DFFPOSX1 _14171_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5847_),
    .CLK(clk_bF$buf10),
    .Q(\genblk1[7].u_ce.Ycalc [11])
);

DFFPOSX1 _8906_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_904_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Ain12b [7])
);

FILL FILL_1__7863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12619_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5375_),
    .Y(_5376_)
);

FILL FILL_1_BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2822_),
    .B(_2826_),
    .C(_2827_),
    .Y(_2828_)
);

FILL FILL_1__8648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8228_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_293_),
    .Y(_6_)
);

INVX1 _11296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .Y(_3934_)
);

FILL FILL_0__12792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7758_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2611_),
    .C(_2612_),
    .Y(_2613_)
);

FILL FILL_0__7338_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2248_),
    .C(_1903_),
    .Y(_2255_)
);

NAND2X1 _9024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_1853_)
);

FILL FILL_2__8717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13997_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6227_),
    .Y(_6228_)
);

FILL FILL_0__13577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13157_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13442_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5042_),
    .CLK(clk_bF$buf62),
    .Q(\genblk1[6].u_ce.Xcalc [1])
);

NAND2X1 _13022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [2]),
    .B(_5174__bF$buf1),
    .Y(_5488_)
);

FILL FILL_2__13904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10084_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(_6875_),
    .Y(_6771_)
);

OAI21X1 _14227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(_6543_),
    .C(_6544_),
    .Y(_7071_[3])
);

FILL FILL_0__7091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12296_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7930_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Xcalc [1])
);

NAND2X1 _7510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [10]),
    .Y(_496_)
);

FILL FILL_1__11289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3628_),
    .B(_3635_),
    .C(_3638_),
    .Y(_3639_)
);

FILL FILL_0__8296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2668_),
    .Y(_3278_)
);

OAI21X1 _10147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2880_),
    .C(_2878_),
    .Y(_2881_)
);

FILL FILL_1__12650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(_1598_),
    .Y(_1599_)
);

FILL FILL_1__7672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12848_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5193_)
);

FILL FILL_0__12428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8037_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6281_),
    .B(_6264_),
    .Y(_6282_)
);

FILL FILL_2__7741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .B(_2467_),
    .Y(_2468_)
);

FILL FILL_0__7147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2070_),
    .B(_2071_),
    .Y(_2072_)
);

FILL FILL_1__11921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14393_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6022_),
    .B(_6039_),
    .C(_6040_),
    .Y(_6045_)
);

FILL FILL_0__13386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5704_),
    .Y(_5706_)
);

FILL FILL_2__13713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9713_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14876_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6767_),
    .CLK(clk_bF$buf67),
    .Q(\u_pa.acc_reg [0])
);

OAI21X1 _14456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6731_),
    .B(_6733_),
    .C(_6735_),
    .Y(_6517_)
);

INVX1 _14036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6394_)
);

FILL FILL_1__7728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [6]),
    .B(_3441_),
    .Y(_3458_)
);

OAI21X1 _10376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3012_),
    .C(_3099_),
    .Y(_3100_)
);

FILL FILL_2__10418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x86550 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [10]),
    .Y(_1778_)
);

INVX1 _8524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .Y(_1420_)
);

NAND2X1 _8104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [4]),
    .Y(_1019_)
);

FILL FILL_1__7481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12657_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5410_),
    .B(_5411_),
    .Y(_5412_)
);

FILL FILL_0__12237_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .B(_4997_),
    .Y(_4263_)
);

OR2X2 _12102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4658_),
    .B(_4636_),
    .Y(_4660_)
);

OAI21X1 _9729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1952_),
    .B(_2486_),
    .C(_2502_),
    .Y(_1732_)
);

NAND2X1 _9309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2125_)
);

FILL FILL_1__8686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6095_),
    .B(_6098_),
    .Y(_6099_)
);

NAND2X1 _13307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5758_),
    .B(_5759_),
    .Y(_5760_)
);

FILL FILL_0__14803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2290_),
    .C(_2278_),
    .Y(_2291_)
);

AOI21X1 _9062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1885_),
    .C(_1888_),
    .Y(_1889_)
);

FILL FILL_1__11730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13195_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13480_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5080_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Yin1 [1])
);

NAND3X1 _13060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5196_),
    .B(_5522_),
    .C(_5521_),
    .Y(_5525_)
);

FILL FILL_2__13942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9102_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6905_),
    .B(_6909_),
    .Y(_6910_)
);

OR2X2 _14265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_6570_),
    .Y(_6572_)
);

FILL FILL_1__7537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14727_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2894_),
    .C(_2873_),
    .Y(_2918_)
);

FILL FILL_2__10647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11261_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [11]),
    .B(_996__bF$buf2),
    .Y(_1633_)
);

AOI21X1 _8333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1206_),
    .B(_1215_),
    .C(_1237_),
    .Y(_1238_)
);

FILL FILL_1__7290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12886_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5225_),
    .C(_5228_),
    .Y(_5229_)
);

FILL FILL_0__12466_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(vdd),
    .Y(_4876_)
);

FILL FILL_0__12046_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2693_),
    .S(_2648__bF$buf3),
    .Y(_2701_)
);

NAND2X1 _9538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2339_),
    .B(_2342_),
    .Y(_2343_)
);

OAI21X1 _9118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1942_),
    .C(_1939_),
    .Y(_1943_)
);

FILL FILL_1__8495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .B(_6317_),
    .C(_6315_),
    .Y(_6318_)
);

NAND2X1 _13536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5916_),
    .B(_5915_),
    .Y(\genblk1[7].u_ce.X_ [0])
);

INVX1 _13116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5575_),
    .Y(_5578_)
);

FILL FILL_0__14612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7185_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_2108_)
);

FILL FILL_0__10952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10112_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_498_),
    .C(_585_),
    .Y(_586_)
);

FILL FILL_2__13751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[4] [1]),
    .B(_4162_),
    .Y(_3427_)
);

NAND2X1 _14494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.Y_ [0]),
    .Y(_6757_)
);

OAI21X1 _14074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6348_),
    .C(_6376_),
    .Y(_6430_)
);

OAI21X1 _8809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_921_),
    .C(_1666_),
    .Y(_896_)
);

FILL FILL_1__7766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13109_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5282_),
    .C(_5279_),
    .Y(_5283_)
);

FILL FILL_2__10456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9912_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_1812_)
);

OAI22X1 _8562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1456_),
    .D(_1454_),
    .Y(_859_)
);

OAI21X1 _8142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_1025_),
    .C(_1010__bF$buf4),
    .Y(_1055_)
);

FILL FILL_1__10810_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3841_),
    .B(_3840_),
    .Y(_3842_)
);

FILL FILL_2__7415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13282_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5448_)
);

FILL FILL_0__12695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12275_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12560_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4214_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [11])
);

OAI21X1 _12140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4689_),
    .B(_4692_),
    .C(_4694_),
    .Y(_4696_)
);

DFFPOSX1 _9767_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1679_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Ycalc [2])
);

OAI21X1 _9347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2161_),
    .C(_2158_),
    .Y(_2162_)
);

FILL FILL_0__8602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14067_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [8]),
    .Y(_6135_)
);

NAND2X1 _13345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5106_),
    .B(_5109_),
    .Y(_5795_)
);

FILL FILL_0__14841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10341_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_92_),
    .Y(_798_)
);

NAND3X1 _7413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_380_),
    .C(_359_),
    .Y(_404_)
);

FILL FILL_2__13980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11546_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .S(vdd),
    .Y(_4400_)
);

FILL FILL_0__9140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11126_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4040_),
    .B(_4041_),
    .Y(_4042_)
);

INVX1 _8618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .Y(_1508_)
);

FILL FILL_1__7575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13338_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5102_)
);

FILL FILL_2__10685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9301_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1249_),
    .B(_1637_),
    .C(_1656_),
    .Y(_888_)
);

MUX2X1 _8371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(_1271_),
    .S(_973__bF$buf2),
    .Y(_1274_)
);

FILL FILL_2__7644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12831_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2721_),
    .B(_2736_),
    .Y(_2737_)
);

OAI21X1 _9576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .B(_2377_),
    .C(_2376_),
    .Y(_2378_)
);

NAND2X1 _9156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1977_),
    .B(_1978_),
    .Y(_1979_)
);

FILL FILL_1__11824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14296_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6352_),
    .C(_6353_),
    .Y(_6354_)
);

MUX2X1 _13574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(\genblk1[7].u_ce.Xin12b [6]),
    .S(vdd),
    .Y(_5952_)
);

FILL FILL_0__13289_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5614_),
    .C(_5171_),
    .Y(_5615_)
);

FILL FILL_0__14650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9616_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6994_),
    .B(_6996_),
    .C(_6833__bF$buf1),
    .Y(_6997_)
);

NOR2X1 _14359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .Y(_6654_)
);

FILL FILL_0__10990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10150_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_539_),
    .C(_585_),
    .Y(_622_)
);

INVX1 _7222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .Y(_221_)
);

DFFPOSX1 _10699_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2525_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [10])
);

OAI21X1 _10279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672__bF$buf4),
    .B(_3007_),
    .C(_2986_),
    .Y(_2529_)
);

FILL FILL_1__12782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11355_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11640_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3380_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[4].u_ce.Acalc [3])
);

NAND2X1 _11220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3861_),
    .B(_3860_),
    .Y(_3862_)
);

DFFPOSX1 _8847_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_845_),
    .CLK(clk_bF$buf14),
    .Q(\genblk1[1].u_ce.Ycalc [6])
);

NOR2X1 _8427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1327_),
    .B(_1326_),
    .Y(_1328_)
);

OAI21X1 _8007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .B(_925_),
    .C(_928_),
    .Y(_929_)
);

FILL FILL_1__7384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5317_),
    .B(_5318_),
    .Y(_5319_)
);

OAI21X1 _12425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4963_),
    .B(_4907_),
    .C(_4962_),
    .Y(_4964_)
);

NAND3X1 _12005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4560_),
    .B(_4566_),
    .C(_4564_),
    .Y(_4567_)
);

FILL FILL_0__13921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9110_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1067_),
    .B(_996__bF$buf0),
    .C(_1091_),
    .D(_1068_),
    .Y(_842_)
);

FILL FILL_0__14706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .B(_2119_),
    .C(_2136_),
    .Y(_2198_)
);

FILL FILL_2_BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8658_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3547_),
    .B(_3522_),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_3566_)
);

FILL FILL_2__8238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13098_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5818_)
);

FILL FILL_2__13425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9005_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [19]),
    .Y(_6829_)
);

DFFPOSX1 _14168_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5844_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Ycalc [8])
);

FILL FILL_1__8801_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_821_)
);

NAND2X1 _7451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf1),
    .B(_435_),
    .Y(_440_)
);

OAI21X1 _10088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .B(_2768_),
    .C(_2824_),
    .Y(_2825_)
);

FILL FILL_1__12171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11164_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .B(_1543_),
    .Y(_1544_)
);

NAND3X1 _8236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .B(_1143_),
    .C(_1144_),
    .Y(_1145_)
);

FILL FILL_1__7193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12789_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [4]),
    .Y(_5137_)
);

FILL FILL_0__12369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4772_),
    .B(_4762_),
    .C(_4785_),
    .Y(_4786_)
);

FILL FILL257550x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [5]),
    .Y(_6225_)
);

DFFPOSX1 _13439_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5039_),
    .CLK(clk_bF$buf77),
    .Q(\genblk1[6].u_ce.Ycalc [10])
);

OR2X2 _13019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .B(_5462_),
    .Y(_5486_)
);

OAI21X1 _14800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7015_),
    .B(_6867_),
    .C(_7016_),
    .Y(_7017_)
);

FILL FILL_2__7682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2012_),
    .B(_2015_),
    .C(_1903_),
    .Y(_2016_)
);

FILL FILL_1__11862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8467_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10720_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2546_),
    .CLK(clk_bF$buf4),
    .Q(\genblk1[3].u_ce.Acalc [7])
);

FILL FILL_0__10435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10015_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2640_),
    .B(_2672__bF$buf2),
    .C(_3027_),
    .D(_2670_),
    .Y(_2530_)
);

INVX1 _13192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5643_),
    .Y(_5650_)
);

DFFPOSX1 _7927_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.Ycalc [10])
);

OAI21X1 _7507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158__bF$buf3),
    .B(_493_),
    .C(_472_),
    .Y(_15_)
);

FILL FILL_2__13234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9654_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf0),
    .B(_4489_),
    .C(_4486_),
    .Y(_4490_)
);

FILL FILL_0__9234_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4127_),
    .B(_4129_),
    .C(_4115_),
    .Y(_3385_)
);

INVX1 _14397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [8]),
    .Y(_6686_)
);

FILL FILL_1__7669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8610_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_172__bF$buf3),
    .C(_414_),
    .Y(_658_)
);

NAND2X1 _7260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_257_)
);

FILL FILL_2__10779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11393_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8885_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_883_),
    .CLK(clk_bF$buf54),
    .Q(\genblk1[1].u_ce.Xin1 [0])
);

OAI21X1 _8465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1363_),
    .C(_1359_),
    .Y(_1364_)
);

AOI22X1 _8045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Xcalc [0]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Xcalc [2]),
    .Y(_963_)
);

FILL FILL_0__7720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .B(_5355_),
    .C(_5243_),
    .Y(_5356_)
);

FILL FILL_0__12178_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [1]),
    .Y(_4995_)
);

NAND2X1 _12043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4600_),
    .B(_4602_),
    .Y(_4603_)
);

FILL FILL_1__11918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8505_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6042_),
    .B(_6023_),
    .C(_5951_),
    .Y(_6043_)
);

INVX1 _13248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5702_),
    .Y(_5703_)
);

FILL FILL_0__14744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [4]),
    .B(_158__bF$buf4),
    .Y(_709_)
);

OAI21X1 _7316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_254_),
    .C(_310_),
    .Y(_311_)
);

FILL FILL_2__13043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11449_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [8]),
    .Y(_4308_)
);

FILL FILL_0__9043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11029_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3933_),
    .B(_3510__bF$buf4),
    .C(_3951_),
    .D(_3948_),
    .Y(_3372_)
);

FILL FILL_0__12810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5401_),
    .B(_5408_),
    .Y(_5409_)
);

OAI21X1 _12519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5025_),
    .B(_4993_),
    .C(_5026_),
    .Y(_4254_)
);

FILL FILL_1__14602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x248550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1578_),
    .Y(_1579_)
);

OAI21X1 _8274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1153_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1181_),
    .Y(_846_)
);

FILL FILL_1__10942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10102_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 )
);

FILL FILL_2__7127_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 )
);

OAI21X1 _12692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5167_),
    .B(_5169_),
    .C(_5172_),
    .Y(_5173_)
);

BUFX2 BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .Y(_6833__bF$buf4)
);

OAI21X1 _12272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4820_),
    .B(_4811_),
    .C(_4346_),
    .Y(_4822_)
);

OAI21X1 _9899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2641_),
    .B(_2642_),
    .C(_2643_),
    .Y(_2644_)
);

NAND3X1 _9479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf0),
    .B(_2282_),
    .C(_2280_),
    .Y(_2288_)
);

MUX2X1 _9059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .S(gnd),
    .Y(_1886_)
);

FILL FILL_1__11727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8314_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6261_),
    .B(_6260_),
    .C(_5951_),
    .Y(_6262_)
);

DFFPOSX1 _13477_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5077_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [4])
);

OAI21X1 _13057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .B(_5518_),
    .C(_5520_),
    .Y(_5522_)
);

FILL FILL_2__13939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10800_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7965_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_49_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Yin12b [10])
);

NAND3X1 _7545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_529_),
    .C(_528_),
    .Y(_530_)
);

OAI21X1 _7125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(\genblk1[0].u_ce.Xcalc [9]),
    .C(_86_),
    .Y(_128_)
);

FILL FILL_2__13692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9692_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4526_),
    .Y(_4527_)
);

FILL FILL_0__9272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11258_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(_4159_),
    .Y(_4160_)
);

NAND2X1 _11123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3767_),
    .B(_3768_),
    .Y(_3769_)
);

FILL FILL257250x158550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7287_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .S(gnd),
    .Y(_5226_)
);

INVX1 _12328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4873_)
);

FILL FILL_1__14831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9013_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_992_),
    .Y(_998_)
);

FILL FILL_1__10331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4639_)
);

NOR2X1 _9288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1840_),
    .Y(_2105_)
);

FILL FILL_1__11956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8543_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [6]),
    .B(_3441_),
    .Y(_3474_)
);

FILL FILL_0__8123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10109_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _13286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5113_),
    .B(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .C(_5737_),
    .D(_5739_),
    .Y(_5055_)
);

FILL FILL_0__14782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8704_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(\genblk1[0].u_ce.Ain12b [6]),
    .Y(_745_)
);

AOI21X1 _7354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_320_),
    .C(_345_),
    .Y(_347_)
);

FILL FILL_2__13081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11487_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf4),
    .B(_4325__bF$buf4),
    .Y(_4344_)
);

FILL FILL_0__9081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11067_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3981_),
    .C(_3986_),
    .Y(_3987_)
);

FILL FILL_1__9909_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .Y(_1809_)
);

INVX1 _8559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .Y(_1454_)
);

AOI21X1 _8139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(_1008_),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_1052_)
);

FILL FILL_1__7096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7814_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2663_),
    .B(_2656_),
    .S(_2648__bF$buf4),
    .Y(_2664_)
);

FILL FILL_1__13699_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2306_),
    .B(_2297_),
    .C(_1832_),
    .Y(_2308_)
);

FILL FILL_1__13279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5180_),
    .Y(_5445_)
);

DFFPOSX1 _12557_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4211_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xcalc [8])
);

OR2X2 _12137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4689_),
    .B(_4692_),
    .Y(_4693_)
);

FILL FILL_1__14640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14418_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [9]),
    .Y(_6927_)
);

FILL FILL_2__7165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12772_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1921_),
    .C(_1922_),
    .Y(_1923_)
);

FILL FILL_1__11765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8352_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_3324_)
);

FILL FILL_0__10338_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(_2934_),
    .C(_2741_),
    .Y(_2935_)
);

INVX1 _13095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .Y(_5558_)
);

FILL FILL_0__14591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9557_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4342_),
    .B(_4389_),
    .C(_4387_),
    .Y(_4397_)
);

FILL FILL_0__9137_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .B(vdd),
    .S(_4037_),
    .Y(_4039_)
);

FILL FILL_1__13911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8513_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_560_),
    .C(_563_),
    .Y(_566_)
);

INVX2 _7163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_164_)
);

OAI21X1 _11581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(_3435_),
    .C(_4180_),
    .Y(_3410_)
);

FILL FILL_0__11296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3805_)
);

FILL FILL_1__9718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11203_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1637_),
    .Y(_1655_)
);

OAI21X1 _8368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1133_),
    .C(_1270_),
    .Y(_1271_)
);

FILL FILL_1__10616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5261_),
    .C(_5262_),
    .Y(_5263_)
);

OAI21X1 _12366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4906_),
    .B(_4907_),
    .C(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .Y(_4909_)
);

FILL FILL_0__13862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14227_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14512_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6500_),
    .CLK(clk_bF$buf9),
    .Q(\u_ot.Ycalc [0])
);

FILL FILL_1__11994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8581_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3484_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3509_),
    .Y(_3352_)
);

FILL FILL_2__8179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10147_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3071_),
    .C(_3099_),
    .Y(_3153_)
);

NAND2X1 _10012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf0),
    .B(_2703_),
    .Y(_2752_)
);

NAND2X1 _7639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xcalc [9]),
    .B(_158__bF$buf0),
    .Y(_619_)
);

NAND2X1 _7219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_217_),
    .Y(_218_)
);

FILL FILL_1__12779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9366_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11637_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3377_),
    .CLK(clk_bF$buf69),
    .Q(\genblk1[4].u_ce.Acalc [0])
);

AOI21X1 _11217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3857_),
    .B(_3858_),
    .C(_3532_),
    .Y(_3859_)
);

FILL FILL_1__13720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8322_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_382_),
    .C(_230_),
    .Y(_384_)
);

FILL FILL_0__13918_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4015_),
    .Y(_4022_)
);

FILL FILL_1__9947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11012_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1488_),
    .B(_1489_),
    .Y(_1490_)
);

NAND2X1 _8177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1086_),
    .B(_1088_),
    .Y(_1089_)
);

FILL FILL_1__10845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7432_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12595_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4249_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin0 [0])
);

AOI21X1 _12175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf0),
    .B(_4687_),
    .C(_4728_),
    .Y(_4729_)
);

FILL FILL_0__13671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8637_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3486__bF$buf3),
    .Y(_3563_)
);

FILL FILL_0__8217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14456_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6957_),
    .B(_6916_),
    .C(_6961_),
    .Y(_6962_)
);

FILL FILL_0__14036_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6620_),
    .B(_6619_),
    .Y(_6621_)
);

FILL FILL_1__11383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8390_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2685_),
    .C(_3344_),
    .Y(_2574_)
);

FILL FILL_0__10376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2790_),
    .C(_2970_),
    .Y(_2971_)
);

INVX1 _7868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(_819_)
);

NAND2X1 _7448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_436_),
    .Y(_437_)
);

FILL FILL_1__12168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9595_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4433_),
    .C(_4424_),
    .Y(_4434_)
);

FILL FILL_0__9175_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3780_),
    .B(_3593_),
    .C(_3524__bF$buf2),
    .Y(_4074_)
);

INVX1 _11026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3676_)
);

FILL FILL_2__11908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8026_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10717_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2543_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Acalc [4])
);

FILL FILL_1__12800_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5646_),
    .B(_5637_),
    .C(_5172_),
    .Y(_5648_)
);

FILL FILL_2__9405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14685_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14550_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\u_ot.LoadCtl [1]),
    .CLK(clk_bF$buf38),
    .Q(\u_ot.LoadCtl [2])
);

FILL FILL_0__14265_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5974_),
    .C(_6472_),
    .Y(_5871_)
);

FILL FILL_1__7822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11192_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3546_),
    .B(_3543_),
    .S(_3486__bF$buf0),
    .Y(_3547_)
);

FILL FILL_0__10185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_3176_),
    .C(_2686__bF$buf1),
    .Y(_3188_)
);

AOI22X1 _10050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2672__bF$buf0),
    .C(_2788_),
    .D(_2744_),
    .Y(_2519_)
);

FILL FILL_1__8607_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_648_),
    .C(_654_),
    .Y(_655_)
);

AOI21X1 _7257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_248_),
    .C(_249_),
    .Y(_254_)
);

FILL FILL_1__12397_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11675_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3415_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[4].u_ce.Ain12b [8])
);

NAND3X1 _11255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf5),
    .B(_3894_),
    .C(_3889_),
    .Y(_3895_)
);

FILL FILL_2__11717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7717_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9823_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1735_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Yin0 [0])
);

AOI21X1 _9403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf1),
    .B(_2173_),
    .C(_2214_),
    .Y(_2215_)
);

FILL FILL_1__8780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13956_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6184_),
    .B(_6188_),
    .Y(_6189_)
);

FILL FILL_0__13536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13116_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5187_),
    .C(_5827_),
    .Y(_5082_)
);

FILL FILL_1__9985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10043_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[0]),
    .B(\u_pa.acc_reg [0]),
    .Y(_6838_)
);

FILL FILL_0__7890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8675_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3585_),
    .B(_3596_),
    .C(_3599_),
    .Y(_3600_)
);

FILL FILL_0__8255_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3239_),
    .B(_3235_),
    .Y(_3240_)
);

NAND3X1 _10106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2841_),
    .C(_2837_),
    .Y(_2842_)
);

FILL FILL_2__9634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8416_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_467_),
    .C(_465_),
    .Y(_473_)
);

FILL FILL_0__11199_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4109_),
    .Y(_4110_)
);

AOI21X1 _11064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3699_),
    .B(_3712_),
    .C(_3512_),
    .Y(_3713_)
);

FILL FILL_2__11946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7526_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf3),
    .B(_2347_),
    .Y(_2430_)
);

FILL FILL_0__7106_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2028_),
    .C(_2026_),
    .Y(_2033_)
);

NAND2X1 _12689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf3),
    .B(_5151__bF$buf1),
    .Y(_5170_)
);

NAND2X1 _12269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4425_),
    .B(_4818_),
    .Y(_4819_)
);

FILL FILL_1__14772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13765_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6004_),
    .B(_6005_),
    .Y(_6006_)
);

FILL FILL_0__13345_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5666_),
    .B(_5667_),
    .Y(_5668_)
);

FILL FILL_1__9374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10272_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7037_),
    .B(_7042_),
    .C(_7048_),
    .Y(_7049_)
);

INVX1 _14415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [10]),
    .Y(_6702_)
);

FILL FILL_2__12484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8064_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10755_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2581_),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[3].u_ce.Ain12b [4])
);

NAND2X1 _10335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3055_),
    .B(_3060_),
    .Y(_3061_)
);

FILL FILL_0__11831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13689_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8903_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_901_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Ain12b [8])
);

FILL FILL_1__7860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5368_),
    .C(_5366_),
    .Y(_5373_)
);

FILL FILL_0__12616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14408_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_275_),
    .B(_290_),
    .Y(_291_)
);

NAND2X1 _11293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .B(_3931_),
    .Y(_3932_)
);

FILL FILL_2__11755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7755_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2608_),
    .C(_2609_),
    .Y(_2610_)
);

FILL FILL_0__7335_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2244_),
    .B(_2226_),
    .C(_2224_),
    .Y(_2252_)
);

NAND2X1 _9021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_1850_)
);

NAND2X1 _12498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_5000_),
    .Y(_5015_)
);

NOR2X1 _12078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4336_),
    .B(_4633_),
    .Y(_4636_)
);

FILL FILL_1__14581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6872_),
    .B(_6871_),
    .Y(_6873_)
);

OAI21X1 _14224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_6541_),
    .C(_6542_),
    .Y(_7071_[2])
);

FILL FILL_1__11286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _10984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3614_),
    .C(_3586_),
    .Y(_3636_)
);

FILL FILL_0__8293_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3274_),
    .C(_2672__bF$buf1),
    .Y(_3276_)
);

FILL FILL_0__10279_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2877_),
    .B(_2849_),
    .Y(_2878_)
);

FILL FILL_2__9672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11220_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1595_),
    .Y(_1596_)
);

FILL FILL_0__9498_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4323_),
    .B(_4340_),
    .Y(_4341_)
);

FILL FILL_0__9078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3984_),
    .B(_3983_),
    .C(_3971_),
    .Y(_3374_)
);

FILL FILL_1__13852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12845_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5190_)
);

FILL FILL_0__12425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12005_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(vdd),
    .Y(_2661_)
);

FILL FILL_1__8454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x241350 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6278_),
    .Y(_6279_)
);

FILL FILL_1__9659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x208950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7564_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .Y(_2465_)
);

FILL FILL_0__7144_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2068_),
    .Y(_2069_)
);

FILL FILL_2__8943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9710_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14873_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6764_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [4])
);

FILL FILL_0__14588_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [6]),
    .B(_6733_),
    .Y(_6734_)
);

OAI21X1 _14033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .B(_6386_),
    .C(_6382_),
    .Y(_6391_)
);

FILL FILL_1__7725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11095_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(\genblk1[4].u_ce.Ycalc [8]),
    .C(_3438_),
    .Y(_3455_)
);

FILL FILL_0__10088_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3073_),
    .B(_3075_),
    .Y(_3097_)
);

FILL FILL_2__9481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1772_),
    .B(_1775_),
    .C(_1768_),
    .Y(_1776_)
);

NAND2X1 _8521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .B(_1417_),
    .Y(_1418_)
);

OAI21X1 _8101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1014_),
    .C(_1015_),
    .Y(_1016_)
);

INVX1 _11998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_4560_)
);

OAI21X1 _11578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_4179_)
);

OAI21X1 _11158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3523_),
    .C(_3801_),
    .Y(_3802_)
);

FILL FILL_1__13661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2486_),
    .Y(_2501_)
);

NOR2X1 _9306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .B(_2119_),
    .Y(_2122_)
);

FILL FILL_1__8683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13859_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf1),
    .B(_6092_),
    .C(_6087_),
    .Y(_6096_)
);

FILL FILL_0__13019_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [7]),
    .Y(_5757_)
);

FILL FILL_0__14800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10366_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14509_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6497_),
    .CLK(clk_bF$buf46),
    .Q(\u_ot.Xcalc [9])
);

FILL FILL_0__7793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8578_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3506_),
    .C(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_3507_)
);

FILL FILL_0__8158_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3128_),
    .Y(_3150_)
);

INVX1 _10009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .Y(_2749_)
);

FILL FILL_1__12932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6907_)
);

OAI21X1 _14262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf2),
    .B(_6568_),
    .C(_6569_),
    .Y(_6489_)
);

FILL FILL_1__7534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13717_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2873_),
    .B(_2895_),
    .C(_2881_),
    .Y(_2915_)
);

FILL FILL_1__8739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10644_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_380_),
    .Y(_381_)
);

AND2X2 _8750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1626_),
    .B(_1630_),
    .Y(_1631_)
);

NAND3X1 _8330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .B(_1229_),
    .C(_1234_),
    .Y(_1235_)
);

NAND2X1 _11387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [0]),
    .B(_3510__bF$buf2),
    .Y(_4020_)
);

FILL FILL_2__7603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7849_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2698_)
);

FILL FILL_0__7429_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain0 [0]),
    .Y(_2340_)
);

OAI21X1 _9115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1910_),
    .C(_1848__bF$buf4),
    .Y(_1940_)
);

FILL FILL_1__8492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13668_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6314_),
    .B(_6312_),
    .Y(_6315_)
);

FILL FILL_0_BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13248_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(_5912_),
    .C(_5913_),
    .Y(_5914_)
);

FILL FILL_0_BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5494_),
    .C(_5574_),
    .Y(_5575_)
);

FILL FILL_0_BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10175_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6949_),
    .Y(_6959_)
);

INVX1 _14318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xcalc [9]),
    .Y(_6618_)
);

FILL FILL_0__7182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_561_),
    .Y(_583_)
);

FILL FILL_0__8387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.Y_ [0]),
    .Y(_3343_)
);

OAI21X1 _10238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2836_),
    .C(_2967_),
    .Y(_2968_)
);

FILL FILL_1__12741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11314_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6740_),
    .C(_6755_),
    .Y(_6532_)
);

NOR2X1 _14071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6405_),
    .Y(_6427_)
);

OAI21X1 _8806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1665_)
);

FILL FILL_1__7763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12939_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5259_),
    .B(_5250_),
    .C(_5188__bF$buf5),
    .Y(_5280_)
);

FILL FILL_0__12519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10453_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_188_),
    .C(_196_),
    .Y(_199_)
);

NAND3X1 _11196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(_3838_),
    .C(_3836_),
    .Y(_3839_)
);

FILL FILL_2__7832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7658_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9764_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1676_),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Ycalc [0])
);

FILL FILL_0__7238_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .Y(_2159_)
);

FILL FILL_2__8617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13897_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6132_),
    .Y(_6133_)
);

OAI21X1 _13342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5791_),
    .B(_5787_),
    .C(_5790_),
    .Y(_5793_)
);

FILL FILL_0__13057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9086_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14547_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6535_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Yin0 [1])
);

NAND2X1 _14127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.X_ [0]),
    .Y(_6471_)
);

FILL FILL_1__7819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_788_),
    .C(_791_),
    .Y(_796_)
);

NAND3X1 _7410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(_381_),
    .C(_367_),
    .Y(_401_)
);

FILL FILL_1__11189_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .S(gnd),
    .Y(_3544_)
);

FILL FILL_0__8196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_3185_)
);

NAND2X1 _10047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2785_),
    .B(_2782_),
    .Y(_2786_)
);

FILL FILL_1__12970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11123_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [0]),
    .B(_996__bF$buf2),
    .Y(_1506_)
);

FILL FILL_1__7572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12748_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12613_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl [3]),
    .CLK(clk_bF$buf32),
    .Q(\genblk1[5].u_ce.LoadCtl [4])
);

FILL FILL_0__12328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10682_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6180_),
    .B(_5963__bF$buf3),
    .Y(_6186_)
);

FILL FILL_2__7641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7887_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .B(_2729_),
    .C(_2732_),
    .Y(_2734_)
);

FILL FILL_0__7467_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1811__bF$buf0),
    .Y(_2375_)
);

NAND3X1 _9153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf4),
    .B(_1975_),
    .C(_1972_),
    .Y(_1976_)
);

FILL FILL_1__11821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14293_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf5),
    .B(_6350_),
    .C(_6347_),
    .Y(_6351_)
);

INVX4 _13571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Vld ),
    .Y(_5949_)
);

FILL FILL_0__13286_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5598_),
    .B(_5588_),
    .C(_5611_),
    .Y(_5612_)
);

FILL FILL_2__13613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9613_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6983_),
    .B(_6980_),
    .C(_6988_),
    .Y(_6994_)
);

INVX1 _14356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin1 [0]),
    .Y(_6651_)
);

FILL FILL_1__7628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7208_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10696_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2522_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Ycalc [7])
);

AND2X2 _10276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3004_),
    .B(_2987_),
    .Y(_3005_)
);

FILL FILL_0__11772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11352_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8844_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_842_),
    .CLK(clk_bF$buf12),
    .Q(\genblk1[1].u_ce.Ycalc [3])
);

NAND3X1 _8424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(_1324_),
    .C(_1322_),
    .Y(_1325_)
);

INVX2 _8004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_926_)
);

FILL FILL_1__7381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12977_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf5),
    .B(_5315_),
    .C(_5312_),
    .Y(_5316_)
);

FILL FILL_0__12137_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4950_),
    .B(_4936_),
    .Y(_4961_)
);

NAND3X1 _12002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4563_),
    .C(_4562_),
    .Y(_4564_)
);

INVX1 _9629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [7]),
    .Y(_2427_)
);

OAI21X1 _9209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2028_),
    .C(_2029_),
    .Y(_2030_)
);

FILL FILL_1__8586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _13627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6002_),
    .B(_5953_),
    .C(_6001_),
    .D(_5945_),
    .Y(_6003_)
);

NAND2X1 _13207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5664_),
    .B(_5661_),
    .Y(_5665_)
);

FILL FILL_0__14703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2194_),
    .Y(_2195_)
);

FILL FILL_1__11210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13095_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5816_)
);

FILL FILL_2__13842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9002_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [5]),
    .Y(_6826_)
);

DFFPOSX1 _14165_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5841_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Ycalc [5])
);

FILL FILL_1__7857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2818_),
    .B(_2821_),
    .Y(_2822_)
);

FILL FILL_2__10967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11161_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1540_),
    .Y(_1541_)
);

NAND3X1 _8233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(_1138_),
    .C(_1141_),
    .Y(_1142_)
);

FILL FILL_1__7190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12786_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [8]),
    .Y(_5134_)
);

FILL FILL_0__12366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4776_),
    .B(_4779_),
    .Y(_4783_)
);

OAI21X1 _9858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(_2597_),
    .C(_2607_),
    .Y(\a[4] [0])
);

AND2X2 _9438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2241_),
    .B(_2242_),
    .Y(_2249_)
);

INVX1 _9018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_1847_)
);

FILL FILL_1__8395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14158_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf2),
    .B(_6218_),
    .C(_6221_),
    .Y(_6222_)
);

DFFPOSX1 _13436_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5036_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [7])
);

NAND3X1 _13016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5199_),
    .B(_5480_),
    .C(_5477_),
    .Y(_5483_)
);

FILL FILL_1__10498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7085_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2012_),
    .Y(_2013_)
);

FILL FILL_0__10852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7924_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf13),
    .Q(\genblk1[0].u_ce.Ycalc [7])
);

AND2X2 _7504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_473_),
    .Y(_491_)
);

FILL FILL_2__13651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9651_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4448_),
    .B(_4325__bF$buf1),
    .C(_4469_),
    .Y(_4487_)
);

FILL FILL_0__9231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11217_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4121_),
    .B(_4126_),
    .Y(_4127_)
);

NAND3X1 _14394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6682_),
    .B(_6683_),
    .C(_6677_),
    .Y(_6684_)
);

OR2X2 _8709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1509_),
    .B(_1010__bF$buf4),
    .Y(_1593_)
);

FILL FILL257550x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13009_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5187_)
);

FILL FILL_2__10356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11390_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8882_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_880_),
    .CLK(clk_bF$buf48),
    .Q(\genblk1[1].u_ce.Xin12b [7])
);

OAI21X1 _8462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1341_),
    .B(_1360_),
    .C(_1010__bF$buf2),
    .Y(_1361_)
);

NAND2X1 _8042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [6]),
    .B(_927_),
    .Y(_960_)
);

INVX1 _11099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .Y(_3746_)
);

FILL FILL_2__7315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13182_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .Y(_5353_)
);

FILL FILL_0__12175_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4988_),
    .B(_4275_),
    .Y(_4993_)
);

NAND2X1 _12040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .B(_4514_),
    .Y(_4600_)
);

FILL FILL_2__12922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2456_),
    .C(_2445_),
    .Y(_2462_)
);

NAND2X1 _9247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_2065_),
    .Y(_2066_)
);

FILL FILL_1__11915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14387_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6038_),
    .B(_6035_),
    .C(_6024_),
    .Y(_6040_)
);

NAND2X1 _13245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain1 [0]),
    .B(_5699_),
    .Y(_5700_)
);

FILL FILL_0__14741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10241_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .B(_697_),
    .C(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .Y(_707_)
);

NAND2X1 _7313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_307_),
    .Y(_308_)
);

FILL FILL_2__13880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11446_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4302_),
    .B(_4305_),
    .C(_4282_),
    .Y(_4306_)
);

FILL FILL_0__9040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3934_),
    .B(_3924_),
    .Y(_3949_)
);

INVX1 _8938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [5]),
    .Y(_1773_)
);

OAI21X1 _8518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1413_),
    .C(_1414_),
    .Y(_1415_)
);

FILL FILL_1__7895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf1),
    .B(_5405_),
    .Y(_5406_)
);

OAI21X1 _12516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5023_),
    .B(_4993_),
    .C(_5024_),
    .Y(_4253_)
);

FILL FILL_2__10585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9201_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1555_),
    .C(_1575_),
    .Y(_1576_)
);

OAI21X1 _8271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf5),
    .B(_1065_),
    .C(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .Y(_1179_)
);

BUFX2 BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf3 )
);

FILL FILL_2__7544_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf2 )
);

FILL FILL_2__7124_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf5)
);

BUFX2 BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf4)
);

BUFX2 BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf3)
);

BUFX2 BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf2)
);

BUFX2 BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf1)
);

BUFX2 BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .Y(_1848__bF$buf0)
);

FILL FILL_2__12731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert384 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Xcalc [11]),
    .Y(_2641_)
);

OAI21X1 _9476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2259_),
    .C(_1848__bF$buf0),
    .Y(_2285_)
);

FILL FILL_2_CLKBUF1_insert387 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1828_),
    .B(_1875_),
    .C(_1873_),
    .Y(_1883_)
);

FILL FILL_2_CLKBUF1_insert389 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8329_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6257_),
    .B(_6258_),
    .Y(_6259_)
);

FILL FILL_0__13189_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13474_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5074_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [9])
);

OR2X2 _13054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .B(_5518_),
    .Y(_5519_)
);

FILL FILL_0__14130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9516_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6902_),
    .B(_6903_),
    .C(_6904_),
    .Y(_6774_)
);

OAI21X1 _14259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6561_),
    .C(_6566_),
    .Y(_6567_)
);

FILL FILL_0__10890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10050_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7962_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_46_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin1 [1])
);

NAND3X1 _7542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(_526_),
    .C(_524_),
    .Y(_527_)
);

NAND2X1 _7122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(_124_),
    .Y(\genblk1[0].u_ce.X_ [0])
);

OAI21X1 _10599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3306_),
    .B(_3302_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_3308_)
);

NAND2X1 _10179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2907_),
    .B(_2911_),
    .Y(_2912_)
);

FILL FILL_1__12682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12262_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4517_),
    .B(_4520_),
    .Y(_4524_)
);

FILL FILL_0__11255_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Xin12b [9]),
    .Y(_4158_)
);

INVX1 _11120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .Y(_3766_)
);

NAND2X1 _8747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1627_),
    .Y(_1628_)
);

INVX1 _8327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .Y(_1232_)
);

FILL FILL_1__7284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13047_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5168_),
    .B(_5215_),
    .C(_5213_),
    .Y(_5223_)
);

NAND2X1 _12325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4860_),
    .B(_4869_),
    .Y(_4871_)
);

FILL FILL_0__13821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9010_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_995_),
    .Y(_838_)
);

FILL FILL_0__14606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2100_),
    .C(_2101_),
    .Y(_2102_)
);

FILL FILL_1__11953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8558_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Xcalc [10]),
    .C(_3438_),
    .Y(_3471_)
);

FILL FILL_0__8120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10106_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5736_),
    .B(_5727_),
    .Y(_5737_)
);

FILL FILL_1__12738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9325_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [5]),
    .B(_6737_),
    .Y(_6754_)
);

INVX1 _14068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [10]),
    .Y(_6424_)
);

FILL FILL_1__8701_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_699_),
    .C(_172__bF$buf3),
    .Y(_742_)
);

INVX1 _7351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [8]),
    .Y(_344_)
);

FILL FILL_1__12491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9906_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Xcalc [1]),
    .C(_1806_),
    .D(_1768_),
    .Y(_1807_)
);

NAND2X1 _8556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1445_),
    .B(_1447_),
    .Y(_1451_)
);

NAND2X1 _8136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_972__bF$buf2),
    .Y(_1049_)
);

FILL FILL_1__7093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13276_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5440_),
    .C(_5441_),
    .Y(_5442_)
);

FILL FILL_0__12689_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12554_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4208_),
    .CLK(clk_bF$buf70),
    .Q(\genblk1[5].u_ce.Xcalc [5])
);

FILL FILL_0__12269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4431_),
    .B(_4638_),
    .Y(_4690_)
);

FILL FILL_0__13630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6099_),
    .B(_6103_),
    .C(_6098_),
    .Y(_6130_)
);

NAND2X1 _13339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [10]),
    .B(_5188__bF$buf4),
    .Y(_5790_)
);

FILL FILL_0__14835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6919_),
    .B(_6916_),
    .C(_6917_),
    .Y(_6924_)
);

FILL FILL_2__7582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf1),
    .B(_1919_),
    .C(_1910_),
    .Y(_1920_)
);

FILL FILL_1__11762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3316_),
    .B(_3321_),
    .C(_3322_),
    .Y(_2555_)
);

FILL FILL_0__10335_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .Y(_2932_)
);

AOI21X1 _13092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf4),
    .B(_5513_),
    .C(_5554_),
    .Y(_5555_)
);

OAI21X1 _7827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_788_),
    .C(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .Y(_794_)
);

NAND2X1 _7407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_397_),
    .Y(_398_)
);

FILL FILL_2__13134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9554_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(\genblk1[4].u_ce.ISout ),
    .Y(_4395_)
);

FILL FILL_0__9134_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4035_),
    .B(_4028_),
    .C(_4033_),
    .Y(_4036_)
);

NAND2X1 _14297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6598_),
    .B(_6599_),
    .Y(_6600_)
);

FILL FILL_0__12901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8510_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_561_),
    .C(_562_),
    .Y(_563_)
);

MUX2X1 _7160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(\genblk1[0].u_ce.Xin12b [6]),
    .S(gnd),
    .Y(_161_)
);

FILL FILL_0__11293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9715_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_984_),
    .C(_1653_),
    .Y(_885_)
);

AOI22X1 _8365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .B(_1266_),
    .C(_1267_),
    .D(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1268_)
);

FILL FILL_1__10613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13085_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf0),
    .B(_5259_),
    .C(_5250_),
    .Y(_5260_)
);

FILL FILL_0__12498_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4905_),
    .B(_4904_),
    .Y(_4906_)
);

FILL FILL_0__12078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8405_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf3),
    .B(_6307_),
    .C(_6329_),
    .Y(_6348_)
);

INVX2 _13568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5946_),
    .Y(_5947_)
);

NAND2X1 _13148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5602_),
    .B(_5605_),
    .Y(_5609_)
);

FILL FILL_0__14644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10144_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_614_),
    .Y(_617_)
);

NAND2X1 _7216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .B(_214_),
    .Y(_215_)
);

FILL FILL_2__13363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11349_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11634_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3374_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [9])
);

OAI21X1 _11214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3835_),
    .B(_3826_),
    .C(_3524__bF$buf1),
    .Y(_3856_)
);

FILL FILL_0__12710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7378_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5274_),
    .B(_5151__bF$buf2),
    .C(_5295_),
    .Y(_5313_)
);

AOI21X1 _12419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4955_),
    .B(_4891_),
    .C(\genblk1[5].u_ce.Ain12b [8]),
    .Y(_4958_)
);

FILL FILL_0__13915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(_1483_),
    .Y(_1487_)
);

NAND3X1 _8174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1071_),
    .B(_1082_),
    .C(_1085_),
    .Y(_1086_)
);

FILL FILL_1__10842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x158550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10002_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12592_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4246_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Yin12b [5])
);

OAI21X1 _12172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4721_),
    .B(_4704_),
    .C(_4717_),
    .Y(_4726_)
);

DFFPOSX1 _9799_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1711_),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[2].u_ce.Acalc [10])
);

OAI21X1 _9379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2061_),
    .C(_2191_),
    .Y(_2192_)
);

FILL FILL_1__11207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8634_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(\genblk1[4].u_ce.Xin12b [8]),
    .S(gnd),
    .Y(_3560_)
);

FILL FILL_0__8214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14099_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6164_),
    .Y(_6166_)
);

OAI21X1 _13377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5401_),
    .B(_5796_),
    .C(_5814_),
    .Y(_5071_)
);

FILL FILL_2__13839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10373_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_799_),
    .C(_817_),
    .Y(_49_)
);

NAND2X1 _7445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_434_)
);

FILL FILL_2__13172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11578_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_4431_)
);

FILL FILL_0__9172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4071_),
    .B(_4070_),
    .C(_4061_),
    .Y(_3381_)
);

AOI21X1 _11023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3672_),
    .B(_3656_),
    .C(_3668_),
    .Y(_3673_)
);

FILL FILL_2__11905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7905_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5128_),
    .B(_5131_),
    .C(_5109_),
    .Y(_5132_)
);

NAND2X1 _12228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4778_),
    .B(_4779_),
    .Y(_4780_)
);

FILL FILL_1__14731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10231_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_2006_),
    .Y(_2010_)
);

FILL FILL_1__11856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8023_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10714_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2540_),
    .CLK(clk_bF$buf4),
    .Q(\genblk1[3].u_ce.Acalc [1])
);

FILL FILL_0__10429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10009_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5251_),
    .B(_5644_),
    .Y(_5645_)
);

FILL FILL_0__14682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9648_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [6]),
    .Y(_4484_)
);

FILL FILL_0__9228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8604_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_158__bF$buf0),
    .C(_652_),
    .D(_156_),
    .Y(_23_)
);

AOI21X1 _7254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_232_),
    .C(_160_),
    .Y(_252_)
);

FILL FILL_1__12394_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11672_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3412_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Yin0 [1])
);

FILL FILL_0__11387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf2),
    .B(_3811_),
    .Y(_3892_)
);

FILL FILL_2__11714_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8879_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_877_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Xin12b [8])
);

OAI21X1 _8459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1274_),
    .C(_1357_),
    .Y(_1358_)
);

OAI21X1 _8039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Xcalc [10]),
    .C(_924_),
    .Y(_957_)
);

FILL FILL_0__7714_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9820_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1732_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Yin12b [5])
);

FILL FILL_1__13599_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2190_),
    .C(_2203_),
    .Y(_2212_)
);

FILL FILL_1__13179_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5343_),
    .B(_5346_),
    .Y(_5350_)
);

NAND2X1 _12457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_4989_),
    .Y(_4991_)
);

AOI22X1 _12037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4292_),
    .B(_4348__bF$buf4),
    .C(_4597_),
    .D(_4420_),
    .Y(_4201_)
);

FILL FILL_1__14120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14318_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[0]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .Y(_6836_)
);

FILL FILL_1__11245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8672_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3586_),
    .Y(_3597_)
);

FILL FILL_0__8252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10658_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .C(_2668_),
    .Y(_3237_)
);

FILL FILL_0__10238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf2),
    .B(_2838_),
    .Y(_2839_)
);

FILL FILL257250x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9457_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [5]),
    .Y(_4303_)
);

FILL FILL_0__9037_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3525_),
    .B(_3944_),
    .C(_3945_),
    .Y(_3946_)
);

FILL FILL_1__13811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8413_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_469_),
    .C(_160_),
    .Y(_471_)
);

FILL FILL_0__11196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4023_),
    .B(_3524__bF$buf4),
    .Y(_4107_)
);

NAND3X1 _11061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .B(_3709_),
    .C(_3708_),
    .Y(_3710_)
);

FILL FILL_1__9618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11103_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1572_),
    .Y(_1573_)
);

NOR2X1 _8268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1159_),
    .Y(_1176_)
);

FILL FILL_1__10936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7103_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5149_),
    .B(_5166_),
    .Y(_5167_)
);

OR2X2 _12266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4814_),
    .B(_4813_),
    .Y(_4816_)
);

FILL FILL_0__13762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9371_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6760_),
    .Y(_7046_)
);

FILL FILL_0__14127_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .Y(_6699_)
);

FILL FILL_1__11894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10467_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10752_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2578_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Ain12b [9])
);

FILL FILL_0__10047_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3016_),
    .B(_3013_),
    .Y(_3058_)
);

DFFPOSX1 _7959_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_43_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Xin12b [4])
);

OR2X2 _7539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_521_),
    .Y(_524_)
);

OAI21X1 _7119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_121_),
    .C(_122_),
    .Y(_123_)
);

DFFPOSX1 _8900_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_898_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Yin0 [1])
);

FILL FILL_1__12679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9686_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4519_),
    .B(_4520_),
    .Y(_4521_)
);

FILL FILL_0__9266_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_4156_)
);

INVX1 _11117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_3763_)
);

FILL FILL_1__13620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14405_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_283_),
    .C(_276_),
    .Y(_288_)
);

FILL FILL_0__13818_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3866_),
    .B(_3927_),
    .C(_3928_),
    .Y(_3929_)
);

FILL FILL_1__9847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1380_),
    .C(_1363_),
    .Y(_1394_)
);

OAI21X1 _8077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_992_),
    .C(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_993_)
);

FILL FILL_1__10325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7332_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5009_),
    .B(_4997_),
    .C(_5013_),
    .Y(_4243_)
);

OAI21X1 _12075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4336_),
    .B(_4633_),
    .C(_4346_),
    .Y(_4634_)
);

FILL FILL_2__12957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8537_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Ycalc [1]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3469_)
);

FILL FILL_0__8117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6868_),
    .B(_6869_),
    .C(_6867_),
    .Y(_6870_)
);

OAI21X1 _14221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_6539_),
    .C(_6540_),
    .Y(_7071_[1])
);

FILL FILL_1__7913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486__bF$buf4),
    .B(_3543_),
    .Y(_3633_)
);

FILL FILL_0__8290_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .B(_3270_),
    .Y(_3273_)
);

FILL FILL_0__10276_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2861_),
    .B(_2874_),
    .C(_2875_),
    .Y(_2876_)
);

OAI21X1 _7768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_164_),
    .C(_134__bF$buf2),
    .Y(_739_)
);

INVX1 _7348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .Y(_342_)
);

FILL FILL_1__12488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9495_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4336_),
    .C(_4337_),
    .Y(_4338_)
);

FILL FILL_0__9075_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3979_),
    .B(_3981_),
    .Y(_3982_)
);

FILL FILL_0__12842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2658_)
);

FILL FILL_1__8451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14634_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6222_),
    .B(_6228_),
    .C(_6254_),
    .Y(_6276_)
);

FILL FILL_0__13627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x169350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8346_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_3317_),
    .C(_3320_),
    .Y(_2554_)
);

FILL FILL_1__12700_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5547_),
    .B(_5530_),
    .C(_5543_),
    .Y(_5552_)
);

FILL FILL_2__9305_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14870_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6761_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.RdyCtl [1])
);

FILL FILL_0__14585_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [9]),
    .B(_6729_),
    .Y(_6732_)
);

INVX1 _14030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6386_),
    .Y(_6389_)
);

FILL FILL_1__7722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11092_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.Acalc [1]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Acalc [3]),
    .Y(_3453_)
);

FILL FILL_0__10085_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3069_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3094_),
    .Y(_2533_)
);

FILL FILL_1__8927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8507_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _7997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_919_)
);

NAND3X1 _7577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf4),
    .B(_559_),
    .C(_556_),
    .Y(_560_)
);

INVX8 _7157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .Y(_158_)
);

FILL FILL_1__12297_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4502_),
    .B(_4556_),
    .C(_4554_),
    .Y(_4557_)
);

OAI21X1 _11575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3607_),
    .B(_4162_),
    .C(_4177_),
    .Y(_3407_)
);

NAND2X1 _11155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3799_)
);

FILL FILL_0__12651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7617_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .B(_2483_),
    .C(_2499_),
    .Y(_1729_)
);

OAI21X1 _9303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .B(_2119_),
    .C(_1832_),
    .Y(_2120_)
);

FILL FILL_1__8680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13856_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6073_),
    .B(_6068_),
    .C(_5963__bF$buf4),
    .Y(_6093_)
);

FILL FILL_0__13016_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5753_),
    .B(_5744_),
    .Y(_5754_)
);

FILL FILL_1__9885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10363_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14506_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6494_),
    .CLK(clk_bF$buf73),
    .Q(\u_ot.Xcalc [6])
);

FILL FILL_0__7790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8575_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3485_),
    .B(_3502_),
    .Y(_3504_)
);

FILL FILL_0__8155_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [10]),
    .Y(_3147_)
);

INVX1 _10006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2745_),
    .Y(_2746_)
);

FILL FILL_0__11922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14919_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf1),
    .B(_375_),
    .C(_372_),
    .Y(_378_)
);

FILL FILL_0__11099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_4014_),
    .Y(_4017_)
);

FILL FILL_2__11846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7846_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [4]),
    .Y(_2695_)
);

FILL FILL_0__7426_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2336_),
    .C(_2329_),
    .Y(_1700_)
);

NAND2X1 _9112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf4),
    .B(_1839_),
    .Y(_1937_)
);

DFFPOSX1 _12589_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4243_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Yin12b [6])
);

NAND2X1 _12169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4723_),
    .B(_4722_),
    .Y(_4724_)
);

FILL FILL_1__14672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6311_),
    .Y(_6312_)
);

FILL FILL_0__13665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(_5909_),
    .C(_5910_),
    .Y(_5911_)
);

FILL FILL_0_BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5537_),
    .B(_5558_),
    .C(_5541_),
    .Y(_5572_)
);

FILL FILL_0_BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6919_),
    .B(_6929_),
    .Y(_6956_)
);

NAND2X1 _14315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6615_),
    .B(_6614_),
    .Y(_6616_)
);

FILL FILL_2__12384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8384_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3333_),
    .B(_2597_),
    .C(_3341_),
    .Y(_2571_)
);

MUX2X1 _10235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2964_),
    .B(_2962_),
    .S(_2649__bF$buf0),
    .Y(_2965_)
);

FILL FILL_2__9763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13589_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1093_),
    .B(_1648_),
    .C(_1663_),
    .Y(_893_)
);

FILL FILL_1__7760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12936_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf2),
    .B(_5179_),
    .Y(_5277_)
);

FILL FILL_0__12516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14308_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_170_),
    .C(_195_),
    .Y(_196_)
);

NAND3X1 _11193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf1),
    .B(_3835_),
    .C(_3826_),
    .Y(_3836_)
);

FILL FILL_1__10648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10228_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf13)
);

FILL FILL_0__7655_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf12)
);

OAI21X1 _9761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2340_),
    .C(_1754_),
    .Y(_1747_)
);

FILL FILL_0__7235_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf11)
);

NAND2X1 _9341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_1916_),
    .Y(_2156_)
);

CLKBUF1 CLKBUF1_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert98 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert99 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf8)
);

NAND2X1 _12398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4937_),
    .B(_4928_),
    .Y(_4939_)
);

FILL FILL_1__14481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14679_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14544_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6532_),
    .CLK(clk_bF$buf19),
    .Q(\u_ot.Yin1 [0])
);

FILL FILL_0__14259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_5887_),
    .C(_6469_),
    .Y(_5868_)
);

FILL FILL_1__7816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11186_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .S(gnd),
    .Y(_3541_)
);

FILL FILL_0__8193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672__bF$buf1),
    .B(_3181_),
    .C(_3182_),
    .Y(_2539_)
);

NOR2X1 _10044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2777_),
    .B(_2778_),
    .Y(_2783_)
);

FILL FILL_0__11960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1500_),
    .Y(_1503_)
);

FILL FILL_0__9398_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11669_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3409_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Yin1 [0])
);

NAND2X1 _11249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3873_),
    .B(_3877_),
    .Y(_3889_)
);

FILL FILL_1__13752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12325_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12610_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .CLK(clk_bF$buf45),
    .Q(\genblk1[5].u_ce.LoadCtl [1])
);

DFFPOSX1 _9817_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1729_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Yin12b [6])
);

FILL FILL_1__8774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14117_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6179_),
    .B(_6181_),
    .C(_6182_),
    .Y(_6183_)
);

FILL FILL_1__9979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7884_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2664_),
    .B(_2701_),
    .C(_2686__bF$buf0),
    .Y(_2731_)
);

FILL FILL_0__7464_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2369_),
    .Y(_2372_)
);

AOI21X1 _9150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1934_),
    .B(_1811__bF$buf1),
    .C(_1955_),
    .Y(_1973_)
);

FILL FILL_0__10811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14488_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6991_)
);

FILL FILL_0__14068_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6647_),
    .B(_6565_),
    .C(_6648_),
    .Y(_6649_)
);

FILL FILL_1__7625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13808_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10693_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2519_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[3].u_ce.Ycalc [4])
);

INVX1 _10273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3001_),
    .Y(_3002_)
);

FILL FILL_2__10315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9381_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8841_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_839_),
    .CLK(clk_bF$buf71),
    .Q(\genblk1[1].u_ce.Ycalc [1])
);

NAND3X1 _8421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf2),
    .B(_1321_),
    .C(_1312_),
    .Y(_1322_)
);

INVX4 _8001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .Y(_923_)
);

AOI22X1 _11898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4295_),
    .B(_4348__bF$buf4),
    .C(_4464_),
    .D(_4420_),
    .Y(_4195_)
);

NAND2X1 _11478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4101_),
    .Y(_4104_)
);

NAND3X1 _11058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3700_),
    .B(_3706_),
    .C(_3703_),
    .Y(_3707_)
);

FILL FILL_1__13981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12134_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .B(_2414_),
    .Y(_2425_)
);

NAND3X1 _9206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf5),
    .B(_2026_),
    .C(_2025_),
    .Y(_2027_)
);

FILL FILL_1__8583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13759_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5999_),
    .B(_5952_),
    .S(vdd),
    .Y(_6000_)
);

FILL FILL_0__13339_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5658_),
    .B(_5656_),
    .Y(_5662_)
);

FILL FILL_0__14700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7039_),
    .B(_7043_),
    .Y(_7044_)
);

AOI21X1 _14409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .B(_6694_),
    .C(_6562__bF$buf1),
    .Y(_6697_)
);

FILL FILL_2_BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x108150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8058_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10749_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2575_),
    .CLK(clk_bF$buf25),
    .Q(\genblk1[3].u_ce.Ain12b [10])
);

OAI21X1 _10329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf1),
    .B(_3053_),
    .C(_3054_),
    .Y(_3055_)
);

FILL FILL_1__12832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14297_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [1]),
    .B(_6821_),
    .C(_6823_),
    .Y(_6824_)
);

DFFPOSX1 _14162_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5838_),
    .CLK(clk_bF$buf75),
    .Q(\genblk1[7].u_ce.Ycalc [2])
);

FILL FILL_1__7854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf2),
    .B(_2815_),
    .C(_2810_),
    .Y(_2819_)
);

FILL FILL_1__8639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10544_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .Y(_285_)
);

OAI21X1 _8650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf1),
    .B(_1537_),
    .C(_1010__bF$buf5),
    .Y(_1538_)
);

INVX1 _8230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .Y(_1139_)
);

AND2X2 _11287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3879_),
    .B(_3882_),
    .Y(_3926_)
);

FILL FILL_2__7503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7749_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .B(_2601_),
    .C(_2604_),
    .Y(_2605_)
);

FILL FILL_0__7329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2190_),
    .C(_2245_),
    .Y(_2246_)
);

NAND3X1 _9015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(gnd),
    .C(_1811__bF$buf0),
    .Y(_1844_)
);

FILL FILL_1__8392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13988_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .Y(_6219_)
);

FILL FILL_0__13568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13148_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13433_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5033_),
    .CLK(clk_bF$buf41),
    .Q(\genblk1[6].u_ce.Ycalc [4])
);

OAI21X1 _13013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5459_),
    .C(_5479_),
    .Y(_5480_)
);

FILL FILL_1__9597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10075_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6864_),
    .B(_6866_),
    .Y(_6867_)
);

OAI21X1 _14218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(_6537_),
    .C(_6538_),
    .Y(_7071_[0])
);

FILL FILL_0__7082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8041_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7921_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[0].u_ce.Ycalc [4])
);

INVX1 _7501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .Y(_488_)
);

NAND2X1 _10978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3630_)
);

FILL FILL_0__8287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3268_),
    .B(_3269_),
    .Y(_3270_)
);

AND2X2 _10138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869_),
    .B(_2872_),
    .Y(_2873_)
);

FILL FILL_1__12641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11214_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(\u_ot.Yin12b [7]),
    .C(_6680_),
    .Y(_6681_)
);

NAND2X1 _8706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1587_),
    .Y(_1590_)
);

FILL FILL_1__7663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12839_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(gnd),
    .C(_5151__bF$buf0),
    .Y(_5184_)
);

FILL FILL_0__12419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10353_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_102_),
    .C(_103_),
    .Y(_104_)
);

AOI21X1 _13909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6269_),
    .B(vdd),
    .C(_6272_),
    .Y(_6273_)
);

NAND2X1 _11096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3738_),
    .Y(_3743_)
);

FILL FILL_2__7732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x93750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7558_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _9664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_2459_),
    .D(_2458_),
    .Y(_1710_)
);

FILL FILL_0__7138_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2062_),
    .Y(_2063_)
);

FILL FILL_1__11912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13797_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6034_),
    .Y(_6037_)
);

FILL FILL_0__13377_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5180_),
    .B(_5151__bF$buf1),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5697_)
);

FILL FILL_0__9704_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [18]),
    .B(_6833__bF$buf0),
    .C(En_bF$buf3),
    .Y(_7070_)
);

NAND2X1 _14447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [8]),
    .B(_6729_),
    .Y(_6730_)
);

NAND2X1 _14027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6382_),
    .B(_6385_),
    .Y(_6386_)
);

FILL FILL_1__7719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_702_),
    .Y(_704_)
);

NAND3X1 _7310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf2),
    .B(_301_),
    .C(_296_),
    .Y(_305_)
);

FILL FILL_1__11089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [7]),
    .B(_3441_),
    .Y(_3450_)
);

FILL FILL_0__8096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3087_),
    .B(_3091_),
    .Y(_3092_)
);

FILL FILL_1__12870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11023_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [9]),
    .Y(_1770_)
);

AND2X2 _8515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1368_),
    .Y(_1412_)
);

FILL FILL_1__7892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5402_),
    .Y(_5403_)
);

FILL FILL_0__12648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12228_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf5),
    .B(_4989_),
    .C(_5022_),
    .Y(_4252_)
);

FILL FILL_1__8677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10582_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf0),
    .B(_6088_),
    .C(_6089_),
    .Y(_6090_)
);

BUFX2 BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 )
);

FILL FILL_2__7541_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf4 )
);

BUFX2 BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf3 )
);

BUFX2 BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf2 )
);

BUFX2 BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf1 )
);

BUFX2 BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf0 )
);

BUFX2 BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2648__bF$buf4)
);

FILL FILL_0__7787_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.Xcalc [0]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Xcalc [2]),
    .Y(_2639_)
);

FILL FILL_0__7367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2281_),
    .C(_2261_),
    .Y(_2282_)
);

NAND2X1 _9053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(\genblk1[1].u_ce.ISout ),
    .Y(_1881_)
);

FILL FILL_1__11721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8746_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6252_),
    .B(_6255_),
    .C(_5974_),
    .Y(_6256_)
);

FILL FILL_0__13186_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13471_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5071_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Yin12b [10])
);

NAND2X1 _13051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5257_),
    .B(_5464_),
    .Y(_5516_)
);

FILL FILL_2__13513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6898_),
    .B(_6901_),
    .Y(_6902_)
);

NAND3X1 _14256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Xin0 [0]),
    .C(\u_ot.Xin0 [1]),
    .Y(_6564_)
);

FILL FILL_1__7528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7108_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .B(_2686__bF$buf0),
    .Y(_3305_)
);

AND2X2 _10176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2903_),
    .B(_2686__bF$buf4),
    .Y(_2909_)
);

FILL FILL_2__10218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11252_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .Y(_1625_)
);

NAND2X1 _8324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1224_),
    .Y(_1229_)
);

FILL FILL_1__7281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12877_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .B(\genblk1[5].u_ce.ISout ),
    .Y(_5221_)
);

FILL FILL_0__12457_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4863_),
    .B(_4865_),
    .C(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4868_)
);

FILL FILL_0__12037_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2690_),
    .C(_2691_),
    .Y(_2692_)
);

NOR2X1 _9529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2334_),
    .B(_2333_),
    .Y(_2335_)
);

OAI21X1 _9109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1932_),
    .C(_1933_),
    .Y(_1934_)
);

FILL FILL_1__8486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6267_),
    .C(_6308_),
    .Y(_6309_)
);

FILL FILL_0_BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5908_),
    .B(_5907_),
    .Y(\genblk1[7].u_ce.Y_ [1])
);

FILL FILL_0_BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5568_),
    .B(_5569_),
    .C(_5172_),
    .Y(_5570_)
);

FILL FILL_0_BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7176_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [0]),
    .B(_1834__bF$buf0),
    .Y(_2099_)
);

FILL FILL_1__11950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10103_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5728_),
    .B(_5732_),
    .Y(_5734_)
);

FILL FILL_2__13742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11308_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6749_),
    .B(_6733_),
    .C(_6752_),
    .Y(_6529_)
);

AND2X2 _14065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6412_),
    .B(_6421_),
    .Y(_6422_)
);

FILL FILL_1__7757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9903_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(\genblk1[2].u_ce.Xcalc [9]),
    .C(_1762_),
    .Y(_1804_)
);

NAND2X1 _8553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1444_),
    .B(_1447_),
    .Y(_1448_)
);

MUX2X1 _8133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(\genblk1[1].u_ce.Xin12b [8]),
    .S(vdd),
    .Y(_1046_)
);

FILL FILL_1__7090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13273_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [0]),
    .B(_5174__bF$buf3),
    .Y(_5439_)
);

FILL FILL_0__12686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12266_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12551_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4205_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xcalc [2])
);

OAI21X1 _12131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4560_),
    .C(_4686_),
    .Y(_4687_)
);

OAI21X1 _9758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_1753_)
);

NAND2X1 _9338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf3),
    .B(_2109_),
    .Y(_2153_)
);

FILL FILL_1__8295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14058_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6123_),
    .B(_6126_),
    .Y(_6127_)
);

AOI21X1 _13336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5777_),
    .B(_5786_),
    .C(_5784_),
    .Y(_5787_)
);

FILL FILL_0__14832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .Y(_1917_)
);

FILL FILL_2__8784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .B(_172__bF$buf5),
    .Y(_791_)
);

AND2X2 _7404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_172__bF$buf1),
    .Y(_395_)
);

FILL FILL_2__13551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11537_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4392_),
    .B(_4391_),
    .C(_4350_),
    .Y(_4393_)
);

FILL FILL_0__9131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11117_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .B(_4033_),
    .Y(_4034_)
);

NAND3X1 _14294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(\u_ot.Xin12b [6]),
    .C(_6596_),
    .Y(_6597_)
);

OAI21X1 _8609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_973__bF$buf3),
    .C(_992_),
    .Y(_1500_)
);

FILL FILL_1__7566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13329_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12607_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4261_),
    .CLK(clk_bF$buf51),
    .Q(\genblk1[5].u_ce.Ain0 [0])
);

FILL FILL_2__10256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9712_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1652_)
);

NAND2X1 _8362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1264_),
    .Y(_1265_)
);

FILL FILL_1__10610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(vdd),
    .Y(_5257_)
);

FILL FILL_0__12495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12075_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4862_),
    .C(_4902_),
    .Y(_4903_)
);

FILL FILL_2__12822_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2709_),
    .B(_2684_),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_2728_)
);

NAND2X1 _9567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .B(_2369_),
    .Y(_2370_)
);

INVX1 _9147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [6]),
    .Y(_1970_)
);

FILL FILL_1__11815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14287_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6326_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6345_),
    .Y(_5853_)
);

INVX1 _13565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5943_),
    .Y(_5944_)
);

NAND2X1 _13145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5604_),
    .B(_5605_),
    .Y(_5606_)
);

FILL FILL_0__14641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10141_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_612_),
    .C(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_614_)
);

OAI22X1 _7213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_162_),
    .C(_210_),
    .D(_154_),
    .Y(_212_)
);

FILL FILL_2__13780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11346_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11631_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3371_),
    .CLK(clk_bF$buf36),
    .Q(\genblk1[4].u_ce.Xcalc [6])
);

NAND2X1 _11211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .B(_3592_),
    .Y(_3853_)
);

NAND2X1 _8838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[1] [1]),
    .Y(_917_)
);

NAND2X1 _8418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1317_),
    .B(_1318_),
    .Y(_1319_)
);

FILL FILL_1__7795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13138_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [6]),
    .Y(_5310_)
);

INVX1 _12416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4954_),
    .Y(_4955_)
);

FILL FILL_0__13912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9101_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(_1478_),
    .Y(_1484_)
);

INVX1 _8171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .Y(_1083_)
);

FILL FILL_2__12631_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9796_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1708_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[2].u_ce.Acalc [7])
);

AOI22X1 _9376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1834__bF$buf3),
    .C(_2189_),
    .D(_1832_),
    .Y(_1692_)
);

FILL FILL_1__11204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8631_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(_3556_),
    .C(_3557_),
    .Y(_3354_)
);

FILL FILL_0__8211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14096_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6162_),
    .Y(_6163_)
);

FILL FILL_0__13089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.X_ [1]),
    .Y(_5813_)
);

FILL FILL257550x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(_6815_),
    .C(_6820_),
    .Y(_6821_)
);

DFFPOSX1 _14159_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5835_),
    .CLK(clk_bF$buf49),
    .Q(\genblk1[7].u_ce.Ycalc [0])
);

FILL FILL_0__10790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10370_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(gnd),
    .Y(_816_)
);

NAND3X1 _7442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf4),
    .B(_427_),
    .C(_430_),
    .Y(_431_)
);

OAI21X1 _10499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_3215_)
);

OAI21X1 _10079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2796_),
    .B(_2791_),
    .C(_2686__bF$buf2),
    .Y(_2816_)
);

FILL FILL_1__12162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11575_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf1),
    .B(_4379_),
    .Y(_4428_)
);

FILL FILL_0__11155_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4048_),
    .B(_4056_),
    .C(_4055_),
    .Y(_4069_)
);

NAND3X1 _11020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .B(_3641_),
    .C(_3669_),
    .Y(_3670_)
);

INVX1 _8647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .Y(_1535_)
);

NAND2X1 _8227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf3),
    .B(_1047_),
    .Y(_1136_)
);

FILL FILL_1__7184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13367_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [5]),
    .Y(_5129_)
);

NAND3X1 _12225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf2),
    .B(_4776_),
    .C(_4773_),
    .Y(_4777_)
);

FILL FILL_0__13721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2005_),
    .B(_2006_),
    .Y(_2007_)
);

FILL FILL_1__11853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8038_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10711_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2537_),
    .CLK(clk_bF$buf21),
    .Q(\genblk1[3].u_ce.Xcalc [10])
);

FILL FILL_0__10426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10006_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5640_),
    .B(_5639_),
    .Y(_5642_)
);

DFFPOSX1 _7918_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf9),
    .Q(\genblk1[0].u_ce.ISout )
);

FILL FILL_1__12638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9645_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4480_),
    .B(_4465_),
    .C(_4417_),
    .Y(_4482_)
);

FILL FILL_0__9225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6675_),
    .C(_6678_),
    .Y(_6679_)
);

FILL FILL_1__8601_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_649_),
    .Y(_650_)
);

AOI21X1 _7251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_244_),
    .C(_233_),
    .Y(_249_)
);

FILL FILL_1__12391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11384_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8876_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_874_),
    .CLK(clk_bF$buf68),
    .Q(\genblk1[1].u_ce.Acalc [11])
);

NAND2X1 _8456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1354_),
    .Y(_1355_)
);

AOI22X1 _8036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.Ycalc [1]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_955_)
);

FILL FILL_0__7711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13176_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5345_),
    .B(_5346_),
    .Y(_5347_)
);

FILL FILL_0__12169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4987_),
    .B(_4988_),
    .Y(_4989_)
);

OAI21X1 _12034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4594_),
    .B(_4537_),
    .C(_4590_),
    .Y(_4595_)
);

FILL FILL_0__13950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11909_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf2),
    .B(_6030_),
    .C(_6033_),
    .Y(_6034_)
);

OAI21X1 _13239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5692_),
    .B(_5694_),
    .C(_5681_),
    .Y(_5053_)
);

FILL FILL_0__14735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14315_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(En_bF$buf3),
    .B(_6804_),
    .Y(_6765_)
);

FILL FILL_2__7482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3534_),
    .B(_3593_),
    .C(_3592_),
    .D(_3530_),
    .Y(_3594_)
);

FILL FILL_2__8267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10655_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3231_),
    .C(_3228_),
    .Y(_3234_)
);

FILL FILL_0__10235_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2836_)
);

OAI21X1 _7727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_701_)
);

OAI21X1 _7307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_277_),
    .C(_172__bF$buf2),
    .Y(_302_)
);

FILL FILL_2__13034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9454_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [9]),
    .Y(_4300_)
);

FILL FILL_0__9034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(_3939_),
    .C(_3942_),
    .Y(_3943_)
);

DFFPOSX1 _14197_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5873_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Yin12b [11])
);

FILL FILL_0__12801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8410_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _7480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_467_),
    .Y(_468_)
);

FILL FILL_0__11193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11520_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _8685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .C(_1568_),
    .D(_1570_),
    .Y(_868_)
);

NAND3X1 _8265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(_1171_),
    .C(_1172_),
    .Y(_1173_)
);

FILL FILL_1__10933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7520_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_134__bF$buf3)
);

FILL FILL_0__7100_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_134__bF$buf2)
);

BUFX2 BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_134__bF$buf1)
);

BUFX2 BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_134__bF$buf0)
);

BUFX2 BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf5)
);

BUFX2 BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf4)
);

BUFX2 BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf3)
);

BUFX2 BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf2)
);

BUFX2 BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf1)
);

OAI21X1 _12683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5162_),
    .C(_5163_),
    .Y(_5164_)
);

FILL FILL_0__12398_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_172__bF$buf0)
);

INVX1 _12263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4812_),
    .Y(_4813_)
);

FILL FILL257250x165750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8305_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6248_),
    .B(_6245_),
    .S(_5926__bF$buf1),
    .Y(_6253_)
);

DFFPOSX1 _13468_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5068_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Xin1 [1])
);

OAI21X1 _13048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5386_),
    .C(_5512_),
    .Y(_5513_)
);

FILL FILL_0__14124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10044_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7956_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_40_),
    .CLK(clk_bF$buf15),
    .Q(\genblk1[0].u_ce.Xin12b [9])
);

INVX1 _7536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .Y(_521_)
);

AOI21X1 _7116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_118_),
    .C(_119_),
    .Y(_120_)
);

FILL FILL_1__12676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9683_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4517_),
    .C(_4513_),
    .Y(_4518_)
);

FILL FILL_0__9263_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3676_),
    .B(_4151_),
    .C(_4153_),
    .Y(_3390_)
);

FILL FILL_0__11249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [11]),
    .B(_3510__bF$buf1),
    .Y(_3760_)
);

FILL FILL_1__7698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14468_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5218_),
    .B(_5217_),
    .C(_5176_),
    .Y(_5219_)
);

AND2X2 _12319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4864_),
    .B(_4862_),
    .Y(_4865_)
);

FILL FILL_1__14822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9004_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1390_),
    .B(_1391_),
    .C(_994_),
    .Y(_1392_)
);

NAND2X1 _8074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_988_),
    .Y(_990_)
);

FILL FILL_1__10322_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_5012_)
);

NAND2X1 _12072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4623_),
    .Y(_4631_)
);

FILL FILL_2__12534_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_2486_)
);

OAI21X1 _9279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2093_),
    .B(_2096_),
    .C(_1903_),
    .Y(_2097_)
);

FILL FILL_1__11947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8534_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [7]),
    .B(_3441_),
    .Y(_3466_)
);

FILL FILL_0__8114_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6069_),
    .Y(_6070_)
);

OR2X2 _13277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5730_),
    .B(_5188__bF$buf0),
    .Y(_5731_)
);

FILL FILL_2__13739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10273_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_728_),
    .C(_726_),
    .Y(_736_)
);

OAI21X1 _7345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_312_),
    .C(_307_),
    .Y(_339_)
);

FILL FILL_2__13072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11478_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4333_),
    .C(_4334_),
    .Y(_4335_)
);

FILL FILL_0__9072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11058_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(_3977_),
    .C(_3978_),
    .Y(_3979_)
);

FILL FILL_2__11805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2653_),
    .C(_2654_),
    .Y(_2655_)
);

OAI21X1 _12968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5433_),
    .B(_5436_),
    .C(_5243_),
    .Y(_5437_)
);

DFFPOSX1 _12548_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4202_),
    .CLK(clk_bF$buf5),
    .Q(\genblk1[5].u_ce.Ycalc [11])
);

OAI21X1 _12128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4679_),
    .B(_4663_),
    .C(_4677_),
    .Y(_4684_)
);

FILL FILL_1__14631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811__bF$buf4),
    .B(_1865_),
    .Y(_1914_)
);

FILL FILL_1__11756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8343_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3316_),
    .B(_3317_),
    .C(_3318_),
    .Y(_2553_)
);

FILL FILL_0__10329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .B(_5548_),
    .Y(_5550_)
);

FILL FILL_2__9722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9548_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4388_),
    .B(_4389_),
    .Y(_4390_)
);

FILL FILL_0__9128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8504_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7994_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl [4]),
    .CLK(clk_bF$buf27),
    .Q(\genblk1[0].u_ce.LoadCtl [5])
);

AOI21X1 _7574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf2),
    .B(_516_),
    .C(_538_),
    .Y(_557_)
);

INVX2 _7154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .Y(_156_)
);

FILL FILL257550x144150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12294_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4553_),
    .B(_4525_),
    .Y(_4554_)
);

FILL FILL_0__11287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(_4159_),
    .Y(_4176_)
);

OAI21X1 _11152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3791_),
    .C(_3775_),
    .Y(_3365_)
);

FILL FILL_1__9709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1648_),
    .C(_1650_),
    .Y(_882_)
);

INVX1 _8359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1262_)
);

FILL FILL_1__10607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7614_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2498_)
);

NAND2X1 _9300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2109_),
    .Y(_2117_)
);

FILL FILL_1__13079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf2),
    .B(_5205_),
    .Y(_5254_)
);

INVX1 _12357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [4]),
    .Y(_4900_)
);

FILL FILL_1__14860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14638_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14503_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6491_),
    .CLK(clk_bF$buf46),
    .Q(\u_ot.Xcalc [3])
);

FILL FILL_0__14218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8572_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3500_),
    .B(_3497_),
    .S(_3487__bF$buf3),
    .Y(_3501_)
);

FILL FILL_0__8152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10138_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3135_),
    .B(_3144_),
    .Y(_3145_)
);

INVX1 _10003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2743_)
);

FILL FILL_2__9531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9357_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11628_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3368_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xcalc [3])
);

MUX2X1 _11208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3849_),
    .B(_3806_),
    .S(gnd),
    .Y(_3850_)
);

FILL FILL_1__13711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14916_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .Y(_375_)
);

FILL FILL_0__13909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11096_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3487__bF$buf4),
    .C(_3506_),
    .Y(_4014_)
);

FILL FILL_1__9938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11003_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(_1480_),
    .Y(_1481_)
);

AOI22X1 _8168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1020_),
    .B(_1079_),
    .C(_1078_),
    .D(_1016_),
    .Y(_1080_)
);

FILL FILL_1__10836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7423_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12586_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4240_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Yin12b [11])
);

NAND2X1 _12166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4717_),
    .B(_4720_),
    .Y(_4721_)
);

FILL FILL_0__13662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14447_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [11]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf1),
    .Y(_6954_)
);

FILL FILL_0__14027_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6583_),
    .B(_6612_),
    .C(\u_ot.ISreg_bF$buf4 ),
    .Y(_6613_)
);

FILL FILL_1__11794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8381_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3324_),
    .Y(_3340_)
);

FILL FILL_0__10367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2747_),
    .C(_2961_),
    .Y(_2962_)
);

FILL FILL_2__9760_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_83_),
    .C(_814_),
    .Y(_46_)
);

NOR2X1 _7439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_428_)
);

FILL FILL_1__12999_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(_1645_),
    .Y(_1662_)
);

FILL FILL_1__12159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9586_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .Y(_4425_)
);

FILL FILL_0__9166_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4065_),
    .B(_4062_),
    .Y(_4066_)
);

INVX1 _11017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ycalc [7]),
    .Y(_3667_)
);

FILL FILL_1__13940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14305_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(\genblk1[0].u_ce.Xin0 [1]),
    .S(gnd),
    .Y(_193_)
);

FILL FILL_0__13718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3831_),
    .B(_3832_),
    .Y(_3833_)
);

FILL FILL_1__9747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11232_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf5),
    .B(_1298_),
    .C(_1276_),
    .Y(_1299_)
);

FILL FILL_1__10645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10225_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf43)
);

FILL FILL_0__7652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7232_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf38)
);

NAND2X1 _12395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4934_),
    .B(_4935_),
    .Y(_4936_)
);

FILL FILL_2__12857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8017_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10708_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2534_),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.Xcalc [7])
);

FILL FILL_1__9080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14676_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14541_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6529_),
    .CLK(clk_bF$buf47),
    .Q(\u_ot.Yin12b [7])
);

FILL FILL_0__14256_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [1]),
    .B(_6466_),
    .Y(_6468_)
);

FILL FILL_1__7813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11183_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3537_),
    .B(_3534_),
    .S(_3487__bF$buf3),
    .Y(_3538_)
);

FILL FILL_0__8190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10596_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3178_),
    .B(_3179_),
    .Y(_3180_)
);

FILL FILL_0__10176_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2748_),
    .Y(_2780_)
);

NOR2X1 _7668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_642_),
    .Y(_647_)
);

INVX1 _7248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .Y(_246_)
);

FILL FILL_1__12388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9395_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11666_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3406_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Yin12b [7])
);

AOI22X1 _11246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3510__bF$buf4),
    .C(_3886_),
    .D(_3508_),
    .Y(_3369_)
);

FILL FILL_0__12742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7708_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9814_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1726_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Yin12b [11])
);

FILL FILL_1__8771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13947_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6166_),
    .B(_6178_),
    .C(_6162_),
    .Y(_6180_)
);

FILL FILL_0__13527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8666_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf1),
    .B(_3589_),
    .C(_3590_),
    .Y(_3591_)
);

FILL FILL_0__8246_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3231_),
    .B(_3230_),
    .Y(_3232_)
);

FILL FILL_2__9205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14485_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6988_)
);

FILL FILL_0__14065_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .C(\u_ot.ISreg_bF$buf2 ),
    .Y(_6646_)
);

FILL FILL_1__7622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13805_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10690_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2516_),
    .CLK(clk_bF$buf38),
    .Q(\genblk1[3].u_ce.ISout )
);

AOI21X1 _10270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2945_),
    .B(_2951_),
    .C(_2977_),
    .Y(_2999_)
);

FILL FILL_1__8827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8407_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [1]),
    .Y(_835_)
);

AOI21X1 _7477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_464_),
    .C(_183_),
    .Y(_465_)
);

FILL FILL_1__12197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4461_),
    .B(_4458_),
    .Y(_4462_)
);

NAND2X1 _11475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4101_),
    .Y(_4102_)
);

NOR2X1 _11055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .B(_3675_),
    .Y(_3704_)
);

FILL FILL256950x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7517_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .B(_2421_),
    .Y(_2422_)
);

INVX1 _9203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2024_)
);

FILL FILL_1__8580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ycalc [2]),
    .B(_5949__bF$buf2),
    .Y(_5997_)
);

NAND2X1 _13201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5656_),
    .B(_5658_),
    .Y(_5659_)
);

FILL FILL_1__9365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7033_),
    .Y(_7041_)
);

INVX1 _14406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [9]),
    .Y(_6694_)
);

FILL FILL_0__7690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8055_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10746_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2572_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin1 [1])
);

NOR2X1 _10326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf1),
    .B(_2925_),
    .Y(_3052_)
);

FILL FILL_2__9854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert221 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert223 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert224 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf3),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

NAND2X1 _11284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .B(_3922_),
    .Y(_3923_)
);

FILL FILL_0__12780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7746_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _9852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_2602_)
);

FILL FILL_0__7326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2242_),
    .B(_2241_),
    .Y(_2243_)
);

NAND2X1 _9012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(_1840_),
    .Y(_1841_)
);

OAI21X1 _12489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_5010_)
);

AND2X2 _12069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4621_),
    .B(_4627_),
    .Y(_4628_)
);

FILL FILL_2__8705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13985_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6216_)
);

FILL FILL_0__13565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13145_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13430_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5030_),
    .CLK(clk_bF$buf47),
    .Q(\genblk1[6].u_ce.ISout )
);

NAND3X1 _13010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf3),
    .B(_5476_),
    .C(_5454_),
    .Y(_5477_)
);

FILL FILL_1__9594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10072_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .B(_6851_),
    .C(_6859_),
    .Y(_6864_)
);

DFFPOSX1 _14215_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.Vld )
);

FILL FILL_1__7907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11277_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3624_),
    .B(_3606_),
    .C(_3623_),
    .Y(_3627_)
);

FILL FILL_0__8284_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .Y(_3267_)
);

NAND3X1 _10135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf4),
    .B(_2867_),
    .C(_2863_),
    .Y(_2870_)
);

FILL FILL_2__9243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1587_),
    .Y(_1588_)
);

FILL FILL_1__7660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12836_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(_5180_),
    .Y(_5181_)
);

FILL FILL_0__12416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2650_),
    .C(_2651_),
    .Y(_2652_)
);

FILL FILL_1__8445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14628_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_100_),
    .Y(\a[1] [1])
);

NAND2X1 _13906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(_6217_),
    .Y(_6270_)
);

AOI21X1 _11093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3723_),
    .B(_3727_),
    .C(_3739_),
    .Y(_3740_)
);

FILL FILL_1__10968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7555_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2455_),
    .Y(_2457_)
);

FILL FILL_0__7135_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2060_),
    .Y(_1686_)
);

NAND2X1 _12298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf5),
    .B(_4833_),
    .Y(_4846_)
);

FILL FILL_0__10902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14579_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [17]),
    .B(_6833__bF$buf0),
    .C(En_bF$buf2),
    .Y(_7068_)
);

INVX1 _14444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.X_ [0]),
    .Y(_6727_)
);

NAND3X1 _14024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf5),
    .B(_6379_),
    .C(_6374_),
    .Y(_6383_)
);

FILL FILL_1__7716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11086_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [11]),
    .C(_3438_),
    .Y(_3447_)
);

FILL FILL_0__8093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3064_),
    .B(_3088_),
    .C(_3063_),
    .Y(_3089_)
);

FILL FILL_0__11860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1768_)
);

NAND2X1 _8512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1408_),
    .Y(_1409_)
);

OAI21X1 _11989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4537_),
    .B(_4550_),
    .C(_4551_),
    .Y(_4552_)
);

FILL FILL_0__9298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(_4155_),
    .C(_4174_),
    .Y(_3404_)
);

NAND2X1 _11149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3792_),
    .B(_3793_),
    .Y(_3794_)
);

FILL FILL_1__13652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13232_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5126_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5400_),
    .Y(_5038_)
);

FILL FILL_0__12645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[5] [0]),
    .B(_4989_),
    .Y(_5021_)
);

OAI21X1 _9717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2496_)
);

FILL FILL_1__8674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14017_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6054_),
    .B(_6076_),
    .C(_6057_),
    .Y(_6087_)
);

FILL FILL_1__9879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7784_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [6]),
    .B(_2603_),
    .Y(_2636_)
);

FILL FILL_0__7364_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2279_)
);

AOI21X1 _9050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1877_),
    .C(_1836_),
    .Y(_1879_)
);

FILL FILL_0__13183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14388_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6899_)
);

INVX8 _14253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .Y(_6562_)
);

FILL FILL_1__7525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x108150 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3288_),
    .B(_3301_),
    .C(_3299_),
    .Y(_3302_)
);

OAI21X1 _10173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2902_),
    .B(_2904_),
    .C(_2905_),
    .Y(_2906_)
);

FILL FILL_2__10635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9281_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Acalc [10]),
    .B(_996__bF$buf2),
    .Y(_1622_)
);

AOI21X1 _8321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1209_),
    .B(_1213_),
    .C(_1225_),
    .Y(_1226_)
);

MUX2X1 _11798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4368_),
    .B(_4365_),
    .S(_4325__bF$buf4),
    .Y(_4369_)
);

AND2X2 _11378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(_4011_),
    .Y(_4012_)
);

FILL FILL_1__13881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x201750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12034_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2687_),
    .C(_2688_),
    .Y(_2689_)
);

NAND2X1 _9526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf2),
    .B(_2319_),
    .Y(_2332_)
);

INVX1 _9106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_1931_)
);

FILL FILL_1__8483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13659_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [11]),
    .Y(_6306_)
);

FILL FILL_0_BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13239_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(_5904_),
    .C(_5905_),
    .Y(_5906_)
);

FILL FILL_0_BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5565_),
    .Y(_5567_)
);

FILL FILL_0_BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10166_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6950_),
    .Y(_6951_)
);

INVX1 _14309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [8]),
    .Y(_6610_)
);

FILL FILL_0__7593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3335_),
    .B(_3321_),
    .C(_3338_),
    .Y(_2568_)
);

NAND2X1 _10229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [1]),
    .B(_2672__bF$buf4),
    .Y(_2959_)
);

FILL FILL_1__12732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11305_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [6]),
    .B(_6733_),
    .Y(_6751_)
);

NAND2X1 _14062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6416_),
    .B(_6417_),
    .Y(_6419_)
);

FILL FILL_1__7754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9900_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .S(gnd),
    .Y(_190_)
);

NAND2X1 _8970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1801_),
    .B(_1800_),
    .Y(\genblk1[2].u_ce.X_ [0])
);

INVX1 _8550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1444_),
    .Y(_1445_)
);

OAI21X1 _8130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .B(_1042_),
    .C(_1043_),
    .Y(_840_)
);

OAI21X1 _11187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487__bF$buf0),
    .B(_3828_),
    .C(_3829_),
    .Y(_3830_)
);

FILL FILL_2__7403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7649_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2486_),
    .C(_1751_),
    .Y(_1744_)
);

FILL FILL_0__7229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2119_),
    .B(_2136_),
    .Y(_2150_)
);

FILL FILL_1__8292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13888_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf1),
    .B(_6120_),
    .C(_6114_),
    .Y(_6124_)
);

FILL FILL_0__13048_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5781_),
    .B(_5769_),
    .C(_5780_),
    .Y(_5784_)
);

FILL FILL_1__9497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10395_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14538_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6526_),
    .CLK(clk_bF$buf51),
    .Q(\u_ot.Yin12b [8])
);

AND2X2 _14118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .B(\genblk1[7].u_ce.LoadCtl [2]),
    .Y(_6466_)
);

AOI21X1 _7821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_787_),
    .C(_785_),
    .Y(_788_)
);

OAI21X1 _7401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .B(_390_),
    .C(_391_),
    .Y(_392_)
);

INVX1 _10878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .Y(_3535_)
);

FILL FILL_0__8187_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_3176_),
    .C(\genblk1[3].u_ce.Ain0 [0]),
    .Y(_3177_)
);

INVX2 _10038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2776_),
    .Y(_2777_)
);

FILL FILL_1__12961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11114_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6590_),
    .B(_6562__bF$buf0),
    .C(_6594_),
    .D(_6592_),
    .Y(_6493_)
);

AND2X2 _8606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1493_),
    .B(_1497_),
    .Y(_1498_)
);

FILL FILL_1__7563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12739_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12604_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4258_),
    .CLK(clk_bF$buf51),
    .Q(\genblk1[5].u_ce.Ain12b [5])
);

FILL FILL_0__12319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10253_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6088_),
    .C(_6117_),
    .Y(_6177_)
);

FILL FILL_2__7632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7878_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_2648__bF$buf3),
    .Y(_2725_)
);

FILL FILL_0__7458_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2366_),
    .Y(_2367_)
);

OAI21X1 _9144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1966_),
    .B(_1951_),
    .C(_1903_),
    .Y(_1968_)
);

FILL FILL_1__11812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6342_),
    .B(_6327_),
    .Y(_6343_)
);

FILL FILL_0__13697_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5940_),
    .B(_5933_),
    .S(_5925__bF$buf1),
    .Y(_5941_)
);

FILL FILL_0__13277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf2),
    .B(_5602_),
    .C(_5599_),
    .Y(_5603_)
);

FILL FILL_0__9604_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6985_),
    .B(_6984_),
    .Y(_6986_)
);

NAND2X1 _14347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6632_),
    .B(_6644_),
    .Y(_6499_)
);

FILL FILL_1__7619_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_610_),
    .B(_608_),
    .C(_603_),
    .Y(_611_)
);

MUX2X1 _7210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_161_),
    .S(gnd),
    .Y(_209_)
);

OAI21X1 _10687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3197_),
    .C(_2593_),
    .Y(_2586_)
);

AOI21X1 _10267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .B(gnd),
    .C(_2995_),
    .Y(_2996_)
);

FILL FILL_1__12770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11343_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_921_),
    .C(_915_),
    .Y(_908_)
);

OAI21X1 _8415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf2),
    .B(_1314_),
    .C(_1315_),
    .Y(_1316_)
);

FILL FILL_1__7792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12968_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5306_),
    .B(_5291_),
    .C(_5243_),
    .Y(_5308_)
);

AOI22X1 _12413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4941_),
    .B(_4348__bF$buf3),
    .C(_4951_),
    .D(_4952_),
    .Y(_4222_)
);

FILL FILL_0__12128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10482_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.ISout ),
    .Y(_5995_)
);

FILL FILL_2__7861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7687_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9793_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1705_),
    .CLK(clk_bF$buf37),
    .Q(\genblk1[2].u_ce.Acalc [4])
);

FILL FILL_2_BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7267_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _9373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2186_),
    .B(_2171_),
    .Y(_2187_)
);

FILL FILL_2_BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14093_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6158_),
    .B(_6146_),
    .C(_6159_),
    .Y(_6160_)
);

FILL FILL_0__13086_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5802_),
    .B(_5104_),
    .C(_5811_),
    .Y(_5068_)
);

FILL FILL_2__13413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9413_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [7]),
    .Y(_6818_)
);

OAI21X1 _14156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5962_),
    .C(_6486_),
    .Y(_5883_)
);

FILL FILL_1__7848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert190 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert192 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert193 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert195 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert197 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert199 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_3212_)
);

OAI21X1 _10076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf2),
    .B(_2811_),
    .C(_2812_),
    .Y(_2813_)
);

FILL FILL_2__10958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11152_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _8644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .C(_1530_),
    .D(_1532_),
    .Y(_865_)
);

INVX1 _8224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1133_)
);

FILL FILL_1__7181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12777_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [9]),
    .Y(_5126_)
);

FILL FILL_0__12357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf4),
    .B(_4601_),
    .Y(_4774_)
);

INVX4 _9849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .Y(_2599_)
);

NAND2X1 _9429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2236_),
    .B(_2239_),
    .Y(_2240_)
);

MUX2X1 _9009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .B(\genblk1[2].u_ce.Xin12b [4]),
    .S(gnd),
    .Y(_1838_)
);

FILL FILL257550x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6199_),
    .B(_6213_),
    .Y(_5847_)
);

OAI21X1 _13427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5695_),
    .C(_5101_),
    .Y(_5094_)
);

NAND2X1 _13007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151__bF$buf3),
    .B(_5473_),
    .Y(_5474_)
);

FILL FILL_2__7670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf4),
    .B(_2003_),
    .C(_1999_),
    .Y(_2004_)
);

FILL FILL_1__11850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10003_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5638_),
    .Y(_5639_)
);

OAI21X1 _7915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_683_),
    .C(_79_),
    .Y(_72_)
);

FILL FILL_2__13642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9642_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4478_),
    .Y(_4479_)
);

FILL FILL_0__9222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11208_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [6]),
    .Y(_6676_)
);

FILL FILL_1__7657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11381_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8873_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_871_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Acalc [8])
);

AOI21X1 _8453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1332_),
    .B(_1347_),
    .C(_1345_),
    .Y(_1352_)
);

NAND2X1 _8033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [7]),
    .B(_927_),
    .Y(_952_)
);

FILL FILL_1__13593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13173_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf5),
    .B(_5343_),
    .C(_5339_),
    .Y(_5344_)
);

FILL FILL_0__12166_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348__bF$buf3),
    .B(_4986_),
    .C(_4985_),
    .Y(_4226_)
);

AOI21X1 _12031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4591_),
    .B(_4590_),
    .C(_4588_),
    .Y(_4592_)
);

AOI21X1 _9658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2450_),
    .B(_2445_),
    .C(_2443_),
    .Y(_2454_)
);

AND2X2 _9238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2045_),
    .B(_2057_),
    .Y(_2058_)
);

FILL FILL_1__8195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5926__bF$buf4),
    .Y(_6031_)
);

NOR2X1 _13236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5682_),
    .B(_5691_),
    .Y(_5692_)
);

FILL FILL_0__14732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10232_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_698_)
);

OAI21X1 _7304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf3),
    .B(_297_),
    .C(_298_),
    .Y(_299_)
);

FILL FILL_2__13031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11437_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4294_),
    .B(_4297_),
    .C(_4282_),
    .Y(_4298_)
);

FILL FILL_0__9031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11017_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .Y(_3940_)
);

DFFPOSX1 _14194_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5870_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin0 [0])
);

AND2X2 _8929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1764_),
    .B(\genblk1[2].u_ce.LoadCtl [3]),
    .Y(_1765_)
);

AOI21X1 _8509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1366_),
    .B(_1367_),
    .C(_977_),
    .Y(_1406_)
);

FILL FILL_1__7886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13229_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5385_),
    .B(_5397_),
    .Y(_5398_)
);

OAI21X1 _12507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4323_),
    .C(_5019_),
    .Y(_4249_)
);

FILL FILL_2__10996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9612_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1558_),
    .Y(_1568_)
);

NAND3X1 _8262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1160_),
    .B(_1166_),
    .C(_1169_),
    .Y(_1170_)
);

FILL FILL_1__10930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10510_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .Y(_3510__bF$buf2)
);

BUFX2 BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .Y(_3510__bF$buf1)
);

FILL FILL_2__7115_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .Y(_3510__bF$buf0)
);

BUFX2 BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .Y(_3486__bF$buf4)
);

BUFX2 BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .Y(_3486__bF$buf3)
);

OAI21X1 _12680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5159_),
    .C(_5160_),
    .Y(_5161_)
);

FILL FILL_0__12395_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4807_),
    .B(_4792_),
    .Y(_4810_)
);

FILL FILL_2__12722_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Xcalc [10]),
    .C(_2600_),
    .Y(_2633_)
);

OAI21X1 _9467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2241_),
    .B(_2271_),
    .C(_2267_),
    .Y(_2276_)
);

AND2X2 _9047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1874_),
    .B(_1875_),
    .Y(_1876_)
);

FILL FILL_1__11715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8302_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926__bF$buf1),
    .B(_6246_),
    .C(_6249_),
    .Y(_6250_)
);

DFFPOSX1 _13465_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5065_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[6].u_ce.Xin12b [4])
);

OAI21X1 _13045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .B(_5489_),
    .C(_5503_),
    .Y(_5510_)
);

FILL FILL_2__13927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10041_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7953_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .CLK(clk_bF$buf31),
    .Q(\genblk1[0].u_ce.Xin12b [10])
);

OAI21X1 _7533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_476_),
    .C(_517_),
    .Y(_518_)
);

NAND2X1 _7113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_116_),
    .Y(\genblk1[0].u_ce.Y_ [1])
);

FILL FILL_2__13680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9680_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324__bF$buf1),
    .B(_4514_),
    .Y(_4515_)
);

FILL FILL_0__9260_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4151_),
    .Y(_4152_)
);

FILL FILL_0__11246_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3755_),
    .B(_3757_),
    .C(_3579_),
    .Y(_3758_)
);

AND2X2 _8738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(_1619_),
    .Y(_1620_)
);

INVX1 _8318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .Y(_1223_)
);

FILL FILL_1__7695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13038_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5214_),
    .B(_5215_),
    .Y(_5216_)
);

AOI21X1 _12316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4619_),
    .B(vdd),
    .C(_4861_),
    .Y(_4862_)
);

FILL FILL_0__13812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9001_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1387_),
    .Y(_1389_)
);

MUX2X1 _8071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_983_),
    .S(_973__bF$buf3),
    .Y(_987_)
);

OAI21X1 _9696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2483_),
    .C(_2484_),
    .Y(_1717_)
);

INVX1 _9276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2093_),
    .Y(_2094_)
);

FILL FILL_1__11944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8531_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Ycalc [11]),
    .C(_3438_),
    .Y(_3463_)
);

FILL FILL_0__8111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8129_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [5]),
    .Y(_6067_)
);

INVX1 _13274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [5]),
    .Y(_5728_)
);

FILL FILL_0__14770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9316_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14899_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6790_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.Atmp [3])
);

INVX1 _14479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Y_ [1]),
    .Y(_6749_)
);

NAND2X1 _14059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6414_),
    .B(_6415_),
    .Y(_6416_)
);

FILL FILL_0__10270_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [6]),
    .B(_158__bF$buf4),
    .Y(_733_)
);

NAND2X1 _7342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_335_),
    .Y(_336_)
);

NAND3X1 _10399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686__bF$buf5),
    .B(_3121_),
    .C(_3118_),
    .Y(_3122_)
);

FILL FILL_1__12482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11475_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4331_),
    .B(_4328_),
    .S(_4325__bF$buf4),
    .Y(_4332_)
);

FILL FILL_0__11055_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .B(_3956_),
    .C(_3524__bF$buf5),
    .Y(_3976_)
);

OAI21X1 _8967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1764_),
    .B(_1797_),
    .C(_1798_),
    .Y(_1799_)
);

NAND3X1 _8547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .B(_1426_),
    .C(_1399_),
    .Y(_1442_)
);

OAI21X1 _8127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996__bF$buf0),
    .B(_1041_),
    .C(_997_),
    .Y(_839_)
);

FILL FILL_1__7084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13267_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5433_),
    .Y(_5434_)
);

DFFPOSX1 _12545_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4199_),
    .CLK(clk_bF$buf53),
    .Q(\genblk1[5].u_ce.Ycalc [8])
);

NOR2X1 _12125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4663_),
    .B(_4680_),
    .Y(_4682_)
);

FILL FILL_0__13621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7399_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .Y(_1911_)
);

FILL FILL_1__11753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8340_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.X_ [0]),
    .Y(_3316_)
);

FILL FILL_0__10326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5543_),
    .B(_5546_),
    .Y(_5547_)
);

OAI21X1 _7818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_766_),
    .C(_780_),
    .Y(_785_)
);

FILL FILL_1__12958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9545_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4386_),
    .B(_4378_),
    .C(_4361_),
    .Y(_4387_)
);

FILL FILL_0__9125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [5]),
    .B(_6591_),
    .Y(_6592_)
);

FILL FILL_1__8921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8501_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7991_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[0].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf78),
    .Q(\genblk1[0].u_ce.LoadCtl [2])
);

OAI21X1 _7571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_554_),
    .Y(_18_)
);

INVX1 _7151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .Y(_153_)
);

FILL FILL_1__12291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11611_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1648_),
    .Y(_1649_)
);

OAI21X1 _8356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_1259_),
    .C(_1068_),
    .Y(_1260_)
);

FILL FILL_1__10604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13076_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .Y(_5251_)
);

FILL FILL_0__12489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12069_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4887_),
    .B(_4896_),
    .C(_4897_),
    .Y(_4898_)
);

FILL FILL_0__13850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8816_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6339_),
    .Y(_6340_)
);

NAND2X1 _13559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .B(vdd),
    .Y(_5938_)
);

NOR2X1 _13139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf4),
    .B(_5427_),
    .Y(_5600_)
);

FILL FILL_0__14635_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl_6_bF$buf1 ),
    .Y(Vld)
);

DFFPOSX1 _14500_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6488_),
    .CLK(clk_bF$buf9),
    .Q(\u_ot.Xcalc [0])
);

FILL FILL_2__7382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x165750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10975_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .Y(_3498_)
);

FILL FILL_2__8167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10555_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3139_),
    .B(_3140_),
    .Y(_3142_)
);

FILL FILL_0__10135_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2674_),
    .Y(_2741_)
);

NAND3X1 _7627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf0),
    .B(_607_),
    .C(_604_),
    .Y(_608_)
);

NAND2X1 _7207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ycalc [2]),
    .B(_158__bF$buf2),
    .Y(_206_)
);

FILL FILL_1__12767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9354_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11625_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3365_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xcalc [0])
);

INVX1 _11205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3846_),
    .Y(_3847_)
);

OAI21X1 _14097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6450_),
    .B(_6446_),
    .C(_5947_),
    .Y(_6452_)
);

FILL FILL_0__12701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14913_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .Y(_372_)
);

FILL FILL_0__13906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11420_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .Y(_1478_)
);

OAI21X1 _8165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf1),
    .B(_1075_),
    .C(_1076_),
    .Y(_1077_)
);

FILL FILL_1__10833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7420_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12583_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4237_),
    .CLK(clk_bF$buf6),
    .Q(\genblk1[5].u_ce.Xin0 [0])
);

FILL FILL_0__12298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _12163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4713_),
    .B(_4710_),
    .Y(_4718_)
);

FILL FILL_2__12205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8205_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6123_),
    .B(_6126_),
    .C(_6156_),
    .Y(_6157_)
);

OAI21X1 _13368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5810_)
);

FILL FILL_0__14864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10364_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_813_)
);

NAND2X1 _7436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_425_)
);

FILL FILL_1__12996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11569_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4421_),
    .Y(_4422_)
);

FILL FILL_0__9163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(vdd),
    .C(_3524__bF$buf4),
    .Y(_4063_)
);

AOI21X1 _11014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3664_),
    .B(_3660_),
    .C(_3512_),
    .Y(_3665_)
);

FILL FILL_0__12930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5120_),
    .B(_5123_),
    .C(_5109_),
    .Y(_5124_)
);

INVX1 _12219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [7]),
    .Y(_4771_)
);

FILL FILL_1__14722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x241350 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf1),
    .B(_1295_),
    .Y(_1296_)
);

FILL FILL_1__10642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10222_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf75)
);

CLKBUF1 CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf73)
);

FILL FILL_2__7667_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf68)
);

NAND2X1 _12392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4932_),
    .B(_4931_),
    .Y(_4933_)
);

FILL FILL256950x208950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12434_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(vdd),
    .C(_1830_),
    .Y(_2399_)
);

NOR2X1 _9179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf3),
    .B(_2000_),
    .Y(_2001_)
);

FILL FILL_1__11847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8014_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10705_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2531_),
    .CLK(clk_bF$buf66),
    .Q(\genblk1[3].u_ce.Xcalc [4])
);

NAND2X1 _13597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_5975_)
);

NOR2X1 _13177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5633_),
    .B(_5618_),
    .Y(_5636_)
);

FILL FILL_2__13639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10920_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_640_),
    .Y(_644_)
);

OAI21X1 _7245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134__bF$buf4),
    .B(_239_),
    .C(_242_),
    .Y(_243_)
);

FILL FILL_1__12385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9392_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11663_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3403_),
    .CLK(clk_bF$buf22),
    .Q(\genblk1[4].u_ce.Yin12b [8])
);

FILL FILL_0__11378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3866_),
    .B(_3883_),
    .Y(_3884_)
);

FILL FILL_2__11705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7705_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9811_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1723_),
    .CLK(clk_bF$buf1),
    .Q(\genblk1[2].u_ce.Xin0 [0])
);

NOR2X1 _12868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf4),
    .B(_5340_),
    .Y(_5341_)
);

OAI21X1 _12448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4984_),
    .B(_4983_),
    .C(_4974_),
    .Y(_4225_)
);

AOI21X1 _12028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4564_),
    .B(_4566_),
    .C(_4560_),
    .Y(_4589_)
);

FILL FILL_1__14111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8663_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3588_)
);

FILL FILL_0__8243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10649_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3224_),
    .B(_3227_),
    .Y(_3229_)
);

FILL FILL_0__10229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9448_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [4]),
    .Y(_4295_)
);

FILL FILL_0__9028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8404_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [0]),
    .Y(_833_)
);

MUX2X1 _7474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_454_),
    .S(_135__bF$buf1),
    .Y(_462_)
);

FILL FILL_1__12194_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4453_),
    .B(_4454_),
    .Y(_4459_)
);

FILL FILL_0__11187_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4098_),
    .Y(_4099_)
);

OR2X2 _11052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .B(_3679_),
    .Y(_3701_)
);

FILL FILL_1__9609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11934_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1559_),
    .B(_1563_),
    .Y(_1565_)
);

INVX1 _8259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .Y(_1167_)
);

FILL FILL_1__10927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7514_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2418_),
    .B(_2417_),
    .Y(_2419_)
);

FILL FILL_1__13399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1983_),
    .B(_2012_),
    .C(_2011_),
    .Y(_2021_)
);

MUX2X1 _12677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5157_),
    .B(_5154_),
    .S(_5151__bF$buf0),
    .Y(_5158_)
);

OAI21X1 _12257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4807_),
    .B(_4792_),
    .C(_4346_),
    .Y(_4808_)
);

FILL FILL_1__14760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10260_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7037_),
    .B(_7036_),
    .Y(_7038_)
);

FILL FILL_0__14118_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6691_),
    .B(_6690_),
    .Y(_6692_)
);

FILL FILL_2__12472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10458_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10743_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2569_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin12b [4])
);

FILL FILL_0__10038_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [5]),
    .Y(_3049_)
);

FILL FILL_2__9431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9677_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4512_)
);

FILL FILL_0__9257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [5]),
    .B(_3437_),
    .Y(_4149_)
);

AND2X2 _11108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3749_),
    .B(_3745_),
    .Y(_3755_)
);

FILL FILL_1__13611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14816_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .Y(_279_)
);

FILL FILL_0__13809_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3880_),
    .B(_3881_),
    .C(_3491_),
    .Y(_3920_)
);

FILL FILL_1__9418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11743_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(_1385_),
    .C(_1014_),
    .Y(_1386_)
);

INVX1 _8068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .Y(_984_)
);

FILL FILL_1__10316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7323_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_4989_),
    .Y(_5008_)
);

OAI21X1 _12066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4445_),
    .C(_4624_),
    .Y(_4625_)
);

FILL FILL_2__12948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14347_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6857_),
    .B(_6858_),
    .C(_6861_),
    .Y(_6862_)
);

DFFPOSX1 _14212_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[7].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf23),
    .Q(\genblk1[7].u_ce.LoadCtl [3])
);

FILL FILL_1__7904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11274_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(_3624_),
    .C(_3512_),
    .Y(_3625_)
);

FILL FILL_0__8281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10687_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3262_),
    .B(_3264_),
    .C(_3247_),
    .Y(_2545_)
);

FILL FILL_0__10267_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2864_),
    .Y(_2867_)
);

FILL FILL_2__9660_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_720_),
    .Y(_731_)
);

NAND3X1 _7339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf2),
    .B(_329_),
    .C(_323_),
    .Y(_333_)
);

FILL FILL_1__12899_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .Y(_1585_)
);

FILL FILL256950x176550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9486_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .Y(_4329_)
);

FILL FILL_0__9066_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3972_),
    .Y(_3973_)
);

FILL FILL_1__13840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12413_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _9905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_2649_)
);

FILL FILL_1__8442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14625_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_97_),
    .C(_98_),
    .Y(_99_)
);

OAI21X1 _13903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [8]),
    .C(_6266_),
    .Y(_6267_)
);

FILL FILL_0__13618_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .Y(_3737_)
);

FILL FILL_1__9647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11132_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1145_),
    .Y(_1203_)
);

FILL FILL_1__10965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7132_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [11]),
    .B(_4348__bF$buf2),
    .Y(_4843_)
);

FILL FILL_2__8931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2770_),
    .B(_3313_),
    .C(_3314_),
    .Y(_2551_)
);

AOI21X1 _14861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6818_),
    .B(_6833__bF$buf3),
    .C(_7066_),
    .Y(_6794_)
);

FILL FILL_0__14576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14156_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6628_),
    .B(_6724_),
    .C(_6725_),
    .Y(_6512_)
);

OAI21X1 _14021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6353_),
    .B(_6347_),
    .C(_5963__bF$buf5),
    .Y(_6380_)
);

FILL FILL_1__7713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11083_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.Acalc [0]),
    .C(_3443_),
    .D(_3444_),
    .Y(_3445_)
);

FILL FILL_0__8090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3081_),
    .B(_3085_),
    .Y(_3086_)
);

FILL FILL_2__10403_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7988_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_72_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Ain0 [1])
);

NOR2X1 _7568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_536_),
    .Y(_552_)
);

MUX2X1 _7148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_142_),
    .S(_134__bF$buf2),
    .Y(_150_)
);

FILL FILL_1__12288_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4545_),
    .B(_4548_),
    .Y(_4549_)
);

FILL FILL_0__9295_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4171_),
    .B(_4155_),
    .C(_4172_),
    .Y(_3403_)
);

NOR2X1 _11146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .B(_3790_),
    .Y(_3791_)
);

FILL FILL_2__11608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7608_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2475_),
    .Y(_2494_)
);

FILL FILL_1__8671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13427_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5904_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6084_),
    .Y(_5841_)
);

FILL FILL_0__13007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10354_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[7]),
    .Y(Dout[7])
);

FILL FILL_0__7781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8566_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3495_)
);

FILL FILL_0__8146_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3137_),
    .B(_3138_),
    .Y(_3139_)
);

FILL FILL_1__12920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14385_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [6]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf1),
    .Y(_6897_)
);

NAND2X1 _14250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [11]),
    .Y(_6560_)
);

FILL FILL_1__7522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13705_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3295_),
    .B(_3280_),
    .C(_3294_),
    .Y(_3299_)
);

NAND3X1 _10170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2889_),
    .B(_2901_),
    .C(_2885_),
    .Y(_2903_)
);

FILL FILL_1__8727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10632_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [8]),
    .B(_701_),
    .C(_765_),
    .Y(_766_)
);

AOI21X1 _7377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_355_),
    .C(_368_),
    .Y(_369_)
);

FILL FILL_1__12097_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4366_)
);

NOR2X1 _11375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .B(_4008_),
    .Y(_4009_)
);

FILL FILL_0__12871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7837_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _9943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_2686_)
);

FILL FILL_0__7417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [11]),
    .B(_1834__bF$buf4),
    .Y(_2329_)
);

OAI21X1 _9103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1908_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_)
);

FILL FILL_1__8480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6303_),
    .B(_6302_),
    .Y(_6304_)
);

FILL FILL_0__13656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13236_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(_5901_),
    .C(_5902_),
    .Y(_5903_)
);

FILL FILL_0_BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5559_),
    .B(_5563_),
    .C(_5192_),
    .Y(_5564_)
);

FILL FILL_0_BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10163_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6948_)
);

NAND3X1 _14306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6606_),
    .B(_6607_),
    .C(_6599_),
    .Y(_6608_)
);

FILL FILL_0__7590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8375_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .B(_3321_),
    .Y(_3337_)
);

OAI21X1 _10226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf0),
    .B(_2956_),
    .C(_2945_),
    .Y(_2957_)
);

FILL FILL_0__11722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14719_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _7186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_179_),
    .S(_134__bF$buf1),
    .Y(_187_)
);

NAND2X1 _11184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3722_),
    .Y(_3827_)
);

FILL FILL_2__7820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7646_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[2] [0]),
    .B(_2486_),
    .Y(_1750_)
);

FILL FILL_0__7226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834__bF$buf0),
    .B(_2147_),
    .C(_2121_),
    .Y(_1690_)
);

NOR2X1 _12389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4889_),
    .Y(_4930_)
);

FILL FILL_2__8605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13885_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6090_),
    .B(_6087_),
    .C(_5963__bF$buf1),
    .Y(_6121_)
);

FILL FILL_0__13045_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5778_),
    .B(_5781_),
    .Y(_5782_)
);

FILL FILL_1__9494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10392_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14535_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6523_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin0 [1])
);

OAI21X1 _14115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_6463_),
    .C(_6464_),
    .Y(_5864_)
);

FILL FILL_1__7807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11177_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3532_)
);

FILL FILL_0__8184_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3173_),
    .B(_3169_),
    .C(_2670_),
    .Y(_3175_)
);

OAI21X1 _10035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf3),
    .B(_2772_),
    .C(_2773_),
    .Y(_2774_)
);

FILL FILL_2__10917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(_1494_),
    .Y(_1495_)
);

FILL FILL_1__7560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12316_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12601_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4255_),
    .CLK(clk_bF$buf30),
    .Q(\genblk1[5].u_ce.Ain12b [6])
);

DFFPOSX1 _9808_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1720_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin12b [5])
);

FILL FILL_1__8765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14108_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6174_),
    .B(_6173_),
    .C(_6021_),
    .Y(_6175_)
);

FILL FILL_1__10868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7875_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(\genblk1[3].u_ce.Xin12b [8]),
    .S(vdd),
    .Y(_2722_)
);

FILL FILL_0__7455_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain1 [0]),
    .B(_2363_),
    .Y(_2364_)
);

INVX1 _9141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1964_),
    .Y(_1965_)
);

NOR3X1 _12198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4710_),
    .B(_4731_),
    .C(_4735_),
    .Y(_4751_)
);

FILL FILL_2__8834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14479_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6981_),
    .B(_6982_),
    .Y(_6983_)
);

FILL FILL_0__14059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6641_),
    .B(_6639_),
    .C(_6613_),
    .Y(_6642_)
);

FILL FILL_1__7616_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[3] [0]),
    .Y(_2592_)
);

FILL FILL_0__10399_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2755_),
    .B(_2940_),
    .Y(_2993_)
);

FILL FILL_0__11760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13198_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_914_)
);

NAND2X1 _8412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_1208_),
    .Y(_1313_)
);

NOR2X1 _11889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .B(_4424_),
    .Y(_4456_)
);

FILL FILL_0__9198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [6]),
    .B(_4095_),
    .Y(_4096_)
);

NOR2X1 _11049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3660_),
    .B(_3688_),
    .Y(_3698_)
);

FILL FILL_1__13972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12965_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5304_),
    .Y(_5305_)
);

FILL FILL_0__12125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4949_),
    .B(_4948_),
    .Y(_4950_)
);

FILL FILL256950x108150 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2375_),
    .Y(_2416_)
);

FILL FILL_1__8994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5991_),
    .B(_5943_),
    .Y(_5993_)
);

FILL FILL_1__9359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x201750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9790_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1702_),
    .CLK(clk_bF$buf24),
    .Q(\genblk1[2].u_ce.Acalc [1])
);

FILL FILL_0__7264_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2183_),
    .Y(_2184_)
);

FILL FILL_2_BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.Atmp [5]),
    .Y(_6815_)
);

NAND2X1 _14153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6485_)
);

FILL FILL_1__7845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert161 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert162 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert164 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert166 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert168 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert169 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [3]),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .Y(_3209_)
);

NAND3X1 _10073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2777_),
    .B(_2799_),
    .C(_2780_),
    .Y(_2810_)
);

FILL FILL_2__10955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9181_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _8641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_1522_),
    .Y(_1530_)
);

OAI21X1 _8221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1130_),
    .B(_1129_),
    .C(_1068_),
    .Y(_1131_)
);

NOR2X1 _11698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.LoadCtl [3]),
    .Y(_4276_)
);

NAND2X1 _11278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(_3916_),
    .Y(_3917_)
);

FILL FILL_1__13781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12354_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2595_),
    .Y(_2596_)
);

NOR3X1 _9426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .B(_2217_),
    .C(_2221_),
    .Y(_2237_)
);

NAND2X1 _9006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [1]),
    .B(_1834__bF$buf0),
    .Y(_1835_)
);

FILL FILL_1__8383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13559_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6196_),
    .B(_6194_),
    .C(_6200_),
    .Y(_6211_)
);

FILL FILL_0__13139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\a[6] [0]),
    .Y(_5100_)
);

INVX1 _13004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5471_)
);

FILL FILL_0__14920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10066_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6858_),
    .B(_6857_),
    .Y(_6859_)
);

DFFPOSX1 _14209_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .CLK(clk_bF$buf65),
    .Q(\genblk1[7].u_ce.LoadCtl [0])
);

FILL FILL_0__7493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12698_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[0] [0]),
    .Y(_78_)
);

FILL FILL_0__8698_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3616_),
    .B(_3615_),
    .Y(_3622_)
);

FILL FILL_0__8278_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .B(_3252_),
    .Y(_3262_)
);

OAI21X1 _10129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2774_),
    .C(_2840_),
    .Y(_2864_)
);

FILL FILL_1__12632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4474_),
    .C(_4475_),
    .Y(_4476_)
);

FILL FILL_0__11205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Yin12b [4]),
    .B(\u_ot.Yin12b [5]),
    .Y(_6673_)
);

FILL FILL_1__7654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10344_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_94_),
    .C(_95_),
    .Y(_96_)
);

DFFPOSX1 _8870_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_868_),
    .CLK(clk_bF$buf46),
    .Q(\genblk1[1].u_ce.Acalc [5])
);

NAND2X1 _8450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1333_),
    .B(_1348_),
    .Y(_1350_)
);

OAI21X1 _8030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Ycalc [11]),
    .C(_924_),
    .Y(_949_)
);

OAI21X1 _11087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3733_),
    .B(_3721_),
    .C(_3579_),
    .Y(_3735_)
);

FILL FILL_2__7303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7549_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2450_),
    .Y(_2452_)
);

FILL FILL_0__7129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2047_),
    .C(_2049_),
    .Y(_2055_)
);

FILL FILL_1__8192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13788_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6026_),
    .C(_6027_),
    .Y(_6028_)
);

FILL FILL_0__13368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5688_),
    .B(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5689_)
);

FILL FILL_1__9397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10295_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [14]),
    .B(_6833__bF$buf3),
    .C(En_bF$buf4),
    .Y(_7065_)
);

NOR2X1 _14438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [3]),
    .B(_6722_),
    .Y(_6723_)
);

OAI21X1 _14018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6289_),
    .C(_6376_),
    .Y(_6377_)
);

NOR2X1 _7721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [3]),
    .B(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .Y(_695_)
);

NAND3X1 _7301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_285_),
    .C(_266_),
    .Y(_296_)
);

AOI22X1 _10778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.Acalc [4]),
    .C(_3441_),
    .D(\genblk1[4].u_ce.Acalc [6]),
    .Y(_3442_)
);

FILL FILL_0__8087_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3082_),
    .B(_3062_),
    .Y(_3083_)
);

FILL FILL_1__12861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11014_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14191_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5867_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin12b [5])
);

NOR2X1 _8926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.LoadCtl [3]),
    .Y(_1762_)
);

NAND2X1 _8506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(_1402_),
    .Y(_1403_)
);

FILL FILL_1__7883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12639_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5387_),
    .C(_5389_),
    .Y(_5395_)
);

FILL FILL_0__12219_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_5018_)
);

FILL FILL_1__8668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10153_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6066_),
    .B(_6081_),
    .Y(_6082_)
);

BUFX2 BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1811__bF$buf3)
);

FILL FILL_2__7532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7112_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert211 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1811__bF$buf2)
);

BUFX2 BUFX2_insert212 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1811__bF$buf1)
);

BUFX2 BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1811__bF$buf0)
);

BUFX2 BUFX2_insert214 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert216 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert217 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf1 )
);

FILL FILL_2__11358_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf0 )
);

FILL FILL_0__12392_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert219 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .Y(_2672__bF$buf4)
);

FILL FILL_0__7778_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _9884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[3].u_ce.Ycalc [1]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2631_)
);

FILL FILL_0__7358_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .Y(_2274_)
);

AOI21X1 _9044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_1864_),
    .C(_1847_),
    .Y(_1873_)
);

FILL FILL_1__11712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13597_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [6]),
    .Y(_6247_)
);

FILL FILL_0__13177_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13462_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5062_),
    .CLK(clk_bF$buf52),
    .Q(\genblk1[6].u_ce.Xin12b [9])
);

NOR2X1 _13042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489_),
    .B(_5506_),
    .Y(_5508_)
);

FILL FILL257250x79350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9504_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6890_),
    .Y(_6894_)
);

NAND2X1 _14247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(\u_ot.Xcalc [10]),
    .Y(_6558_)
);

FILL FILL_1__7519_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7950_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Acalc [9])
);

NAND2X1 _7530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_515_)
);

OAI21X1 _7110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_113_),
    .C(_114_),
    .Y(_115_)
);

OAI21X1 _10587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3295_),
    .B(_3292_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_3297_)
);

OAI21X1 _10167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2811_),
    .C(_2840_),
    .Y(_2900_)
);

FILL FILL_1__12670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11243_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010__bF$buf5),
    .B(\genblk1[1].u_ce.Ain12b [9]),
    .Y(_1617_)
);

OAI21X1 _8315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .B(_1207_),
    .C(_1065_),
    .Y(_1221_)
);

FILL FILL_1__7692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12868_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5212_),
    .B(_5204_),
    .C(_5187_),
    .Y(_5213_)
);

FILL FILL_0__12448_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [1]),
    .B(_4348__bF$buf1),
    .Y(_4859_)
);

FILL FILL_0__12028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10382_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .B(_6299_),
    .Y(_6301_)
);

NAND2X1 _13518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5900_),
    .B(_5899_),
    .Y(\genblk1[7].u_ce.Y_ [0])
);

FILL FILL_2__7341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7587_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .B(_2479_),
    .C(_2482_),
    .Y(_1716_)
);

FILL FILL_0__7167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2090_),
    .B(_2066_),
    .Y(_2091_)
);

FILL FILL_1__11941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6063_),
    .C(_6064_),
    .Y(_6065_)
);

NAND2X1 _13271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5724_),
    .B(_5723_),
    .Y(_5725_)
);

FILL FILL_2__13313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9313_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14896_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6787_),
    .CLK(clk_bF$buf34),
    .Q(\u_pa.Atmp [0])
);

INVX1 _14476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Y_ [0]),
    .Y(_6747_)
);

OAI21X1 _14056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6330_),
    .C(_6376_),
    .Y(_6413_)
);

FILL FILL_1__7748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7328_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3119_)
);

FILL FILL_2__10858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11052_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _8964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1794_),
    .C(_1795_),
    .Y(_1796_)
);

NOR2X1 _8544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1433_),
    .Y(_1439_)
);

OAI21X1 _8124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .B(_1008_),
    .C(_1038_),
    .Y(_1039_)
);

FILL FILL_1__7081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13264_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5430_),
    .B(_5406_),
    .Y(_5431_)
);

FILL FILL_0__12677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12257_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12542_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4196_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ycalc [5])
);

AOI21X1 _12122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4674_),
    .B(_4676_),
    .C(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4679_)
);

OAI21X1 _9749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_2483_),
    .C(_2513_),
    .Y(_1741_)
);

NAND2X1 _9329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2144_),
    .Y(_2145_)
);

FILL FILL_1__8286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_6030_),
    .C(_6117_),
    .Y(_6118_)
);

OR2X2 _13327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf4),
    .B(\genblk1[6].u_ce.Ain12b [9]),
    .Y(_5779_)
);

FILL FILL_0__14823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7396_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .Y(_1908_)
);

FILL FILL_1__11750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10323_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _13080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .B(_5536_),
    .Y(_5544_)
);

OAI21X1 _7815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_778_),
    .C(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .Y(_783_)
);

FILL FILL_2__13122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11528_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4383_),
    .B(_4382_),
    .S(_4325__bF$buf4),
    .Y(_4384_)
);

FILL FILL_0__9122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11108_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf0),
    .B(_6588_),
    .C(_6589_),
    .Y(_6492_)
);

FILL FILL_1__7557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(_1645_),
    .Y(_1647_)
);

NOR3X1 _8353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1256_),
    .C(_1240_),
    .Y(_1257_)
);

FILL FILL_1__10601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13073_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5247_),
    .Y(_5248_)
);

FILL FILL_0__12486_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4894_),
    .Y(_4895_)
);

FILL FILL_0__12066_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_2718_),
    .C(_2719_),
    .Y(_2516_)
);

OAI21X1 _9558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .B(_1811__bF$buf0),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_2361_)
);

OAI21X1 _9138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1960_),
    .C(_1961_),
    .Y(_1962_)
);

FILL FILL_1__8095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14278_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6311_),
    .B(_6336_),
    .C(_5963__bF$buf2),
    .Y(_6337_)
);

NAND2X1 _13556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_5935_)
);

INVX1 _13136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [7]),
    .Y(_5597_)
);

FILL FILL_0__14632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10132_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .Y(_605_)
);

INVX1 _7204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.ISout ),
    .Y(_204_)
);

FILL FILL_2__13351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9369_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11622_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3362_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[4].u_ce.Ycalc [9])
);

FILL FILL_0__11337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3844_),
    .B(_3843_),
    .C(_3579_),
    .Y(_3845_)
);

AOI21X1 _14094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6434_),
    .B(_5963__bF$buf0),
    .C(_6205_),
    .Y(_6449_)
);

OAI21X1 _8829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1548_),
    .B(_1648_),
    .C(_912_),
    .Y(_905_)
);

NAND2X1 _8409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xcalc [2]),
    .B(_996__bF$buf1),
    .Y(_1310_)
);

FILL FILL_1__7786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5300_),
    .C(_5301_),
    .Y(_5302_)
);

NOR2X1 _12407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4943_),
    .B(_4946_),
    .Y(_4947_)
);

FILL FILL_1__14910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1465_),
    .B(_1467_),
    .C(_1474_),
    .Y(_1475_)
);

NAND2X1 _8162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1074_)
);

FILL FILL_1__10830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10410_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12580_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4234_),
    .CLK(clk_bF$buf33),
    .Q(\genblk1[5].u_ce.Xin12b [5])
);

FILL FILL_0__12295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4693_),
    .B(_4712_),
    .Y(_4715_)
);

DFFPOSX1 _9787_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1699_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Xcalc [10])
);

OR2X2 _9367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2180_),
    .B(_2179_),
    .Y(_2181_)
);

FILL FILL_0__8622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14087_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .B(_6123_),
    .Y(_6154_)
);

OAI21X1 _13365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5155_),
    .B(_5807_),
    .C(_5808_),
    .Y(_5065_)
);

FILL FILL_2__13827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10361_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_810_),
    .C(_811_),
    .Y(_43_)
);

NAND2X1 _7433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_422_),
    .Y(_12_)
);

FILL FILL_2__13580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11566_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4419_)
);

FILL FILL_0__9160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11146_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4047_),
    .B(_4060_),
    .Y(_3380_)
);

NOR2X1 _11011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3661_),
    .B(_3640_),
    .Y(_3662_)
);

OR2X2 _8638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_1527_)
);

NAND2X1 _8218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1127_),
    .Y(_1128_)
);

FILL FILL_1__7595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13358_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [4]),
    .Y(_5121_)
);

OAI21X1 _12216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4768_),
    .B(_4762_),
    .C(_4417_),
    .Y(_4769_)
);

FILL FILL_0__13712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9321_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1292_),
    .Y(_1293_)
);

FILL FILL_0__14917_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2393_),
    .C(_2390_),
    .Y(_2396_)
);

INVX1 _9176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_1998_)
);

FILL FILL_1__11844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8011_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10702_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2528_),
    .CLK(clk_bF$buf8),
    .Q(\genblk1[3].u_ce.Xcalc [1])
);

FILL FILL_0__10417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Xin12b [4]),
    .Y(_5972_)
);

OAI21X1 _13174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5633_),
    .B(_5618_),
    .C(_5172_),
    .Y(_5634_)
);

OAI21X1 _7909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_83_),
    .C(_76_),
    .Y(_69_)
);

FILL FILL_0__14670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9636_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf0),
    .B(_4472_),
    .C(_4467_),
    .Y(_4473_)
);

FILL FILL_0__9216_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7014_),
    .B(_6886_),
    .C(_6913_),
    .Y(_7016_)
);

OR2X2 _14379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6670_),
    .B(_6669_),
    .Y(_6671_)
);

FILL FILL_0__10590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10170_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_606_),
    .Y(_641_)
);

NOR2X1 _7242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_135__bF$buf1),
    .Y(_240_)
);

NAND2X1 _10299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3026_),
    .B(_3025_),
    .Y(_3027_)
);

FILL FILL_1__12382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11375_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11660_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3400_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin0 [1])
);

OAI21X1 _11240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3877_),
    .C(_3872_),
    .Y(_3881_)
);

DFFPOSX1 _8867_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_865_),
    .CLK(clk_bF$buf55),
    .Q(\genblk1[1].u_ce.Acalc [2])
);

NAND3X1 _8447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1018_),
    .B(_1344_),
    .C(_1343_),
    .Y(_1347_)
);

AOI22X1 _8027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.Ycalc [0]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Ycalc [2]),
    .Y(_947_)
);

FILL FILL_0__7702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13167_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5338_)
);

NAND2X1 _12445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4980_),
    .B(_4981_),
    .Y(_4982_)
);

NAND2X1 _12025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4584_),
    .B(_4585_),
    .Y(_4586_)
);

FILL FILL_2__12907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8660_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3585_)
);

FILL FILL_0__8240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10646_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2943_),
    .C(_3225_),
    .Y(_3226_)
);

FILL FILL_0__10226_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_684_),
    .Y(_693_)
);

FILL FILL_1__12858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ycalc [10]),
    .Y(_4292_)
);

FILL FILL_0__9025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14188_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5864_),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[7].u_ce.Xin12b [6])
);

FILL FILL_1__8821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8401_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .B(_799_),
    .C(_831_),
    .Y(_61_)
);

OAI21X1 _7471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135__bF$buf1),
    .B(_455_),
    .C(_458_),
    .Y(_459_)
);

FILL FILL_1__12191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11511_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _8676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(_1010__bF$buf4),
    .Y(_1562_)
);

INVX1 _8256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1163_),
    .Y(_1164_)
);

FILL FILL_1__10924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10504_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert180 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .Y(_2649__bF$buf0)
);

FILL FILL_2__7529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7511_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert181 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf4 )
);

FILL FILL_1__13396_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert183 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert185 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert186 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_158__bF$buf4)
);

BUFX2 BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_158__bF$buf3)
);

BUFX2 BUFX2_insert188 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_158__bF$buf2)
);

INVX1 _12674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .Y(_5155_)
);

FILL FILL_0__12389_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_158__bF$buf1)
);

OAI21X1 _12254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4804_),
    .C(_4792_),
    .Y(_4805_)
);

FILL FILL_0__13750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8716_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6244_)
);

DFFPOSX1 _13459_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5059_),
    .CLK(clk_bF$buf56),
    .Q(\genblk1[6].u_ce.Xin12b [10])
);

AOI21X1 _13039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .B(_5502_),
    .C(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5505_)
);

INVX1 _14820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[18]),
    .Y(_7035_)
);

FILL FILL_0__14115_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6663_),
    .B(_6688_),
    .C(\u_ot.ISreg_bF$buf1 ),
    .Y(_6689_)
);

FILL FILL256650x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8067_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10740_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2566_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Yin12b [9])
);

FILL FILL_0__10455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3045_),
    .B(_3028_),
    .Y(_3047_)
);

DFFPOSX1 _7947_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Acalc [6])
);

NAND2X1 _7527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_511_),
    .Y(_513_)
);

AOI21X1 _7107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_110_),
    .C(_111_),
    .Y(_112_)
);

FILL FILL_1__12667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9674_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4499_),
    .B(_4477_),
    .C(_4478_),
    .Y(_4509_)
);

FILL FILL_0__9254_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Acalc [11]),
    .B(_3510__bF$buf2),
    .Y(_4147_)
);

AOI21X1 _11105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3720_),
    .B(_3729_),
    .C(_3751_),
    .Y(_3752_)
);

FILL FILL_1__7689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14813_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_276_)
);

FILL FILL_0__13806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11320_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _8485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1320_),
    .B(_1382_),
    .C(_1323_),
    .Y(_1383_)
);

INVX1 _8065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_981_)
);

FILL FILL_1__10313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12198_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4373_),
    .C(_5006_),
    .Y(_4238_)
);

NAND2X1 _12063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4622_)
);

FILL FILL_2__12525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8105_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6060_),
    .B(_6061_),
    .C(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6062_)
);

OAI21X1 _13268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5684_),
    .C(_5721_),
    .Y(_5722_)
);

FILL FILL_0__14764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10264_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(_726_),
    .Y(_728_)
);

OAI21X1 _7336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_296_),
    .C(_172__bF$buf2),
    .Y(_330_)
);

FILL FILL_1__12896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11469_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_4326_)
);

FILL FILL_0__9063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _11334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3470_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_3970_),
    .D(_3968_),
    .Y(_3373_)
);

FILL FILL_0__12830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14268_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [0]),
    .Y(_2646_)
);

NAND2X1 _12959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .B(_5427_),
    .Y(_5428_)
);

DFFPOSX1 _12539_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4193_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ycalc [2])
);

OAI21X1 _12119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4675_),
    .C(_4672_),
    .Y(_4676_)
);

FILL FILL_1__14622_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6237_),
    .B(_6258_),
    .C(_6256_),
    .Y(_6264_)
);

FILL FILL_0__13615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9224_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _8294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1182_),
    .B(_996__bF$buf4),
    .C(_1200_),
    .D(_1180_),
    .Y(_847_)
);

FILL FILL_1__10962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x151350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4839_),
    .B(_4828_),
    .Y(_4841_)
);

FILL FILL_2__12334_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2297_),
    .B(_2306_),
    .Y(_2307_)
);

INVX1 _9079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1905_)
);

FILL FILL_1__11747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x118950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2600_),
    .B(_2606_),
    .Y(_3312_)
);

DFFPOSX1 _13497_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[6].u_ce.LoadCtl [1]),
    .CLK(clk_bF$buf29),
    .Q(\genblk1[6].u_ce.LoadCtl [2])
);

NOR2X1 _13077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5519_),
    .B(_5538_),
    .Y(_5541_)
);

FILL FILL_2__9713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10073_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7985_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_69_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Ain1 [0])
);

INVX1 _7565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .Y(_549_)
);

NAND2X1 _7145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(gnd),
    .Y(_147_)
);

FILL FILL_1__12285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11698_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4543_),
    .C(_4539_),
    .Y(_4546_)
);

FILL FILL_0__9292_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_4151_),
    .C(_4170_),
    .Y(_3402_)
);

FILL FILL_0__11278_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3787_),
    .B(_3785_),
    .S(_3487__bF$buf0),
    .Y(_3788_)
);

FILL FILL_2__14497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7605_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1859_),
    .C(_2492_),
    .Y(_1724_)
);

INVX1 _12768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5245_)
);

OAI21X1 _12348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4354_),
    .B(_4891_),
    .C(_4890_),
    .Y(_4892_)
);

FILL FILL_1__14851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10351_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[4]),
    .Y(Dout[4])
);

FILL FILL_0__14629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8563_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3492_)
);

FILL FILL_0__8143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3053_),
    .C(_3099_),
    .Y(_3136_)
);

FILL FILL_0__11910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9348_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11619_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3359_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[4].u_ce.Ycalc [6])
);

FILL FILL_1__13702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256350x201750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Acalc [8]),
    .B(_158__bF$buf3),
    .Y(_763_)
);

NAND3X1 _7374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_335_),
    .C(_365_),
    .Y(_366_)
);

FILL FILL256950x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12094_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4363_)
);

FILL FILL_0__11087_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3997_),
    .Y(_4006_)
);

FILL FILL_1__9929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11834_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1828_),
    .Y(_1829_)
);

INVX1 _8579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1465_),
    .Y(_1472_)
);

INVX1 _8159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1071_)
);

FILL FILL_1__10827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7834_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648__bF$buf4),
    .B(_2682_),
    .C(_2681_),
    .Y(_2683_)
);

FILL FILL_0__7414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2314_),
    .Y(_2327_)
);

FILL FILL_1__13299_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .Y(_1926_)
);

OAI21X1 _12997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_5249_),
    .C(_5463_),
    .Y(_5464_)
);

DFFPOSX1 _12577_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4231_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Xin12b [6])
);

NAND3X1 _12157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .B(_4633_),
    .C(_4650_),
    .Y(_4712_)
);

FILL FILL_1__14660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert200 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert202 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert204 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert205 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert207 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert209 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14438_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6944_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(_6945_),
    .Y(_6777_)
);

FILL FILL_0__14018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(\u_ot.Xin12b [7]),
    .C(_6604_),
    .Y(_6605_)
);

FILL FILL_2__12372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8372_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [1]),
    .Y(_3335_)
);

FILL FILL_0__10358_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649__bF$buf0),
    .B(_2949_),
    .Y(_2954_)
);

FILL FILL_2__9751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9577_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4350_),
    .Y(_4417_)
);

FILL FILL_0__9157_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4055_),
    .B(_4057_),
    .Y(_4058_)
);

NAND3X1 _11008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .B(_3657_),
    .C(_3658_),
    .Y(_3659_)
);

FILL FILL_1__13931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x104550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x183750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14716_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_184_)
);

FILL FILL_0__13709_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Xcalc [2]),
    .B(_3510__bF$buf3),
    .Y(_3824_)
);

FILL FILL_1__9738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9318_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972__bF$buf0),
    .B(_1289_),
    .Y(_1290_)
);

FILL FILL_1__10636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7223_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4926_),
    .Y(_4927_)
);

FILL FILL_2__12848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14667_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14532_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6520_),
    .CLK(clk_bF$buf38),
    .Q(\u_ot.Xin1 [0])
);

FILL FILL_0__14247_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6461_),
    .B(_6459_),
    .C(_6462_),
    .Y(_5863_)
);

FILL FILL_1__7804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11174_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_3529_)
);

FILL FILL_0__8181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10167_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3157_),
    .B(_2686__bF$buf4),
    .C(_2928_),
    .Y(_3172_)
);

NAND2X1 _10032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2771_)
);

FILL FILL_2__9560_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_637_),
    .C(_635_),
    .Y(_638_)
);

OAI21X1 _7239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_235_),
    .C(_236_),
    .Y(_237_)
);

FILL FILL_2__13386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12799_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1483_),
    .Y(_1492_)
);

FILL FILL_1__12379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9386_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11657_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3397_),
    .CLK(clk_bF$buf59),
    .Q(\genblk1[4].u_ce.Xin1 [0])
);

OAI21X1 _11237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3877_),
    .C(_3873_),
    .Y(_3878_)
);

FILL FILL_1__13740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12313_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9805_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1717_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin12b [6])
);

FILL FILL_1__8762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13938_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6168_),
    .B(_6171_),
    .Y(_6172_)
);

FILL FILL_0__13518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11032_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _8197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1101_),
    .Y(_1108_)
);

FILL FILL_1__10865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7452_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4747_),
    .Y(_4748_)
);

FILL FILL_2__12657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8657_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _10928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3580_),
    .Y(_3582_)
);

FILL FILL_0__8237_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Acalc [4]),
    .B(_2672__bF$buf3),
    .Y(_3223_)
);

FILL FILL_0__14476_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6962_),
    .B(_6977_),
    .C(_6979_),
    .Y(_6980_)
);

FILL FILL_0__14056_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Xin12b [10]),
    .Y(_6639_)
);

FILL FILL_1__7613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3347_),
    .B(_2597_),
    .C(_2590_),
    .Y(_2583_)
);

FILL FILL_0__10396_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .C(_2989_),
    .Y(_2990_)
);

FILL FILL_1__8818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10303_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(gnd),
    .Y(_830_)
);

NAND2X1 _7468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_456_)
);

FILL FILL_1__12188_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _11886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4452_),
    .Y(_4453_)
);

FILL FILL_0__9195_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4092_),
    .Y(_4093_)
);

OAI21X1 _11046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3667_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3695_),
    .Y(_3360_)
);

FILL FILL_0__12962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7508_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2412_),
    .Y(_2413_)
);

FILL FILL_1__8991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13747_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5962_),
    .B(_5979_),
    .C(_5987_),
    .Y(_5990_)
);

FILL FILL_0__13327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7012_),
    .B(_7028_),
    .Y(_7032_)
);

FILL FILL_2_BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8046_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10737_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2563_),
    .CLK(clk_bF$buf7),
    .Q(\genblk1[3].u_ce.Yin12b [10])
);

NAND3X1 _10317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .B(_3043_),
    .C(_3042_),
    .Y(_3044_)
);

FILL FILL_1__12820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14285_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.RdyCtl [1]),
    .B(_6810_),
    .C(_6812_),
    .Y(_6813_)
);

OAI21X1 _14150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6475_),
    .B(_5887_),
    .C(_6483_),
    .Y(_5880_)
);

FILL FILL_1__7842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert130 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert131 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert133 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert135 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert136 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert138 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3198_),
    .Y(_3207_)
);

OAI21X1 _10070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2627_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_2807_),
    .Y(_2520_)
);

FILL FILL_1__8627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10532_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _7697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_672_),
    .Y(_673_)
);

OAI21X1 _7277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_272_),
    .C(_273_),
    .Y(_274_)
);

INVX2 _11695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4272_),
    .Y(_4273_)
);

INVX1 _11275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3911_),
    .Y(_3914_)
);

FILL FILL_2__7911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7737_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9843_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl [5]),
    .CLK(clk_bF$buf63),
    .Q(\genblk1[2].u_ce.Vld )
);

FILL FILL_0__7317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2233_),
    .Y(_2234_)
);

OAI21X1 _9003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1829_),
    .C(_1832_),
    .Y(_1833_)
);

FILL FILL_1__8380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6206_),
    .B(_6207_),
    .Y(_6208_)
);

FILL FILL_0__13136_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5830_),
    .B(_5104_),
    .C(_5098_),
    .Y(_5091_)
);

NAND2X1 _13001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5150__bF$buf1),
    .B(_5467_),
    .Y(_5468_)
);

FILL FILL_1__9585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10063_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [3]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf0),
    .Y(_6856_)
);

DFFPOSX1 _14206_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5882_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[7].u_ce.Yin0 [0])
);

FILL FILL_0__7490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8695_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3618_),
    .C(_3615_),
    .Y(_3619_)
);

FILL FILL_0__8275_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3257_),
    .B(\genblk1[3].u_ce.Ain12b [6]),
    .Y(_3259_)
);

AOI21X1 _10126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2860_),
    .B(_2834_),
    .C(_2859_),
    .Y(_2861_)
);

FILL FILL_2__9234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_83_),
    .C(_93_),
    .Y(\a[1] [0])
);

NAND3X1 _11084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .B(_3731_),
    .C(_3730_),
    .Y(_3732_)
);

FILL FILL_2__7720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7546_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2405_),
    .C(_2447_),
    .Y(_2449_)
);

FILL FILL_0__7126_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2047_),
    .C(_2051_),
    .Y(_2052_)
);

FILL FILL_1__11900_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4837_),
    .B(_4836_),
    .C(_4446_),
    .Y(_4838_)
);

FILL FILL_2__8505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13785_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5961_),
    .B(_5986_),
    .C(_6004_),
    .Y(_6025_)
);

FILL FILL_0__13365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5445_),
    .B(_5678_),
    .C(_5188__bF$buf4),
    .Y(_5686_)
);

FILL FILL_1__9394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10292_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6799_),
    .B(_6833__bF$buf3),
    .C(_7063_),
    .Y(_6791_)
);

AND2X2 _14435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6719_),
    .B(_6718_),
    .Y(_6720_)
);

NAND2X1 _14015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6350_),
    .B(_6352_),
    .Y(_6374_)
);

FILL FILL_1__7707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3437_),
    .B(\genblk1[4].u_ce.Acalc [8]),
    .C(_3438_),
    .Y(_3439_)
);

FILL FILL_0__8084_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2650_),
    .B(_3074_),
    .C(_3077_),
    .Y(_3080_)
);

FILL FILL_2__10817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13289_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _8923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1758_),
    .Y(_1759_)
);

INVX1 _8503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .Y(_1400_)
);

FILL FILL_1__7880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5387_),
    .C(_5391_),
    .Y(_5392_)
);

FILL FILL_0__12636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12216_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4466_),
    .B(_5000_),
    .C(_5016_),
    .Y(_4246_)
);

NAND2X1 _9708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.X_ [0]),
    .Y(_2491_)
);

FILL FILL_1__8665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14008_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6077_),
    .B(_6074_),
    .C(_6067_),
    .Y(_6079_)
);

FILL FILL_1__10768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7775_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [7]),
    .B(_2603_),
    .Y(_2628_)
);

FILL FILL_0__7355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2267_),
    .B(_2270_),
    .Y(_2271_)
);

MUX2X1 _9041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1869_),
    .B(_1868_),
    .S(_1811__bF$buf2),
    .Y(_1870_)
);

INVX1 _12098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4655_),
    .Y(_4656_)
);

FILL FILL_2__8734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .B(_6890_),
    .Y(_6891_)
);

NAND2X1 _14244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [9]),
    .Y(_6556_)
);

FILL FILL_1__7516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b [9]),
    .B(_2686__bF$buf1),
    .Y(_3294_)
);

FILL FILL_0__10299_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2897_),
    .B(_2896_),
    .C(_2744_),
    .Y(_2898_)
);

FILL FILL_2__10206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1614_),
    .Y(_1615_)
);

NAND3X1 _8312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .B(_1217_),
    .C(_1216_),
    .Y(_1218_)
);

OAI22X1 _11789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4356_),
    .B(_4359_),
    .C(_4324__bF$buf0),
    .D(_4353_),
    .Y(_4360_)
);

FILL FILL_0__9098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4002_),
    .B(_4003_),
    .Y(_4004_)
);

FILL FILL_1__13872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12865_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5209_),
    .B(_5208_),
    .S(_5151__bF$buf0),
    .Y(_5210_)
);

FILL FILL_0__12445_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4853_),
    .B(_4856_),
    .Y(_4857_)
);

FILL FILL_0__12025_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _9937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2679_),
    .B(_2658_),
    .C(_2649__bF$buf4),
    .Y(_2680_)
);

OAI21X1 _9517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2323_),
    .B(_2322_),
    .C(_1932_),
    .Y(_2324_)
);

FILL FILL_1__8474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert171 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert173 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6296_),
    .B(_6297_),
    .C(_5971_),
    .Y(_6298_)
);

FILL FILL_0_BUFX2_insert174 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(_5896_),
    .C(_5897_),
    .Y(_5898_)
);

FILL FILL_0_BUFX2_insert176 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert178 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7584_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2479_),
    .C(_2480_),
    .Y(_1715_)
);

FILL FILL_0__7164_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .B(_2087_),
    .Y(_2088_)
);

FILL FILL_0__10931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257250x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9310_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14893_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6784_),
    .CLK(clk_bF$buf72),
    .Q(\u_pa.acc_reg [17])
);

OAI21X1 _14473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6702_),
    .B(_6724_),
    .C(_6745_),
    .Y(_6524_)
);

NAND2X1 _14053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xcalc [9]),
    .B(_5949__bF$buf0),
    .Y(_6410_)
);

FILL FILL_1__7745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13508_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3115_),
    .B(_3091_),
    .C(_3114_),
    .Y(_3116_)
);

FILL FILL_2__10855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9081_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1793_),
    .B(_1792_),
    .Y(\genblk1[2].u_ce.Y_ [1])
);

AOI21X1 _8541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1435_),
    .B(_1436_),
    .C(_993_),
    .Y(_1437_)
);

INVX1 _8121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1035_),
    .Y(_1036_)
);

NAND2X1 _11598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .B(_4159_),
    .Y(_3425_)
);

OR2X2 _11178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3820_),
    .B(_3798_),
    .Y(_3822_)
);

FILL FILL_1__13681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12254_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Ain12b [9]),
    .Y(_2512_)
);

INVX1 _9326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .Y(_2142_)
);

FILL FILL_1__8283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13879_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6115_)
);

FILL FILL_0__13039_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5740_),
    .B(_5736_),
    .C(_5774_),
    .Y(_5776_)
);

FILL FILL_0__14820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10386_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14529_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6517_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin12b [7])
);

OAI21X1 _14109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_6459_),
    .C(_6460_),
    .Y(_5862_)
);

FILL FILL_0__7393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10320_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Ain12b [9]),
    .B(_172__bF$buf3),
    .Y(_780_)
);

FILL FILL_0__8598_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3526_)
);

FILL FILL_0__8178_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3152_),
    .B(_3162_),
    .C(_3168_),
    .Y(_3169_)
);

AOI21X1 _10029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2745_),
    .B(_2762_),
    .C(_2763_),
    .Y(_2768_)
);

FILL FILL_1__12952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11525_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _11810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4380_),
    .B(_4379_),
    .S(_4325__bF$buf4),
    .Y(_4381_)
);

FILL FILL_0__11105_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6586_),
    .C(_6585_),
    .Y(_6587_)
);

FILL FILL_1__7554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9700_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(_927_),
    .Y(_1645_)
);

NAND2X1 _8350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(_1233_),
    .Y(_1254_)
);

FILL FILL_2__7203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7869_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672__bF$buf4),
    .B(_2717_),
    .C(_2673_),
    .Y(_2515_)
);

FILL FILL_0__7449_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2356_),
    .B(_2358_),
    .C(_2345_),
    .Y(_1702_)
);

NAND3X1 _9135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf4),
    .B(_1958_),
    .C(_1953_),
    .Y(_1959_)
);

FILL FILL_1__8092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14275_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf2),
    .B(_6333_),
    .C(_6328_),
    .Y(_6334_)
);

FILL FILL_0__13688_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5930_),
    .C(_5931_),
    .Y(_5932_)
);

FILL FILL_0__13268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5594_),
    .B(_5588_),
    .C(_5243_),
    .Y(_5595_)
);

FILL FILL_1__9297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6965_),
    .B(_6973_),
    .Y(_6977_)
);

NAND2X1 _14338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [11]),
    .B(_6635_),
    .Y(_6636_)
);

AOI21X1 _7621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_577_),
    .C(_600_),
    .Y(_602_)
);

OR2X2 _7201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_152_),
    .Y(_202_)
);

NAND2X1 _10678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[3] [1]),
    .B(_3324_),
    .Y(_2589_)
);

AOI21X1 _10258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2960_),
    .B(_2981_),
    .C(_2979_),
    .Y(_2987_)
);

FILL FILL_1__12761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11334_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6429_),
    .B(_6439_),
    .C(_6445_),
    .Y(_6446_)
);

NAND2X1 _8826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .B(_1645_),
    .Y(_911_)
);

OR2X2 _8406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1306_),
    .B(_1284_),
    .Y(_1308_)
);

FILL FILL_1__7783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12959_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf5),
    .B(_5298_),
    .C(_5293_),
    .Y(_5299_)
);

FILL FILL_0__12119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf4),
    .B(_4861_),
    .Y(_4944_)
);

FILL FILL_0__13900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10053_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5961_),
    .C(_5986_),
    .Y(_5987_)
);

FILL FILL_2__7432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7258_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9784_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1696_),
    .CLK(clk_bF$buf42),
    .Q(\genblk1[2].u_ce.Xcalc [7])
);

NAND2X1 _9364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .B(_2177_),
    .Y(_2178_)
);

FILL FILL_2__8217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14084_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6138_),
    .B(_6151_),
    .C(_5951_),
    .Y(_6152_)
);

FILL FILL_0__13077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5802_),
    .B(_5804_),
    .C(_5806_),
    .Y(_5064_)
);

FILL FILL_1__12817_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf3)
);

FILL FILL_0__9404_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert105 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert106 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert107 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf0)
);

OAI21X1 _14567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6799_),
    .B(_6800_),
    .C(_6809_),
    .Y(_6810_)
);

NAND2X1 _14147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Y_ [1]),
    .B(_6466_),
    .Y(_6482_)
);

FILL FILL_1__7839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7419_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_807_),
    .C(_809_),
    .Y(_42_)
);

AOI21X1 _7430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_403_),
    .C(_409_),
    .Y(_420_)
);

NAND2X1 _10487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3202_),
    .B(_3203_),
    .Y(_3204_)
);

AND2X2 _10067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2789_),
    .B(_2804_),
    .Y(_2805_)
);

FILL FILL_1__12990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11143_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .C(gnd),
    .Y(_1524_)
);

NAND3X1 _8215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1114_),
    .B(_1121_),
    .C(_1124_),
    .Y(_1125_)
);

FILL FILL_1__7592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12768_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ycalc [10]),
    .Y(_5118_)
);

FILL FILL_0__12348_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4758_),
    .B(_4740_),
    .C(_4738_),
    .Y(_4766_)
);

FILL FILL_1__8797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10282_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6204_),
    .Y(_6205_)
);

NAND2X1 _13418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[6] [1]),
    .B(_5807_),
    .Y(_5097_)
);

FILL FILL_0__14914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7487_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _9593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2393_),
    .B(_2392_),
    .Y(_2394_)
);

AOI21X1 _9173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .B(_1963_),
    .C(_1964_),
    .Y(_1995_)
);

FILL FILL_1__11841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10414_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5967_),
    .C(_5968_),
    .Y(_5969_)
);

OAI21X1 _13171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5630_),
    .C(_5618_),
    .Y(_5631_)
);

NAND2X1 _7906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\a[0] [1]),
    .B(_810_),
    .Y(_75_)
);

FILL FILL_1__12626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9633_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4427_),
    .B(_4325__bF$buf1),
    .C(_4469_),
    .Y(_4470_)
);

FILL FILL_0__9213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7012_),
    .B(_7009_),
    .Y(_7013_)
);

OAI21X1 _14376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6545_),
    .B(\u_ot.LoadCtl_6_bF$buf1 ),
    .C(_6668_),
    .Y(_6504_)
);

FILL FILL_1__7648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14418_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3023_),
    .B(_3022_),
    .Y(_3024_)
);

FILL FILL_0__11792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11372_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8864_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_862_),
    .CLK(clk_bF$buf61),
    .Q(\genblk1[1].u_ce.Xcalc [11])
);

OAI21X1 _8444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(_1340_),
    .C(_1342_),
    .Y(_1344_)
);

NAND2X1 _8024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ycalc [6]),
    .B(_927_),
    .Y(_944_)
);

FILL FILL_2__14591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12997_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_5303_),
    .C(_5304_),
    .Y(_5335_)
);

FILL FILL_0__12157_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .Y(_4979_)
);

NAND2X1 _12022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4575_),
    .B(_4582_),
    .Y(_4583_)
);

OAI21X1 _9649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .B(_2436_),
    .C(_2434_),
    .Y(_2446_)
);

OAI21X1 _9229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1956_),
    .C(_2002_),
    .Y(_2049_)
);

FILL FILL_1__8186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6010_),
    .B(_5998_),
    .C(_6011_),
    .Y(_6022_)
);

NOR2X1 _13227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(gnd),
    .Y(_5683_)
);

FILL FILL_0__14723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10223_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(_689_),
    .Y(_690_)
);

FILL FILL_2__13022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11428_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4286_),
    .B(_4289_),
    .C(_4282_),
    .Y(_4290_)
);

FILL FILL_0__9022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11008_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14185_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5861_),
    .CLK(clk_bF$buf0),
    .Q(\genblk1[7].u_ce.Xin12b [11])
);

FILL FILL_1__7877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7457_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5296_),
    .C(_5342_),
    .Y(_5389_)
);

FILL FILL_0__11181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9603_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b [5]),
    .Y(_1559_)
);

NAND3X1 _8253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(_1139_),
    .C(_1122_),
    .Y(_1161_)
);

FILL FILL_1__10921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10501_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert150 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .Y(_135__bF$buf0)
);

BUFX2 BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .Y(_5151__bF$buf4)
);

FILL FILL_1__13393_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert152 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .Y(_5151__bF$buf3)
);

BUFX2 BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .Y(_5151__bF$buf2)
);

BUFX2 BUFX2_insert154 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .Y(_5151__bF$buf1)
);

BUFX2 BUFX2_insert155 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .Y(_5151__bF$buf0)
);

BUFX2 BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .Y(_4325__bF$buf4)
);

BUFX2 BUFX2_insert157 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .Y(_4325__bF$buf3)
);

BUFX2 BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .Y(_4325__bF$buf2)
);

INVX1 _12671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5152_)
);

FILL FILL_0__12386_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert159 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .Y(_4325__bF$buf1)
);

NAND3X1 _12251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf2),
    .B(_4796_),
    .C(_4794_),
    .Y(_4802_)
);

OAI21X1 _9878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Ycalc [11]),
    .C(_2600_),
    .Y(_2625_)
);

NAND3X1 _9458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848__bF$buf0),
    .B(_2264_),
    .C(_2259_),
    .Y(_2268_)
);

MUX2X1 _9038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_1865_),
    .S(_1811__bF$buf4),
    .Y(_1867_)
);

FILL FILL_1__11706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5962_),
    .C(_6240_),
    .Y(_6241_)
);

DFFPOSX1 _13456_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5056_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Acalc [7])
);

OAI21X1 _13036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5501_),
    .C(_5498_),
    .Y(_5502_)
);

FILL FILL_2__13918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10032_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7944_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .CLK(clk_bF$buf58),
    .Q(\genblk1[0].u_ce.Acalc [3])
);

NAND2X1 _7524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .B(_508_),
    .Y(_510_)
);

NAND2X1 _7104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_108_),
    .Y(\genblk1[0].u_ce.Y_ [0])
);

FILL FILL_2__13251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9689_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4493_),
    .B(_4490_),
    .C(_4485_),
    .Y(_4506_)
);

FILL FILL_2__9269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11237_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _11522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4140_),
    .B(_4144_),
    .Y(_4145_)
);

NAND3X1 _11102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .B(_3743_),
    .C(_3748_),
    .Y(_3749_)
);

OAI21X1 _8729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1611_),
    .B(_1555_),
    .C(_1610_),
    .Y(_1612_)
);

NAND3X1 _8309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1214_),
    .C(_1212_),
    .Y(_1215_)
);

FILL FILL_1__7686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13029_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5206_),
    .B(_5205_),
    .S(_5151__bF$buf0),
    .Y(_5207_)
);

INVX1 _12307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Ain0 [0]),
    .Y(_4854_)
);

FILL FILL_1__14810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9412_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1379_),
    .Y(_1380_)
);

NAND2X1 _8062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_978_)
);

FILL FILL_1__10310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12195_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.X_ [0]),
    .Y(_5005_)
);

NOR2X1 _12060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4354_),
    .Y(_4619_)
);

FILL FILL_2__12522_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.X_ [0]),
    .Y(_2478_)
);

INVX1 _9267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .Y(_2085_)
);

FILL FILL_1__11935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10508_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6046_),
    .B(_6058_),
    .C(_6056_),
    .Y(_6059_)
);

INVX1 _13265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Ain12b [4]),
    .Y(_5719_)
);

FILL FILL_2__13727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10261_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_724_),
    .Y(_725_)
);

OAI21X1 _7333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_239_),
    .C(_326_),
    .Y(_327_)
);

FILL FILL_2__13060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11466_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .Y(_4323_)
);

FILL FILL_0__9060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11046_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .Y(_3968_)
);

OAI21X1 _8958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1764_),
    .B(_1789_),
    .C(_1790_),
    .Y(_1791_)
);

OAI21X1 _8538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1410_),
    .C(_1433_),
    .Y(_1434_)
);

MUX2X1 _8118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1032_),
    .B(_1029_),
    .S(_972__bF$buf2),
    .Y(_1033_)
);

FILL FILL_1__7495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13258_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5413_),
    .Y(_5425_)
);

DFFPOSX1 _12536_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4190_),
    .CLK(clk_bF$buf20),
    .Q(\genblk1[5].u_ce.Ycalc [0])
);

INVX1 _12116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .Y(_4673_)
);

FILL FILL_0__13612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9221_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .Y(_1198_)
);

FILL FILL_1_CLKBUF1_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert98 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert99 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2301_),
    .B(_2302_),
    .Y(_2304_)
);

INVX2 _9076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1836_),
    .Y(_1903_)
);

FILL FILL_1__11744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8331_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3306_),
    .B(_3302_),
    .C(_3305_),
    .Y(_3310_)
);

FILL FILL_0__10317_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _13494_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5094_),
    .CLK(clk_bF$buf44),
    .Q(\genblk1[6].u_ce.Ain0 [1])
);

NAND3X1 _13074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .B(_5459_),
    .C(_5476_),
    .Y(_5538_)
);

FILL FILL_2__9710_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_777_),
    .C(_763_),
    .Y(_33_)
);

FILL FILL_2__13956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9536_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf5),
    .B(_4340_),
    .C(_4377_),
    .Y(_4378_)
);

FILL FILL_0__9116_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6922_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(_6923_),
    .Y(_6775_)
);

NAND3X1 _14279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(\u_ot.Xin12b [4]),
    .C(_6583_),
    .Y(_6584_)
);

FILL FILL_0__10490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10070_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7982_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_66_),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[0].u_ce.Ain12b [7])
);

OAI21X1 _7562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_545_),
    .C(_172__bF$buf4),
    .Y(_546_)
);

NAND2X1 _7142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_144_)
);

NAND2X1 _10199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2929_),
    .B(_2930_),
    .Y(_2931_)
);

FILL FILL_1__12282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x172950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11695_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4540_),
    .Y(_4543_)
);

NAND2X1 _11560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4151_),
    .Y(_4169_)
);

FILL FILL_0__11275_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_3647_),
    .C(_3784_),
    .Y(_3785_)
);

INVX1 _8767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.X_ [1]),
    .Y(_1643_)
);

NAND2X1 _8347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1248_),
    .B(_1250_),
    .Y(_1251_)
);

FILL FILL_2__14494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13067_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5176_),
    .Y(_5243_)
);

NOR2X1 _12345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4325__bF$buf3),
    .Y(_4889_)
);

FILL FILL_2__12807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14626_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[11]),
    .Y(Dout[11])
);

FILL FILL_0__7199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8560_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3489_)
);

FILL FILL_0__8140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10126_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xcalc [9]),
    .B(_2672__bF$buf2),
    .Y(_3133_)
);

FILL FILL257250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _7618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_158__bF$buf0),
    .C(_599_),
    .D(_596_),
    .Y(_20_)
);

FILL FILL_2__13765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9345_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11616_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3356_),
    .CLK(clk_bF$buf74),
    .Q(\genblk1[4].u_ce.Ycalc [3])
);

AOI22X1 _14088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6424_),
    .B(_5949__bF$buf0),
    .C(_6443_),
    .D(_5947_),
    .Y(_5858_)
);

FILL FILL_1__8721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8301_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _7791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_760_),
    .Y(_761_)
);

NAND2X1 _7371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_332_),
    .Y(_363_)
);

FILL FILL_1__12091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11831_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _8996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1818_),
    .S(_1810__bF$buf0),
    .Y(_1826_)
);

OAI21X1 _8576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1468_),
    .B(_1459_),
    .C(_994_),
    .Y(_1470_)
);

INVX2 _8156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .Y(_1068_)
);

FILL FILL_1__10824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xcalc [1]),
    .B(_5174__bF$buf3),
    .Y(_5461_)
);

FILL FILL_0__12289_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _12574_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4228_),
    .CLK(clk_bF$buf60),
    .Q(\genblk1[5].u_ce.Xin12b [11])
);

NAND2X1 _12154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4708_),
    .Y(_4709_)
);

FILL FILL_0__13650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8616_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Yin12b [8]),
    .B(_6148_),
    .C(_6147_),
    .Y(_6149_)
);

NAND2X1 _13359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(_5804_),
    .Y(_5805_)
);

FILL FILL_0__14855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14435_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6938_),
    .B(_6941_),
    .Y(_6943_)
);

FILL FILL_0__14015_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6562__bF$buf1),
    .B(_6601_),
    .C(_6602_),
    .Y(_6494_)
);

FILL FILL_1__11782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10775_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Y_ [0]),
    .Y(_3333_)
);

FILL FILL_0__10355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _10220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2950_),
    .Y(_2951_)
);

NAND2X1 _7847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(_807_),
    .Y(_808_)
);

NAND2X1 _7427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_416_),
    .Y(_417_)
);

FILL FILL_2__13994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9574_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4413_),
    .Y(_4414_)
);

FILL FILL_0__9154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4050_),
    .B(_4054_),
    .Y(_4055_)
);

NAND3X1 _11005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3647_),
    .B(_3652_),
    .C(_3655_),
    .Y(_3656_)
);

FILL FILL_0__12921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14713_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Xin12b [4]),
    .Y(_181_)
);

FILL FILL_0__13706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11220_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1287_)
);

FILL FILL_1__10633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7220_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4906_),
    .Y(_4924_)
);

FILL FILL_0__12098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8005_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5964_),
    .C(_5965_),
    .Y(_5966_)
);

NAND3X1 _13168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5188__bF$buf2),
    .B(_5622_),
    .C(_5620_),
    .Y(_5628_)
);

FILL FILL_0__14664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10164_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _7656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_629_),
    .C(_634_),
    .Y(_635_)
);

NAND3X1 _7236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_195_),
    .C(_213_),
    .Y(_234_)
);

FILL FILL_1__12796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9383_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _11654_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3394_),
    .CLK(clk_bF$buf17),
    .Q(\genblk1[4].u_ce.Xin12b [7])
);

FILL FILL_0__11369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3855_),
    .B(_3874_),
    .C(_3524__bF$buf1),
    .Y(_3875_)
);

FILL FILL_0__12730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7398_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9802_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1714_),
    .CLK(clk_bF$buf16),
    .Q(\genblk1[2].u_ce.Xin12b [11])
);

AOI21X1 _12859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5319_),
    .B(_5316_),
    .C(_5311_),
    .Y(_5332_)
);

NAND3X1 _12439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4969_),
    .B(_4970_),
    .C(_4959_),
    .Y(_4976_)
);

NAND2X1 _12019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362__bF$buf3),
    .B(_4579_),
    .Y(_4580_)
);

FILL FILL_1__14102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13935_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5963__bF$buf3),
    .B(_6166_),
    .C(_6163_),
    .Y(_6169_)
);

FILL FILL_0__13515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9124_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1104_),
    .C(_1101_),
    .Y(_1105_)
);

FILL FILL256650x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7467_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xcalc [6]),
    .Y(_4745_)
);

FILL FILL_2__12234_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [5]),
    .Y(_2211_)
);

FILL FILL_1__11227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8654_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3579_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_3580_)
);

FILL FILL_0__8234_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_3211_),
    .C(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .Y(_3221_)
);

OAI21X1 _13397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5104_),
    .C(_5825_),
    .Y(_5080_)
);

FILL FILL_2__13019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8815_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_83_),
    .C(_828_),
    .Y(_58_)
);

NAND2X1 _7465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_453_)
);

FILL FILL_1__12185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325__bF$buf1),
    .B(_4448_),
    .C(_4449_),
    .Y(_4450_)
);

FILL FILL_0__9192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11178_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4087_),
    .B(_4069_),
    .C(_4089_),
    .Y(_4090_)
);

OAI21X1 _11043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524__bF$buf2),
    .B(_3579_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_3693_)
);

FILL FILL_1__10918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7505_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .Y(_2410_)
);

FILL FILL256650x201750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .Y(_5149_)
);

OAI21X1 _12248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4776_),
    .B(_4773_),
    .C(_4362__bF$buf2),
    .Y(_4799_)
);

FILL FILL_1__14751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10251_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7025_),
    .B(_7028_),
    .C(_6833__bF$buf0),
    .Y(_7030_)
);

FILL FILL_0__14109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8043_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _10734_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2560_),
    .CLK(clk_bF$buf28),
    .Q(\genblk1[3].u_ce.Xin1 [1])
);

FILL FILL_0__10449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _10314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(_3040_),
    .C(_3038_),
    .Y(_3041_)
);

FILL FILL_0__11810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9668_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4498_),
    .B(_4502_),
    .C(_4503_),
    .Y(_4504_)
);

FILL FILL_0__9248_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4141_),
    .Y(_4142_)
);

FILL FILL_1__13602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8204_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .Y(_670_)
);

FILL FILL_1__14807_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_270_),
    .C(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_271_)
);

INVX1 _11692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [2]),
    .Y(_4270_)
);

OAI21X1 _11272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_3830_),
    .C(_3910_),
    .Y(_3911_)
);

FILL FILL_1__9409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11734_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _8899_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_897_),
    .CLK(clk_bF$buf3),
    .Q(\genblk1[1].u_ce.Yin0 [0])
);

AOI21X1 _8479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973__bF$buf0),
    .B(_1335_),
    .C(_1376_),
    .Y(_1377_)
);

NAND2X1 _8059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_975_)
);

FILL FILL_1__10307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL257550x104550 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9840_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(\genblk1[2].u_ce.LoadCtl [2]),
    .CLK(clk_bF$buf43),
    .Q(\genblk1[2].u_ce.LoadCtl [3])
);

FILL FILL_0__7314_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _9420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xcalc [6]),
    .Y(_2231_)
);

FILL FILL256950x183750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf1),
    .B(_1811__bF$buf2),
    .Y(_1830_)
);

INVX1 _12897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5366_),
    .Y(_5369_)
);

OAI21X1 _12477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4992_),
    .B(_4273_),
    .C(_5003_),
    .Y(_4235_)
);

OAI21X1 _12057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4614_),
    .C(_4615_),
    .Y(_4616_)
);

FILL FILL_1__14560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14338_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .B(_6851_),
    .C(_6853_),
    .Y(_6854_)
);

DFFPOSX1 _14203_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5879_),
    .CLK(clk_bF$buf39),
    .Q(\genblk1[7].u_ce.Yin12b [5])
);

FILL FILL_2__12272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8692_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3586_),
    .C(_3524__bF$buf3),
    .Y(_3616_)
);

FILL FILL_0__8272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10678_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .B(_3213_),
    .C(_2686__bF$buf1),
    .Y(_3256_)
);

FILL FILL_0__10258_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ycalc [8]),
    .Y(_2858_)
);

FILL FILL_2__9651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9477_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Xcalc [1]),
    .C(_4320_),
    .D(_4282_),
    .Y(_4321_)
);

FILL FILL_0__9057_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3959_),
    .B(_3961_),
    .Y(_3965_)
);

FILL FILL_1__13831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14616_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _7083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_87_),
    .C(_90_),
    .Y(_91_)
);

FILL FILL_0__13609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3722_),
    .B(_3728_),
    .C(_3726_),
    .Y(_3729_)
);

FILL FILL_1__9638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1190_),
    .C(_1188_),
    .Y(_1195_)
);

FILL FILL_1__10956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x86550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin12b [10]),
    .B(_4833_),
    .C(_4834_),
    .Y(_4835_)
);

FILL FILL_2__12748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14567_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_pa.acc_reg [11]),
    .B(_6833__bF$buf4),
    .C(En_bF$buf4),
    .Y(_7062_)
);

FILL FILL_0__14147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6706_),
    .B(_6717_),
    .Y(_6511_)
);

OAI21X1 _14012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6346_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6371_),
    .Y(_5854_)
);

FILL FILL_1__7704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11074_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _10772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [10]),
    .Y(_3436_)
);

FILL FILL_0__8081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10067_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3075_),
    .C(_3076_),
    .Y(_3077_)
);

FILL FILL_2__9460_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _7979_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_63_),
    .CLK(clk_bF$buf11),
    .Q(\genblk1[0].u_ce.Ain12b [8])
);

FILL FILL_2__9040_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _7559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172__bF$buf4),
    .B(_542_),
    .C(_537_),
    .Y(_543_)
);

OAI21X1 _7139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_139_),
    .C(_140_),
    .Y(_141_)
);

FILL FILL_2__13286_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Acalc [2]),
    .Y(_1756_)
);

FILL FILL_1__12699_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_1316_),
    .C(_1396_),
    .Y(_1397_)
);

FILL FILL_1__12279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_4450_),
    .C(_4516_),
    .Y(_4540_)
);

FILL FILL_0__9286_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _11557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3498_),
    .C(_4167_),
    .Y(_3399_)
);

AOI22X1 _11137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .B(_3780_),
    .C(_3781_),
    .D(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3782_)
);

FILL FILL_1__13640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12213_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_1759_),
    .C(_2489_),
    .Y(_1721_)
);

FILL FILL_1__8662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13838_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6073_),
    .Y(_6076_)
);

FILL FILL_0__13418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11772_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _8097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1012_)
);

FILL FILL_1__10345_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _14908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7071_[0]),
    .Y(Dout[0])
);

FILL FILL_0__7772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7352_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _12095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4652_),
    .B(_4641_),
    .S(vdd),
    .Y(_4653_)
);

FILL FILL_2__12977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8557_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _10828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .Y(_3486_)
);

FILL FILL_0__8137_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _10408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3128_),
    .Y(_3131_)
);

FILL FILL_1__12911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14376_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6871_),
    .B(_6887_),
    .C(_6886_),
    .Y(_6888_)
);

NAND2X1 _14241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [8]),
    .Y(_6554_)
);

FILL FILL_1__7513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256650x136950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3289_),
    .B(_3291_),
    .C(_3277_),
    .Y(_2547_)
);

FILL FILL_0__10296_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _10161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2894_),
    .Y(_2895_)
);

FILL FILL_1__8718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10203_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _7788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .Y(_758_)
);

AOI21X1 _7368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_360_),
    .C(_160_),
    .Y(_361_)
);

FILL FILL_1__12088_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .B(_4354_),
    .C(_4325__bF$buf3),
    .Y(_4357_)
);

FILL FILL_0__9095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4000_),
    .B(_3997_),
    .Y(_4001_)
);

FILL FILL_0__12862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7828_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .B(_2675_),
    .S(_2649__bF$buf2),
    .Y(_2677_)
);

FILL FILL_0__7408_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _9514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Xin12b [10]),
    .B(_2319_),
    .C(_2320_),
    .Y(_2321_)
);

FILL FILL_1__8471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert140 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert142 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert143 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13647_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6274_),
    .B(_6265_),
    .C(_5963__bF$buf2),
    .Y(_6295_)
);

FILL FILL_0_BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13227_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_5893_),
    .C(_5894_),
    .Y(_5895_)
);

FILL FILL_0_BUFX2_insert145 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert147 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert149 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6940_)
);

FILL FILL_0__7581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__12786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8366_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2899_),
    .B(_3313_),
    .C(_3331_),
    .Y(_2563_)
);

NAND2X1 _10217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_2948_)
);

FILL FILL_1__12720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11713_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14890_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6781_),
    .CLK(clk_bF$buf40),
    .Q(\u_pa.acc_reg [14])
);

NAND2X1 _14470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.X_ [1]),
    .Y(_6744_)
);

OR2X2 _14050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6405_),
    .Y(_6408_)
);

FILL FILL_1__7742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12918_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3095_),
    .B(_2672__bF$buf2),
    .C(_3113_),
    .D(_3110_),
    .Y(_2534_)
);

FILL FILL_1__8947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10432_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _7597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .B(_579_),
    .Y(_580_)
);

OAI21X1 _7177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_176_),
    .C(_177_),
    .Y(_178_)
);

OAI21X1 _11595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4187_),
    .B(_4155_),
    .C(_4188_),
    .Y(_3416_)
);

NAND3X1 _11175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3535_),
    .B(_3816_),
    .C(_3813_),
    .Y(_3819_)
);

FILL FILL_2__11217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7637_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Ain12b [8]),
    .Y(_2510_)
);

FILL FILL_0__7217_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _9323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2127_),
    .S(gnd),
    .Y(_2139_)
);

FILL FILL_1__8280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13876_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6111_),
    .B(_6095_),
    .C(_6107_),
    .Y(_6112_)
);

FILL FILL_0__13036_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5750_),
    .B(_5764_),
    .C(_5762_),
    .Y(_5773_)
);

FILL FILL_1__9485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10383_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _14526_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6514_),
    .CLK(clk_bF$buf64),
    .Q(\u_ot.Xin12b [8])
);

INVX1 _14106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[6].u_ce.X_ [0]),
    .Y(_6458_)
);

FILL FILL_0__7390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__8595_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _10866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3523_)
);

FILL FILL_0__8175_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _10446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3147_),
    .B(_2672__bF$buf2),
    .C(_3166_),
    .D(_2670_),
    .Y(_2537_)
);

AOI21X1 _10026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2765_),
    .B(_2746_),
    .C(_2674_),
    .Y(_2766_)
);

FILL FILL_2__10908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__7200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__11446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7866_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _9972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .B(_2684_),
    .C(_2714_),
    .Y(_2715_)
);

FILL FILL_0__7446_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _9552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .B(_2355_),
    .Y(_2356_)
);

AOI21X1 _9132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1913_),
    .B(_1811__bF$buf1),
    .C(_1955_),
    .Y(_1956_)
);

FILL FILL_1__11800_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4726_),
    .B(_4741_),
    .Y(_4743_)
);

FILL FILL_2__8825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__8405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14272_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5925__bF$buf3),
    .B(_6250_),
    .Y(_6331_)
);

FILL FILL_0__13685_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(_5927_),
    .C(_5928_),
    .Y(_5929_)
);

FILL FILL_0__13265_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5584_),
    .B(_5566_),
    .C(_5564_),
    .Y(_5592_)
);

FILL FILL256950x115350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__9294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10192_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6970_),
    .B(_6973_),
    .C(_6833__bF$buf2),
    .Y(_6975_)
);

INVX1 _14335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ot.Xin12b [11]),
    .Y(_6633_)
);

FILL FILL_1__7607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__11397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _10675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3349_),
    .B(_3321_),
    .C(_2587_),
    .Y(_2580_)
);

AOI21X1 _10255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2984_),
    .B(_2983_),
    .C(_2674_),
    .Y(_2985_)
);

FILL FILL_0__11751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _8823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1641_),
    .C(_1674_),
    .Y(_902_)
);

NAND3X1 _8403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1021_),
    .B(_1302_),
    .C(_1299_),
    .Y(_1305_)
);

FILL FILL_1__7780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__14130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__13123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__12956_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5253_),
    .B(_5151__bF$buf2),
    .C(_5295_),
    .Y(_5296_)
);

INVX1 _12401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[5].u_ce.Acalc [7]),
    .Y(_4941_)
);

FILL FILL_0__12116_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _9608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_2407_),
    .Y(_2408_)
);

FILL FILL_1__8985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__8145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14328_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _13606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(\genblk1[7].u_ce.Xin0 [1]),
    .S(vdd),
    .Y(_5984_)
);

FILL FILL_1__10668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__10248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__7255_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _9781_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1693_),
    .CLK(clk_bF$buf2),
    .Q(\genblk1[2].u_ce.Xcalc [4])
);

NOR2X1 _9361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810__bF$buf3),
    .B(_2174_),
    .Y(_2175_)
);

FILL FILL_2__8634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__10602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__14081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__13074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL256950x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__13401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__12814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__9401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__14279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6802_),
    .B(_6806_),
    .Y(_6807_)
);

OAI21X1 _14144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6477_),
    .B(_6463_),
    .C(_6480_),
    .Y(_5877_)
);

FILL FILL_1__7836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__7416_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _10484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .B(gnd),
    .S(_3199_),
    .Y(_3201_)
);

FILL FILL_0__10199_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _10064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .B(_2797_),
    .C(_2790_),
    .Y(_2802_)
);

FILL FILL_2__10946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__10106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__9172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__11140_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _8632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1521_)
);

NOR3X1 _8212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1081_),
    .B(_1100_),
    .C(_1072_),
    .Y(_1122_)
);

endmodule
