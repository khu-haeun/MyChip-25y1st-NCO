magic
tech scmos
magscale 1 2
timestamp 1740657676
<< metal1 >>
rect -62 5778 -2 6018
rect 5910 6002 6002 6018
rect 4067 5937 4093 5943
rect 2487 5857 2513 5863
rect -62 5762 30 5778
rect -62 5298 -2 5762
rect 5942 5538 6002 6002
rect 5910 5522 6002 5538
rect 4187 5457 4213 5463
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 5507 5177 5573 5183
rect 5447 5137 5513 5143
rect 5942 5058 6002 5522
rect 5910 5042 6002 5058
rect 3167 4917 3253 4923
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 2947 4637 2973 4643
rect 5942 4578 6002 5042
rect 5910 4562 6002 4578
rect 5157 4497 5173 4503
rect 5157 4427 5163 4497
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 5737 4143 5743 4173
rect 5737 4137 5773 4143
rect 5942 4098 6002 4562
rect 5910 4082 6002 4098
rect 5727 4017 5763 4023
rect 5757 3967 5763 4017
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 2687 3697 2713 3703
rect 5197 3703 5203 3753
rect 5187 3697 5203 3703
rect 2307 3677 2333 3683
rect 5942 3618 6002 4082
rect 5910 3602 6002 3618
rect 5427 3517 5473 3523
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 647 3197 693 3203
rect 5942 3138 6002 3602
rect 5910 3122 6002 3138
rect 4427 3057 4473 3063
rect 3187 3037 3233 3043
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 1867 2777 1913 2783
rect 5942 2658 6002 3122
rect 5910 2642 6002 2658
rect 4347 2497 4373 2503
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 5942 2178 6002 2642
rect 5910 2162 6002 2178
rect 287 2117 313 2123
rect 5447 2117 5493 2123
rect 5717 2077 5733 2083
rect 147 2017 213 2023
rect 5717 2003 5723 2077
rect 5717 1997 5733 2003
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 1567 1777 1593 1783
rect 5942 1698 6002 2162
rect 5910 1682 6002 1698
rect 1067 1617 1093 1623
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 2927 1357 2953 1363
rect 5942 1218 6002 1682
rect 5910 1202 6002 1218
rect 5247 1137 5263 1143
rect 5257 1127 5263 1137
rect -62 962 30 978
rect -62 498 -2 962
rect 3847 857 3933 863
rect 4727 857 4773 863
rect 5942 738 6002 1202
rect 5910 722 6002 738
rect 4267 657 4333 663
rect -62 482 30 498
rect -62 18 -2 482
rect 2747 377 2813 383
rect 5942 258 6002 722
rect 5910 242 6002 258
rect 1947 197 1993 203
rect -62 2 30 18
rect 5942 2 6002 242
<< m2contact >>
rect 4053 5933 4067 5947
rect 4093 5933 4107 5947
rect 2473 5853 2487 5867
rect 2513 5853 2527 5867
rect 4173 5453 4187 5467
rect 4213 5453 4227 5467
rect 5493 5173 5507 5187
rect 5573 5173 5587 5187
rect 5433 5133 5447 5147
rect 5513 5133 5527 5147
rect 3153 4913 3167 4927
rect 3253 4913 3267 4927
rect 2933 4633 2947 4647
rect 2973 4633 2987 4647
rect 5173 4493 5187 4507
rect 5153 4413 5167 4427
rect 5733 4173 5747 4187
rect 5773 4133 5787 4147
rect 5713 4013 5727 4027
rect 5753 3953 5767 3967
rect 5193 3753 5207 3767
rect 2673 3693 2687 3707
rect 2713 3693 2727 3707
rect 5173 3693 5187 3707
rect 2293 3673 2307 3687
rect 2333 3673 2347 3687
rect 5413 3513 5427 3527
rect 5473 3513 5487 3527
rect 633 3193 647 3207
rect 693 3193 707 3207
rect 4413 3053 4427 3067
rect 4473 3053 4487 3067
rect 3173 3033 3187 3047
rect 3233 3033 3247 3047
rect 1853 2773 1867 2787
rect 1913 2773 1927 2787
rect 4333 2493 4347 2507
rect 4373 2493 4387 2507
rect 273 2113 287 2127
rect 313 2113 327 2127
rect 5433 2113 5447 2127
rect 5493 2113 5507 2127
rect 133 2013 147 2027
rect 213 2013 227 2027
rect 5733 2073 5747 2087
rect 5733 1993 5747 2007
rect 1553 1773 1567 1787
rect 1593 1773 1607 1787
rect 1053 1613 1067 1627
rect 1093 1613 1107 1627
rect 2913 1353 2927 1367
rect 2953 1353 2967 1367
rect 5233 1133 5247 1147
rect 5253 1113 5267 1127
rect 3833 853 3847 867
rect 3933 853 3947 867
rect 4713 853 4727 867
rect 4773 853 4787 867
rect 4253 653 4267 667
rect 4333 653 4347 667
rect 2733 373 2747 387
rect 2813 373 2827 387
rect 1933 193 1947 207
rect 1993 193 2007 207
<< metal2 >>
rect 4436 6056 4463 6063
rect 96 5936 123 5943
rect 116 5887 123 5936
rect 216 5896 223 5913
rect 596 5887 603 5923
rect 956 5916 983 5923
rect 16 5847 23 5873
rect 76 5387 83 5873
rect 236 5667 243 5883
rect 976 5883 983 5916
rect 1007 5916 1023 5923
rect 216 5636 243 5643
rect 116 5587 123 5603
rect 116 5436 123 5473
rect 156 5443 163 5573
rect 156 5436 183 5443
rect 96 5416 103 5433
rect 136 5363 143 5413
rect 176 5407 183 5436
rect 136 5356 163 5363
rect 136 5176 143 5193
rect 156 5167 163 5356
rect 76 4956 103 4963
rect 96 4907 103 4956
rect 116 4887 123 4923
rect 56 4696 83 4703
rect 116 4696 143 4703
rect 56 4507 63 4696
rect 56 4443 63 4493
rect 56 4436 83 4443
rect 116 4367 123 4443
rect 16 3907 23 4253
rect 136 4227 143 4696
rect 96 4196 103 4213
rect 96 4016 123 4023
rect 16 1347 23 3853
rect 116 3703 123 4016
rect 136 3923 143 4193
rect 156 3947 163 4933
rect 176 4927 183 5193
rect 196 5187 203 5433
rect 216 5427 223 5636
rect 256 5467 263 5623
rect 276 5436 283 5673
rect 316 5443 323 5873
rect 676 5867 683 5873
rect 716 5807 723 5883
rect 816 5847 823 5883
rect 856 5787 863 5883
rect 976 5876 1003 5883
rect 416 5636 423 5673
rect 556 5636 563 5653
rect 316 5436 343 5443
rect 336 5427 343 5436
rect 196 4947 203 5173
rect 216 5156 223 5373
rect 256 5207 263 5423
rect 296 5407 303 5423
rect 256 5127 263 5143
rect 256 4967 263 5113
rect 276 5087 283 5123
rect 256 4936 263 4953
rect 176 4207 183 4913
rect 296 4907 303 5393
rect 436 5147 443 5453
rect 456 5407 463 5633
rect 536 5423 543 5603
rect 556 5436 563 5453
rect 596 5436 603 5473
rect 616 5467 623 5673
rect 696 5656 723 5663
rect 716 5607 723 5656
rect 836 5656 843 5673
rect 516 5416 543 5423
rect 516 5387 523 5416
rect 456 5123 463 5373
rect 536 5156 563 5163
rect 456 5116 483 5123
rect 396 4936 403 5073
rect 356 4923 363 4933
rect 436 4923 443 4973
rect 456 4947 463 5073
rect 356 4916 383 4923
rect 416 4916 443 4923
rect 476 4923 483 5116
rect 516 5087 523 5123
rect 556 4987 563 5156
rect 576 4963 583 5413
rect 616 5167 623 5453
rect 656 5436 663 5473
rect 676 5456 683 5593
rect 796 5396 823 5403
rect 596 5156 613 5163
rect 636 5156 643 5173
rect 676 5143 683 5213
rect 796 5176 803 5396
rect 656 5136 683 5143
rect 556 4956 583 4963
rect 536 4927 543 4943
rect 476 4916 503 4923
rect 196 4487 203 4873
rect 216 4696 223 4893
rect 256 4487 263 4703
rect 276 4487 283 4683
rect 356 4476 363 4493
rect 396 4476 423 4483
rect 256 4456 283 4463
rect 276 4427 283 4456
rect 316 4456 343 4463
rect 196 4187 203 4413
rect 296 4407 303 4433
rect 216 4216 223 4393
rect 296 4227 303 4353
rect 136 3916 163 3923
rect 96 3696 123 3703
rect 96 3607 103 3696
rect 116 3516 143 3523
rect 116 3323 123 3516
rect 116 3316 143 3323
rect 76 3147 83 3223
rect 96 3087 103 3203
rect 116 3167 123 3223
rect 136 3127 143 3316
rect 56 3036 63 3073
rect 156 3067 163 3916
rect 176 3547 183 3973
rect 216 3587 223 4013
rect 236 3987 243 4173
rect 256 4016 263 4193
rect 276 4127 283 4203
rect 296 4167 303 4213
rect 296 4003 303 4153
rect 316 4127 323 4456
rect 356 4216 363 4433
rect 376 4327 383 4463
rect 416 4447 423 4476
rect 376 4167 383 4193
rect 396 4187 403 4213
rect 416 4127 423 4203
rect 436 4147 443 4693
rect 496 4667 503 4916
rect 616 4907 623 5113
rect 676 4956 683 5073
rect 696 4907 703 4923
rect 536 4663 543 4893
rect 516 4656 543 4663
rect 476 4447 483 4463
rect 496 4227 503 4493
rect 516 4287 523 4656
rect 536 4427 543 4633
rect 576 4627 583 4663
rect 636 4483 643 4683
rect 696 4667 703 4893
rect 716 4647 723 5173
rect 736 5127 743 5163
rect 776 4923 783 5133
rect 816 4936 823 4953
rect 776 4916 803 4923
rect 756 4676 763 4693
rect 776 4687 783 4916
rect 796 4676 823 4683
rect 816 4667 823 4676
rect 836 4643 843 4913
rect 856 4787 863 5393
rect 896 5227 903 5433
rect 916 5407 923 5653
rect 956 5647 963 5673
rect 996 5627 1003 5876
rect 936 5587 943 5623
rect 976 5607 983 5623
rect 1016 5607 1023 5916
rect 1456 5916 1483 5923
rect 1496 5916 1523 5923
rect 1476 5907 1483 5916
rect 1196 5887 1203 5903
rect 1196 5647 1203 5773
rect 1056 5616 1083 5623
rect 976 5436 983 5573
rect 1076 5467 1083 5616
rect 1016 5436 1043 5443
rect 996 5187 1003 5423
rect 1036 5407 1043 5436
rect 1156 5436 1163 5613
rect 1196 5436 1203 5573
rect 1056 5156 1063 5433
rect 1216 5427 1223 5623
rect 1136 5327 1143 5423
rect 1176 5387 1183 5423
rect 1116 5156 1143 5163
rect 916 5107 923 5143
rect 1016 5103 1023 5143
rect 1116 5127 1123 5156
rect 1216 5143 1223 5313
rect 1236 5187 1243 5633
rect 1256 5587 1263 5873
rect 1316 5867 1323 5883
rect 1356 5807 1363 5883
rect 1336 5647 1343 5793
rect 1296 5407 1303 5423
rect 1336 5387 1343 5633
rect 1356 5607 1363 5623
rect 1396 5567 1403 5793
rect 1436 5707 1443 5893
rect 1516 5867 1523 5916
rect 1876 5916 1903 5923
rect 1516 5623 1523 5673
rect 1556 5636 1563 5653
rect 1596 5647 1603 5673
rect 1516 5616 1543 5623
rect 1636 5623 1643 5633
rect 1616 5616 1643 5623
rect 1476 5467 1483 5613
rect 1476 5403 1483 5453
rect 1556 5403 1563 5553
rect 1656 5436 1663 5893
rect 1696 5507 1703 5903
rect 1796 5896 1823 5903
rect 1796 5887 1803 5896
rect 1896 5887 1903 5916
rect 2016 5916 2043 5923
rect 2036 5867 2043 5916
rect 2276 5916 2283 5933
rect 2316 5916 2323 6013
rect 3376 5936 3403 5943
rect 3476 5936 3503 5943
rect 2516 5916 2543 5923
rect 2576 5916 2603 5923
rect 2656 5916 2663 5933
rect 3376 5927 3383 5936
rect 1996 5643 2003 5693
rect 1976 5636 2003 5643
rect 1736 5616 1763 5623
rect 1736 5607 1743 5616
rect 1696 5436 1703 5493
rect 1476 5396 1503 5403
rect 1536 5396 1563 5403
rect 1616 5416 1643 5423
rect 1616 5383 1623 5416
rect 1616 5376 1643 5383
rect 1556 5176 1583 5183
rect 1196 5136 1223 5143
rect 996 5096 1023 5103
rect 996 4967 1003 5096
rect 1016 5087 1023 5096
rect 1156 5087 1163 5123
rect 916 4956 943 4963
rect 916 4907 923 4956
rect 1076 4923 1083 4973
rect 1116 4936 1123 4953
rect 1076 4916 1103 4923
rect 1136 4916 1143 4953
rect 896 4647 903 4703
rect 916 4667 923 4683
rect 1036 4663 1043 4773
rect 1176 4727 1183 5113
rect 1236 5107 1243 5153
rect 1276 5136 1303 5143
rect 1236 4956 1243 5093
rect 1276 4927 1283 5136
rect 1336 4967 1343 5143
rect 1416 5127 1423 5143
rect 1476 5007 1483 5163
rect 1556 5147 1563 5176
rect 1636 5167 1643 5376
rect 1676 5187 1683 5423
rect 1676 5116 1703 5123
rect 1456 4956 1483 4963
rect 1436 4927 1443 4943
rect 1076 4676 1083 4713
rect 1036 4656 1063 4663
rect 816 4636 843 4643
rect 636 4476 663 4483
rect 276 3996 303 4003
rect 296 3947 303 3996
rect 476 3976 483 3993
rect 496 3943 503 4133
rect 476 3936 503 3943
rect 236 3736 243 3933
rect 276 3727 283 3743
rect 216 3507 223 3523
rect 196 3143 203 3393
rect 236 3267 243 3593
rect 256 3507 263 3573
rect 256 3307 263 3493
rect 236 3167 243 3253
rect 176 3136 203 3143
rect 96 3036 103 3053
rect 56 2523 63 2753
rect 76 2723 83 2763
rect 156 2743 163 3013
rect 136 2736 163 2743
rect 76 2716 103 2723
rect 96 2536 103 2716
rect 56 2516 83 2523
rect 76 1987 83 2516
rect 96 2276 103 2473
rect 116 2367 123 2523
rect 136 2243 143 2273
rect 116 2236 143 2243
rect 96 2027 103 2043
rect 136 2027 143 2043
rect 156 1783 163 2713
rect 176 2367 183 3136
rect 216 3087 223 3133
rect 216 3036 223 3073
rect 236 3003 243 3153
rect 256 3127 263 3223
rect 296 3167 303 3723
rect 316 3607 323 3733
rect 416 3687 423 3733
rect 316 3516 323 3533
rect 336 3483 343 3503
rect 336 3476 363 3483
rect 356 3447 363 3476
rect 336 3216 343 3313
rect 236 2996 263 3003
rect 216 2527 223 2543
rect 256 2467 263 2996
rect 276 2727 283 2743
rect 96 1596 103 1783
rect 136 1776 163 1783
rect 36 1327 43 1573
rect 116 1563 123 1573
rect 96 1556 123 1563
rect 96 1363 103 1556
rect 76 1356 103 1363
rect 76 1343 83 1356
rect 56 1336 83 1343
rect 116 1336 123 1533
rect 56 1107 63 1336
rect 156 1327 163 1776
rect 176 1547 183 2353
rect 196 2263 203 2453
rect 276 2276 283 2293
rect 196 2256 223 2263
rect 236 2056 243 2113
rect 256 2107 263 2243
rect 296 2127 303 3133
rect 316 3067 323 3113
rect 316 2727 323 3053
rect 356 2767 363 3433
rect 416 3247 423 3673
rect 396 3063 403 3153
rect 416 3087 423 3233
rect 436 3207 443 3933
rect 456 3447 463 3793
rect 476 3707 483 3936
rect 516 3747 523 4183
rect 536 4127 543 4193
rect 536 4007 543 4113
rect 556 4027 563 4473
rect 596 4327 603 4443
rect 636 4403 643 4443
rect 616 4396 643 4403
rect 616 4207 623 4396
rect 656 4267 663 4476
rect 716 4456 723 4473
rect 696 4216 703 4413
rect 496 3667 503 3723
rect 596 3707 603 3973
rect 656 3967 663 4213
rect 716 4207 723 4313
rect 556 3696 583 3703
rect 476 3447 483 3483
rect 516 3476 543 3483
rect 496 3236 503 3253
rect 396 3056 423 3063
rect 416 2747 423 3056
rect 436 3007 443 3043
rect 516 3036 523 3053
rect 376 2523 383 2693
rect 436 2587 443 2993
rect 476 2756 483 3013
rect 536 2987 543 3476
rect 556 3107 563 3653
rect 576 3587 583 3696
rect 616 3667 623 3953
rect 696 3867 703 3983
rect 636 3527 643 3703
rect 576 3516 603 3523
rect 576 3483 583 3516
rect 576 3476 603 3483
rect 576 3007 583 3273
rect 596 3267 603 3476
rect 616 3247 623 3493
rect 636 3207 643 3233
rect 616 3187 623 3203
rect 616 2967 623 3153
rect 456 2707 463 2743
rect 476 2556 483 2613
rect 496 2607 503 2743
rect 516 2556 523 2573
rect 356 2516 383 2523
rect 316 2127 323 2493
rect 376 2327 383 2516
rect 536 2523 543 2953
rect 576 2776 603 2783
rect 636 2776 643 2993
rect 556 2527 563 2713
rect 576 2707 583 2776
rect 516 2516 543 2523
rect 416 2276 443 2283
rect 256 2023 263 2043
rect 236 2016 263 2023
rect 216 1787 223 2013
rect 196 1563 203 1593
rect 236 1576 243 2016
rect 276 1587 283 2113
rect 336 2096 343 2273
rect 356 2207 363 2263
rect 396 2227 403 2243
rect 396 2107 403 2213
rect 436 2187 443 2276
rect 436 2096 443 2113
rect 456 2107 463 2313
rect 316 2076 323 2093
rect 356 2076 373 2083
rect 376 2027 383 2073
rect 196 1556 223 1563
rect 176 1147 183 1513
rect 76 1116 83 1133
rect 96 1087 103 1093
rect 156 863 163 1113
rect 136 856 163 863
rect 136 823 143 856
rect 176 827 183 1133
rect 276 887 283 1083
rect 296 1027 303 1973
rect 336 1796 363 1803
rect 356 1647 363 1796
rect 356 1607 363 1633
rect 376 1627 383 2013
rect 396 1667 403 2093
rect 456 1867 463 2053
rect 476 1847 483 2513
rect 496 2276 503 2293
rect 496 1827 503 2093
rect 516 2067 523 2516
rect 576 2207 583 2673
rect 596 2567 603 2733
rect 656 2687 663 3653
rect 716 3647 723 3993
rect 676 3227 683 3553
rect 736 3516 743 4273
rect 756 4143 763 4633
rect 776 4407 783 4633
rect 816 4443 823 4636
rect 856 4456 863 4473
rect 916 4447 923 4653
rect 996 4476 1003 4613
rect 1036 4496 1043 4513
rect 816 4436 843 4443
rect 776 4216 803 4223
rect 776 4167 783 4216
rect 816 4167 823 4203
rect 756 4136 783 4143
rect 776 3727 783 4136
rect 756 3687 763 3703
rect 776 3543 783 3683
rect 776 3536 803 3543
rect 796 3507 803 3536
rect 816 3523 823 3673
rect 836 3667 843 3983
rect 876 3787 883 4253
rect 1016 4227 1023 4463
rect 1056 4327 1063 4463
rect 916 3987 923 4163
rect 1047 4156 1063 4163
rect 976 3996 983 4133
rect 1036 3987 1043 4153
rect 1056 4007 1063 4073
rect 856 3536 863 3573
rect 876 3547 883 3733
rect 896 3583 903 3973
rect 916 3736 923 3753
rect 896 3576 923 3583
rect 816 3516 843 3523
rect 876 3516 903 3523
rect 696 3496 723 3503
rect 696 3287 703 3496
rect 816 3487 823 3516
rect 696 3207 703 3223
rect 676 2747 683 3193
rect 756 3167 763 3453
rect 776 3187 783 3473
rect 816 3236 823 3253
rect 796 3207 803 3223
rect 696 3043 703 3093
rect 696 3036 723 3043
rect 696 2727 703 3036
rect 736 3007 743 3023
rect 736 2723 743 2763
rect 736 2716 763 2723
rect 616 2327 623 2543
rect 676 2527 683 2543
rect 696 2527 703 2573
rect 696 2283 703 2333
rect 676 2276 703 2283
rect 607 2256 623 2263
rect 596 2107 603 2253
rect 716 2127 723 2593
rect 736 2547 743 2613
rect 756 2543 763 2716
rect 796 2627 803 2743
rect 816 2603 823 3173
rect 856 3147 863 3243
rect 876 3227 883 3473
rect 896 3267 903 3516
rect 856 2987 863 3003
rect 916 2967 923 3576
rect 936 3007 943 3673
rect 956 3507 963 3573
rect 1016 3516 1023 3753
rect 1056 3567 1063 3993
rect 1076 3747 1083 4453
rect 1096 3727 1103 4673
rect 1216 4647 1223 4663
rect 1116 4407 1123 4443
rect 1156 4423 1163 4433
rect 1136 4416 1163 4423
rect 1116 4147 1123 4393
rect 1136 4216 1143 4416
rect 1176 4187 1183 4223
rect 1196 4167 1203 4203
rect 1156 3996 1163 4013
rect 1176 3967 1183 3983
rect 1196 3923 1203 4153
rect 1196 3916 1223 3923
rect 1116 3703 1123 3773
rect 1076 3647 1083 3703
rect 1096 3696 1123 3703
rect 1056 3516 1063 3553
rect 1096 3543 1103 3696
rect 1096 3536 1123 3543
rect 976 3496 1003 3503
rect 976 3467 983 3496
rect 796 2596 823 2603
rect 796 2556 803 2596
rect 836 2556 843 2613
rect 756 2536 783 2543
rect 756 2487 763 2536
rect 816 2523 823 2543
rect 796 2516 823 2523
rect 736 2267 743 2293
rect 796 2287 803 2516
rect 676 2047 683 2093
rect 756 2076 763 2273
rect 856 2267 863 2953
rect 896 2687 903 2723
rect 916 2556 923 2573
rect 896 2527 903 2543
rect 936 2507 943 2993
rect 956 2583 963 3293
rect 976 3256 983 3293
rect 1096 3283 1103 3536
rect 1156 3527 1163 3733
rect 1216 3707 1223 3916
rect 1236 3867 1243 4853
rect 1256 4667 1263 4913
rect 1276 4663 1283 4693
rect 1276 4656 1303 4663
rect 1276 4456 1283 4633
rect 1336 4447 1343 4643
rect 1356 4547 1363 4633
rect 1356 4456 1363 4533
rect 1396 4467 1403 4673
rect 1416 4663 1423 4913
rect 1476 4887 1483 4956
rect 1636 4947 1643 4973
rect 1596 4936 1623 4943
rect 1616 4927 1623 4936
rect 1676 4936 1683 5116
rect 1736 4947 1743 5593
rect 1756 5436 1763 5553
rect 1876 5427 1883 5633
rect 1896 5456 1903 5613
rect 1916 5567 1923 5623
rect 1956 5527 1963 5623
rect 2036 5607 2043 5853
rect 2076 5616 2103 5623
rect 2016 5436 2043 5443
rect 2076 5436 2083 5616
rect 2136 5607 2143 5623
rect 2216 5616 2243 5623
rect 1776 5407 1783 5423
rect 1996 5347 2003 5433
rect 1956 5176 1983 5183
rect 1456 4676 1463 4693
rect 1416 4656 1443 4663
rect 1456 4636 1483 4643
rect 1456 4447 1463 4636
rect 1476 4627 1483 4636
rect 1636 4587 1643 4933
rect 1656 4567 1663 4913
rect 1696 4907 1703 4923
rect 1696 4627 1703 4893
rect 1716 4627 1723 4663
rect 1736 4647 1743 4913
rect 1776 4667 1783 4933
rect 1816 4787 1823 5163
rect 1836 5127 1843 5143
rect 1916 5143 1923 5153
rect 1956 5147 1963 5176
rect 1916 5136 1943 5143
rect 1916 4956 1923 5136
rect 2016 5127 2023 5436
rect 2056 5147 2063 5423
rect 2136 5407 2143 5593
rect 2236 5483 2243 5616
rect 2216 5476 2243 5483
rect 2216 5456 2223 5476
rect 2176 5423 2183 5433
rect 2176 5416 2203 5423
rect 2196 5407 2203 5416
rect 2096 5156 2103 5393
rect 2256 5367 2263 5613
rect 2276 5427 2283 5873
rect 2356 5636 2363 5653
rect 2396 5636 2403 5673
rect 2436 5647 2443 5883
rect 2516 5867 2523 5916
rect 2596 5883 2603 5916
rect 2876 5916 2893 5923
rect 2576 5876 2603 5883
rect 2476 5663 2483 5853
rect 2576 5667 2583 5876
rect 2456 5656 2483 5663
rect 2456 5623 2463 5656
rect 2296 5436 2303 5573
rect 2376 5436 2383 5473
rect 2416 5467 2423 5623
rect 2436 5616 2463 5623
rect 2236 5156 2263 5163
rect 2136 4976 2163 4983
rect 1896 4927 1903 4943
rect 2116 4923 2123 4953
rect 2136 4927 2143 4976
rect 2216 4927 2223 4943
rect 2096 4916 2123 4923
rect 1896 4887 1903 4913
rect 1836 4656 1843 4693
rect 1536 4456 1543 4473
rect 1576 4467 1583 4513
rect 1676 4476 1683 4573
rect 1736 4487 1743 4633
rect 1836 4476 1843 4613
rect 1876 4476 1883 4673
rect 1296 4347 1303 4443
rect 1296 4216 1303 4313
rect 1316 4127 1323 4193
rect 1336 4187 1343 4223
rect 1316 4016 1323 4113
rect 1336 3996 1343 4013
rect 1356 3987 1363 4203
rect 1196 3667 1203 3703
rect 1236 3696 1263 3703
rect 1196 3587 1203 3653
rect 1256 3516 1263 3696
rect 1156 3503 1163 3513
rect 1076 3276 1103 3283
rect 1136 3496 1163 3503
rect 1016 3256 1043 3263
rect 1036 3187 1043 3256
rect 1016 3036 1023 3173
rect 1056 3043 1063 3093
rect 1076 3047 1083 3276
rect 1136 3236 1143 3496
rect 1236 3447 1243 3503
rect 1096 3067 1103 3193
rect 1116 3087 1123 3223
rect 1156 3187 1163 3223
rect 1196 3216 1203 3333
rect 1236 3187 1243 3233
rect 1036 3036 1063 3043
rect 1036 2743 1043 3036
rect 1116 2783 1123 3033
rect 1236 3023 1243 3173
rect 1256 3063 1263 3333
rect 1276 3207 1283 3223
rect 1296 3067 1303 3713
rect 1316 3187 1323 3223
rect 1256 3056 1283 3063
rect 1256 3047 1263 3056
rect 1316 3023 1323 3053
rect 1156 3007 1163 3023
rect 1216 3016 1243 3023
rect 1296 3016 1323 3023
rect 976 2707 983 2743
rect 1016 2736 1043 2743
rect 1096 2776 1123 2783
rect 1156 2776 1163 2813
rect 956 2576 983 2583
rect 976 2567 983 2576
rect 956 2467 963 2543
rect 996 2527 1003 2713
rect 776 2227 783 2263
rect 436 1816 463 1823
rect 436 1767 443 1816
rect 536 1787 543 1813
rect 416 1563 423 1593
rect 396 1556 423 1563
rect 336 1347 343 1353
rect 336 1316 343 1333
rect 436 1327 443 1613
rect 496 1596 503 1753
rect 536 1607 543 1773
rect 356 1163 363 1313
rect 496 1303 503 1553
rect 516 1527 523 1583
rect 476 1296 503 1303
rect 476 1283 483 1296
rect 456 1276 483 1283
rect 336 1156 363 1163
rect 336 1116 343 1156
rect 376 1116 383 1253
rect 356 1087 363 1103
rect 76 743 83 813
rect 56 736 83 743
rect 56 663 63 736
rect 36 656 63 663
rect 36 367 43 656
rect 96 623 103 813
rect 116 807 123 823
rect 136 816 163 823
rect 396 803 403 853
rect 356 796 403 803
rect 236 656 243 673
rect 76 616 103 623
rect 176 636 203 643
rect 76 407 83 616
rect 176 347 183 636
rect 356 636 363 796
rect 96 307 103 343
rect 176 323 183 333
rect 176 316 203 323
rect 96 156 103 233
rect 116 176 123 313
rect 236 176 243 613
rect 256 567 263 623
rect 336 567 343 623
rect 376 616 383 673
rect 416 647 423 1113
rect 536 907 543 1083
rect 556 867 563 1853
rect 616 1796 623 1833
rect 596 1747 603 1783
rect 676 1767 683 2033
rect 696 1827 703 2053
rect 796 1783 803 1813
rect 596 1567 603 1733
rect 616 1596 623 1633
rect 656 1596 663 1653
rect 736 1647 743 1783
rect 776 1776 803 1783
rect 816 1767 823 1793
rect 836 1767 843 2113
rect 896 2107 903 2313
rect 916 2287 923 2313
rect 996 2263 1003 2473
rect 916 2256 943 2263
rect 976 2256 1003 2263
rect 876 2056 883 2073
rect 916 2067 923 2256
rect 1016 2227 1023 2673
rect 1096 2587 1103 2776
rect 1096 2556 1123 2563
rect 1136 2556 1163 2563
rect 1116 2487 1123 2556
rect 1136 2307 1143 2333
rect 1036 2283 1043 2293
rect 1036 2276 1063 2283
rect 1136 2263 1143 2293
rect 1116 2256 1143 2263
rect 1156 2263 1163 2556
rect 1176 2307 1183 2613
rect 1156 2256 1183 2263
rect 996 2127 1003 2173
rect 936 2076 963 2083
rect 996 2076 1003 2113
rect 896 2027 903 2043
rect 896 1847 903 2013
rect 936 2007 943 2076
rect 856 1796 863 1813
rect 876 1747 883 1763
rect 916 1647 923 1783
rect 716 1547 723 1613
rect 756 1603 763 1633
rect 936 1627 943 1833
rect 736 1596 763 1603
rect 576 1167 583 1293
rect 616 1267 623 1303
rect 456 603 463 833
rect 496 647 503 843
rect 556 827 563 853
rect 596 827 603 1153
rect 636 1096 643 1173
rect 696 1116 703 1253
rect 716 943 723 1133
rect 736 1107 743 1596
rect 816 1563 823 1613
rect 936 1596 943 1613
rect 796 1556 823 1563
rect 796 1336 803 1513
rect 836 1343 843 1593
rect 976 1347 983 2053
rect 996 1827 1003 1993
rect 996 1796 1003 1813
rect 1116 1787 1123 2093
rect 1156 2076 1163 2213
rect 1176 2147 1183 2256
rect 1196 2227 1203 2993
rect 1216 2827 1223 3016
rect 1216 2727 1223 2813
rect 1296 2783 1303 3016
rect 1336 3003 1343 3953
rect 1376 3763 1383 4333
rect 1396 4147 1403 4413
rect 1496 4187 1503 4193
rect 1416 4023 1423 4173
rect 1436 4087 1443 4183
rect 1476 4147 1483 4183
rect 1396 4016 1423 4023
rect 1396 3967 1403 4016
rect 1356 3756 1383 3763
rect 1356 3347 1363 3756
rect 1376 3736 1393 3743
rect 1376 3687 1383 3736
rect 1436 3736 1443 3893
rect 1456 3547 1463 3993
rect 1496 3587 1503 4073
rect 1516 3987 1523 4113
rect 1536 4007 1543 4413
rect 1616 4227 1623 4473
rect 1616 4196 1623 4213
rect 1576 3996 1583 4173
rect 1636 4167 1643 4453
rect 1676 4436 1703 4443
rect 1596 4127 1603 4163
rect 1556 3976 1563 3993
rect 1556 3747 1563 3813
rect 1636 3787 1643 4013
rect 1676 3947 1683 4436
rect 1736 4207 1743 4223
rect 1716 4167 1723 4203
rect 1707 3996 1723 4003
rect 1716 3927 1723 3996
rect 1556 3716 1563 3733
rect 1636 3716 1643 3773
rect 1536 3523 1543 3703
rect 1576 3687 1583 3693
rect 1516 3516 1543 3523
rect 1556 3516 1563 3573
rect 1376 3447 1383 3483
rect 1276 2776 1303 2783
rect 1316 2996 1343 3003
rect 1276 2756 1283 2776
rect 1296 2727 1303 2743
rect 1216 2556 1243 2563
rect 1216 2427 1223 2556
rect 1236 2263 1243 2273
rect 1316 2267 1323 2996
rect 1336 2687 1343 2773
rect 1356 2527 1363 3073
rect 1376 3027 1383 3433
rect 1416 3407 1423 3483
rect 1456 3256 1483 3263
rect 1516 3256 1523 3333
rect 1456 3247 1463 3256
rect 1596 3223 1603 3553
rect 1656 3523 1663 3613
rect 1636 3516 1663 3523
rect 1636 3223 1643 3516
rect 1596 3216 1623 3223
rect 1636 3216 1663 3223
rect 1396 3036 1403 3053
rect 1436 3036 1443 3173
rect 1416 3007 1423 3013
rect 1536 2987 1543 3003
rect 1416 2776 1443 2783
rect 1436 2727 1443 2776
rect 1496 2776 1523 2783
rect 1436 2627 1443 2713
rect 1216 2256 1243 2263
rect 1356 2263 1363 2473
rect 1376 2427 1383 2523
rect 1456 2487 1463 2773
rect 1496 2747 1503 2776
rect 1496 2567 1503 2733
rect 1536 2687 1543 2763
rect 1596 2556 1603 3053
rect 1336 2256 1363 2263
rect 1316 2147 1323 2193
rect 1276 2076 1303 2083
rect 1316 2076 1323 2133
rect 1136 2056 1143 2073
rect 1176 1947 1183 2063
rect 1256 2027 1263 2073
rect 1296 2047 1303 2076
rect 1056 1627 1063 1783
rect 1156 1767 1163 1833
rect 1256 1807 1263 2013
rect 1296 1827 1303 2033
rect 1376 1967 1383 2263
rect 1416 2087 1423 2453
rect 1436 2287 1443 2413
rect 1456 2227 1463 2263
rect 1196 1796 1223 1803
rect 996 1607 1003 1613
rect 996 1563 1003 1593
rect 1036 1576 1043 1593
rect 996 1556 1023 1563
rect 1056 1483 1063 1563
rect 1036 1476 1063 1483
rect 836 1336 863 1343
rect 756 1147 763 1333
rect 856 1287 863 1336
rect 956 1316 963 1333
rect 976 1287 983 1303
rect 1036 1267 1043 1476
rect 1096 1407 1103 1613
rect 1176 1587 1183 1773
rect 1216 1687 1223 1796
rect 1236 1767 1243 1783
rect 1276 1627 1283 1653
rect 1216 1596 1243 1603
rect 1056 1307 1063 1323
rect 1096 1316 1103 1393
rect 1136 1327 1143 1583
rect 1216 1347 1223 1596
rect 1316 1583 1323 1813
rect 1376 1783 1383 1953
rect 1376 1776 1403 1783
rect 1436 1727 1443 2043
rect 1456 1767 1463 2213
rect 1476 1827 1483 2553
rect 1516 2427 1523 2543
rect 1576 2387 1583 2543
rect 1496 2276 1503 2333
rect 1536 2287 1543 2313
rect 1576 2203 1583 2373
rect 1576 2196 1603 2203
rect 1496 1807 1503 2053
rect 1516 2043 1523 2073
rect 1516 2036 1543 2043
rect 1556 1787 1563 2013
rect 1576 2007 1583 2043
rect 1596 2027 1603 2196
rect 1616 1987 1623 2263
rect 1636 2147 1643 2993
rect 1676 2787 1683 3533
rect 1696 3527 1703 3703
rect 1736 3647 1743 3873
rect 1756 3563 1763 4013
rect 1796 3887 1803 4473
rect 1856 4447 1863 4463
rect 1896 4327 1903 4873
rect 2256 4867 2263 5156
rect 2276 4967 2283 5413
rect 2316 5387 2323 5423
rect 2356 5407 2363 5423
rect 2416 5367 2423 5433
rect 2436 5407 2443 5616
rect 2456 5436 2463 5493
rect 2536 5436 2543 5473
rect 2556 5467 2563 5633
rect 2556 5427 2563 5453
rect 2476 5387 2483 5423
rect 2316 4936 2323 5353
rect 2336 5143 2343 5173
rect 2496 5156 2503 5393
rect 2576 5147 2583 5653
rect 2676 5607 2683 5623
rect 2816 5603 2823 5613
rect 2896 5607 2903 5913
rect 2956 5887 2963 5923
rect 3196 5916 3223 5923
rect 3216 5907 3223 5916
rect 3036 5707 3043 5873
rect 3216 5687 3223 5873
rect 2816 5596 2843 5603
rect 2616 5347 2623 5453
rect 2636 5436 2643 5533
rect 2796 5456 2803 5513
rect 2656 5367 2663 5423
rect 2696 5327 2703 5423
rect 2716 5387 2723 5453
rect 2776 5327 2783 5423
rect 2656 5156 2663 5173
rect 2336 5136 2363 5143
rect 2396 5067 2403 5143
rect 2476 5116 2493 5123
rect 2416 4956 2423 5053
rect 2276 4923 2283 4933
rect 2276 4916 2303 4923
rect 1976 4643 1983 4693
rect 2196 4676 2203 4693
rect 1956 4636 1983 4643
rect 2056 4627 2063 4663
rect 2116 4647 2123 4663
rect 1856 4167 1863 4203
rect 1876 4187 1883 4223
rect 1916 4216 1923 4553
rect 1936 4436 1963 4443
rect 1936 4407 1943 4436
rect 1996 4427 2003 4433
rect 1996 4403 2003 4413
rect 1976 4396 2003 4403
rect 1796 3727 1803 3743
rect 1776 3687 1783 3723
rect 1756 3556 1783 3563
rect 1776 3487 1783 3556
rect 1796 3507 1803 3713
rect 1856 3667 1863 3993
rect 1916 3943 1923 3963
rect 1896 3936 1923 3943
rect 1896 3847 1903 3936
rect 1936 3907 1943 4393
rect 1876 3727 1883 3773
rect 1856 3516 1863 3633
rect 1876 3496 1883 3513
rect 1696 3036 1703 3333
rect 1776 3236 1783 3473
rect 1896 3407 1903 3833
rect 1956 3767 1963 4153
rect 1976 3967 1983 4396
rect 2016 4203 2023 4533
rect 2136 4483 2143 4653
rect 2176 4627 2183 4643
rect 2256 4483 2263 4493
rect 2136 4476 2163 4483
rect 2236 4476 2263 4483
rect 1996 4196 2023 4203
rect 1996 4027 2003 4196
rect 2136 4183 2143 4476
rect 2056 4176 2083 4183
rect 2136 4176 2163 4183
rect 2056 4167 2063 4176
rect 2156 4087 2163 4176
rect 2196 4067 2203 4183
rect 2276 4167 2283 4713
rect 2296 4667 2303 4713
rect 1996 4007 2003 4013
rect 2016 3996 2023 4053
rect 2156 4016 2183 4023
rect 2036 3967 2043 3983
rect 1976 3736 1983 3933
rect 1916 3427 1923 3723
rect 1936 3567 1943 3733
rect 1916 3287 1923 3413
rect 1876 3236 1883 3273
rect 1756 3207 1763 3223
rect 1756 3036 1763 3073
rect 1796 3023 1803 3213
rect 1856 3203 1863 3213
rect 1856 3196 1883 3203
rect 1716 3016 1743 3023
rect 1776 3016 1803 3023
rect 1696 2756 1703 2813
rect 1716 2727 1723 2733
rect 1696 2536 1703 2573
rect 1676 2487 1683 2523
rect 1736 2503 1743 3016
rect 1816 2807 1823 3193
rect 1836 3043 1843 3093
rect 1836 3036 1863 3043
rect 1876 3036 1883 3196
rect 1896 3067 1903 3223
rect 1856 2907 1863 3036
rect 1756 2727 1763 2773
rect 1776 2747 1783 2763
rect 1756 2527 1763 2553
rect 1776 2527 1783 2733
rect 1796 2707 1803 2753
rect 1816 2687 1823 2763
rect 1856 2727 1863 2773
rect 1876 2747 1883 2953
rect 1836 2543 1843 2593
rect 1716 2496 1743 2503
rect 1676 2263 1683 2293
rect 1656 2256 1683 2263
rect 1716 2167 1723 2496
rect 1796 2427 1803 2543
rect 1836 2536 1863 2543
rect 1736 2307 1743 2313
rect 1776 2296 1803 2303
rect 1796 2227 1803 2296
rect 1856 2263 1863 2513
rect 1856 2256 1883 2263
rect 1716 2076 1723 2153
rect 1636 2007 1643 2053
rect 1576 1787 1583 1973
rect 1636 1796 1643 1833
rect 1356 1687 1363 1693
rect 1256 1547 1263 1583
rect 1296 1576 1323 1583
rect 1316 1567 1323 1576
rect 1356 1563 1363 1673
rect 1356 1556 1383 1563
rect 1236 1307 1243 1313
rect 1056 1187 1063 1293
rect 936 1116 943 1153
rect 1076 1123 1083 1303
rect 1116 1267 1123 1303
rect 1176 1267 1183 1303
rect 776 1087 783 1103
rect 716 936 743 943
rect 636 823 643 833
rect 736 827 743 936
rect 776 843 783 1073
rect 1016 1067 1023 1123
rect 1056 1116 1083 1123
rect 836 867 843 1013
rect 976 856 983 893
rect 776 836 803 843
rect 836 836 843 853
rect 616 816 643 823
rect 796 823 803 836
rect 796 816 823 823
rect 596 807 603 813
rect 616 647 623 673
rect 656 636 663 693
rect 456 596 483 603
rect 536 567 543 613
rect 416 363 423 393
rect 716 387 723 603
rect 456 367 463 383
rect 496 376 523 383
rect 416 356 443 363
rect 476 347 483 363
rect 296 247 303 323
rect 316 147 323 343
rect 516 327 523 376
rect 736 343 743 413
rect 716 336 743 343
rect 576 247 583 323
rect 336 136 343 213
rect 356 156 363 233
rect 396 156 403 233
rect 456 147 463 193
rect 496 176 503 213
rect 576 147 583 233
rect 696 163 703 323
rect 696 156 723 163
rect 467 136 483 143
rect 656 127 663 143
rect 716 127 723 156
rect 776 147 783 813
rect 816 727 823 816
rect 796 427 803 673
rect 816 607 823 653
rect 856 647 863 733
rect 876 636 883 673
rect 836 407 843 633
rect 856 616 863 633
rect 796 227 803 393
rect 876 356 883 593
rect 796 136 803 213
rect 816 116 823 233
rect 856 227 863 343
rect 936 327 943 373
rect 836 136 843 193
rect 916 127 923 173
rect 956 167 963 713
rect 996 647 1003 673
rect 1036 647 1043 753
rect 1056 523 1063 1116
rect 1176 1116 1203 1123
rect 1076 847 1083 1093
rect 1096 887 1103 1033
rect 1156 1027 1163 1103
rect 1096 856 1103 873
rect 1136 867 1143 1013
rect 1196 887 1203 1116
rect 1196 847 1203 873
rect 1156 667 1163 673
rect 1216 667 1223 1303
rect 1256 867 1263 1333
rect 1316 1283 1323 1533
rect 1416 1527 1423 1563
rect 1316 1276 1343 1283
rect 1416 1116 1423 1493
rect 1436 1347 1443 1573
rect 1456 1316 1463 1633
rect 1476 1627 1483 1783
rect 1676 1783 1683 1993
rect 1576 1596 1583 1613
rect 1496 1387 1503 1593
rect 1596 1587 1603 1773
rect 1616 1587 1623 1783
rect 1656 1776 1683 1783
rect 1696 1767 1703 2063
rect 1716 1947 1723 2033
rect 1636 1596 1643 1633
rect 1576 1303 1583 1513
rect 1716 1507 1723 1933
rect 1736 1647 1743 1783
rect 1756 1727 1763 2093
rect 1776 1847 1783 2133
rect 1856 2076 1863 2213
rect 1836 2047 1843 2063
rect 1856 1827 1863 2033
rect 1836 1796 1863 1803
rect 1776 1747 1783 1753
rect 1736 1527 1743 1633
rect 1616 1316 1623 1393
rect 1736 1336 1743 1513
rect 1776 1336 1783 1733
rect 1816 1616 1823 1633
rect 1436 1287 1443 1303
rect 1336 1083 1343 1113
rect 1436 1087 1443 1103
rect 1316 1076 1343 1083
rect 1436 1067 1443 1073
rect 1236 787 1243 803
rect 1276 727 1283 833
rect 1136 607 1143 623
rect 1256 616 1263 633
rect 1276 607 1283 713
rect 1296 616 1303 853
rect 1316 836 1343 843
rect 1316 767 1323 836
rect 1356 747 1363 803
rect 1036 516 1063 523
rect 956 143 963 153
rect 936 136 963 143
rect 976 136 983 213
rect 996 163 1003 363
rect 1036 247 1043 516
rect 1056 347 1063 493
rect 1107 376 1123 383
rect 1076 327 1083 343
rect 1096 307 1103 373
rect 996 156 1023 163
rect 1016 87 1023 156
rect 1076 143 1083 213
rect 1236 207 1243 603
rect 1436 596 1443 793
rect 1456 787 1463 1073
rect 1456 616 1463 773
rect 1476 667 1483 1303
rect 1576 1296 1603 1303
rect 1576 1287 1583 1296
rect 1636 1167 1643 1303
rect 1596 1083 1603 1113
rect 1576 1076 1603 1083
rect 1496 843 1503 873
rect 1496 836 1523 843
rect 1536 643 1543 823
rect 1516 636 1543 643
rect 1576 636 1603 643
rect 1356 356 1383 363
rect 1276 307 1283 323
rect 1376 227 1383 356
rect 1396 327 1403 593
rect 1436 307 1443 353
rect 1536 347 1543 393
rect 1596 387 1603 636
rect 1616 387 1623 1133
rect 1716 1116 1723 1133
rect 1836 1116 1843 1713
rect 1856 1627 1863 1796
rect 1896 1687 1903 3033
rect 1936 3007 1943 3273
rect 1956 3047 1963 3653
rect 1976 3536 1983 3553
rect 2016 3547 2023 3733
rect 1996 3263 2003 3273
rect 2036 3267 2043 3753
rect 2096 3736 2123 3743
rect 2116 3707 2123 3736
rect 1976 3256 2003 3263
rect 1976 3227 1983 3256
rect 1956 2807 1963 3013
rect 1976 2987 1983 3193
rect 2056 3003 2063 3053
rect 2036 2996 2063 3003
rect 2036 2827 2043 2853
rect 1927 2776 1943 2783
rect 1916 2567 1923 2753
rect 1916 2527 1923 2553
rect 1936 2287 1943 2733
rect 1996 2727 2003 2763
rect 2016 2707 2023 2753
rect 1976 2427 1983 2523
rect 2036 2407 2043 2813
rect 2076 2807 2083 3493
rect 2136 3467 2143 3483
rect 2136 3287 2143 3453
rect 2156 3387 2163 3953
rect 2176 3767 2183 4016
rect 2216 3996 2243 4003
rect 2216 3927 2223 3996
rect 2316 3827 2323 4613
rect 2336 4476 2343 4513
rect 2356 4496 2363 4633
rect 2376 4547 2383 4663
rect 2376 4476 2383 4533
rect 2396 4243 2403 4953
rect 2436 4696 2443 4713
rect 2496 4687 2503 5113
rect 2596 4956 2603 4973
rect 2576 4936 2583 4953
rect 2616 4867 2623 4943
rect 2656 4887 2663 4973
rect 2676 4967 2683 5143
rect 2696 4927 2703 5153
rect 2416 4527 2423 4673
rect 2576 4567 2583 4663
rect 2656 4587 2663 4693
rect 2516 4476 2543 4483
rect 2536 4467 2543 4476
rect 2436 4456 2463 4463
rect 2396 4236 2423 4243
rect 2416 4203 2423 4236
rect 2436 4207 2443 4456
rect 2496 4427 2503 4463
rect 2476 4227 2483 4233
rect 2516 4216 2523 4413
rect 2396 4196 2423 4203
rect 2256 3716 2263 3753
rect 2296 3707 2303 3733
rect 2336 3687 2343 4183
rect 2376 4167 2383 4183
rect 2356 3727 2363 3973
rect 2376 3727 2383 3753
rect 2096 3087 2103 3253
rect 2096 3047 2103 3073
rect 2116 3027 2123 3273
rect 2156 3236 2163 3273
rect 2136 3067 2143 3223
rect 2196 3047 2203 3533
rect 2236 3427 2243 3503
rect 2276 3487 2283 3533
rect 2296 3467 2303 3673
rect 2396 3527 2403 4173
rect 2556 4167 2563 4533
rect 2656 4523 2663 4573
rect 2696 4567 2703 4913
rect 2716 4867 2723 5173
rect 2856 5147 2863 5493
rect 2956 5463 2963 5613
rect 2976 5507 2983 5623
rect 3016 5607 3023 5623
rect 3176 5623 3183 5653
rect 3216 5636 3223 5673
rect 3256 5636 3283 5643
rect 3176 5616 3203 5623
rect 3276 5607 3283 5636
rect 2956 5456 2983 5463
rect 2936 5387 2943 5423
rect 2976 5407 2983 5456
rect 2876 5176 2903 5183
rect 2936 5176 2963 5183
rect 2736 4967 2743 5143
rect 2776 5127 2783 5143
rect 2756 5107 2763 5123
rect 2876 5107 2883 5176
rect 2756 4936 2763 4953
rect 2736 4703 2743 4793
rect 2716 4696 2743 4703
rect 2716 4627 2723 4696
rect 2636 4516 2663 4523
rect 2636 4227 2643 4516
rect 2656 4443 2663 4493
rect 2696 4456 2703 4553
rect 2736 4443 2743 4493
rect 2656 4436 2683 4443
rect 2716 4436 2743 4443
rect 2596 4147 2603 4183
rect 2436 4007 2443 4013
rect 2436 3976 2443 3993
rect 2496 3987 2503 4013
rect 2516 3947 2523 4013
rect 2596 3996 2603 4113
rect 2576 3967 2583 3983
rect 2636 3967 2643 4183
rect 2656 3967 2663 4213
rect 2476 3736 2483 3933
rect 2536 3707 2543 3723
rect 2556 3687 2563 3733
rect 2316 3467 2323 3483
rect 2236 3267 2243 3373
rect 2296 3263 2303 3333
rect 2376 3267 2383 3493
rect 2396 3367 2403 3493
rect 2276 3256 2303 3263
rect 2256 3087 2263 3243
rect 2296 3207 2303 3256
rect 2336 3223 2343 3253
rect 2396 3236 2403 3353
rect 2336 3216 2363 3223
rect 2256 3036 2283 3043
rect 2156 2967 2163 3023
rect 2056 2527 2063 2773
rect 2136 2756 2143 2773
rect 2176 2743 2183 2773
rect 2116 2563 2123 2743
rect 2156 2736 2183 2743
rect 2236 2743 2243 3033
rect 2256 3007 2263 3036
rect 2296 2967 2303 3023
rect 2336 3016 2343 3073
rect 2356 2967 2363 3216
rect 2376 3203 2383 3223
rect 2416 3207 2423 3223
rect 2376 3196 2403 3203
rect 2296 2767 2303 2783
rect 2236 2736 2263 2743
rect 2096 2556 2123 2563
rect 2076 2276 2083 2433
rect 2096 2303 2103 2556
rect 2136 2536 2143 2573
rect 2176 2536 2203 2543
rect 2156 2516 2163 2533
rect 2196 2487 2203 2536
rect 2236 2527 2243 2713
rect 2256 2567 2263 2736
rect 2276 2707 2283 2763
rect 2316 2756 2343 2763
rect 2336 2747 2343 2756
rect 2256 2503 2263 2533
rect 2256 2496 2283 2503
rect 2096 2296 2123 2303
rect 1916 2256 1943 2263
rect 1916 1647 1923 2133
rect 1936 1767 1943 2256
rect 1996 2187 2003 2233
rect 1976 2076 1983 2093
rect 1996 2063 2003 2173
rect 2016 2167 2023 2263
rect 2056 2147 2063 2263
rect 2036 2076 2063 2083
rect 1996 2056 2023 2063
rect 1956 1816 1963 2053
rect 2056 1947 2063 2076
rect 2116 1867 2123 2296
rect 2136 2076 2143 2193
rect 2156 2107 2163 2473
rect 2236 2276 2243 2453
rect 2276 2267 2283 2496
rect 2316 2327 2323 2523
rect 2336 2327 2343 2733
rect 2356 2367 2363 2933
rect 2376 2547 2383 3133
rect 2396 3127 2403 3196
rect 2436 3147 2443 3513
rect 2516 3507 2523 3553
rect 2536 3487 2543 3533
rect 2536 3256 2543 3273
rect 2556 3227 2563 3673
rect 2576 3567 2583 3953
rect 2596 3703 2603 3953
rect 2676 3807 2683 4413
rect 2696 4127 2703 4193
rect 2716 4183 2723 4313
rect 2796 4243 2803 4993
rect 2816 4927 2823 4973
rect 2896 4956 2923 4963
rect 2816 4627 2823 4913
rect 2836 4667 2843 4913
rect 2916 4907 2923 4956
rect 2936 4923 2943 5133
rect 2956 5127 2963 5176
rect 2976 5007 2983 5373
rect 3016 5227 3023 5593
rect 3236 5587 3243 5603
rect 3056 5383 3063 5403
rect 3056 5376 3083 5383
rect 3076 5307 3083 5376
rect 3016 5156 3023 5173
rect 2956 4976 2983 4983
rect 2956 4947 2963 4976
rect 2936 4916 2963 4923
rect 2876 4647 2883 4683
rect 2916 4676 2923 4693
rect 2896 4647 2903 4663
rect 2956 4647 2963 4916
rect 2996 4867 3003 4943
rect 2976 4647 2983 4693
rect 3016 4667 3023 4993
rect 3036 4676 3043 4713
rect 2836 4456 2843 4633
rect 2816 4427 2823 4443
rect 2856 4407 2863 4443
rect 2796 4236 2823 4243
rect 2716 4176 2743 4183
rect 2776 4007 2783 4153
rect 2796 4087 2803 4133
rect 2696 3887 2703 3963
rect 2616 3736 2623 3773
rect 2596 3696 2623 3703
rect 2576 3516 2583 3533
rect 2616 3516 2623 3696
rect 2636 3687 2643 3723
rect 2676 3707 2683 3723
rect 2696 3687 2703 3753
rect 2716 3736 2743 3743
rect 2776 3736 2783 3753
rect 2716 3707 2723 3736
rect 2796 3707 2803 4073
rect 2716 3647 2723 3693
rect 2596 3267 2603 3503
rect 2636 3496 2643 3513
rect 2616 3256 2623 3353
rect 2656 3287 2663 3533
rect 2656 3263 2663 3273
rect 2656 3256 2683 3263
rect 2396 3027 2403 3043
rect 2436 2827 2443 3113
rect 2476 3043 2483 3173
rect 2456 3036 2483 3043
rect 2456 2947 2463 3036
rect 2596 3027 2603 3253
rect 2396 2776 2403 2793
rect 2436 2776 2443 2813
rect 2496 2807 2503 3013
rect 2416 2447 2423 2543
rect 2476 2527 2483 2543
rect 2336 2296 2343 2313
rect 2176 2247 2183 2263
rect 2116 1847 2123 1853
rect 1996 1816 2023 1823
rect 1856 1547 1863 1593
rect 1856 1147 1863 1493
rect 1876 1303 1883 1613
rect 1976 1587 1983 1633
rect 1896 1567 1903 1583
rect 1876 1296 1903 1303
rect 1876 1267 1883 1296
rect 1856 1067 1863 1103
rect 1936 887 1943 1293
rect 1956 1207 1963 1373
rect 1996 1307 2003 1753
rect 2016 1727 2023 1816
rect 2016 1247 2023 1373
rect 2036 1347 2043 1833
rect 2076 1576 2083 1833
rect 2116 1796 2123 1813
rect 2156 1807 2163 2093
rect 2096 1627 2103 1783
rect 2136 1707 2143 1763
rect 2096 1583 2103 1613
rect 2096 1576 2123 1583
rect 2136 1567 2143 1593
rect 2056 1387 2063 1563
rect 2096 1343 2103 1453
rect 2176 1387 2183 1953
rect 2196 1803 2203 2073
rect 2216 1827 2223 2263
rect 2256 2127 2263 2253
rect 2236 2063 2243 2113
rect 2316 2076 2323 2253
rect 2236 2056 2263 2063
rect 2396 2027 2403 2393
rect 2496 2307 2503 2793
rect 2576 2776 2583 2793
rect 2516 2747 2523 2763
rect 2616 2727 2623 3213
rect 2636 3007 2643 3243
rect 2676 3227 2683 3256
rect 2696 3247 2703 3293
rect 2676 3207 2683 3213
rect 2716 3207 2723 3633
rect 2736 3516 2743 3553
rect 2796 3496 2803 3593
rect 2756 3483 2763 3493
rect 2736 3476 2763 3483
rect 2736 3287 2743 3476
rect 2776 3347 2783 3353
rect 2736 3256 2743 3273
rect 2776 3256 2783 3333
rect 2816 3267 2823 4236
rect 2876 4196 2883 4213
rect 2856 4127 2863 4163
rect 2856 3996 2863 4033
rect 2896 3996 2903 4013
rect 2876 3887 2883 3983
rect 2856 3736 2863 3833
rect 2836 3507 2843 3733
rect 2876 3607 2883 3723
rect 2916 3607 2923 4513
rect 2936 4427 2943 4633
rect 2976 4476 2983 4613
rect 3056 4607 3063 4643
rect 3076 4523 3083 5293
rect 3096 4956 3103 5153
rect 3116 5147 3123 5273
rect 3156 5207 3163 5433
rect 3196 5416 3203 5433
rect 3236 5407 3243 5433
rect 3176 5387 3183 5403
rect 3216 5367 3223 5403
rect 3136 5156 3163 5163
rect 3136 5127 3143 5156
rect 3196 5123 3203 5153
rect 3176 5116 3203 5123
rect 3136 4976 3143 5113
rect 3236 4976 3243 5093
rect 3256 4987 3263 5593
rect 3336 5587 3343 5623
rect 3356 5607 3363 5893
rect 3416 5747 3423 5903
rect 3476 5767 3483 5936
rect 3796 5936 3823 5943
rect 3616 5916 3643 5923
rect 3556 5667 3563 5673
rect 3516 5636 3523 5653
rect 3556 5636 3563 5653
rect 3596 5627 3603 5733
rect 3616 5727 3623 5916
rect 3696 5887 3703 5903
rect 3816 5867 3823 5936
rect 3836 5923 3843 5933
rect 3916 5923 3923 5933
rect 3836 5916 3863 5923
rect 3896 5916 3923 5923
rect 3836 5907 3843 5916
rect 3916 5887 3923 5916
rect 3776 5667 3783 5753
rect 3796 5656 3803 5673
rect 3836 5656 3843 5693
rect 3536 5607 3543 5623
rect 3616 5587 3623 5633
rect 3296 5416 3303 5493
rect 3336 5167 3343 5573
rect 3476 5436 3483 5493
rect 3616 5467 3623 5573
rect 3456 5187 3463 5423
rect 3556 5387 3563 5433
rect 3596 5416 3603 5433
rect 3576 5307 3583 5403
rect 3616 5343 3623 5403
rect 3596 5336 3623 5343
rect 3536 5156 3543 5253
rect 3596 5143 3603 5336
rect 3696 5267 3703 5403
rect 3736 5367 3743 5403
rect 3756 5367 3763 5653
rect 3576 5136 3603 5143
rect 3576 5123 3583 5136
rect 3276 4956 3303 4963
rect 3096 4687 3103 4833
rect 3116 4667 3123 4943
rect 3156 4927 3163 4943
rect 3136 4607 3143 4683
rect 3196 4567 3203 4663
rect 3216 4527 3223 4933
rect 3256 4927 3263 4943
rect 3276 4903 3283 4913
rect 3256 4896 3283 4903
rect 3256 4667 3263 4896
rect 3296 4867 3303 4956
rect 3316 4907 3323 4953
rect 3336 4923 3343 5123
rect 3456 5116 3483 5123
rect 3556 5116 3583 5123
rect 3396 4956 3403 4973
rect 3336 4916 3363 4923
rect 3296 4703 3303 4853
rect 3356 4827 3363 4916
rect 3376 4887 3383 4943
rect 3296 4696 3323 4703
rect 3316 4676 3323 4696
rect 3276 4647 3283 4673
rect 3356 4663 3363 4813
rect 3336 4656 3363 4663
rect 3396 4663 3403 4713
rect 3396 4656 3423 4663
rect 3056 4516 3083 4523
rect 2996 4443 3003 4453
rect 2996 4436 3023 4443
rect 2936 4216 2963 4223
rect 2936 4167 2943 4216
rect 3016 4147 3023 4436
rect 3056 4087 3063 4516
rect 3087 4476 3103 4483
rect 2996 3996 3003 4033
rect 2976 3547 2983 3993
rect 3056 3667 3063 3693
rect 2976 3523 2983 3533
rect 2956 3516 2983 3523
rect 2856 3227 2863 3493
rect 2916 3236 2923 3273
rect 2756 3007 2763 3213
rect 2796 3067 2803 3133
rect 2736 2807 2743 3003
rect 2796 3003 2803 3053
rect 2876 3047 2883 3053
rect 2876 3003 2883 3033
rect 2796 2996 2823 3003
rect 2856 2996 2883 3003
rect 2896 2983 2903 3193
rect 2936 3067 2943 3213
rect 2956 3043 2963 3473
rect 2976 3187 2983 3516
rect 3036 3487 3043 3523
rect 2996 3236 3023 3243
rect 2996 3227 3003 3236
rect 2936 3036 2963 3043
rect 2936 3003 2943 3036
rect 2936 2996 2963 3003
rect 2876 2976 2903 2983
rect 2696 2776 2723 2783
rect 2416 2096 2423 2273
rect 2456 2263 2463 2293
rect 2516 2267 2523 2713
rect 2676 2707 2683 2763
rect 2716 2707 2723 2776
rect 2736 2747 2743 2773
rect 2756 2743 2763 2953
rect 2816 2776 2843 2783
rect 2756 2736 2783 2743
rect 2556 2556 2583 2563
rect 2616 2556 2643 2563
rect 2716 2556 2723 2573
rect 2736 2563 2743 2733
rect 2736 2556 2763 2563
rect 2576 2447 2583 2556
rect 2436 2243 2443 2263
rect 2456 2256 2483 2263
rect 2436 2236 2463 2243
rect 2436 2047 2443 2063
rect 2196 1796 2223 1803
rect 2276 1796 2283 2013
rect 2456 1967 2463 2236
rect 2536 2227 2543 2273
rect 2576 2263 2583 2313
rect 2596 2303 2603 2543
rect 2636 2487 2643 2556
rect 2736 2547 2743 2556
rect 2596 2296 2623 2303
rect 2556 2167 2563 2263
rect 2576 2256 2603 2263
rect 2476 1783 2483 1833
rect 2496 1787 2503 2153
rect 2556 2056 2563 2073
rect 2596 2047 2603 2073
rect 2536 1887 2543 2033
rect 2576 1947 2583 2043
rect 2616 1827 2623 2296
rect 2636 2087 2643 2353
rect 2756 2263 2763 2433
rect 2736 2256 2763 2263
rect 2776 2247 2783 2736
rect 2836 2687 2843 2776
rect 2696 2147 2703 2243
rect 2636 1807 2643 2013
rect 2676 2007 2683 2043
rect 2696 2027 2703 2133
rect 2776 2056 2783 2213
rect 2796 2207 2803 2573
rect 2816 2467 2823 2573
rect 2856 2556 2863 2573
rect 2876 2447 2883 2976
rect 2956 2927 2963 2996
rect 2956 2743 2963 2813
rect 2976 2756 2983 2773
rect 3016 2747 3023 3053
rect 3056 2967 3063 3593
rect 3076 3227 3083 4473
rect 3256 4456 3263 4493
rect 3296 4443 3303 4473
rect 3316 4447 3323 4633
rect 3356 4456 3363 4656
rect 3456 4567 3463 4663
rect 3476 4647 3483 5116
rect 3556 4956 3563 5033
rect 3636 4967 3643 5253
rect 3656 5143 3663 5213
rect 3656 5136 3683 5143
rect 3676 4967 3683 5136
rect 3716 5047 3723 5143
rect 3736 5063 3743 5353
rect 3776 5167 3783 5653
rect 3796 5403 3803 5433
rect 3916 5423 3923 5873
rect 4056 5867 4063 5933
rect 4096 5916 4103 5933
rect 4256 5916 4263 5933
rect 4416 5916 4443 5923
rect 4456 5916 4463 6056
rect 4476 6027 4483 6063
rect 4436 5887 4443 5916
rect 4696 5887 4703 5923
rect 3936 5627 3943 5693
rect 3996 5656 4023 5663
rect 3956 5456 3963 5613
rect 3976 5607 3983 5643
rect 3996 5436 4003 5453
rect 3916 5416 3943 5423
rect 3796 5396 3823 5403
rect 3936 5287 3943 5416
rect 3976 5387 3983 5423
rect 3836 5176 3863 5183
rect 3836 5107 3843 5176
rect 3996 5156 4003 5173
rect 4016 5167 4023 5656
rect 4056 5607 4063 5853
rect 4116 5603 4123 5633
rect 4296 5623 4303 5713
rect 4336 5656 4363 5663
rect 4096 5596 4123 5603
rect 4196 5507 4203 5623
rect 4296 5616 4323 5623
rect 4336 5507 4343 5656
rect 4436 5647 4443 5873
rect 4816 5767 4823 5883
rect 4496 5636 4503 5713
rect 4776 5667 4783 5753
rect 4476 5507 4483 5623
rect 4516 5607 4523 5623
rect 4136 5456 4173 5463
rect 4136 5436 4143 5456
rect 4176 5436 4193 5443
rect 4116 5416 4123 5433
rect 4196 5407 4203 5433
rect 4216 5387 4223 5453
rect 4236 5436 4243 5453
rect 4296 5436 4323 5443
rect 4236 5176 4263 5183
rect 4116 5156 4123 5173
rect 3736 5056 3763 5063
rect 3696 4956 3703 4973
rect 3516 4936 3543 4943
rect 3516 4847 3523 4936
rect 3556 4707 3563 4873
rect 3576 4807 3583 4943
rect 3596 4696 3623 4703
rect 3616 4587 3623 4696
rect 3636 4687 3643 4893
rect 3656 4627 3663 4643
rect 3756 4547 3763 5056
rect 3856 4963 3863 5093
rect 3816 4927 3823 4963
rect 3856 4956 3883 4963
rect 4016 4843 4023 5113
rect 4096 5107 4103 5123
rect 4176 4987 4183 5173
rect 4256 5127 4263 5176
rect 4296 5143 4303 5233
rect 4316 5187 4323 5436
rect 4476 5423 4483 5453
rect 4516 5427 4523 5533
rect 4536 5467 4543 5633
rect 4616 5607 4623 5623
rect 4556 5443 4563 5493
rect 4536 5436 4563 5443
rect 4596 5436 4603 5453
rect 4696 5443 4703 5653
rect 4676 5436 4703 5443
rect 4456 5416 4483 5423
rect 4336 5156 4343 5193
rect 4296 5136 4323 5143
rect 4216 4956 4223 4973
rect 4136 4936 4163 4943
rect 4136 4907 4143 4936
rect 4196 4887 4203 4943
rect 4336 4923 4343 4973
rect 4316 4916 4343 4923
rect 4016 4836 4043 4843
rect 3936 4676 3943 4693
rect 3816 4656 3843 4663
rect 3236 4427 3243 4443
rect 3276 4436 3303 4443
rect 3096 4196 3103 4213
rect 3156 4167 3163 4213
rect 3176 4187 3183 4213
rect 3216 4196 3223 4293
rect 3236 4207 3243 4413
rect 3276 4307 3283 4436
rect 3296 4187 3303 4253
rect 3116 4156 3143 4163
rect 3116 3967 3123 4003
rect 3136 3967 3143 4156
rect 3176 4163 3183 4173
rect 3176 4156 3203 4163
rect 3156 4027 3163 4153
rect 3316 4147 3323 4433
rect 3336 4267 3343 4443
rect 3336 4167 3343 4203
rect 3416 4187 3423 4213
rect 3236 4016 3243 4133
rect 3196 3996 3223 4003
rect 3196 3927 3203 3996
rect 3316 3987 3323 3993
rect 3356 3976 3363 4133
rect 3396 4047 3403 4183
rect 3196 3747 3203 3913
rect 3096 3207 3103 3593
rect 3156 3587 3163 3703
rect 3156 3543 3163 3573
rect 3136 3536 3163 3543
rect 3136 3236 3143 3536
rect 3196 3516 3203 3533
rect 3216 3447 3223 3873
rect 3256 3703 3263 3733
rect 3256 3696 3283 3703
rect 3236 3627 3243 3693
rect 3296 3523 3303 3593
rect 3276 3516 3303 3523
rect 3096 3187 3103 3193
rect 3216 3107 3223 3433
rect 3316 3407 3323 3973
rect 3396 3963 3403 4013
rect 3376 3956 3403 3963
rect 3436 3867 3443 4513
rect 3456 4496 3483 4503
rect 3456 4427 3463 4496
rect 3796 4496 3803 4553
rect 3836 4507 3843 4656
rect 3916 4647 3923 4663
rect 3676 4476 3703 4483
rect 3656 4447 3663 4463
rect 3376 3727 3383 3753
rect 3256 3227 3263 3393
rect 3356 3263 3363 3693
rect 3376 3516 3383 3713
rect 3396 3687 3403 3703
rect 3396 3487 3403 3503
rect 3436 3267 3443 3493
rect 3456 3387 3463 4393
rect 3696 4387 3703 4476
rect 3756 4476 3783 4483
rect 3756 4427 3763 4476
rect 3496 4196 3503 4213
rect 3476 4067 3483 4193
rect 3596 4167 3603 4203
rect 3476 3996 3483 4033
rect 3516 3996 3523 4053
rect 3476 3703 3483 3733
rect 3476 3696 3503 3703
rect 3556 3667 3563 3723
rect 3556 3647 3563 3653
rect 3476 3516 3503 3523
rect 3476 3507 3483 3516
rect 3516 3483 3523 3533
rect 3516 3476 3543 3483
rect 3356 3256 3383 3263
rect 3276 3127 3283 3233
rect 3336 3207 3343 3223
rect 3116 3036 3123 3053
rect 3236 3047 3243 3073
rect 2936 2736 2963 2743
rect 2916 2556 2943 2563
rect 2936 2547 2943 2556
rect 2836 2263 2843 2333
rect 2896 2307 2903 2543
rect 2956 2283 2963 2433
rect 2876 2276 2903 2283
rect 2936 2276 2963 2283
rect 2836 2256 2863 2263
rect 2896 2243 2903 2276
rect 2896 2236 2923 2243
rect 2876 2096 2883 2113
rect 2816 2043 2823 2053
rect 2576 1796 2603 1803
rect 2236 1727 2243 1783
rect 2296 1727 2303 1783
rect 2236 1707 2243 1713
rect 2256 1596 2263 1633
rect 2196 1576 2203 1593
rect 2076 1336 2103 1343
rect 1956 1116 1963 1193
rect 1976 1103 1983 1153
rect 2016 1116 2023 1233
rect 1976 1096 2003 1103
rect 1756 856 1783 863
rect 1756 807 1763 856
rect 1796 787 1803 843
rect 1796 767 1803 773
rect 1636 603 1643 673
rect 1656 647 1663 673
rect 1776 667 1783 733
rect 1816 727 1823 863
rect 1836 827 1843 843
rect 1796 656 1803 673
rect 1776 636 1783 653
rect 1816 636 1823 653
rect 1716 603 1723 633
rect 1636 596 1663 603
rect 1696 596 1723 603
rect 1076 136 1103 143
rect 1116 123 1123 133
rect 1176 123 1183 173
rect 1116 116 1183 123
rect 1236 156 1263 163
rect 1236 107 1243 156
rect 1376 147 1383 213
rect 1556 207 1563 373
rect 1576 327 1583 343
rect 1636 287 1643 363
rect 1396 156 1403 173
rect 1456 167 1463 193
rect 1556 143 1563 193
rect 1656 183 1663 373
rect 1696 327 1703 573
rect 1756 356 1763 393
rect 1636 176 1663 183
rect 1556 136 1583 143
rect 1636 27 1643 176
rect 1656 156 1683 163
rect 1716 156 1723 353
rect 1736 327 1743 343
rect 1736 247 1743 313
rect 1656 127 1663 156
rect 1736 136 1763 143
rect 1756 127 1763 136
rect 1756 107 1763 113
rect 1776 107 1783 343
rect 1796 287 1803 363
rect 1816 147 1823 313
rect 1856 283 1863 873
rect 1896 387 1903 853
rect 1916 627 1923 813
rect 1936 807 1943 813
rect 1976 707 1983 813
rect 1956 607 1963 623
rect 1956 356 1963 533
rect 1976 367 1983 593
rect 1876 323 1883 333
rect 1876 316 1903 323
rect 1836 276 1863 283
rect 1696 -24 1703 13
rect 1736 -24 1743 33
rect 1836 27 1843 276
rect 1916 267 1923 343
rect 1856 156 1863 253
rect 1936 247 1943 313
rect 1916 203 1923 233
rect 1996 223 2003 1033
rect 2016 907 2023 993
rect 2056 907 2063 1103
rect 2096 1047 2103 1336
rect 1976 216 2003 223
rect 1916 196 1933 203
rect 1876 87 1883 143
rect 1936 123 1943 173
rect 1927 116 1943 123
rect 1876 -24 1883 13
rect 1976 -17 1983 216
rect 1996 176 2003 193
rect 2016 183 2023 893
rect 2096 856 2123 863
rect 2036 687 2043 843
rect 2056 663 2063 853
rect 2116 787 2123 856
rect 2036 656 2063 663
rect 2036 427 2043 613
rect 2056 447 2063 613
rect 2036 363 2043 413
rect 2136 403 2143 1373
rect 2196 1316 2203 1333
rect 2216 1203 2223 1303
rect 2216 1196 2243 1203
rect 2156 1136 2163 1153
rect 2176 887 2183 1103
rect 2196 836 2203 853
rect 2156 647 2163 833
rect 2216 827 2223 1133
rect 2236 1047 2243 1196
rect 2296 1116 2303 1693
rect 2416 1647 2423 1783
rect 2456 1776 2483 1783
rect 2556 1747 2563 1783
rect 2596 1647 2603 1796
rect 2656 1787 2663 1813
rect 2676 1763 2683 1933
rect 2736 1816 2743 1873
rect 2756 1807 2763 2043
rect 2796 2036 2823 2043
rect 2656 1756 2683 1763
rect 2356 1616 2383 1623
rect 2376 1607 2383 1616
rect 2316 1527 2323 1593
rect 2416 1427 2423 1633
rect 2456 1616 2463 1633
rect 2476 1596 2503 1603
rect 2496 1567 2503 1596
rect 2496 1547 2503 1553
rect 2356 1287 2363 1303
rect 2276 1047 2283 1103
rect 2176 747 2183 803
rect 2236 687 2243 853
rect 2316 847 2323 893
rect 2296 787 2303 823
rect 2156 603 2163 633
rect 2236 603 2243 673
rect 2296 643 2303 773
rect 2356 747 2363 843
rect 2376 787 2383 1413
rect 2516 1227 2523 1633
rect 2556 1576 2563 1593
rect 2536 1336 2563 1343
rect 2596 1336 2623 1343
rect 2536 1307 2543 1336
rect 2536 1143 2543 1293
rect 2616 1187 2623 1336
rect 2516 1136 2543 1143
rect 2396 1083 2403 1113
rect 2396 1076 2423 1083
rect 2516 847 2523 1136
rect 2616 1127 2623 1173
rect 2636 1147 2643 1673
rect 2656 1307 2663 1756
rect 2776 1727 2783 1813
rect 2856 1807 2863 2073
rect 2896 2047 2903 2063
rect 2676 1547 2683 1573
rect 2756 1527 2763 1563
rect 2776 1503 2783 1713
rect 2756 1496 2783 1503
rect 2756 1307 2763 1496
rect 2736 1187 2743 1303
rect 2736 1167 2743 1173
rect 2636 1116 2643 1133
rect 2676 1116 2683 1133
rect 2556 1047 2563 1103
rect 2736 1087 2743 1123
rect 2776 1107 2783 1313
rect 2796 1287 2803 1793
rect 2836 1767 2843 1783
rect 2896 1576 2903 1633
rect 2916 1567 2923 2236
rect 2956 2147 2963 2276
rect 2976 2267 2983 2713
rect 2996 2707 3003 2743
rect 2996 2647 3003 2693
rect 3036 2583 3043 2913
rect 3076 2827 3083 2973
rect 3076 2763 3083 2813
rect 3016 2576 3043 2583
rect 3056 2756 3083 2763
rect 3016 2567 3023 2576
rect 3036 2467 3043 2543
rect 3056 2407 3063 2756
rect 3076 2556 3083 2573
rect 3116 2543 3123 2733
rect 3156 2687 3163 2743
rect 3176 2583 3183 3033
rect 3196 3023 3203 3033
rect 3196 3016 3223 3023
rect 3196 3007 3203 3016
rect 3236 2996 3243 3033
rect 3296 3003 3303 3193
rect 3356 3147 3363 3233
rect 3356 3087 3363 3133
rect 3376 3043 3383 3256
rect 3396 3243 3403 3253
rect 3396 3236 3423 3243
rect 3456 3236 3463 3293
rect 3356 3036 3383 3043
rect 3276 2996 3303 3003
rect 3196 2747 3203 2993
rect 3096 2536 3123 2543
rect 3156 2576 3183 2583
rect 3096 2527 3103 2536
rect 2996 2263 3003 2373
rect 3036 2276 3043 2293
rect 3096 2276 3123 2283
rect 2996 2256 3023 2263
rect 2936 1847 2943 2113
rect 2976 2076 2983 2193
rect 3036 1767 3043 2213
rect 2936 1576 2943 1613
rect 2876 1547 2883 1563
rect 2976 1387 2983 1573
rect 2996 1527 3003 1573
rect 3016 1563 3023 1633
rect 3056 1607 3063 2273
rect 3116 2267 3123 2276
rect 3136 2087 3143 2393
rect 3156 2327 3163 2576
rect 3216 2563 3223 2773
rect 3236 2587 3243 2793
rect 3276 2743 3283 2893
rect 3276 2736 3303 2743
rect 3196 2556 3223 2563
rect 3256 2556 3263 2593
rect 3176 2447 3183 2543
rect 3156 2227 3163 2263
rect 3176 2027 3183 2043
rect 3196 2007 3203 2053
rect 3216 2007 3223 2373
rect 3236 2207 3243 2543
rect 3276 2323 3283 2593
rect 3296 2567 3303 2736
rect 3336 2587 3343 3033
rect 3356 2607 3363 3036
rect 3396 3016 3403 3153
rect 3416 3047 3423 3236
rect 3496 3227 3503 3453
rect 3476 3207 3483 3223
rect 3516 3203 3523 3476
rect 3576 3467 3583 3993
rect 3596 3827 3603 4153
rect 3616 3996 3623 4073
rect 3636 4016 3643 4033
rect 3656 4027 3663 4183
rect 3776 4183 3783 4213
rect 3756 4176 3783 4183
rect 3716 3747 3723 4173
rect 3836 4167 3843 4493
rect 3856 4443 3863 4473
rect 3896 4456 3903 4593
rect 3856 4436 3883 4443
rect 3756 3963 3763 4073
rect 3796 3996 3803 4053
rect 3756 3956 3783 3963
rect 3776 3707 3783 3723
rect 3636 3647 3643 3693
rect 3696 3647 3703 3683
rect 3556 3236 3563 3253
rect 3496 3196 3523 3203
rect 3436 3047 3443 3193
rect 3496 3167 3503 3196
rect 3376 2987 3383 3003
rect 3376 2756 3383 2953
rect 3416 2867 3423 2993
rect 3436 2987 3443 3033
rect 3396 2707 3403 2723
rect 3296 2387 3303 2553
rect 3336 2327 3343 2573
rect 3396 2556 3403 2613
rect 3416 2523 3423 2753
rect 3436 2727 3443 2973
rect 3456 2763 3463 2833
rect 3516 2807 3523 3173
rect 3536 3067 3543 3223
rect 3556 3056 3583 3063
rect 3576 3007 3583 3056
rect 3596 3007 3603 3233
rect 3616 3027 3623 3253
rect 3636 3227 3643 3553
rect 3656 3487 3663 3513
rect 3676 3496 3683 3573
rect 3696 3516 3703 3613
rect 3776 3607 3783 3693
rect 3796 3647 3803 3743
rect 3836 3736 3843 3813
rect 3736 3527 3743 3533
rect 3656 3227 3663 3473
rect 3696 3243 3703 3293
rect 3696 3236 3723 3243
rect 3656 3036 3663 3113
rect 3636 3016 3643 3033
rect 3576 2776 3603 2783
rect 3636 2776 3643 2793
rect 3516 2767 3523 2773
rect 3456 2756 3483 2763
rect 3396 2516 3423 2523
rect 3256 2316 3283 2323
rect 3256 2243 3263 2316
rect 3336 2296 3363 2303
rect 3256 2236 3283 2243
rect 3276 2127 3283 2236
rect 3316 2207 3323 2283
rect 3356 2147 3363 2296
rect 3396 2283 3403 2516
rect 3376 2276 3403 2283
rect 3136 1803 3143 1933
rect 3116 1796 3143 1803
rect 3096 1587 3103 1593
rect 3016 1556 3043 1563
rect 3096 1547 3103 1573
rect 2836 1316 2843 1333
rect 2816 1287 2823 1303
rect 2796 1123 2803 1273
rect 2796 1116 2813 1123
rect 2856 1116 2863 1303
rect 2916 1227 2923 1353
rect 2956 1336 2963 1353
rect 2436 807 2443 843
rect 2476 787 2483 843
rect 2376 747 2383 773
rect 2356 727 2363 733
rect 2156 596 2183 603
rect 2216 596 2243 603
rect 2276 636 2303 643
rect 2336 636 2343 693
rect 2276 507 2283 636
rect 2356 616 2363 673
rect 2416 667 2423 773
rect 2416 627 2423 653
rect 2436 636 2443 713
rect 2496 627 2503 793
rect 2556 647 2563 1033
rect 2616 827 2623 843
rect 2136 396 2163 403
rect 2116 376 2143 383
rect 2036 356 2063 363
rect 2136 347 2143 376
rect 2016 176 2043 183
rect 1976 -24 2003 -17
rect 2036 -24 2043 176
rect 2116 156 2123 293
rect 2156 183 2163 396
rect 2176 363 2183 413
rect 2356 387 2363 433
rect 2256 376 2283 383
rect 2176 356 2203 363
rect 2276 307 2283 376
rect 2136 176 2163 183
rect 2136 47 2143 176
rect 2176 156 2183 253
rect 2416 147 2423 473
rect 2496 376 2503 393
rect 2536 387 2543 633
rect 2616 596 2623 713
rect 2656 376 2663 413
rect 2676 407 2683 853
rect 2696 827 2703 873
rect 2716 856 2743 863
rect 2716 787 2723 856
rect 2776 827 2783 863
rect 2716 627 2723 773
rect 2736 616 2743 633
rect 2776 616 2783 693
rect 2836 667 2843 1073
rect 2876 867 2883 1213
rect 2916 1007 2923 1213
rect 2936 1067 2943 1273
rect 2996 1096 3003 1133
rect 3016 1087 3023 1193
rect 3036 1096 3043 1233
rect 3056 1147 3063 1533
rect 3116 1367 3123 1796
rect 3216 1627 3223 1763
rect 3136 1527 3143 1593
rect 3176 1556 3183 1613
rect 3196 1576 3203 1593
rect 3236 1563 3243 1593
rect 3256 1567 3263 1813
rect 3276 1603 3283 1993
rect 3316 1927 3323 2043
rect 3336 1843 3343 2093
rect 3376 2047 3383 2276
rect 3396 2076 3403 2113
rect 3416 2107 3423 2313
rect 3436 2267 3443 2713
rect 3476 2276 3483 2733
rect 3496 2707 3503 2743
rect 3536 2667 3543 2743
rect 3516 2536 3523 2573
rect 3556 2523 3563 2653
rect 3576 2627 3583 2776
rect 3656 2556 3663 2793
rect 3496 2347 3503 2523
rect 3536 2516 3563 2523
rect 3676 2487 3683 2543
rect 3696 2287 3703 2993
rect 3716 2747 3723 3213
rect 3776 3067 3783 3223
rect 3796 3103 3803 3573
rect 3836 3547 3843 3593
rect 3816 3487 3823 3503
rect 3816 3227 3823 3453
rect 3836 3223 3843 3493
rect 3856 3267 3863 4436
rect 3916 4427 3923 4443
rect 3896 4047 3903 4163
rect 3956 4007 3963 4533
rect 3976 4247 3983 4573
rect 4036 4407 4043 4836
rect 4076 4483 4083 4613
rect 4116 4583 4123 4693
rect 4136 4607 4143 4663
rect 4116 4576 4143 4583
rect 4076 4476 4103 4483
rect 4136 4476 4143 4576
rect 4036 4087 4043 4183
rect 4076 4083 4083 4476
rect 4156 4467 4163 4773
rect 4336 4707 4343 4916
rect 4376 4907 4383 5163
rect 4396 5147 4403 5193
rect 4436 5147 4443 5393
rect 4476 5227 4483 5416
rect 4536 5247 4543 5436
rect 4496 5156 4503 5173
rect 4536 5167 4543 5213
rect 4576 5143 4583 5153
rect 4516 5127 4523 5143
rect 4556 5136 4583 5143
rect 4436 4936 4443 5013
rect 4216 4667 4223 4693
rect 4056 4076 4083 4083
rect 4056 4027 4063 4076
rect 4096 4063 4103 4113
rect 4076 4056 4103 4063
rect 4027 3996 4043 4003
rect 4076 3996 4083 4056
rect 3936 3947 3943 3983
rect 3896 3467 3903 3933
rect 3916 3627 3923 3683
rect 3936 3667 3943 3703
rect 4016 3687 4023 3993
rect 4056 3967 4063 3983
rect 3916 3496 3923 3573
rect 3996 3483 4003 3653
rect 4036 3567 4043 3713
rect 4056 3687 4063 3703
rect 4096 3536 4103 3613
rect 4116 3607 4123 3723
rect 4116 3516 4123 3553
rect 4136 3507 4143 3553
rect 3976 3476 4003 3483
rect 3836 3216 3863 3223
rect 3896 3207 3903 3223
rect 3796 3096 3823 3103
rect 3776 3016 3783 3053
rect 3796 3027 3803 3073
rect 3816 3027 3823 3096
rect 3796 2996 3803 3013
rect 3836 2987 3843 3003
rect 3776 2756 3783 2773
rect 3836 2747 3843 2953
rect 3856 2867 3863 3193
rect 3876 3167 3883 3203
rect 3756 2647 3763 2743
rect 3796 2627 3803 2743
rect 3716 2556 3723 2593
rect 3756 2543 3763 2613
rect 3836 2556 3843 2593
rect 3856 2587 3863 2853
rect 3916 2787 3923 3333
rect 3976 3127 3983 3223
rect 3996 3187 4003 3203
rect 3976 3107 3983 3113
rect 3956 3016 3963 3053
rect 4036 3047 4043 3233
rect 3996 3003 4003 3013
rect 3936 2967 3943 3003
rect 3976 2996 4003 3003
rect 3876 2547 3883 2773
rect 3896 2727 3903 2763
rect 3936 2756 3943 2813
rect 3956 2627 3963 2743
rect 3896 2556 3903 2573
rect 3736 2536 3763 2543
rect 3936 2543 3943 2613
rect 3976 2567 3983 2933
rect 3996 2847 4003 2996
rect 4016 2947 4023 3033
rect 3916 2536 3943 2543
rect 3936 2527 3943 2536
rect 3716 2296 3723 2333
rect 3756 2296 3783 2303
rect 3456 2187 3463 2263
rect 3436 2083 3443 2153
rect 3516 2143 3523 2263
rect 3496 2136 3523 2143
rect 3576 2256 3603 2263
rect 3416 2076 3443 2083
rect 3316 1836 3343 1843
rect 3276 1596 3303 1603
rect 3216 1556 3243 1563
rect 3276 1507 3283 1596
rect 3296 1336 3303 1393
rect 3096 1316 3103 1333
rect 3076 1167 3083 1303
rect 3156 1207 3163 1333
rect 3176 1143 3183 1333
rect 3176 1136 3203 1143
rect 2876 836 2883 853
rect 2856 747 2863 823
rect 2896 787 2903 823
rect 2796 447 2803 603
rect 2816 387 2823 653
rect 2936 627 2943 1053
rect 3056 867 3063 1083
rect 3116 843 3123 1133
rect 3196 1123 3203 1136
rect 3196 1116 3223 1123
rect 3116 836 3143 843
rect 2996 647 3003 813
rect 3076 803 3083 813
rect 3136 807 3143 836
rect 3056 796 3083 803
rect 3016 656 3023 713
rect 3156 687 3163 823
rect 3036 636 3043 673
rect 2516 327 2523 363
rect 2696 347 2703 383
rect 2736 363 2743 373
rect 2716 356 2743 363
rect 2756 327 2763 373
rect 2816 356 2823 373
rect 2896 367 2903 613
rect 3096 607 3103 673
rect 3116 603 3123 633
rect 3156 616 3163 653
rect 3216 627 3223 1116
rect 3256 847 3263 1233
rect 3296 1127 3303 1273
rect 3316 1087 3323 1836
rect 3376 1796 3383 1853
rect 3416 1787 3423 2076
rect 3456 2047 3463 2073
rect 3496 2067 3503 2136
rect 3516 1927 3523 2073
rect 3536 2047 3543 2063
rect 3576 1967 3583 2256
rect 3616 2076 3623 2113
rect 3776 2107 3783 2296
rect 3876 2276 3883 2313
rect 3956 2287 3963 2333
rect 3736 2076 3763 2083
rect 3716 2047 3723 2063
rect 3756 2027 3763 2076
rect 3516 1827 3523 1833
rect 3356 1667 3363 1783
rect 3396 1776 3413 1783
rect 3476 1647 3483 1803
rect 3516 1796 3523 1813
rect 3496 1767 3503 1783
rect 3576 1763 3583 1913
rect 3596 1787 3603 2013
rect 3756 1823 3763 1993
rect 3736 1816 3763 1823
rect 3576 1756 3603 1763
rect 3336 1596 3343 1613
rect 3376 1316 3383 1353
rect 3396 1347 3403 1573
rect 3436 1367 3443 1563
rect 3476 1467 3483 1563
rect 3556 1407 3563 1613
rect 3596 1596 3603 1756
rect 3616 1747 3623 1803
rect 3736 1787 3743 1816
rect 3776 1787 3783 1803
rect 3816 1787 3823 2053
rect 3636 1596 3643 1613
rect 3556 1336 3563 1393
rect 3356 1207 3363 1303
rect 3576 1303 3583 1333
rect 3596 1327 3603 1553
rect 3616 1447 3623 1583
rect 3656 1527 3663 1733
rect 3676 1627 3683 1773
rect 3736 1587 3743 1653
rect 3756 1607 3763 1613
rect 3716 1547 3723 1563
rect 3756 1556 3763 1593
rect 3776 1587 3783 1633
rect 3836 1327 3843 2273
rect 3976 2267 3983 2553
rect 4016 2536 4023 2753
rect 4036 2647 4043 3013
rect 4056 2967 4063 3353
rect 4096 3247 4103 3493
rect 4156 3487 4163 4393
rect 4176 3927 4183 4493
rect 4256 4227 4263 4433
rect 4276 4427 4283 4463
rect 4176 3347 4183 3693
rect 4156 3227 4163 3253
rect 4096 3036 4103 3093
rect 4136 3036 4143 3073
rect 4116 2827 4123 3023
rect 4136 2827 4143 2973
rect 4196 2847 4203 4213
rect 4256 4196 4263 4213
rect 4236 4147 4243 4163
rect 4256 4027 4263 4153
rect 4216 3996 4223 4013
rect 4236 3907 4243 3983
rect 4216 3707 4223 3723
rect 4236 3667 4243 3743
rect 4276 3736 4283 3953
rect 4296 3703 4303 4453
rect 4336 4167 4343 4473
rect 4356 4467 4363 4653
rect 4376 4487 4383 4653
rect 4416 4476 4423 4893
rect 4456 4507 4463 4683
rect 4476 4483 4483 4613
rect 4456 4476 4483 4483
rect 4436 4383 4443 4463
rect 4436 4376 4463 4383
rect 4396 4216 4403 4233
rect 4316 3987 4323 4033
rect 4327 3976 4343 3983
rect 4276 3696 4303 3703
rect 4276 3503 4283 3696
rect 4316 3627 4323 3973
rect 4356 3967 4363 4013
rect 4416 3963 4423 4133
rect 4436 4027 4443 4073
rect 4396 3956 4423 3963
rect 4436 3907 4443 4013
rect 4276 3496 4303 3503
rect 4096 2756 4103 2793
rect 4176 2776 4183 2833
rect 4216 2807 4223 3233
rect 4236 3207 4243 3223
rect 4256 3016 4263 3473
rect 4296 3447 4303 3496
rect 4236 2963 4243 3003
rect 4316 2987 4323 3033
rect 4236 2956 4263 2963
rect 4076 2687 4083 2743
rect 3896 2187 3903 2263
rect 4016 2107 4023 2263
rect 4056 2247 4063 2263
rect 3956 2076 3973 2083
rect 4036 2083 4043 2233
rect 4076 2167 4083 2633
rect 4096 2107 4103 2693
rect 4116 2627 4123 2733
rect 4136 2576 4143 2653
rect 4156 2556 4163 2613
rect 4176 2567 4183 2593
rect 4176 2527 4183 2553
rect 4236 2327 4243 2813
rect 4256 2767 4263 2956
rect 4316 2767 4323 2973
rect 4296 2667 4303 2723
rect 4256 2527 4263 2533
rect 4336 2507 4343 3833
rect 4356 3716 4363 3733
rect 4436 3703 4443 3893
rect 4416 3696 4443 3703
rect 4456 3703 4463 4376
rect 4476 4227 4483 4476
rect 4496 4023 4503 5053
rect 4516 4956 4543 4963
rect 4576 4956 4583 4993
rect 4536 4867 4543 4956
rect 4556 4827 4563 4923
rect 4596 4887 4603 5313
rect 4636 4827 4643 4953
rect 4536 4467 4543 4693
rect 4576 4676 4583 4693
rect 4656 4667 4663 5413
rect 4676 5407 4683 5436
rect 4716 5387 4723 5423
rect 4776 5387 4783 5473
rect 4836 5367 4843 5673
rect 4956 5527 4963 5623
rect 4756 5143 4763 5353
rect 4676 5067 4683 5143
rect 4756 5136 4783 5143
rect 4816 4963 4823 5143
rect 4856 4987 4863 5393
rect 4816 4956 4843 4963
rect 4856 4956 4863 4973
rect 4696 4867 4703 4943
rect 4836 4867 4843 4956
rect 4896 4927 4903 5353
rect 4976 5207 4983 5953
rect 5056 5916 5063 6063
rect 5096 5916 5123 5923
rect 5036 5616 5043 5653
rect 5056 5567 5063 5613
rect 5036 5436 5043 5513
rect 4916 5127 4923 5143
rect 4956 5087 4963 5143
rect 5056 5107 5063 5553
rect 5116 5483 5123 5916
rect 5136 5887 5143 5923
rect 5227 5916 5243 5923
rect 5196 5663 5203 5873
rect 5196 5656 5223 5663
rect 5216 5627 5223 5656
rect 5236 5527 5243 5916
rect 5416 5916 5423 6063
rect 5456 5916 5483 5923
rect 5116 5476 5143 5483
rect 5116 5407 5123 5443
rect 5136 5187 5143 5476
rect 5156 5407 5163 5453
rect 4936 4927 4943 4993
rect 4996 4956 5003 4973
rect 4976 4927 4983 4943
rect 4676 4667 4683 4673
rect 4556 4647 4563 4653
rect 4636 4627 4643 4663
rect 4556 4456 4563 4493
rect 4576 4476 4583 4493
rect 4656 4467 4663 4483
rect 4596 4387 4603 4463
rect 4716 4447 4723 4653
rect 4756 4607 4763 4663
rect 4756 4483 4763 4593
rect 4796 4567 4803 4663
rect 4736 4476 4763 4483
rect 4776 4476 4783 4493
rect 4596 4183 4603 4213
rect 4736 4187 4743 4413
rect 4496 4016 4523 4023
rect 4456 3696 4483 3703
rect 4376 3667 4383 3683
rect 4396 3516 4403 3613
rect 4376 3167 4383 3503
rect 4396 3187 4403 3233
rect 4416 3067 4423 3433
rect 4436 3207 4443 3593
rect 4456 3487 4463 3696
rect 4476 3327 4483 3633
rect 4516 3567 4523 4016
rect 4536 4007 4543 4183
rect 4576 4176 4603 4183
rect 4596 4087 4603 4176
rect 4596 3927 4603 4073
rect 4636 4067 4643 4183
rect 4696 4147 4703 4183
rect 4636 3947 4643 4053
rect 4656 3996 4663 4033
rect 4756 3987 4763 4213
rect 4536 3683 4543 3913
rect 4536 3676 4563 3683
rect 4396 2947 4403 3023
rect 4436 2787 4443 3173
rect 4496 3127 4503 3203
rect 4356 2307 4363 2753
rect 4396 2687 4403 2743
rect 4456 2647 4463 2763
rect 4436 2523 4443 2593
rect 4376 2507 4383 2523
rect 4416 2516 4443 2523
rect 4216 2296 4243 2303
rect 4196 2167 4203 2283
rect 4236 2267 4243 2296
rect 4276 2263 4283 2293
rect 4276 2256 4303 2263
rect 4347 2256 4363 2263
rect 4316 2207 4323 2243
rect 4016 2076 4043 2083
rect 3856 1776 3863 1813
rect 3916 1767 3923 2013
rect 3936 1887 3943 2063
rect 3976 2007 3983 2073
rect 4016 1907 4023 2076
rect 3916 1596 3923 1653
rect 3936 1607 3943 1783
rect 3956 1767 3963 1813
rect 3996 1627 4003 1793
rect 4036 1647 4043 2043
rect 4076 2007 4083 2043
rect 4036 1616 4043 1633
rect 3856 1567 3863 1583
rect 3876 1316 3883 1353
rect 3576 1296 3603 1303
rect 3336 1116 3343 1153
rect 3296 847 3303 1073
rect 3356 847 3363 1193
rect 3456 1107 3463 1233
rect 3576 1207 3583 1296
rect 3476 1103 3483 1193
rect 3516 1136 3523 1193
rect 3576 1116 3583 1133
rect 3616 1116 3623 1133
rect 3476 1096 3503 1103
rect 3456 856 3483 863
rect 3416 807 3423 853
rect 3436 787 3443 843
rect 3356 727 3363 753
rect 3316 636 3323 693
rect 3356 636 3363 713
rect 3116 596 3143 603
rect 3476 587 3483 856
rect 3496 623 3503 1073
rect 3536 636 3543 653
rect 3496 616 3523 623
rect 3196 427 3203 433
rect 2916 356 2923 373
rect 2836 267 2843 343
rect 2936 307 2943 313
rect 2976 307 2983 343
rect 3096 327 3103 383
rect 3176 367 3183 413
rect 3196 343 3203 413
rect 3256 376 3263 393
rect 3196 336 3223 343
rect 2336 107 2343 143
rect 2516 116 2523 173
rect 2536 136 2543 193
rect 2596 87 2603 153
rect 2636 123 2643 193
rect 2756 156 2763 213
rect 2776 176 2783 213
rect 2876 156 2883 193
rect 2916 156 2923 193
rect 2936 136 2943 273
rect 3056 207 3063 273
rect 2996 176 3023 183
rect 2996 167 3003 176
rect 3036 156 3043 193
rect 3156 167 3163 213
rect 2896 127 2903 133
rect 2636 116 2663 123
rect 3176 123 3183 173
rect 3216 156 3243 163
rect 3176 116 3203 123
rect 3236 107 3243 156
rect 3296 147 3303 553
rect 3496 463 3503 616
rect 3556 567 3563 1113
rect 3596 1087 3603 1103
rect 3636 1096 3643 1313
rect 3676 1287 3683 1303
rect 3696 867 3703 1193
rect 3816 907 3823 1313
rect 3856 1247 3863 1303
rect 3836 867 3843 1233
rect 3896 1167 3903 1303
rect 3936 1287 3943 1593
rect 3996 1583 4003 1613
rect 3996 1576 4023 1583
rect 4056 1367 4063 1893
rect 4096 1683 4103 2093
rect 4176 2076 4183 2113
rect 4296 2096 4303 2133
rect 4336 2076 4343 2113
rect 4156 2047 4163 2063
rect 4136 1807 4143 2033
rect 4276 2027 4283 2063
rect 4316 2047 4323 2053
rect 4356 1887 4363 2256
rect 4376 1827 4383 2493
rect 4476 2283 4483 3053
rect 4496 3036 4503 3073
rect 4536 3036 4543 3453
rect 4556 3187 4563 3676
rect 4576 3487 4583 3833
rect 4716 3707 4723 3853
rect 4596 3627 4603 3703
rect 4736 3703 4743 3913
rect 4736 3696 4763 3703
rect 4696 3607 4703 3693
rect 4776 3667 4783 4393
rect 4796 4147 4803 4163
rect 4836 4043 4843 4533
rect 4856 4196 4863 4373
rect 4816 4036 4843 4043
rect 4816 3723 4823 4036
rect 4876 3807 4883 4913
rect 4896 4407 4903 4873
rect 4936 4696 4963 4703
rect 4936 4587 4943 4696
rect 4956 4476 4963 4553
rect 4936 4427 4943 4463
rect 4916 3887 4923 4393
rect 4956 4107 4963 4173
rect 4956 4016 4963 4093
rect 4976 3996 4983 4053
rect 4856 3723 4863 3753
rect 4816 3716 4843 3723
rect 4856 3716 4883 3723
rect 4916 3716 4923 3733
rect 4796 3647 4803 3703
rect 4656 3516 4683 3523
rect 4696 3516 4703 3593
rect 4676 3483 4683 3516
rect 4656 3476 4683 3483
rect 4556 3016 4563 3053
rect 4576 2947 4583 3473
rect 4636 3387 4643 3433
rect 4636 3203 4643 3373
rect 4656 3207 4663 3476
rect 4736 3227 4743 3243
rect 4716 3207 4723 3223
rect 4616 3196 4643 3203
rect 4616 3023 4623 3033
rect 4676 3027 4683 3093
rect 4616 3016 4643 3023
rect 4556 2776 4563 2813
rect 4496 2747 4503 2773
rect 4556 2607 4563 2713
rect 4616 2687 4623 3016
rect 4516 2556 4523 2573
rect 4556 2556 4563 2593
rect 4536 2527 4543 2543
rect 4456 2276 4483 2283
rect 4396 2207 4403 2263
rect 4516 2227 4523 2493
rect 4636 2327 4643 2833
rect 4676 2783 4683 2953
rect 4656 2776 4683 2783
rect 4716 2776 4743 2783
rect 4396 2027 4403 2073
rect 4436 2036 4443 2133
rect 4456 2056 4463 2073
rect 4496 2047 4503 2093
rect 4516 2067 4523 2153
rect 4476 2036 4493 2043
rect 4096 1676 4123 1683
rect 4076 1587 4083 1603
rect 3996 1336 4013 1343
rect 3896 1116 3903 1133
rect 3936 1116 3943 1233
rect 3996 1227 4003 1336
rect 4056 1336 4063 1353
rect 4076 1327 4083 1513
rect 4036 1116 4043 1193
rect 4076 1116 4083 1173
rect 4116 1167 4123 1676
rect 4136 1336 4143 1393
rect 4176 1336 4203 1343
rect 4196 1287 4203 1336
rect 4196 1127 4203 1273
rect 3916 1007 3923 1103
rect 4196 987 4203 1113
rect 4216 863 4223 1813
rect 4236 1763 4243 1803
rect 4436 1787 4443 1853
rect 4476 1807 4483 1873
rect 4447 1776 4463 1783
rect 4236 1756 4263 1763
rect 4256 1327 4263 1756
rect 4356 1596 4363 1613
rect 4336 1336 4343 1553
rect 4376 1527 4383 1583
rect 4436 1567 4443 1773
rect 4256 1047 4263 1113
rect 4196 856 4223 863
rect 3696 807 3703 823
rect 3616 636 3643 643
rect 3696 636 3703 793
rect 3796 767 3803 803
rect 3616 607 3623 636
rect 3756 616 3763 673
rect 3776 647 3783 713
rect 3836 687 3843 853
rect 3936 836 3943 853
rect 3656 587 3663 603
rect 3776 596 3783 633
rect 3836 603 3843 633
rect 3856 627 3863 833
rect 3916 727 3923 803
rect 3976 707 3983 853
rect 3816 596 3843 603
rect 3476 456 3503 463
rect 3456 387 3463 393
rect 3336 363 3343 373
rect 3376 367 3383 383
rect 3416 376 3443 383
rect 3336 356 3363 363
rect 3356 227 3363 356
rect 3396 347 3403 363
rect 3316 156 3323 173
rect 3376 136 3383 193
rect 3436 187 3443 376
rect 3456 327 3463 373
rect 3476 207 3483 456
rect 3516 407 3523 473
rect 3916 447 3923 603
rect 3956 596 3963 633
rect 3976 627 3983 693
rect 4056 643 4063 823
rect 4096 647 4103 803
rect 4036 636 4063 643
rect 4036 467 4043 636
rect 4056 603 4063 613
rect 4136 603 4143 793
rect 4196 687 4203 856
rect 4236 787 4243 793
rect 4156 636 4183 643
rect 4156 627 4163 636
rect 4236 627 4243 713
rect 4056 596 4083 603
rect 4116 596 4143 603
rect 4136 427 4143 596
rect 3496 156 3503 273
rect 3476 107 3483 143
rect 3516 136 3523 393
rect 4076 376 4083 413
rect 3896 356 3923 363
rect 3596 327 3603 343
rect 3616 267 3623 353
rect 3676 247 3683 343
rect 3876 307 3883 343
rect 3816 176 3823 213
rect 3616 156 3623 173
rect 3696 127 3703 153
rect 3876 147 3883 293
rect 3916 267 3923 356
rect 3896 156 3903 253
rect 3936 156 3943 293
rect 4016 183 4023 373
rect 4056 347 4063 363
rect 4056 247 4063 333
rect 4096 227 4103 413
rect 4156 363 4163 453
rect 4176 407 4183 593
rect 4196 567 4203 623
rect 4256 547 4263 653
rect 4156 356 4183 363
rect 4216 356 4223 373
rect 4256 343 4263 433
rect 4276 347 4283 833
rect 4116 267 4123 313
rect 4196 267 4203 343
rect 4236 336 4263 343
rect 4296 307 4303 1073
rect 4316 827 4323 1103
rect 4356 967 4363 1373
rect 4416 1327 4423 1433
rect 4436 1116 4443 1133
rect 4376 1087 4383 1113
rect 4376 836 4383 853
rect 4396 807 4403 823
rect 4336 636 4343 653
rect 4376 636 4383 693
rect 4416 636 4423 933
rect 4456 887 4463 1613
rect 4516 1603 4523 1803
rect 4536 1627 4543 2293
rect 4576 2167 4583 2243
rect 4636 2207 4643 2263
rect 4636 2107 4643 2113
rect 4636 2067 4643 2093
rect 4516 1596 4543 1603
rect 4536 1576 4543 1596
rect 4556 1467 4563 1563
rect 4516 1316 4523 1353
rect 4476 1303 4483 1313
rect 4476 1296 4503 1303
rect 4536 1207 4543 1303
rect 4476 1116 4483 1173
rect 4456 867 4463 873
rect 4456 727 4463 823
rect 4476 723 4483 993
rect 4476 716 4503 723
rect 4356 607 4363 623
rect 4316 376 4323 573
rect 4436 427 4443 653
rect 4356 376 4363 413
rect 4016 176 4043 183
rect 3836 127 3843 143
rect 4116 143 4123 253
rect 4156 176 4163 213
rect 4116 136 4143 143
rect 4056 127 4063 133
rect 4276 123 4283 153
rect 4316 136 4323 333
rect 4336 327 4343 363
rect 4356 123 4363 173
rect 4396 127 4403 413
rect 4436 356 4443 373
rect 4456 367 4463 633
rect 4496 627 4503 716
rect 4516 636 4523 693
rect 4476 356 4483 413
rect 4436 176 4443 293
rect 4516 207 4523 353
rect 4416 156 4423 173
rect 4516 147 4523 193
rect 4276 116 4303 123
rect 4336 116 4363 123
rect 4536 27 4543 913
rect 4556 783 4563 1093
rect 4576 807 4583 1813
rect 4596 1027 4603 1613
rect 4656 1607 4663 2776
rect 4736 2727 4743 2776
rect 4756 2707 4763 3373
rect 4796 3067 4803 3553
rect 4836 3327 4843 3716
rect 4976 3687 4983 3873
rect 4996 3847 5003 4473
rect 5016 4407 5023 4493
rect 5036 4183 5043 4593
rect 5056 4547 5063 5093
rect 5116 4936 5123 5013
rect 5136 4956 5143 5053
rect 5176 4967 5183 5393
rect 5156 4927 5163 4943
rect 5076 4507 5083 4913
rect 5156 4587 5163 4663
rect 5156 4483 5163 4573
rect 5176 4507 5183 4673
rect 5196 4587 5203 5373
rect 5216 5127 5223 5173
rect 5236 5123 5243 5453
rect 5256 5427 5263 5653
rect 5316 5636 5323 5653
rect 5296 5607 5303 5623
rect 5276 5427 5283 5573
rect 5316 5407 5323 5423
rect 5256 5147 5263 5163
rect 5296 5156 5303 5173
rect 5276 5127 5283 5143
rect 5236 5116 5263 5123
rect 5256 4967 5263 5116
rect 5156 4476 5183 4483
rect 5016 4176 5043 4183
rect 5016 4047 5023 4176
rect 5056 4016 5063 4233
rect 5096 4227 5103 4413
rect 5096 4176 5103 4213
rect 5136 4187 5143 4473
rect 5156 4447 5163 4476
rect 5167 4416 5183 4423
rect 5156 3987 5163 4393
rect 5176 4363 5183 4416
rect 5196 4387 5203 4463
rect 5276 4407 5283 5033
rect 5296 4963 5303 5073
rect 5316 5047 5323 5143
rect 5336 5063 5343 5413
rect 5376 5187 5383 5893
rect 5396 5636 5423 5643
rect 5456 5636 5463 5693
rect 5476 5687 5483 5916
rect 5396 5487 5403 5636
rect 5496 5627 5503 5913
rect 5556 5887 5563 5903
rect 5476 5607 5483 5623
rect 5396 5367 5403 5433
rect 5416 5407 5423 5473
rect 5436 5447 5443 5553
rect 5456 5456 5463 5473
rect 5496 5443 5503 5613
rect 5516 5607 5523 5653
rect 5536 5583 5543 5633
rect 5556 5623 5563 5673
rect 5636 5663 5643 5873
rect 5636 5656 5663 5663
rect 5616 5636 5623 5653
rect 5556 5616 5603 5623
rect 5476 5436 5503 5443
rect 5496 5407 5503 5436
rect 5516 5576 5543 5583
rect 5356 5087 5363 5173
rect 5376 5107 5383 5143
rect 5336 5056 5363 5063
rect 5296 4956 5323 4963
rect 5336 4956 5343 4973
rect 5296 4607 5303 4663
rect 5316 4607 5323 4956
rect 5356 4927 5363 5056
rect 5376 4687 5383 4693
rect 5376 4656 5383 4673
rect 5296 4403 5303 4573
rect 5376 4447 5383 4473
rect 5316 4427 5323 4443
rect 5356 4436 5373 4443
rect 5296 4396 5323 4403
rect 5176 4356 5203 4363
rect 5176 4147 5183 4333
rect 4996 3683 5003 3693
rect 4996 3676 5023 3683
rect 4876 3487 4883 3503
rect 4816 3203 4823 3273
rect 4856 3247 4863 3273
rect 4816 3196 4843 3203
rect 4816 3036 4823 3093
rect 4836 3087 4843 3196
rect 4776 3016 4803 3023
rect 4776 3007 4783 3016
rect 4796 2756 4803 2793
rect 4776 2727 4783 2743
rect 4696 2263 4703 2673
rect 4716 2556 4723 2573
rect 4816 2263 4823 2293
rect 4676 2256 4703 2263
rect 4676 1827 4683 2256
rect 4756 2247 4763 2263
rect 4796 2256 4823 2263
rect 4756 2127 4763 2233
rect 4776 2227 4783 2243
rect 4796 2076 4823 2083
rect 4676 1747 4683 1783
rect 4696 1707 4703 2073
rect 4796 2067 4803 2076
rect 4556 776 4583 783
rect 4556 636 4563 693
rect 4576 307 4583 776
rect 4596 627 4603 953
rect 4616 927 4623 1593
rect 4696 1587 4703 1693
rect 4756 1596 4763 1653
rect 4836 1607 4843 2573
rect 4856 2287 4863 2993
rect 4876 2587 4883 3033
rect 4896 3007 4903 3653
rect 4936 3047 4943 3673
rect 4956 3243 4963 3533
rect 4996 3496 5003 3676
rect 5036 3487 5043 3513
rect 4976 3467 4983 3483
rect 4956 3236 4983 3243
rect 5016 3236 5023 3293
rect 5036 3207 5043 3223
rect 5056 3183 5063 3973
rect 5076 3547 5083 3983
rect 5196 3976 5203 4356
rect 5276 4196 5283 4213
rect 5216 4167 5223 4183
rect 5216 4007 5223 4153
rect 5236 4007 5243 4153
rect 5256 4147 5263 4183
rect 5176 3783 5183 3963
rect 5216 3867 5223 3963
rect 5176 3776 5203 3783
rect 5196 3767 5203 3776
rect 5196 3723 5203 3733
rect 5176 3716 5203 3723
rect 5096 3696 5123 3703
rect 5156 3696 5173 3703
rect 5096 3667 5103 3696
rect 5096 3536 5103 3653
rect 5096 3467 5103 3493
rect 5076 3223 5083 3253
rect 5116 3236 5123 3273
rect 5136 3267 5143 3533
rect 5156 3227 5163 3243
rect 5076 3216 5103 3223
rect 5136 3207 5143 3223
rect 5036 3176 5063 3183
rect 4976 3083 4983 3113
rect 4956 3076 4983 3083
rect 4956 3056 4963 3076
rect 4896 2736 4903 2853
rect 4976 2647 4983 2743
rect 4996 2587 5003 3053
rect 5036 3047 5043 3176
rect 5076 3036 5083 3053
rect 5136 3043 5143 3153
rect 5176 3087 5183 3673
rect 5196 3103 5203 3633
rect 5216 3523 5223 3813
rect 5236 3687 5243 3973
rect 5276 3827 5283 4153
rect 5296 4087 5303 4183
rect 5316 4167 5323 4396
rect 5396 4347 5403 5113
rect 5416 4867 5423 4953
rect 5416 4627 5423 4853
rect 5436 4667 5443 5133
rect 5476 5127 5483 5393
rect 5496 5067 5503 5173
rect 5516 5147 5523 5576
rect 5576 5387 5583 5403
rect 5576 5156 5583 5173
rect 5516 4887 5523 5113
rect 5476 4676 5483 4693
rect 5456 4643 5463 4663
rect 5536 4647 5543 4663
rect 5436 4636 5463 4643
rect 5416 4247 5423 4613
rect 5336 4127 5343 4213
rect 5296 3847 5303 3963
rect 5276 3727 5283 3753
rect 5256 3667 5263 3683
rect 5216 3516 5243 3523
rect 5216 3387 5223 3516
rect 5256 3387 5263 3503
rect 5296 3387 5303 3793
rect 5316 3467 5323 3753
rect 5356 3547 5363 4233
rect 5436 4087 5443 4636
rect 5456 4476 5463 4613
rect 5536 4403 5543 4613
rect 5556 4423 5563 5093
rect 5596 5087 5603 5143
rect 5616 5107 5623 5593
rect 5636 5507 5643 5623
rect 5636 5447 5643 5493
rect 5636 5047 5643 5433
rect 5636 4947 5643 4953
rect 5576 4663 5583 4693
rect 5576 4656 5603 4663
rect 5576 4443 5583 4656
rect 5636 4627 5643 4933
rect 5656 4727 5663 5656
rect 5716 5607 5723 5933
rect 5756 5916 5763 5953
rect 5796 5916 5823 5923
rect 5676 5436 5683 5453
rect 5696 5163 5703 5513
rect 5716 5436 5723 5573
rect 5696 5156 5723 5163
rect 5676 4703 5683 4943
rect 5716 4703 5723 5156
rect 5656 4696 5683 4703
rect 5696 4696 5723 4703
rect 5656 4663 5663 4696
rect 5656 4656 5683 4663
rect 5656 4607 5663 4656
rect 5576 4436 5603 4443
rect 5556 4416 5583 4423
rect 5536 4396 5563 4403
rect 5516 4183 5523 4213
rect 5536 4196 5543 4233
rect 5496 4176 5523 4183
rect 5476 4127 5483 4163
rect 5456 3996 5463 4033
rect 5376 3967 5383 3993
rect 5396 3707 5403 3743
rect 5436 3736 5443 3853
rect 5416 3687 5423 3723
rect 5396 3483 5403 3513
rect 5336 3447 5343 3483
rect 5376 3476 5403 3483
rect 5216 3127 5223 3293
rect 5256 3236 5263 3293
rect 5236 3203 5243 3223
rect 5236 3196 5263 3203
rect 5236 3187 5243 3196
rect 5196 3096 5223 3103
rect 5116 3036 5143 3043
rect 5036 2723 5043 3033
rect 5016 2716 5043 2723
rect 4876 2556 4903 2563
rect 4916 2556 4923 2573
rect 4936 2563 4943 2573
rect 4936 2556 4963 2563
rect 4876 2267 4883 2513
rect 4896 2347 4903 2556
rect 4876 2076 4883 2093
rect 4876 1796 4883 1833
rect 4896 1827 4903 2093
rect 4896 1767 4903 1783
rect 4876 1616 4903 1623
rect 4816 1576 4843 1583
rect 4636 1467 4643 1563
rect 4676 1527 4683 1563
rect 4676 1367 4683 1513
rect 4676 1336 4683 1353
rect 4636 1127 4643 1273
rect 4696 1247 4703 1313
rect 4716 1116 4723 1133
rect 4696 1027 4703 1103
rect 4736 1007 4743 1103
rect 4796 867 4803 1553
rect 4836 1547 4843 1576
rect 4876 1547 4883 1616
rect 4936 1567 4943 2273
rect 4956 2207 4963 2303
rect 4976 2076 4983 2153
rect 4996 1827 5003 2293
rect 5016 2127 5023 2716
rect 5076 2647 5083 2933
rect 5036 2587 5043 2633
rect 5036 2567 5043 2573
rect 5036 2067 5043 2313
rect 5056 2307 5063 2633
rect 5136 2547 5143 3036
rect 5096 2296 5103 2313
rect 5076 2267 5083 2283
rect 5136 2247 5143 2533
rect 5176 2347 5183 3073
rect 5216 3043 5223 3096
rect 5256 3047 5263 3196
rect 5216 3036 5243 3043
rect 5236 2747 5243 3036
rect 5316 2783 5323 3313
rect 5336 3047 5343 3393
rect 5356 3167 5363 3453
rect 5376 3407 5383 3476
rect 5416 3263 5423 3513
rect 5396 3256 5423 3263
rect 5356 3056 5363 3073
rect 5376 3036 5383 3113
rect 5316 2776 5343 2783
rect 5196 2607 5203 2743
rect 5316 2727 5323 2733
rect 5256 2563 5263 2573
rect 5336 2563 5343 2776
rect 5396 2623 5403 3256
rect 5416 3207 5423 3223
rect 5416 2787 5423 3033
rect 5436 2743 5443 3533
rect 5456 3263 5463 3593
rect 5476 3527 5483 4093
rect 5556 3767 5563 4396
rect 5556 3716 5563 3733
rect 5496 3516 5503 3533
rect 5456 3256 5483 3263
rect 5476 3223 5483 3256
rect 5456 3216 5483 3223
rect 5496 3207 5503 3373
rect 5536 3216 5543 3233
rect 5576 3227 5583 4416
rect 5616 4216 5643 4223
rect 5676 4216 5683 4233
rect 5616 4207 5623 4216
rect 5656 4167 5663 4203
rect 5676 4107 5683 4173
rect 5696 4027 5703 4696
rect 5716 4587 5723 4663
rect 5736 4483 5743 5893
rect 5816 5887 5823 5916
rect 5756 5527 5763 5623
rect 5776 4667 5783 5873
rect 5796 5567 5803 5623
rect 5936 5587 5943 5913
rect 5816 5123 5823 5423
rect 5836 5156 5863 5163
rect 5816 5116 5843 5123
rect 5816 4647 5823 4713
rect 5716 4476 5743 4483
rect 5756 4476 5763 4573
rect 5716 4027 5723 4476
rect 5736 4187 5743 4293
rect 5596 3607 5603 4013
rect 5616 3736 5643 3743
rect 5616 3407 5623 3736
rect 5656 3687 5663 3723
rect 5636 3516 5643 3533
rect 5676 3516 5683 3593
rect 5696 3507 5703 3953
rect 5716 3727 5723 3933
rect 5736 3603 5743 4153
rect 5756 4147 5763 4433
rect 5776 4307 5783 4463
rect 5776 4167 5783 4183
rect 5796 4147 5803 4163
rect 5776 4027 5783 4133
rect 5796 4027 5803 4113
rect 5756 3996 5783 4003
rect 5816 3996 5823 4153
rect 5836 4007 5843 5116
rect 5856 4947 5863 5156
rect 5856 4647 5863 4663
rect 5756 3987 5763 3996
rect 5756 3747 5763 3953
rect 5816 3767 5823 3953
rect 5776 3736 5783 3753
rect 5716 3596 5743 3603
rect 5616 3256 5643 3263
rect 5676 3256 5703 3263
rect 5456 3023 5463 3113
rect 5556 3107 5563 3173
rect 5496 3056 5523 3063
rect 5556 3056 5563 3093
rect 5516 3027 5523 3056
rect 5576 3036 5583 3113
rect 5456 3016 5483 3023
rect 5596 3023 5603 3253
rect 5616 3247 5623 3256
rect 5616 3127 5623 3233
rect 5656 3043 5663 3193
rect 5696 3187 5703 3256
rect 5656 3036 5683 3043
rect 5596 3016 5623 3023
rect 5416 2647 5423 2743
rect 5436 2736 5463 2743
rect 5396 2616 5423 2623
rect 5256 2556 5283 2563
rect 5316 2556 5343 2563
rect 5196 2307 5203 2553
rect 5016 1803 5023 2063
rect 5036 1807 5043 2053
rect 4996 1796 5023 1803
rect 5076 1763 5083 2073
rect 5056 1756 5083 1763
rect 4996 1616 5023 1623
rect 4856 1336 4883 1343
rect 4916 1336 4923 1373
rect 4856 1287 4863 1336
rect 4956 1307 4963 1373
rect 4856 1136 4883 1143
rect 4876 1123 4883 1136
rect 4936 1127 4943 1173
rect 4976 1143 4983 1593
rect 4996 1587 5003 1616
rect 5036 1596 5043 1653
rect 5056 1583 5063 1756
rect 5056 1576 5083 1583
rect 5096 1347 5103 2233
rect 5136 2096 5143 2153
rect 5156 2147 5163 2273
rect 5176 2267 5183 2283
rect 5236 2187 5243 2263
rect 5256 2187 5263 2556
rect 5336 2327 5343 2556
rect 5396 2267 5403 2593
rect 5376 2187 5383 2263
rect 5176 1823 5183 2173
rect 5236 2076 5243 2133
rect 5156 1816 5183 1823
rect 5156 1796 5163 1816
rect 5136 1407 5143 1793
rect 5156 1596 5163 1653
rect 5176 1647 5183 1783
rect 5196 1707 5203 2073
rect 5336 1987 5343 2173
rect 5376 2096 5383 2153
rect 5236 1787 5243 1813
rect 5196 1596 5203 1673
rect 5216 1576 5223 1693
rect 5016 1247 5023 1303
rect 4976 1136 5003 1143
rect 4876 1116 4903 1123
rect 4816 1103 4823 1113
rect 4996 1107 5003 1136
rect 5016 1116 5023 1133
rect 4816 1096 4843 1103
rect 4836 1087 4843 1096
rect 4616 787 4623 843
rect 4636 827 4643 863
rect 4716 827 4723 853
rect 4776 843 4783 853
rect 4747 836 4763 843
rect 4776 836 4803 843
rect 4736 803 4743 833
rect 4736 796 4763 803
rect 4656 643 4663 753
rect 4636 636 4663 643
rect 4596 347 4603 363
rect 4636 356 4643 373
rect 4616 307 4623 343
rect 4656 327 4663 333
rect 4576 176 4583 233
rect 4616 156 4643 163
rect 4596 127 4603 143
rect 4636 127 4643 156
rect 4616 -24 4623 13
rect 4676 -17 4683 673
rect 4696 656 4723 663
rect 4696 567 4703 656
rect 4756 623 4763 796
rect 4776 787 4783 803
rect 4736 616 4763 623
rect 4696 347 4703 553
rect 4796 367 4803 633
rect 4836 623 4843 853
rect 4876 683 4883 973
rect 5076 947 5083 1313
rect 5096 1067 5103 1313
rect 5156 1287 5163 1303
rect 5156 1167 5163 1193
rect 4916 836 4923 873
rect 4896 807 4903 823
rect 5036 807 5043 823
rect 5116 707 5123 1113
rect 5136 1027 5143 1133
rect 5156 1116 5163 1153
rect 5196 1116 5203 1353
rect 5216 1187 5223 1333
rect 5236 1147 5243 1333
rect 5256 1147 5263 1633
rect 5316 1596 5323 1613
rect 5336 1607 5343 1803
rect 5356 1687 5363 2093
rect 5416 1903 5423 2616
rect 5436 2387 5443 2736
rect 5616 2743 5623 2853
rect 5676 2747 5683 3013
rect 5596 2736 5623 2743
rect 5596 2587 5603 2736
rect 5636 2576 5663 2583
rect 5656 2563 5663 2576
rect 5536 2556 5563 2563
rect 5556 2547 5563 2556
rect 5656 2556 5683 2563
rect 5456 2536 5483 2543
rect 5456 2527 5463 2536
rect 5456 2256 5463 2293
rect 5396 1896 5423 1903
rect 5376 1596 5383 1613
rect 5176 1087 5183 1103
rect 5216 1087 5223 1093
rect 5136 847 5143 1013
rect 5116 687 5123 693
rect 4876 676 4903 683
rect 4896 643 4903 676
rect 4996 656 5023 663
rect 5016 643 5023 656
rect 4896 636 4923 643
rect 5016 636 5043 643
rect 4816 616 4843 623
rect 4816 403 4823 616
rect 4876 447 4883 613
rect 4916 407 4923 636
rect 4816 396 4843 403
rect 4816 347 4823 373
rect 4696 156 4703 233
rect 4836 176 4843 396
rect 4896 376 4923 383
rect 5016 376 5023 393
rect 5056 376 5063 433
rect 4856 343 4863 353
rect 4856 336 4883 343
rect 4896 327 4903 376
rect 5036 327 5043 353
rect 4876 143 4883 293
rect 5096 207 5103 673
rect 5116 636 5123 673
rect 5136 607 5143 833
rect 5156 823 5163 1053
rect 5196 836 5203 893
rect 5156 816 5183 823
rect 5176 627 5183 816
rect 5216 647 5223 823
rect 5116 343 5123 393
rect 5196 343 5203 433
rect 5116 336 5143 343
rect 5176 336 5203 343
rect 5236 287 5243 843
rect 4856 136 4883 143
rect 4976 136 4983 173
rect 5096 156 5103 173
rect 5136 156 5143 193
rect 5016 123 5023 133
rect 5216 127 5223 163
rect 5256 127 5263 1113
rect 5276 627 5283 1113
rect 5296 1047 5303 1093
rect 5296 356 5303 373
rect 5316 227 5323 1173
rect 5336 1147 5343 1393
rect 5356 1347 5363 1593
rect 5356 1307 5363 1333
rect 5356 1116 5363 1173
rect 5396 1167 5403 1896
rect 5416 1347 5423 1553
rect 5436 1387 5443 2113
rect 5456 2067 5463 2193
rect 5476 2087 5483 2373
rect 5496 2127 5503 2313
rect 5536 2263 5543 2333
rect 5576 2276 5583 2293
rect 5656 2287 5663 2556
rect 5716 2307 5723 3596
rect 5776 3523 5783 3533
rect 5756 3516 5783 3523
rect 5796 3487 5803 3693
rect 5736 3263 5743 3393
rect 5736 3256 5763 3263
rect 5736 3247 5743 3256
rect 5776 3227 5783 3243
rect 5736 3036 5763 3043
rect 5736 2867 5743 3036
rect 5776 2927 5783 3193
rect 5736 2743 5743 2773
rect 5736 2736 5763 2743
rect 5756 2556 5763 2573
rect 5536 2256 5563 2263
rect 5496 2096 5503 2113
rect 5476 1643 5483 2053
rect 5516 1807 5523 1973
rect 5516 1783 5523 1793
rect 5496 1776 5523 1783
rect 5496 1747 5503 1776
rect 5456 1636 5483 1643
rect 5456 1607 5463 1636
rect 5496 1596 5503 1673
rect 5416 1316 5423 1333
rect 5456 1316 5463 1353
rect 5436 1247 5443 1283
rect 5356 836 5363 933
rect 5376 907 5383 1103
rect 5336 767 5343 803
rect 5376 636 5383 673
rect 5416 427 5423 1133
rect 5456 1116 5463 1193
rect 5496 1116 5503 1313
rect 5516 1307 5523 1753
rect 5536 1627 5543 2256
rect 5576 1847 5583 2233
rect 5596 2107 5603 2263
rect 5616 2076 5643 2083
rect 5576 1776 5603 1783
rect 5536 1527 5543 1613
rect 5596 1607 5603 1776
rect 5616 1603 5623 2076
rect 5636 1767 5643 2033
rect 5656 1867 5663 2253
rect 5676 2247 5683 2273
rect 5696 2127 5703 2263
rect 5756 2243 5763 2283
rect 5736 2236 5763 2243
rect 5676 2067 5683 2093
rect 5696 2087 5703 2113
rect 5616 1596 5643 1603
rect 5636 1563 5643 1596
rect 5616 1556 5643 1563
rect 5556 1316 5563 1333
rect 5476 1027 5483 1103
rect 5516 1087 5523 1103
rect 5476 827 5483 843
rect 5516 836 5523 893
rect 5556 847 5563 1013
rect 5556 823 5563 833
rect 5536 816 5563 823
rect 5576 727 5583 1153
rect 5636 1143 5643 1556
rect 5656 1307 5663 1833
rect 5696 1823 5703 2073
rect 5716 1887 5723 2093
rect 5736 2087 5743 2236
rect 5756 2076 5763 2113
rect 5776 2107 5783 2293
rect 5816 2247 5823 3673
rect 5836 3503 5843 3933
rect 5856 3547 5863 4213
rect 5876 4047 5883 4643
rect 5896 4167 5903 4653
rect 5876 3687 5883 3973
rect 5836 3496 5863 3503
rect 5836 3207 5843 3473
rect 5836 2727 5843 2913
rect 5856 2243 5863 3496
rect 5836 2236 5863 2243
rect 5747 1996 5763 2003
rect 5676 1816 5703 1823
rect 5676 1687 5683 1816
rect 5716 1596 5723 1853
rect 5756 1596 5763 1996
rect 5776 1647 5783 2033
rect 5816 1947 5823 2093
rect 5836 2047 5843 2236
rect 5856 2076 5863 2113
rect 5796 1643 5803 1873
rect 5816 1803 5823 1933
rect 5816 1796 5863 1803
rect 5796 1636 5823 1643
rect 5796 1596 5803 1613
rect 5776 1567 5783 1583
rect 5616 1136 5643 1143
rect 5656 1136 5683 1143
rect 5616 1007 5623 1136
rect 5676 1123 5683 1136
rect 5676 1116 5703 1123
rect 5616 707 5623 993
rect 5696 823 5703 1093
rect 5736 1003 5743 1553
rect 5756 1083 5763 1533
rect 5776 1127 5783 1313
rect 5816 1143 5823 1636
rect 5796 1136 5823 1143
rect 5756 1076 5783 1083
rect 5676 816 5703 823
rect 5716 996 5743 1003
rect 5476 643 5483 653
rect 5456 636 5483 643
rect 5516 627 5523 693
rect 5676 687 5683 816
rect 5536 636 5563 643
rect 5416 407 5423 413
rect 5356 376 5383 383
rect 5356 367 5363 376
rect 5456 287 5463 613
rect 5536 587 5543 636
rect 5636 636 5663 643
rect 5656 627 5663 636
rect 5576 607 5583 623
rect 5536 356 5543 393
rect 5516 307 5523 323
rect 5436 156 5443 173
rect 5516 156 5523 273
rect 5576 243 5583 593
rect 5596 327 5603 573
rect 5556 236 5583 243
rect 5556 147 5563 236
rect 5616 183 5623 613
rect 5696 587 5703 713
rect 5716 667 5723 996
rect 5776 783 5783 1076
rect 5756 776 5783 783
rect 5716 347 5723 363
rect 5656 307 5663 343
rect 5696 327 5703 343
rect 5596 176 5623 183
rect 5496 127 5503 143
rect 5596 127 5603 176
rect 5656 156 5663 193
rect 5756 147 5763 776
rect 5796 643 5803 1136
rect 5836 1083 5843 1753
rect 5856 1316 5863 1796
rect 5876 1767 5883 2233
rect 5916 2107 5923 4933
rect 5896 2076 5923 2083
rect 5916 2047 5923 2076
rect 5876 1127 5883 1173
rect 5776 636 5803 643
rect 5816 1076 5843 1083
rect 5776 607 5783 636
rect 5816 627 5823 1076
rect 5796 587 5803 603
rect 5796 287 5803 353
rect 4956 87 4963 123
rect 4996 116 5023 123
rect 5796 107 5803 213
rect 5816 187 5823 323
rect 5856 167 5863 613
rect 5816 127 5823 153
rect 5836 107 5843 123
rect 4656 -24 4683 -17
<< m3contact >>
rect 2313 6013 2327 6027
rect 73 5893 87 5907
rect 1173 5933 1187 5947
rect 1673 5933 1687 5947
rect 2173 5933 2187 5947
rect 2273 5933 2287 5947
rect 213 5913 227 5927
rect 293 5913 307 5927
rect 333 5913 347 5927
rect 473 5913 487 5927
rect 513 5913 527 5927
rect 313 5893 327 5907
rect 353 5893 367 5907
rect 693 5893 707 5907
rect 833 5893 847 5907
rect 13 5873 27 5887
rect 73 5873 87 5887
rect 113 5873 127 5887
rect 193 5873 207 5887
rect 13 5833 27 5847
rect 313 5873 327 5887
rect 593 5873 607 5887
rect 673 5873 687 5887
rect 993 5913 1007 5927
rect 273 5673 287 5687
rect 233 5653 247 5667
rect 93 5633 107 5647
rect 193 5613 207 5627
rect 113 5573 127 5587
rect 153 5573 167 5587
rect 113 5473 127 5487
rect 93 5433 107 5447
rect 133 5413 147 5427
rect 73 5373 87 5387
rect 193 5433 207 5447
rect 173 5393 187 5407
rect 133 5193 147 5207
rect 93 5173 107 5187
rect 173 5193 187 5207
rect 113 5153 127 5167
rect 153 5153 167 5167
rect 133 4953 147 4967
rect 153 4933 167 4947
rect 93 4893 107 4907
rect 113 4873 127 4887
rect 93 4673 107 4687
rect 53 4493 67 4507
rect 93 4453 107 4467
rect 113 4353 127 4367
rect 13 4253 27 4267
rect 93 4213 107 4227
rect 133 4213 147 4227
rect 133 4193 147 4207
rect 113 4153 127 4167
rect 73 3973 87 3987
rect 13 3893 27 3907
rect 13 3853 27 3867
rect 253 5453 267 5467
rect 233 5433 247 5447
rect 293 5633 307 5647
rect 673 5853 687 5867
rect 813 5833 827 5847
rect 713 5793 727 5807
rect 853 5773 867 5787
rect 413 5673 427 5687
rect 613 5673 627 5687
rect 833 5673 847 5687
rect 953 5673 967 5687
rect 553 5653 567 5667
rect 453 5633 467 5647
rect 393 5613 407 5627
rect 433 5613 447 5627
rect 393 5453 407 5467
rect 433 5453 447 5467
rect 213 5413 227 5427
rect 213 5373 227 5387
rect 193 5173 207 5187
rect 333 5413 347 5427
rect 413 5413 427 5427
rect 293 5393 307 5407
rect 253 5193 267 5207
rect 253 5113 267 5127
rect 273 5073 287 5087
rect 253 4953 267 4967
rect 193 4933 207 4947
rect 213 4933 227 4947
rect 173 4913 187 4927
rect 233 4913 247 4927
rect 273 4913 287 4927
rect 373 5153 387 5167
rect 593 5473 607 5487
rect 553 5453 567 5467
rect 653 5653 667 5667
rect 673 5633 687 5647
rect 793 5653 807 5667
rect 913 5653 927 5667
rect 813 5633 827 5647
rect 673 5593 687 5607
rect 713 5593 727 5607
rect 653 5473 667 5487
rect 613 5453 627 5467
rect 453 5393 467 5407
rect 573 5413 587 5427
rect 453 5373 467 5387
rect 513 5373 527 5387
rect 433 5133 447 5147
rect 353 5113 367 5127
rect 493 5153 507 5167
rect 473 5133 487 5147
rect 393 5073 407 5087
rect 453 5073 467 5087
rect 353 4933 367 4947
rect 433 4973 447 4987
rect 453 4933 467 4947
rect 513 5073 527 5087
rect 513 4973 527 4987
rect 553 4973 567 4987
rect 693 5433 707 5447
rect 893 5433 907 5447
rect 833 5413 847 5427
rect 673 5213 687 5227
rect 633 5173 647 5187
rect 613 5153 627 5167
rect 713 5173 727 5187
rect 753 5173 767 5187
rect 853 5393 867 5407
rect 613 5113 627 5127
rect 493 4933 507 4947
rect 213 4893 227 4907
rect 293 4893 307 4907
rect 193 4873 207 4887
rect 233 4673 247 4687
rect 433 4693 447 4707
rect 473 4693 487 4707
rect 353 4673 367 4687
rect 373 4633 387 4647
rect 353 4493 367 4507
rect 193 4473 207 4487
rect 253 4473 267 4487
rect 273 4473 287 4487
rect 213 4453 227 4467
rect 193 4433 207 4447
rect 233 4433 247 4447
rect 293 4433 307 4447
rect 193 4413 207 4427
rect 273 4413 287 4427
rect 173 4193 187 4207
rect 213 4393 227 4407
rect 293 4393 307 4407
rect 293 4353 307 4367
rect 253 4213 267 4227
rect 293 4213 307 4227
rect 233 4193 247 4207
rect 253 4193 267 4207
rect 193 4173 207 4187
rect 233 4173 247 4187
rect 193 4013 207 4027
rect 213 4013 227 4027
rect 173 3973 187 3987
rect 153 3933 167 3947
rect 133 3713 147 3727
rect 73 3673 87 3687
rect 93 3593 107 3607
rect 93 3513 107 3527
rect 73 3133 87 3147
rect 113 3153 127 3167
rect 133 3113 147 3127
rect 53 3073 67 3087
rect 93 3073 107 3087
rect 293 4153 307 4167
rect 273 4113 287 4127
rect 353 4433 367 4447
rect 413 4433 427 4447
rect 373 4313 387 4327
rect 393 4213 407 4227
rect 373 4193 387 4207
rect 393 4173 407 4187
rect 373 4153 387 4167
rect 533 4913 547 4927
rect 673 5073 687 5087
rect 533 4893 547 4907
rect 613 4893 627 4907
rect 693 4893 707 4907
rect 453 4653 467 4667
rect 493 4653 507 4667
rect 593 4673 607 4687
rect 453 4493 467 4507
rect 493 4493 507 4507
rect 473 4433 487 4447
rect 533 4633 547 4647
rect 613 4653 627 4667
rect 573 4613 587 4627
rect 553 4473 567 4487
rect 693 4653 707 4667
rect 773 5153 787 5167
rect 773 5133 787 5147
rect 733 5113 747 5127
rect 733 4953 747 4967
rect 813 4953 827 4967
rect 753 4693 767 4707
rect 833 4913 847 4927
rect 773 4673 787 4687
rect 733 4653 747 4667
rect 813 4653 827 4667
rect 713 4633 727 4647
rect 753 4633 767 4647
rect 773 4633 787 4647
rect 953 5633 967 5647
rect 993 5613 1007 5627
rect 1073 5913 1087 5927
rect 1333 5893 1347 5907
rect 1433 5893 1447 5907
rect 1473 5893 1487 5907
rect 1193 5873 1207 5887
rect 1253 5873 1267 5887
rect 1193 5773 1207 5787
rect 1153 5633 1167 5647
rect 1193 5633 1207 5647
rect 1233 5633 1247 5647
rect 973 5593 987 5607
rect 1013 5593 1027 5607
rect 933 5573 947 5587
rect 973 5573 987 5587
rect 933 5433 947 5447
rect 1153 5613 1167 5627
rect 1173 5613 1187 5627
rect 1073 5453 1087 5467
rect 953 5413 967 5427
rect 913 5393 927 5407
rect 893 5213 907 5227
rect 1053 5433 1067 5447
rect 1113 5433 1127 5447
rect 1193 5573 1207 5587
rect 1033 5393 1047 5407
rect 993 5173 1007 5187
rect 1213 5413 1227 5427
rect 1173 5373 1187 5387
rect 1133 5313 1147 5327
rect 1213 5313 1227 5327
rect 873 5133 887 5147
rect 893 5113 907 5127
rect 993 5113 1007 5127
rect 913 5093 927 5107
rect 1173 5153 1187 5167
rect 1313 5853 1327 5867
rect 1333 5793 1347 5807
rect 1353 5793 1367 5807
rect 1393 5793 1407 5807
rect 1333 5633 1347 5647
rect 1313 5613 1327 5627
rect 1253 5573 1267 5587
rect 1273 5453 1287 5467
rect 1293 5393 1307 5407
rect 1353 5593 1367 5607
rect 1573 5913 1587 5927
rect 1833 5913 1847 5927
rect 1653 5893 1667 5907
rect 1513 5853 1527 5867
rect 1433 5693 1447 5707
rect 1513 5673 1527 5687
rect 1593 5673 1607 5687
rect 1433 5613 1447 5627
rect 1473 5613 1487 5627
rect 1553 5653 1567 5667
rect 1593 5633 1607 5647
rect 1633 5633 1647 5647
rect 1573 5613 1587 5627
rect 1393 5553 1407 5567
rect 1553 5553 1567 5567
rect 1413 5453 1427 5467
rect 1473 5453 1487 5467
rect 1393 5413 1407 5427
rect 1513 5413 1527 5427
rect 1853 5893 1867 5907
rect 1973 5913 1987 5927
rect 1793 5873 1807 5887
rect 1893 5873 1907 5887
rect 2093 5913 2107 5927
rect 2553 5933 2567 5947
rect 2653 5933 2667 5947
rect 2193 5893 2207 5907
rect 2453 5893 2467 5907
rect 2273 5873 2287 5887
rect 2033 5853 2047 5867
rect 1993 5693 2007 5707
rect 1873 5633 1887 5647
rect 1933 5633 1947 5647
rect 1713 5613 1727 5627
rect 1833 5613 1847 5627
rect 1733 5593 1747 5607
rect 1693 5493 1707 5507
rect 1333 5373 1347 5387
rect 1233 5173 1247 5187
rect 1233 5153 1247 5167
rect 1433 5153 1447 5167
rect 1113 5113 1127 5127
rect 1173 5113 1187 5127
rect 1013 5073 1027 5087
rect 1153 5073 1167 5087
rect 1073 4973 1087 4987
rect 993 4953 1007 4967
rect 973 4913 987 4927
rect 1113 4953 1127 4967
rect 1133 4953 1147 4967
rect 1153 4933 1167 4947
rect 913 4893 927 4907
rect 853 4773 867 4787
rect 1033 4773 1047 4787
rect 873 4673 887 4687
rect 933 4693 947 4707
rect 913 4653 927 4667
rect 1233 5093 1247 5107
rect 1313 5113 1327 5127
rect 1453 5133 1467 5147
rect 1413 5113 1427 5127
rect 1613 5173 1627 5187
rect 1673 5173 1687 5187
rect 1593 5153 1607 5167
rect 1633 5153 1647 5167
rect 1713 5153 1727 5167
rect 1553 5133 1567 5147
rect 1473 4993 1487 5007
rect 1633 4973 1647 4987
rect 1293 4953 1307 4967
rect 1333 4953 1347 4967
rect 1413 4953 1427 4967
rect 1393 4933 1407 4947
rect 1253 4913 1267 4927
rect 1273 4913 1287 4927
rect 1413 4913 1427 4927
rect 1433 4913 1447 4927
rect 1233 4853 1247 4867
rect 1073 4713 1087 4727
rect 1173 4713 1187 4727
rect 1173 4693 1187 4707
rect 1093 4673 1107 4687
rect 533 4413 547 4427
rect 513 4273 527 4287
rect 493 4213 507 4227
rect 493 4193 507 4207
rect 533 4193 547 4207
rect 473 4173 487 4187
rect 433 4133 447 4147
rect 493 4133 507 4147
rect 313 4113 327 4127
rect 413 4113 427 4127
rect 233 3973 247 3987
rect 413 3993 427 4007
rect 453 3993 467 4007
rect 473 3993 487 4007
rect 313 3973 327 3987
rect 433 3973 447 3987
rect 233 3933 247 3947
rect 293 3933 307 3947
rect 433 3933 447 3947
rect 313 3733 327 3747
rect 353 3733 367 3747
rect 393 3733 407 3747
rect 413 3733 427 3747
rect 253 3713 267 3727
rect 273 3713 287 3727
rect 233 3593 247 3607
rect 213 3573 227 3587
rect 173 3533 187 3547
rect 213 3493 227 3507
rect 193 3393 207 3407
rect 253 3573 267 3587
rect 253 3493 267 3507
rect 253 3293 267 3307
rect 233 3253 247 3267
rect 213 3213 227 3227
rect 233 3153 247 3167
rect 93 3053 107 3067
rect 153 3053 167 3067
rect 73 3013 87 3027
rect 113 3013 127 3027
rect 153 3013 167 3027
rect 53 2753 67 2767
rect 113 2753 127 2767
rect 93 2733 107 2747
rect 153 2713 167 2727
rect 93 2473 107 2487
rect 113 2353 127 2367
rect 133 2273 147 2287
rect 113 2053 127 2067
rect 93 2013 107 2027
rect 73 1973 87 1987
rect 213 3133 227 3147
rect 213 3073 227 3087
rect 373 3713 387 3727
rect 413 3673 427 3687
rect 313 3593 327 3607
rect 313 3533 327 3547
rect 353 3513 367 3527
rect 373 3493 387 3507
rect 353 3433 367 3447
rect 333 3313 347 3327
rect 293 3153 307 3167
rect 293 3133 307 3147
rect 253 3113 267 3127
rect 273 3033 287 3047
rect 233 2733 247 2747
rect 233 2573 247 2587
rect 213 2513 227 2527
rect 273 2713 287 2727
rect 193 2453 207 2467
rect 253 2453 267 2467
rect 173 2353 187 2367
rect 133 1593 147 1607
rect 33 1573 47 1587
rect 73 1573 87 1587
rect 113 1573 127 1587
rect 13 1333 27 1347
rect 113 1533 127 1547
rect 33 1313 47 1327
rect 273 2293 287 2307
rect 233 2273 247 2287
rect 233 2113 247 2127
rect 313 3113 327 3127
rect 313 3053 327 3067
rect 413 3233 427 3247
rect 393 3153 407 3167
rect 453 3793 467 3807
rect 533 4113 547 4127
rect 613 4453 627 4467
rect 593 4313 607 4327
rect 713 4473 727 4487
rect 693 4433 707 4447
rect 733 4433 747 4447
rect 693 4413 707 4427
rect 653 4253 667 4267
rect 653 4213 667 4227
rect 713 4313 727 4327
rect 613 4193 627 4207
rect 633 4193 647 4207
rect 553 4013 567 4027
rect 533 3993 547 4007
rect 573 3993 587 4007
rect 613 3993 627 4007
rect 593 3973 607 3987
rect 513 3733 527 3747
rect 473 3693 487 3707
rect 533 3713 547 3727
rect 733 4273 747 4287
rect 673 4193 687 4207
rect 713 4193 727 4207
rect 713 3993 727 4007
rect 613 3953 627 3967
rect 653 3953 667 3967
rect 513 3693 527 3707
rect 493 3653 507 3667
rect 553 3653 567 3667
rect 493 3493 507 3507
rect 453 3433 467 3447
rect 473 3433 487 3447
rect 493 3253 507 3267
rect 453 3233 467 3247
rect 473 3213 487 3227
rect 513 3213 527 3227
rect 433 3193 447 3207
rect 413 3073 427 3087
rect 373 3013 387 3027
rect 353 2753 367 2767
rect 513 3053 527 3067
rect 473 3013 487 3027
rect 433 2993 447 3007
rect 353 2733 367 2747
rect 413 2733 427 2747
rect 313 2713 327 2727
rect 373 2693 387 2707
rect 333 2533 347 2547
rect 313 2513 327 2527
rect 593 3693 607 3707
rect 693 3853 707 3867
rect 613 3653 627 3667
rect 573 3573 587 3587
rect 613 3533 627 3547
rect 673 3693 687 3707
rect 653 3673 667 3687
rect 653 3653 667 3667
rect 633 3513 647 3527
rect 613 3493 627 3507
rect 573 3273 587 3287
rect 553 3093 567 3107
rect 553 3033 567 3047
rect 593 3253 607 3267
rect 593 3233 607 3247
rect 613 3233 627 3247
rect 633 3233 647 3247
rect 613 3173 627 3187
rect 613 3153 627 3167
rect 573 2993 587 3007
rect 533 2973 547 2987
rect 633 2993 647 3007
rect 533 2953 547 2967
rect 613 2953 627 2967
rect 513 2753 527 2767
rect 453 2693 467 2707
rect 473 2613 487 2627
rect 433 2573 447 2587
rect 493 2593 507 2607
rect 513 2573 527 2587
rect 453 2533 467 2547
rect 493 2533 507 2547
rect 313 2493 327 2507
rect 473 2513 487 2527
rect 553 2713 567 2727
rect 613 2753 627 2767
rect 593 2733 607 2747
rect 573 2693 587 2707
rect 573 2673 587 2687
rect 373 2313 387 2327
rect 453 2313 467 2327
rect 333 2273 347 2287
rect 373 2273 387 2287
rect 293 2113 307 2127
rect 253 2093 267 2107
rect 213 2033 227 2047
rect 213 1773 227 1787
rect 193 1593 207 1607
rect 313 2093 327 2107
rect 393 2213 407 2227
rect 353 2193 367 2207
rect 433 2173 447 2187
rect 433 2113 447 2127
rect 393 2093 407 2107
rect 453 2093 467 2107
rect 373 2073 387 2087
rect 373 2013 387 2027
rect 293 1973 307 1987
rect 273 1573 287 1587
rect 253 1553 267 1567
rect 173 1533 187 1547
rect 173 1513 187 1527
rect 93 1313 107 1327
rect 153 1313 167 1327
rect 193 1313 207 1327
rect 73 1133 87 1147
rect 173 1133 187 1147
rect 113 1113 127 1127
rect 153 1113 167 1127
rect 53 1093 67 1107
rect 93 1093 107 1107
rect 133 1093 147 1107
rect 93 1073 107 1087
rect 33 813 47 827
rect 73 813 87 827
rect 93 813 107 827
rect 253 1093 267 1107
rect 233 1073 247 1087
rect 313 1753 327 1767
rect 353 1633 367 1647
rect 453 2053 467 2067
rect 453 1853 467 1867
rect 493 2293 507 2307
rect 493 2093 507 2107
rect 473 1833 487 1847
rect 553 2513 567 2527
rect 533 2253 547 2267
rect 553 2233 567 2247
rect 713 3633 727 3647
rect 673 3553 687 3567
rect 893 4633 907 4647
rect 853 4473 867 4487
rect 893 4453 907 4467
rect 993 4613 1007 4627
rect 1033 4513 1047 4527
rect 873 4433 887 4447
rect 913 4433 927 4447
rect 773 4393 787 4407
rect 873 4253 887 4267
rect 833 4213 847 4227
rect 853 4193 867 4207
rect 773 4153 787 4167
rect 813 4153 827 4167
rect 773 3713 787 3727
rect 793 3693 807 3707
rect 753 3673 767 3687
rect 813 3673 827 3687
rect 773 3513 787 3527
rect 1073 4453 1087 4467
rect 1053 4313 1067 4327
rect 1013 4213 1027 4227
rect 933 4193 947 4207
rect 1033 4193 1047 4207
rect 1033 4153 1047 4167
rect 973 4133 987 4147
rect 1013 3993 1027 4007
rect 1053 4073 1067 4087
rect 1053 3993 1067 4007
rect 893 3973 907 3987
rect 913 3973 927 3987
rect 953 3973 967 3987
rect 993 3973 1007 3987
rect 1033 3973 1047 3987
rect 873 3773 887 3787
rect 873 3733 887 3747
rect 833 3653 847 3667
rect 853 3573 867 3587
rect 913 3753 927 3767
rect 1013 3753 1027 3767
rect 953 3733 967 3747
rect 933 3713 947 3727
rect 933 3673 947 3687
rect 873 3533 887 3547
rect 753 3493 767 3507
rect 793 3493 807 3507
rect 773 3473 787 3487
rect 813 3473 827 3487
rect 873 3473 887 3487
rect 753 3453 767 3467
rect 693 3273 707 3287
rect 673 3213 687 3227
rect 733 3213 747 3227
rect 673 3193 687 3207
rect 713 3193 727 3207
rect 813 3253 827 3267
rect 833 3213 847 3227
rect 793 3193 807 3207
rect 773 3173 787 3187
rect 813 3173 827 3187
rect 753 3153 767 3167
rect 693 3093 707 3107
rect 673 2733 687 2747
rect 753 3033 767 3047
rect 773 3013 787 3027
rect 733 2993 747 3007
rect 693 2713 707 2727
rect 773 2753 787 2767
rect 753 2733 767 2747
rect 653 2673 667 2687
rect 733 2613 747 2627
rect 713 2593 727 2607
rect 693 2573 707 2587
rect 593 2553 607 2567
rect 653 2553 667 2567
rect 673 2513 687 2527
rect 693 2513 707 2527
rect 693 2333 707 2347
rect 613 2313 627 2327
rect 633 2273 647 2287
rect 593 2253 607 2267
rect 653 2253 667 2267
rect 573 2193 587 2207
rect 733 2533 747 2547
rect 793 2613 807 2627
rect 893 3253 907 3267
rect 873 3213 887 3227
rect 853 3133 867 3147
rect 873 3013 887 3027
rect 893 2993 907 3007
rect 853 2973 867 2987
rect 953 3573 967 3587
rect 1033 3693 1047 3707
rect 1073 3733 1087 3747
rect 1153 4653 1167 4667
rect 1213 4633 1227 4647
rect 1133 4453 1147 4467
rect 1153 4433 1167 4447
rect 1113 4393 1127 4407
rect 1153 4193 1167 4207
rect 1173 4173 1187 4187
rect 1193 4153 1207 4167
rect 1113 4133 1127 4147
rect 1153 4013 1167 4027
rect 1113 3973 1127 3987
rect 1173 3953 1187 3967
rect 1213 3993 1227 4007
rect 1113 3773 1127 3787
rect 1093 3713 1107 3727
rect 1153 3733 1167 3747
rect 1073 3633 1087 3647
rect 1053 3553 1067 3567
rect 953 3493 967 3507
rect 1033 3493 1047 3507
rect 973 3453 987 3467
rect 953 3293 967 3307
rect 973 3293 987 3307
rect 933 2993 947 3007
rect 853 2953 867 2967
rect 913 2953 927 2967
rect 833 2613 847 2627
rect 753 2473 767 2487
rect 733 2293 747 2307
rect 753 2273 767 2287
rect 793 2273 807 2287
rect 833 2273 847 2287
rect 733 2253 747 2267
rect 713 2113 727 2127
rect 593 2093 607 2107
rect 673 2093 687 2107
rect 713 2093 727 2107
rect 573 2073 587 2087
rect 613 2073 627 2087
rect 513 2053 527 2067
rect 873 2753 887 2767
rect 893 2673 907 2687
rect 913 2573 927 2587
rect 893 2513 907 2527
rect 1273 4693 1287 4707
rect 1253 4653 1267 4667
rect 1313 4673 1327 4687
rect 1353 4673 1367 4687
rect 1393 4673 1407 4687
rect 1273 4633 1287 4647
rect 1353 4633 1367 4647
rect 1353 4533 1367 4547
rect 1553 4933 1567 4947
rect 1633 4933 1647 4947
rect 1753 5553 1767 5567
rect 1793 5433 1807 5447
rect 1893 5613 1907 5627
rect 1913 5553 1927 5567
rect 2033 5593 2047 5607
rect 1953 5513 1967 5527
rect 1993 5433 2007 5447
rect 2133 5593 2147 5607
rect 1813 5413 1827 5427
rect 1873 5413 1887 5427
rect 1913 5413 1927 5427
rect 1773 5393 1787 5407
rect 1993 5333 2007 5347
rect 1773 4973 1787 4987
rect 1733 4933 1747 4947
rect 1773 4933 1787 4947
rect 1793 4933 1807 4947
rect 1533 4913 1547 4927
rect 1573 4913 1587 4927
rect 1613 4913 1627 4927
rect 1473 4873 1487 4887
rect 1453 4693 1467 4707
rect 1493 4673 1507 4687
rect 1593 4673 1607 4687
rect 1393 4453 1407 4467
rect 1613 4633 1627 4647
rect 1473 4613 1487 4627
rect 1653 4913 1667 4927
rect 1633 4573 1647 4587
rect 1733 4913 1747 4927
rect 1693 4893 1707 4907
rect 1853 5153 1867 5167
rect 1913 5153 1927 5167
rect 1873 5133 1887 5147
rect 1833 5113 1847 5127
rect 1873 4953 1887 4967
rect 1953 5133 1967 5147
rect 1993 5133 2007 5147
rect 2113 5433 2127 5447
rect 2093 5413 2107 5427
rect 2253 5613 2267 5627
rect 2173 5433 2187 5447
rect 2093 5393 2107 5407
rect 2133 5393 2147 5407
rect 2193 5393 2207 5407
rect 2393 5673 2407 5687
rect 2353 5653 2367 5667
rect 2473 5873 2487 5887
rect 2693 5913 2707 5927
rect 2833 5913 2847 5927
rect 2893 5913 2907 5927
rect 2673 5893 2687 5907
rect 2713 5893 2727 5907
rect 2433 5633 2447 5647
rect 2333 5613 2347 5627
rect 2373 5613 2387 5627
rect 2513 5653 2527 5667
rect 2573 5653 2587 5667
rect 2493 5633 2507 5647
rect 2553 5633 2567 5647
rect 2293 5573 2307 5587
rect 2373 5473 2387 5487
rect 2333 5433 2347 5447
rect 2413 5453 2427 5467
rect 2413 5433 2427 5447
rect 2273 5413 2287 5427
rect 2253 5353 2267 5367
rect 2053 5133 2067 5147
rect 2013 5113 2027 5127
rect 2113 4953 2127 4967
rect 1933 4933 1947 4947
rect 2073 4933 2087 4947
rect 1893 4913 1907 4927
rect 2053 4913 2067 4927
rect 2173 4953 2187 4967
rect 2133 4913 2147 4927
rect 2213 4913 2227 4927
rect 1893 4873 1907 4887
rect 1813 4773 1827 4787
rect 1833 4693 1847 4707
rect 1753 4653 1767 4667
rect 1773 4653 1787 4667
rect 1873 4673 1887 4687
rect 1733 4633 1747 4647
rect 1693 4613 1707 4627
rect 1713 4613 1727 4627
rect 1673 4573 1687 4587
rect 1653 4553 1667 4567
rect 1573 4513 1587 4527
rect 1533 4473 1547 4487
rect 1613 4473 1627 4487
rect 1833 4613 1847 4627
rect 1733 4473 1747 4487
rect 1793 4473 1807 4487
rect 1573 4453 1587 4467
rect 1253 4433 1267 4447
rect 1333 4433 1347 4447
rect 1373 4433 1387 4447
rect 1413 4433 1427 4447
rect 1453 4433 1467 4447
rect 1513 4433 1527 4447
rect 1553 4433 1567 4447
rect 1393 4413 1407 4427
rect 1533 4413 1547 4427
rect 1293 4333 1307 4347
rect 1373 4333 1387 4347
rect 1293 4313 1307 4327
rect 1313 4193 1327 4207
rect 1333 4173 1347 4187
rect 1313 4113 1327 4127
rect 1333 4013 1347 4027
rect 1293 3993 1307 4007
rect 1353 3973 1367 3987
rect 1333 3953 1347 3967
rect 1233 3853 1247 3867
rect 1293 3713 1307 3727
rect 1213 3693 1227 3707
rect 1193 3653 1207 3667
rect 1193 3573 1207 3587
rect 1153 3513 1167 3527
rect 1213 3513 1227 3527
rect 993 3233 1007 3247
rect 1013 3173 1027 3187
rect 1033 3173 1047 3187
rect 1053 3093 1067 3107
rect 1093 3233 1107 3247
rect 1273 3493 1287 3507
rect 1233 3433 1247 3447
rect 1193 3333 1207 3347
rect 1253 3333 1267 3347
rect 1093 3193 1107 3207
rect 1233 3233 1247 3247
rect 1153 3173 1167 3187
rect 1233 3173 1247 3187
rect 1113 3073 1127 3087
rect 1093 3053 1107 3067
rect 1073 3033 1087 3047
rect 1113 3033 1127 3047
rect 1133 3033 1147 3047
rect 1193 3033 1207 3047
rect 1273 3193 1287 3207
rect 1313 3173 1327 3187
rect 1293 3053 1307 3067
rect 1313 3053 1327 3067
rect 1253 3033 1267 3047
rect 1153 2993 1167 3007
rect 1193 2993 1207 3007
rect 1153 2813 1167 2827
rect 993 2713 1007 2727
rect 973 2693 987 2707
rect 973 2553 987 2567
rect 933 2493 947 2507
rect 1013 2673 1027 2687
rect 993 2513 1007 2527
rect 993 2473 1007 2487
rect 953 2453 967 2467
rect 893 2313 907 2327
rect 913 2313 927 2327
rect 813 2253 827 2267
rect 853 2253 867 2267
rect 773 2213 787 2227
rect 833 2113 847 2127
rect 693 2053 707 2067
rect 733 2053 747 2067
rect 673 2033 687 2047
rect 553 1853 567 1867
rect 493 1813 507 1827
rect 533 1813 547 1827
rect 473 1793 487 1807
rect 533 1773 547 1787
rect 433 1753 447 1767
rect 493 1753 507 1767
rect 393 1653 407 1667
rect 373 1613 387 1627
rect 433 1613 447 1627
rect 353 1593 367 1607
rect 413 1593 427 1607
rect 373 1573 387 1587
rect 353 1553 367 1567
rect 333 1353 347 1367
rect 333 1333 347 1347
rect 533 1593 547 1607
rect 473 1573 487 1587
rect 493 1553 507 1567
rect 353 1313 367 1327
rect 433 1313 447 1327
rect 513 1513 527 1527
rect 373 1253 387 1267
rect 413 1113 427 1127
rect 393 1093 407 1107
rect 353 1073 367 1087
rect 293 1013 307 1027
rect 273 873 287 887
rect 393 853 407 867
rect 313 833 327 847
rect 173 813 187 827
rect 353 813 367 827
rect 113 793 127 807
rect 233 673 247 687
rect 73 393 87 407
rect 33 353 47 367
rect 73 353 87 367
rect 113 353 127 367
rect 313 633 327 647
rect 373 673 387 687
rect 213 613 227 627
rect 233 613 247 627
rect 213 353 227 367
rect 133 333 147 347
rect 173 333 187 347
rect 113 313 127 327
rect 93 293 107 307
rect 93 233 107 247
rect 513 1093 527 1107
rect 493 1073 507 1087
rect 533 893 547 907
rect 613 1833 627 1847
rect 573 1793 587 1807
rect 633 1773 647 1787
rect 693 1813 707 1827
rect 793 1813 807 1827
rect 813 1793 827 1807
rect 673 1753 687 1767
rect 593 1733 607 1747
rect 653 1653 667 1667
rect 613 1633 627 1647
rect 633 1613 647 1627
rect 913 2273 927 2287
rect 893 2093 907 2107
rect 873 2073 887 2087
rect 953 2233 967 2247
rect 1133 2753 1147 2767
rect 1173 2613 1187 2627
rect 1093 2573 1107 2587
rect 1113 2473 1127 2487
rect 1133 2333 1147 2347
rect 1033 2293 1047 2307
rect 1133 2293 1147 2307
rect 1093 2273 1107 2287
rect 1073 2253 1087 2267
rect 1173 2293 1187 2307
rect 1013 2213 1027 2227
rect 1153 2213 1167 2227
rect 993 2173 1007 2187
rect 993 2113 1007 2127
rect 1113 2093 1127 2107
rect 913 2053 927 2067
rect 853 2033 867 2047
rect 893 2013 907 2027
rect 973 2053 987 2067
rect 1013 2053 1027 2067
rect 933 1993 947 2007
rect 893 1833 907 1847
rect 933 1833 947 1847
rect 853 1813 867 1827
rect 893 1793 907 1807
rect 753 1753 767 1767
rect 813 1753 827 1767
rect 833 1753 847 1767
rect 873 1733 887 1747
rect 733 1633 747 1647
rect 753 1633 767 1647
rect 913 1633 927 1647
rect 713 1613 727 1627
rect 593 1553 607 1567
rect 813 1613 827 1627
rect 933 1613 947 1627
rect 713 1533 727 1547
rect 573 1293 587 1307
rect 613 1253 627 1267
rect 693 1253 707 1267
rect 633 1173 647 1187
rect 573 1153 587 1167
rect 593 1153 607 1167
rect 473 853 487 867
rect 513 853 527 867
rect 553 853 567 867
rect 453 833 467 847
rect 413 633 427 647
rect 653 1113 667 1127
rect 713 1133 727 1147
rect 673 1093 687 1107
rect 773 1573 787 1587
rect 753 1553 767 1567
rect 833 1593 847 1607
rect 893 1593 907 1607
rect 793 1513 807 1527
rect 753 1333 767 1347
rect 873 1573 887 1587
rect 913 1573 927 1587
rect 993 1993 1007 2007
rect 993 1813 1007 1827
rect 1033 1793 1047 1807
rect 1133 2073 1147 2087
rect 1213 2813 1227 2827
rect 1453 4193 1467 4207
rect 1493 4193 1507 4207
rect 1413 4173 1427 4187
rect 1393 4133 1407 4147
rect 1493 4173 1507 4187
rect 1473 4133 1487 4147
rect 1513 4113 1527 4127
rect 1433 4073 1447 4087
rect 1493 4073 1507 4087
rect 1453 3993 1467 4007
rect 1433 3973 1447 3987
rect 1393 3953 1407 3967
rect 1433 3893 1447 3907
rect 1393 3733 1407 3747
rect 1413 3713 1427 3727
rect 1373 3673 1387 3687
rect 1633 4453 1647 4467
rect 1613 4213 1627 4227
rect 1573 4173 1587 4187
rect 1533 3993 1547 4007
rect 1553 3993 1567 4007
rect 1633 4153 1647 4167
rect 1593 4113 1607 4127
rect 1633 4013 1647 4027
rect 1613 3993 1627 4007
rect 1513 3973 1527 3987
rect 1593 3973 1607 3987
rect 1553 3813 1567 3827
rect 1773 4213 1787 4227
rect 1733 4193 1747 4207
rect 1753 4193 1767 4207
rect 1713 4153 1727 4167
rect 1753 4013 1767 4027
rect 1693 3993 1707 4007
rect 1673 3933 1687 3947
rect 1733 3993 1747 4007
rect 1713 3913 1727 3927
rect 1733 3873 1747 3887
rect 1633 3773 1647 3787
rect 1553 3733 1567 3747
rect 1513 3713 1527 3727
rect 1673 3713 1687 3727
rect 1493 3573 1507 3587
rect 1453 3533 1467 3547
rect 1573 3693 1587 3707
rect 1573 3673 1587 3687
rect 1653 3673 1667 3687
rect 1653 3613 1667 3627
rect 1553 3573 1567 3587
rect 1593 3553 1607 3567
rect 1393 3493 1407 3507
rect 1373 3433 1387 3447
rect 1353 3333 1367 3347
rect 1353 3073 1367 3087
rect 1233 2753 1247 2767
rect 1253 2733 1267 2747
rect 1213 2713 1227 2727
rect 1293 2713 1307 2727
rect 1273 2553 1287 2567
rect 1253 2533 1267 2547
rect 1293 2533 1307 2547
rect 1213 2413 1227 2427
rect 1233 2273 1247 2287
rect 1333 2773 1347 2787
rect 1333 2673 1347 2687
rect 1413 3393 1427 3407
rect 1513 3333 1527 3347
rect 1453 3233 1467 3247
rect 1493 3233 1507 3247
rect 1673 3533 1687 3547
rect 1433 3173 1447 3187
rect 1393 3053 1407 3067
rect 1593 3053 1607 3067
rect 1373 3013 1387 3027
rect 1413 3013 1427 3027
rect 1453 3013 1467 3027
rect 1553 3013 1567 3027
rect 1413 2993 1427 3007
rect 1573 2993 1587 3007
rect 1533 2973 1547 2987
rect 1373 2773 1387 2787
rect 1393 2753 1407 2767
rect 1453 2773 1467 2787
rect 1433 2713 1447 2727
rect 1433 2613 1447 2627
rect 1393 2533 1407 2547
rect 1353 2513 1367 2527
rect 1353 2473 1367 2487
rect 1313 2253 1327 2267
rect 1413 2513 1427 2527
rect 1553 2773 1567 2787
rect 1493 2733 1507 2747
rect 1533 2673 1547 2687
rect 1473 2553 1487 2567
rect 1493 2553 1507 2567
rect 1533 2553 1547 2567
rect 1633 2993 1647 3007
rect 1453 2473 1467 2487
rect 1413 2453 1427 2467
rect 1373 2413 1387 2427
rect 1193 2213 1207 2227
rect 1313 2193 1327 2207
rect 1173 2133 1187 2147
rect 1313 2133 1327 2147
rect 1193 2073 1207 2087
rect 1253 2073 1267 2087
rect 1293 2033 1307 2047
rect 1253 2013 1267 2027
rect 1173 1933 1187 1947
rect 1153 1833 1167 1847
rect 1013 1753 1027 1767
rect 1113 1773 1127 1787
rect 1433 2413 1447 2427
rect 1433 2273 1447 2287
rect 1453 2213 1467 2227
rect 1413 2073 1427 2087
rect 1413 2053 1427 2067
rect 1393 2033 1407 2047
rect 1373 1953 1387 1967
rect 1293 1813 1307 1827
rect 1313 1813 1327 1827
rect 1173 1773 1187 1787
rect 1153 1753 1167 1767
rect 993 1613 1007 1627
rect 1113 1613 1127 1627
rect 993 1593 1007 1607
rect 1033 1593 1047 1607
rect 813 1313 827 1327
rect 953 1333 967 1347
rect 973 1333 987 1347
rect 913 1313 927 1327
rect 933 1293 947 1307
rect 853 1273 867 1287
rect 973 1273 987 1287
rect 1253 1793 1267 1807
rect 1233 1753 1247 1767
rect 1213 1673 1227 1687
rect 1273 1653 1287 1667
rect 1273 1613 1287 1627
rect 1093 1393 1107 1407
rect 1173 1573 1187 1587
rect 1353 1773 1367 1787
rect 1513 2413 1527 2427
rect 1573 2373 1587 2387
rect 1493 2333 1507 2347
rect 1533 2313 1547 2327
rect 1533 2273 1547 2287
rect 1513 2253 1527 2267
rect 1513 2073 1527 2087
rect 1493 2053 1507 2067
rect 1473 1813 1487 1827
rect 1553 2053 1567 2067
rect 1553 2013 1567 2027
rect 1493 1793 1507 1807
rect 1593 2013 1607 2027
rect 1573 1993 1587 2007
rect 1733 3633 1747 3647
rect 1813 4453 1827 4467
rect 1853 4433 1867 4447
rect 2353 5393 2367 5407
rect 2313 5373 2327 5387
rect 2453 5493 2467 5507
rect 2533 5473 2547 5487
rect 2493 5433 2507 5447
rect 2553 5453 2567 5467
rect 2433 5393 2447 5407
rect 2513 5413 2527 5427
rect 2553 5413 2567 5427
rect 2493 5393 2507 5407
rect 2473 5373 2487 5387
rect 2313 5353 2327 5367
rect 2413 5353 2427 5367
rect 2273 4953 2287 4967
rect 2273 4933 2287 4947
rect 2333 5173 2347 5187
rect 2853 5633 2867 5647
rect 2633 5613 2647 5627
rect 2753 5613 2767 5627
rect 2813 5613 2827 5627
rect 2673 5593 2687 5607
rect 3233 5913 3247 5927
rect 3313 5913 3327 5927
rect 3373 5913 3387 5927
rect 3053 5893 3067 5907
rect 3213 5893 3227 5907
rect 3353 5893 3367 5907
rect 2953 5873 2967 5887
rect 3033 5873 3047 5887
rect 3073 5873 3087 5887
rect 3213 5873 3227 5887
rect 3033 5693 3047 5707
rect 3213 5673 3227 5687
rect 3173 5653 3187 5667
rect 2953 5613 2967 5627
rect 2893 5593 2907 5607
rect 2633 5533 2647 5547
rect 2613 5453 2627 5467
rect 2793 5513 2807 5527
rect 2673 5453 2687 5467
rect 2713 5453 2727 5467
rect 2853 5493 2867 5507
rect 2653 5353 2667 5367
rect 2613 5333 2627 5347
rect 2833 5433 2847 5447
rect 2713 5373 2727 5387
rect 2813 5413 2827 5427
rect 2693 5313 2707 5327
rect 2773 5313 2787 5327
rect 2653 5173 2667 5187
rect 2713 5173 2727 5187
rect 2613 5153 2627 5167
rect 2693 5153 2707 5167
rect 2573 5133 2587 5147
rect 2633 5133 2647 5147
rect 2493 5113 2507 5127
rect 2393 5053 2407 5067
rect 2413 5053 2427 5067
rect 2393 4953 2407 4967
rect 2453 4953 2467 4967
rect 2333 4913 2347 4927
rect 2253 4853 2267 4867
rect 2273 4713 2287 4727
rect 2293 4713 2307 4727
rect 1973 4693 1987 4707
rect 2073 4693 2087 4707
rect 2193 4693 2207 4707
rect 1933 4673 1947 4687
rect 2133 4653 2147 4667
rect 2113 4633 2127 4647
rect 2053 4613 2067 4627
rect 1913 4553 1927 4567
rect 1893 4313 1907 4327
rect 2013 4533 2027 4547
rect 1973 4453 1987 4467
rect 1993 4433 2007 4447
rect 1993 4413 2007 4427
rect 1933 4393 1947 4407
rect 1893 4193 1907 4207
rect 1873 4173 1887 4187
rect 1853 4153 1867 4167
rect 1853 3993 1867 4007
rect 1793 3873 1807 3887
rect 1833 3733 1847 3747
rect 1793 3713 1807 3727
rect 1813 3713 1827 3727
rect 1773 3673 1787 3687
rect 1753 3533 1767 3547
rect 1693 3513 1707 3527
rect 1733 3493 1747 3507
rect 1893 3973 1907 3987
rect 1873 3953 1887 3967
rect 1953 4153 1967 4167
rect 1933 3893 1947 3907
rect 1893 3833 1907 3847
rect 1873 3773 1887 3787
rect 1873 3713 1887 3727
rect 1853 3653 1867 3667
rect 1853 3633 1867 3647
rect 1813 3513 1827 3527
rect 1873 3513 1887 3527
rect 1793 3493 1807 3507
rect 1833 3493 1847 3507
rect 1773 3473 1787 3487
rect 1693 3333 1707 3347
rect 1733 3233 1747 3247
rect 2113 4473 2127 4487
rect 2173 4613 2187 4627
rect 2253 4493 2267 4507
rect 2033 4153 2047 4167
rect 2053 4153 2067 4167
rect 2153 4073 2167 4087
rect 2313 4673 2327 4687
rect 2353 4673 2367 4687
rect 2293 4653 2307 4667
rect 2333 4653 2347 4667
rect 2353 4633 2367 4647
rect 2313 4613 2327 4627
rect 2273 4153 2287 4167
rect 2013 4053 2027 4067
rect 2193 4053 2207 4067
rect 1993 4013 2007 4027
rect 1993 3993 2007 4007
rect 2053 3993 2067 4007
rect 1993 3973 2007 3987
rect 2133 3973 2147 3987
rect 1973 3953 1987 3967
rect 2033 3953 2047 3967
rect 2153 3953 2167 3967
rect 1973 3933 1987 3947
rect 1953 3753 1967 3767
rect 1933 3733 1947 3747
rect 2033 3753 2047 3767
rect 2013 3733 2027 3747
rect 1953 3713 1967 3727
rect 1953 3653 1967 3667
rect 1933 3553 1947 3567
rect 1913 3413 1927 3427
rect 1893 3393 1907 3407
rect 1873 3273 1887 3287
rect 1913 3273 1927 3287
rect 1933 3273 1947 3287
rect 1913 3233 1927 3247
rect 1793 3213 1807 3227
rect 1853 3213 1867 3227
rect 1753 3193 1767 3207
rect 1753 3073 1767 3087
rect 1813 3193 1827 3207
rect 1693 2813 1707 2827
rect 1673 2773 1687 2787
rect 1653 2753 1667 2767
rect 1673 2733 1687 2747
rect 1713 2733 1727 2747
rect 1713 2713 1727 2727
rect 1693 2573 1707 2587
rect 1713 2513 1727 2527
rect 1833 3093 1847 3107
rect 1893 3053 1907 3067
rect 1893 3033 1907 3047
rect 1873 2953 1887 2967
rect 1853 2893 1867 2907
rect 1813 2793 1827 2807
rect 1753 2773 1767 2787
rect 1793 2773 1807 2787
rect 1833 2773 1847 2787
rect 1793 2753 1807 2767
rect 1773 2733 1787 2747
rect 1753 2713 1767 2727
rect 1753 2553 1767 2567
rect 1793 2693 1807 2707
rect 1873 2733 1887 2747
rect 1853 2713 1867 2727
rect 1813 2673 1827 2687
rect 1833 2593 1847 2607
rect 1813 2553 1827 2567
rect 1873 2553 1887 2567
rect 1753 2513 1767 2527
rect 1773 2513 1787 2527
rect 1673 2473 1687 2487
rect 1673 2293 1687 2307
rect 1853 2513 1867 2527
rect 1793 2413 1807 2427
rect 1733 2313 1747 2327
rect 1733 2293 1747 2307
rect 1753 2273 1767 2287
rect 1793 2213 1807 2227
rect 1853 2213 1867 2227
rect 1713 2153 1727 2167
rect 1633 2133 1647 2147
rect 1653 2073 1667 2087
rect 1773 2133 1787 2147
rect 1753 2093 1767 2107
rect 1633 2053 1647 2067
rect 1633 1993 1647 2007
rect 1673 1993 1687 2007
rect 1573 1973 1587 1987
rect 1613 1973 1627 1987
rect 1633 1833 1647 1847
rect 1593 1793 1607 1807
rect 1453 1753 1467 1767
rect 1433 1713 1447 1727
rect 1353 1693 1367 1707
rect 1353 1673 1367 1687
rect 1313 1553 1327 1567
rect 1453 1633 1467 1647
rect 1393 1573 1407 1587
rect 1433 1573 1447 1587
rect 1253 1533 1267 1547
rect 1313 1533 1327 1547
rect 1213 1333 1227 1347
rect 1253 1333 1267 1347
rect 1133 1313 1147 1327
rect 1193 1313 1207 1327
rect 1233 1313 1247 1327
rect 1053 1293 1067 1307
rect 1033 1253 1047 1267
rect 1053 1173 1067 1187
rect 933 1153 947 1167
rect 753 1133 767 1147
rect 893 1113 907 1127
rect 1113 1253 1127 1267
rect 1173 1253 1187 1267
rect 733 1093 747 1107
rect 773 1073 787 1087
rect 633 833 647 847
rect 553 813 567 827
rect 593 813 607 827
rect 1013 1053 1027 1067
rect 833 1013 847 1027
rect 973 893 987 907
rect 833 853 847 867
rect 1013 853 1027 867
rect 653 813 667 827
rect 733 813 747 827
rect 773 813 787 827
rect 873 833 887 847
rect 993 833 1007 847
rect 593 793 607 807
rect 653 693 667 707
rect 613 673 627 687
rect 493 633 507 647
rect 613 633 627 647
rect 493 613 507 627
rect 533 613 547 627
rect 733 613 747 627
rect 513 593 527 607
rect 253 553 267 567
rect 333 553 347 567
rect 533 553 547 567
rect 413 393 427 407
rect 353 353 367 367
rect 753 593 767 607
rect 733 413 747 427
rect 453 353 467 367
rect 293 233 307 247
rect 133 153 147 167
rect 473 333 487 347
rect 713 373 727 387
rect 593 353 607 367
rect 673 333 687 347
rect 513 313 527 327
rect 353 233 367 247
rect 393 233 407 247
rect 573 233 587 247
rect 333 213 347 227
rect 213 133 227 147
rect 313 133 327 147
rect 493 213 507 227
rect 453 193 467 207
rect 533 153 547 167
rect 633 153 647 167
rect 673 153 687 167
rect 373 133 387 147
rect 453 133 467 147
rect 513 133 527 147
rect 573 133 587 147
rect 693 133 707 147
rect 853 813 867 827
rect 1033 753 1047 767
rect 853 733 867 747
rect 813 713 827 727
rect 793 673 807 687
rect 813 653 827 667
rect 953 713 967 727
rect 873 673 887 687
rect 833 633 847 647
rect 853 633 867 647
rect 913 633 927 647
rect 813 593 827 607
rect 793 413 807 427
rect 893 613 907 627
rect 873 593 887 607
rect 793 393 807 407
rect 833 393 847 407
rect 833 353 847 367
rect 933 373 947 387
rect 813 233 827 247
rect 793 213 807 227
rect 773 133 787 147
rect 653 113 667 127
rect 713 113 727 127
rect 893 333 907 347
rect 933 313 947 327
rect 853 213 867 227
rect 833 193 847 207
rect 913 173 927 187
rect 993 673 1007 687
rect 1013 653 1027 667
rect 993 633 1007 647
rect 1033 633 1047 647
rect 1133 1113 1147 1127
rect 1073 1093 1087 1107
rect 1113 1093 1127 1107
rect 1093 1033 1107 1047
rect 1133 1013 1147 1027
rect 1153 1013 1167 1027
rect 1093 873 1107 887
rect 1193 873 1207 887
rect 1133 853 1147 867
rect 1073 833 1087 847
rect 1113 833 1127 847
rect 1193 833 1207 847
rect 1153 673 1167 687
rect 1233 1293 1247 1307
rect 1413 1513 1427 1527
rect 1413 1493 1427 1507
rect 1353 1313 1367 1327
rect 1333 1113 1347 1127
rect 1433 1333 1447 1347
rect 1513 1773 1527 1787
rect 1573 1773 1587 1787
rect 1473 1613 1487 1627
rect 1573 1613 1587 1627
rect 1493 1593 1507 1607
rect 1533 1593 1547 1607
rect 1713 2033 1727 2047
rect 1713 1933 1727 1947
rect 1693 1753 1707 1767
rect 1633 1633 1647 1647
rect 1673 1593 1687 1607
rect 1513 1573 1527 1587
rect 1553 1573 1567 1587
rect 1593 1573 1607 1587
rect 1613 1573 1627 1587
rect 1653 1573 1667 1587
rect 1693 1573 1707 1587
rect 1573 1513 1587 1527
rect 1493 1373 1507 1387
rect 1493 1313 1507 1327
rect 1813 2073 1827 2087
rect 1873 2053 1887 2067
rect 1833 2033 1847 2047
rect 1853 2033 1867 2047
rect 1773 1833 1787 1847
rect 1853 1813 1867 1827
rect 1773 1773 1787 1787
rect 1773 1753 1787 1767
rect 1773 1733 1787 1747
rect 1753 1713 1767 1727
rect 1733 1633 1747 1647
rect 1733 1513 1747 1527
rect 1713 1493 1727 1507
rect 1613 1393 1627 1407
rect 1833 1713 1847 1727
rect 1813 1633 1827 1647
rect 1793 1573 1807 1587
rect 1653 1313 1667 1327
rect 1753 1313 1767 1327
rect 1433 1273 1447 1287
rect 1453 1113 1467 1127
rect 1293 1093 1307 1107
rect 1273 1073 1287 1087
rect 1393 1093 1407 1107
rect 1433 1073 1447 1087
rect 1453 1073 1467 1087
rect 1433 1053 1447 1067
rect 1253 853 1267 867
rect 1293 853 1307 867
rect 1253 833 1267 847
rect 1273 833 1287 847
rect 1233 773 1247 787
rect 1273 713 1287 727
rect 1153 653 1167 667
rect 1213 653 1227 667
rect 1253 633 1267 647
rect 1373 833 1387 847
rect 1393 813 1407 827
rect 1313 753 1327 767
rect 1433 793 1447 807
rect 1353 733 1367 747
rect 1413 613 1427 627
rect 1133 593 1147 607
rect 973 373 987 387
rect 1013 373 1027 387
rect 973 213 987 227
rect 953 153 967 167
rect 1053 493 1067 507
rect 1093 373 1107 387
rect 1053 333 1067 347
rect 1073 313 1087 327
rect 1133 333 1147 347
rect 1093 293 1107 307
rect 1033 233 1047 247
rect 1073 213 1087 227
rect 853 113 867 127
rect 913 113 927 127
rect 953 113 967 127
rect 993 113 1007 127
rect 1273 593 1287 607
rect 1393 593 1407 607
rect 1453 773 1467 787
rect 1573 1273 1587 1287
rect 1633 1153 1647 1167
rect 1613 1133 1627 1147
rect 1713 1133 1727 1147
rect 1593 1113 1607 1127
rect 1553 1093 1567 1107
rect 1533 1073 1547 1087
rect 1493 873 1507 887
rect 1553 833 1567 847
rect 1473 653 1487 667
rect 1573 813 1587 827
rect 1553 593 1567 607
rect 1253 353 1267 367
rect 1333 313 1347 327
rect 1273 293 1287 307
rect 1533 393 1547 407
rect 1433 353 1447 367
rect 1473 353 1487 367
rect 1513 353 1527 367
rect 1393 313 1407 327
rect 1673 1113 1687 1127
rect 1873 1793 1887 1807
rect 1973 3553 1987 3567
rect 2013 3533 2027 3547
rect 1993 3493 2007 3507
rect 1993 3273 2007 3287
rect 2053 3733 2067 3747
rect 2073 3713 2087 3727
rect 2113 3693 2127 3707
rect 2073 3493 2087 3507
rect 2113 3493 2127 3507
rect 2033 3253 2047 3267
rect 2013 3233 2027 3247
rect 1973 3213 1987 3227
rect 1973 3193 1987 3207
rect 1953 3033 1967 3047
rect 1953 3013 1967 3027
rect 1933 2993 1947 3007
rect 2053 3053 2067 3067
rect 2013 3013 2027 3027
rect 1993 2993 2007 3007
rect 1973 2973 1987 2987
rect 2033 2853 2047 2867
rect 2033 2813 2047 2827
rect 1953 2793 1967 2807
rect 1973 2773 1987 2787
rect 1913 2753 1927 2767
rect 1953 2753 1967 2767
rect 1933 2733 1947 2747
rect 1913 2553 1927 2567
rect 1913 2513 1927 2527
rect 2013 2753 2027 2767
rect 1993 2713 2007 2727
rect 2013 2693 2027 2707
rect 1993 2533 2007 2547
rect 2013 2513 2027 2527
rect 1973 2413 1987 2427
rect 2093 3473 2107 3487
rect 2133 3453 2147 3467
rect 2273 3993 2287 4007
rect 2253 3973 2267 3987
rect 2293 3973 2307 3987
rect 2213 3913 2227 3927
rect 2333 4513 2347 4527
rect 2373 4533 2387 4547
rect 2433 4713 2447 4727
rect 2473 4693 2487 4707
rect 2593 4973 2607 4987
rect 2653 4973 2667 4987
rect 2573 4953 2587 4967
rect 2633 4953 2647 4967
rect 2673 4953 2687 4967
rect 2693 4913 2707 4927
rect 2653 4873 2667 4887
rect 2613 4853 2627 4867
rect 2653 4693 2667 4707
rect 2413 4673 2427 4687
rect 2453 4673 2467 4687
rect 2493 4673 2507 4687
rect 2593 4673 2607 4687
rect 2633 4673 2647 4687
rect 2613 4653 2627 4667
rect 2653 4573 2667 4587
rect 2573 4553 2587 4567
rect 2553 4533 2567 4547
rect 2413 4513 2427 4527
rect 2473 4473 2487 4487
rect 2353 4193 2367 4207
rect 2533 4453 2547 4467
rect 2493 4413 2507 4427
rect 2513 4413 2527 4427
rect 2473 4233 2487 4247
rect 2473 4213 2487 4227
rect 2433 4193 2447 4207
rect 2493 4193 2507 4207
rect 2313 3813 2327 3827
rect 2173 3753 2187 3767
rect 2253 3753 2267 3767
rect 2213 3713 2227 3727
rect 2293 3733 2307 3747
rect 2233 3693 2247 3707
rect 2273 3693 2287 3707
rect 2293 3693 2307 3707
rect 2393 4173 2407 4187
rect 2373 4153 2387 4167
rect 2353 3973 2367 3987
rect 2373 3753 2387 3767
rect 2353 3713 2367 3727
rect 2373 3713 2387 3727
rect 2373 3673 2387 3687
rect 2193 3533 2207 3547
rect 2213 3533 2227 3547
rect 2273 3533 2287 3547
rect 2153 3373 2167 3387
rect 2113 3273 2127 3287
rect 2133 3273 2147 3287
rect 2153 3273 2167 3287
rect 2093 3253 2107 3267
rect 2093 3073 2107 3087
rect 2093 3033 2107 3047
rect 2133 3053 2147 3067
rect 2273 3473 2287 3487
rect 3093 5613 3107 5627
rect 3013 5593 3027 5607
rect 2973 5493 2987 5507
rect 2973 5393 2987 5407
rect 2933 5373 2947 5387
rect 2973 5373 2987 5387
rect 2853 5133 2867 5147
rect 2773 5113 2787 5127
rect 2913 5153 2927 5167
rect 2933 5133 2947 5147
rect 2753 5093 2767 5107
rect 2873 5093 2887 5107
rect 2793 4993 2807 5007
rect 2733 4953 2747 4967
rect 2753 4953 2767 4967
rect 2733 4913 2747 4927
rect 2773 4913 2787 4927
rect 2713 4853 2727 4867
rect 2733 4793 2747 4807
rect 2773 4693 2787 4707
rect 2753 4673 2767 4687
rect 2713 4613 2727 4627
rect 2693 4553 2707 4567
rect 2573 4493 2587 4507
rect 2593 4453 2607 4467
rect 2653 4493 2667 4507
rect 2733 4493 2747 4507
rect 2673 4413 2687 4427
rect 2633 4213 2647 4227
rect 2653 4213 2667 4227
rect 2553 4153 2567 4167
rect 2613 4153 2627 4167
rect 2593 4133 2607 4147
rect 2593 4113 2607 4127
rect 2433 4013 2447 4027
rect 2493 4013 2507 4027
rect 2513 4013 2527 4027
rect 2553 4013 2567 4027
rect 2433 3993 2447 4007
rect 2473 3973 2487 3987
rect 2493 3973 2507 3987
rect 2413 3953 2427 3967
rect 2453 3953 2467 3967
rect 2533 3973 2547 3987
rect 2573 3953 2587 3967
rect 2593 3953 2607 3967
rect 2633 3953 2647 3967
rect 2653 3953 2667 3967
rect 2473 3933 2487 3947
rect 2513 3933 2527 3947
rect 2513 3733 2527 3747
rect 2553 3733 2567 3747
rect 2493 3713 2507 3727
rect 2533 3693 2547 3707
rect 2553 3673 2567 3687
rect 2513 3553 2527 3567
rect 2493 3533 2507 3547
rect 2393 3513 2407 3527
rect 2433 3513 2447 3527
rect 2333 3493 2347 3507
rect 2373 3493 2387 3507
rect 2393 3493 2407 3507
rect 2353 3473 2367 3487
rect 2293 3453 2307 3467
rect 2313 3453 2327 3467
rect 2233 3413 2247 3427
rect 2233 3373 2247 3387
rect 2293 3333 2307 3347
rect 2233 3253 2247 3267
rect 2393 3353 2407 3367
rect 2333 3253 2347 3267
rect 2373 3253 2387 3267
rect 2353 3233 2367 3247
rect 2293 3193 2307 3207
rect 2253 3073 2267 3087
rect 2333 3073 2347 3087
rect 2133 3033 2147 3047
rect 2193 3033 2207 3047
rect 2233 3033 2247 3047
rect 2113 3013 2127 3027
rect 2213 3013 2227 3027
rect 2153 2953 2167 2967
rect 2073 2793 2087 2807
rect 2053 2773 2067 2787
rect 2133 2773 2147 2787
rect 2173 2773 2187 2787
rect 2093 2753 2107 2767
rect 2073 2733 2087 2747
rect 2313 3033 2327 3047
rect 2253 2993 2267 3007
rect 2373 3133 2387 3147
rect 2293 2953 2307 2967
rect 2353 2953 2367 2967
rect 2353 2933 2367 2947
rect 2253 2773 2267 2787
rect 2233 2713 2247 2727
rect 2133 2573 2147 2587
rect 2053 2513 2067 2527
rect 2073 2433 2087 2447
rect 2033 2393 2047 2407
rect 1933 2273 1947 2287
rect 2033 2273 2047 2287
rect 2153 2533 2167 2547
rect 2113 2513 2127 2527
rect 2293 2753 2307 2767
rect 2333 2733 2347 2747
rect 2273 2693 2287 2707
rect 2253 2553 2267 2567
rect 2253 2533 2267 2547
rect 2293 2533 2307 2547
rect 2233 2513 2247 2527
rect 2273 2513 2287 2527
rect 2153 2473 2167 2487
rect 2193 2473 2207 2487
rect 1913 2133 1927 2147
rect 1893 1673 1907 1687
rect 1993 2233 2007 2247
rect 1993 2173 2007 2187
rect 1973 2093 1987 2107
rect 1953 2053 1967 2067
rect 2013 2153 2027 2167
rect 2093 2253 2107 2267
rect 2053 2133 2067 2147
rect 2053 1933 2067 1947
rect 2133 2193 2147 2207
rect 2233 2453 2247 2467
rect 2193 2273 2207 2287
rect 2413 3193 2427 3207
rect 2533 3533 2547 3547
rect 2473 3493 2487 3507
rect 2513 3493 2527 3507
rect 2533 3473 2547 3487
rect 2533 3273 2547 3287
rect 2493 3253 2507 3267
rect 2513 3233 2527 3247
rect 2713 4313 2727 4327
rect 2693 4193 2707 4207
rect 2813 4973 2827 4987
rect 2853 4973 2867 4987
rect 2833 4933 2847 4947
rect 2873 4933 2887 4947
rect 2813 4913 2827 4927
rect 2833 4913 2847 4927
rect 2953 5113 2967 5127
rect 3253 5593 3267 5607
rect 3273 5593 3287 5607
rect 3313 5593 3327 5607
rect 3233 5573 3247 5587
rect 3153 5433 3167 5447
rect 3193 5433 3207 5447
rect 3233 5433 3247 5447
rect 3073 5413 3087 5427
rect 3093 5393 3107 5407
rect 3073 5293 3087 5307
rect 3013 5213 3027 5227
rect 3013 5173 3027 5187
rect 3053 5153 3067 5167
rect 2993 5133 3007 5147
rect 3033 5133 3047 5147
rect 2973 4993 2987 5007
rect 3013 4993 3027 5007
rect 2953 4933 2967 4947
rect 2913 4893 2927 4907
rect 2913 4693 2927 4707
rect 2833 4653 2847 4667
rect 2933 4653 2947 4667
rect 2993 4853 3007 4867
rect 2973 4693 2987 4707
rect 3033 4713 3047 4727
rect 3013 4653 3027 4667
rect 2833 4633 2847 4647
rect 2873 4633 2887 4647
rect 2893 4633 2907 4647
rect 2953 4633 2967 4647
rect 2813 4613 2827 4627
rect 2913 4513 2927 4527
rect 2813 4413 2827 4427
rect 2853 4393 2867 4407
rect 2753 4193 2767 4207
rect 2793 4193 2807 4207
rect 2773 4153 2787 4167
rect 2693 4113 2707 4127
rect 2793 4133 2807 4147
rect 2793 4073 2807 4087
rect 2773 3993 2787 4007
rect 2713 3973 2727 3987
rect 2733 3953 2747 3967
rect 2693 3873 2707 3887
rect 2673 3793 2687 3807
rect 2613 3773 2627 3787
rect 2693 3753 2707 3767
rect 2773 3753 2787 3767
rect 2653 3733 2667 3747
rect 2573 3553 2587 3567
rect 2573 3533 2587 3547
rect 2753 3713 2767 3727
rect 2793 3693 2807 3707
rect 2633 3673 2647 3687
rect 2693 3673 2707 3687
rect 2713 3633 2727 3647
rect 2653 3533 2667 3547
rect 2633 3513 2647 3527
rect 2613 3353 2627 3367
rect 2593 3253 2607 3267
rect 2693 3293 2707 3307
rect 2653 3273 2667 3287
rect 2553 3213 2567 3227
rect 2473 3173 2487 3187
rect 2433 3133 2447 3147
rect 2393 3113 2407 3127
rect 2433 3113 2447 3127
rect 2393 3013 2407 3027
rect 2513 3033 2527 3047
rect 2613 3213 2627 3227
rect 2493 3013 2507 3027
rect 2593 3013 2607 3027
rect 2453 2933 2467 2947
rect 2433 2813 2447 2827
rect 2393 2793 2407 2807
rect 2493 2793 2507 2807
rect 2573 2793 2587 2807
rect 2413 2753 2427 2767
rect 2393 2553 2407 2567
rect 2453 2553 2467 2567
rect 2373 2533 2387 2547
rect 2473 2513 2487 2527
rect 2413 2433 2427 2447
rect 2393 2393 2407 2407
rect 2353 2353 2367 2367
rect 2313 2313 2327 2327
rect 2333 2313 2347 2327
rect 2373 2293 2387 2307
rect 2353 2273 2367 2287
rect 2173 2233 2187 2247
rect 2153 2093 2167 2107
rect 2113 1853 2127 1867
rect 2033 1833 2047 1847
rect 2073 1833 2087 1847
rect 2113 1833 2127 1847
rect 1973 1793 1987 1807
rect 1933 1753 1947 1767
rect 1993 1753 2007 1767
rect 1913 1633 1927 1647
rect 1973 1633 1987 1647
rect 1853 1613 1867 1627
rect 1873 1613 1887 1627
rect 1913 1613 1927 1627
rect 1853 1593 1867 1607
rect 1853 1533 1867 1547
rect 1853 1493 1867 1507
rect 1953 1593 1967 1607
rect 1933 1573 1947 1587
rect 1973 1573 1987 1587
rect 1893 1553 1907 1567
rect 1953 1373 1967 1387
rect 1933 1293 1947 1307
rect 1873 1253 1887 1267
rect 1853 1133 1867 1147
rect 1873 1113 1887 1127
rect 1813 1093 1827 1107
rect 1853 1053 1867 1067
rect 2013 1713 2027 1727
rect 2013 1373 2027 1387
rect 1993 1293 2007 1307
rect 2113 1813 2127 1827
rect 2173 2073 2187 2087
rect 2193 2073 2207 2087
rect 2173 1953 2187 1967
rect 2153 1793 2167 1807
rect 2133 1693 2147 1707
rect 2093 1613 2107 1627
rect 2133 1593 2147 1607
rect 2093 1553 2107 1567
rect 2133 1553 2147 1567
rect 2093 1453 2107 1467
rect 2053 1373 2067 1387
rect 2033 1333 2047 1347
rect 2253 2253 2267 2267
rect 2273 2253 2287 2267
rect 2313 2253 2327 2267
rect 2233 2113 2247 2127
rect 2253 2113 2267 2127
rect 2273 2093 2287 2107
rect 2293 2053 2307 2067
rect 2533 2773 2547 2787
rect 2553 2753 2567 2767
rect 2513 2733 2527 2747
rect 2693 3233 2707 3247
rect 2673 3213 2687 3227
rect 2793 3593 2807 3607
rect 2733 3553 2747 3567
rect 2773 3513 2787 3527
rect 2753 3493 2767 3507
rect 2773 3353 2787 3367
rect 2773 3333 2787 3347
rect 2733 3273 2747 3287
rect 2873 4213 2887 4227
rect 2853 4113 2867 4127
rect 2853 4033 2867 4047
rect 2893 4013 2907 4027
rect 2833 3973 2847 3987
rect 2873 3873 2887 3887
rect 2853 3833 2867 3847
rect 2833 3733 2847 3747
rect 2893 3733 2907 3747
rect 2973 4613 2987 4627
rect 3053 4593 3067 4607
rect 3113 5273 3127 5287
rect 3093 5153 3107 5167
rect 3173 5373 3187 5387
rect 3233 5393 3247 5407
rect 3213 5353 3227 5367
rect 3153 5193 3167 5207
rect 3113 5133 3127 5147
rect 3193 5153 3207 5167
rect 3133 5113 3147 5127
rect 3233 5093 3247 5107
rect 3673 5933 3687 5947
rect 3513 5893 3527 5907
rect 3473 5753 3487 5767
rect 3413 5733 3427 5747
rect 3593 5733 3607 5747
rect 3553 5673 3567 5687
rect 3513 5653 3527 5667
rect 3553 5653 3567 5667
rect 3373 5633 3387 5647
rect 3653 5893 3667 5907
rect 3773 5893 3787 5907
rect 3693 5873 3707 5887
rect 3833 5933 3847 5947
rect 3873 5933 3887 5947
rect 3913 5933 3927 5947
rect 3993 5933 4007 5947
rect 4253 5933 4267 5947
rect 3833 5893 3847 5907
rect 4013 5893 4027 5907
rect 3913 5873 3927 5887
rect 3813 5853 3827 5867
rect 3773 5753 3787 5767
rect 3613 5713 3627 5727
rect 3833 5693 3847 5707
rect 3793 5673 3807 5687
rect 3753 5653 3767 5667
rect 3773 5653 3787 5667
rect 3613 5633 3627 5647
rect 3653 5633 3667 5647
rect 3693 5633 3707 5647
rect 3493 5613 3507 5627
rect 3573 5613 3587 5627
rect 3593 5613 3607 5627
rect 3353 5593 3367 5607
rect 3533 5593 3547 5607
rect 3633 5613 3647 5627
rect 3673 5613 3687 5627
rect 3333 5573 3347 5587
rect 3613 5573 3627 5587
rect 3293 5493 3307 5507
rect 3273 5393 3287 5407
rect 3313 5393 3327 5407
rect 3473 5493 3487 5507
rect 3433 5433 3447 5447
rect 3613 5453 3627 5467
rect 3553 5433 3567 5447
rect 3593 5433 3607 5447
rect 3413 5413 3427 5427
rect 3713 5413 3727 5427
rect 3553 5373 3567 5387
rect 3573 5293 3587 5307
rect 3533 5253 3547 5267
rect 3453 5173 3467 5187
rect 3273 5153 3287 5167
rect 3333 5153 3347 5167
rect 3433 5153 3447 5167
rect 3313 5133 3327 5147
rect 3733 5353 3747 5367
rect 3753 5353 3767 5367
rect 3633 5253 3647 5267
rect 3693 5253 3707 5267
rect 3253 4973 3267 4987
rect 3093 4833 3107 4847
rect 3093 4673 3107 4687
rect 3213 4933 3227 4947
rect 3153 4913 3167 4927
rect 3113 4653 3127 4667
rect 3173 4673 3187 4687
rect 3153 4653 3167 4667
rect 3133 4593 3147 4607
rect 3193 4553 3207 4567
rect 3273 4913 3287 4927
rect 3313 4953 3327 4967
rect 3393 4973 3407 4987
rect 3353 4953 3367 4967
rect 3313 4893 3327 4907
rect 3293 4853 3307 4867
rect 3413 4933 3427 4947
rect 3373 4873 3387 4887
rect 3353 4813 3367 4827
rect 3273 4673 3287 4687
rect 3253 4653 3267 4667
rect 3293 4653 3307 4667
rect 3393 4713 3407 4727
rect 3273 4633 3287 4647
rect 3313 4633 3327 4647
rect 3013 4473 3027 4487
rect 2953 4453 2967 4467
rect 2993 4453 3007 4467
rect 2933 4413 2947 4427
rect 2993 4213 3007 4227
rect 2973 4193 2987 4207
rect 2933 4153 2947 4167
rect 3013 4133 3027 4147
rect 3213 4513 3227 4527
rect 3113 4493 3127 4507
rect 3253 4493 3267 4507
rect 3073 4473 3087 4487
rect 3133 4473 3147 4487
rect 3053 4073 3067 4087
rect 2993 4033 3007 4047
rect 2973 3993 2987 4007
rect 3033 3993 3047 4007
rect 2873 3593 2887 3607
rect 2913 3593 2927 3607
rect 3013 3693 3027 3707
rect 3053 3693 3067 3707
rect 3053 3653 3067 3667
rect 3053 3593 3067 3607
rect 2973 3533 2987 3547
rect 2913 3513 2927 3527
rect 2833 3493 2847 3507
rect 2853 3493 2867 3507
rect 2813 3253 2827 3267
rect 2753 3233 2767 3247
rect 2953 3473 2967 3487
rect 2913 3273 2927 3287
rect 2873 3233 2887 3247
rect 2753 3213 2767 3227
rect 2853 3213 2867 3227
rect 2893 3213 2907 3227
rect 2933 3213 2947 3227
rect 2673 3193 2687 3207
rect 2713 3193 2727 3207
rect 2673 3013 2687 3027
rect 2713 3013 2727 3027
rect 2893 3193 2907 3207
rect 2793 3133 2807 3147
rect 2793 3053 2807 3067
rect 2873 3053 2887 3067
rect 2633 2993 2647 3007
rect 2693 2993 2707 3007
rect 2753 2993 2767 3007
rect 2873 3033 2887 3047
rect 2833 3013 2847 3027
rect 2933 3053 2947 3067
rect 3033 3473 3047 3487
rect 2993 3213 3007 3227
rect 3033 3193 3047 3207
rect 2973 3173 2987 3187
rect 3013 3053 3027 3067
rect 2973 3013 2987 3027
rect 2753 2953 2767 2967
rect 2733 2793 2747 2807
rect 2653 2773 2667 2787
rect 2513 2713 2527 2727
rect 2613 2713 2627 2727
rect 2453 2293 2467 2307
rect 2493 2293 2507 2307
rect 2413 2273 2427 2287
rect 2733 2773 2747 2787
rect 2733 2733 2747 2747
rect 2773 2773 2787 2787
rect 2793 2753 2807 2767
rect 2673 2693 2687 2707
rect 2713 2693 2727 2707
rect 2713 2573 2727 2587
rect 2533 2533 2547 2547
rect 2573 2433 2587 2447
rect 2573 2313 2587 2327
rect 2533 2273 2547 2287
rect 2513 2253 2527 2267
rect 2433 2033 2447 2047
rect 2273 2013 2287 2027
rect 2393 2013 2407 2027
rect 2213 1813 2227 1827
rect 2733 2533 2747 2547
rect 2633 2473 2647 2487
rect 2753 2433 2767 2447
rect 2633 2353 2647 2367
rect 2533 2213 2547 2227
rect 2493 2153 2507 2167
rect 2553 2153 2567 2167
rect 2453 1953 2467 1967
rect 2473 1833 2487 1847
rect 2553 2073 2567 2087
rect 2593 2073 2607 2087
rect 2533 2033 2547 2047
rect 2593 2033 2607 2047
rect 2573 1933 2587 1947
rect 2533 1873 2547 1887
rect 2673 2273 2687 2287
rect 2713 2273 2727 2287
rect 2833 2673 2847 2687
rect 2793 2573 2807 2587
rect 2813 2573 2827 2587
rect 2853 2573 2867 2587
rect 2773 2233 2787 2247
rect 2773 2213 2787 2227
rect 2693 2133 2707 2147
rect 2633 2073 2647 2087
rect 2653 2053 2667 2067
rect 2633 2033 2647 2047
rect 2633 2013 2647 2027
rect 2613 1813 2627 1827
rect 2833 2533 2847 2547
rect 2813 2453 2827 2467
rect 2993 2993 3007 3007
rect 2953 2913 2967 2927
rect 2953 2813 2967 2827
rect 2913 2753 2927 2767
rect 2973 2773 2987 2787
rect 3293 4473 3307 4487
rect 3433 4633 3447 4647
rect 3553 5033 3567 5047
rect 3653 5213 3667 5227
rect 3813 5633 3827 5647
rect 3793 5433 3807 5447
rect 3833 5413 3847 5427
rect 4133 5913 4147 5927
rect 4293 5913 4307 5927
rect 4473 6013 4487 6027
rect 4973 5953 4987 5967
rect 4113 5893 4127 5907
rect 4153 5893 4167 5907
rect 4273 5893 4287 5907
rect 4313 5893 4327 5907
rect 4573 5913 4587 5927
rect 4613 5913 4627 5927
rect 4793 5893 4807 5907
rect 4933 5893 4947 5907
rect 4433 5873 4447 5887
rect 4693 5873 4707 5887
rect 4773 5873 4787 5887
rect 4053 5853 4067 5867
rect 3933 5693 3947 5707
rect 3953 5653 3967 5667
rect 3933 5613 3947 5627
rect 3953 5613 3967 5627
rect 3973 5593 3987 5607
rect 3993 5453 4007 5467
rect 3853 5393 3867 5407
rect 3973 5373 3987 5387
rect 3933 5273 3947 5287
rect 3773 5153 3787 5167
rect 3893 5173 3907 5187
rect 3993 5173 4007 5187
rect 3873 5153 3887 5167
rect 4293 5713 4307 5727
rect 4073 5633 4087 5647
rect 4113 5633 4127 5647
rect 4233 5633 4247 5647
rect 4053 5593 4067 5607
rect 4173 5593 4187 5607
rect 4913 5873 4927 5887
rect 4953 5873 4967 5887
rect 4773 5753 4787 5767
rect 4813 5753 4827 5767
rect 4493 5713 4507 5727
rect 4433 5633 4447 5647
rect 4833 5673 4847 5687
rect 4693 5653 4707 5667
rect 4773 5653 4787 5667
rect 4813 5653 4827 5667
rect 4533 5633 4547 5647
rect 4633 5633 4647 5647
rect 4673 5633 4687 5647
rect 4373 5613 4387 5627
rect 4513 5593 4527 5607
rect 4513 5533 4527 5547
rect 4193 5493 4207 5507
rect 4333 5493 4347 5507
rect 4473 5493 4487 5507
rect 4113 5433 4127 5447
rect 4233 5453 4247 5467
rect 4473 5453 4487 5467
rect 4193 5433 4207 5447
rect 4153 5413 4167 5427
rect 4193 5393 4207 5407
rect 4273 5393 4287 5407
rect 4213 5373 4227 5387
rect 4293 5233 4307 5247
rect 4113 5173 4127 5187
rect 4173 5173 4187 5187
rect 4193 5173 4207 5187
rect 4013 5153 4027 5167
rect 4013 5113 4027 5127
rect 3833 5093 3847 5107
rect 3853 5093 3867 5107
rect 3713 5033 3727 5047
rect 3693 4973 3707 4987
rect 3593 4953 3607 4967
rect 3633 4953 3647 4967
rect 3673 4953 3687 4967
rect 3733 4953 3747 4967
rect 3553 4873 3567 4887
rect 3513 4833 3527 4847
rect 3633 4893 3647 4907
rect 3573 4793 3587 4807
rect 3553 4693 3567 4707
rect 3573 4673 3587 4687
rect 3473 4633 3487 4647
rect 3633 4673 3647 4687
rect 3673 4673 3687 4687
rect 3653 4613 3667 4627
rect 3613 4573 3627 4587
rect 3453 4553 3467 4567
rect 3953 4953 3967 4967
rect 3993 4953 4007 4967
rect 3813 4913 3827 4927
rect 4093 5093 4107 5107
rect 4213 5153 4227 5167
rect 4393 5433 4407 5447
rect 4433 5433 4447 5447
rect 4413 5413 4427 5427
rect 4653 5613 4667 5627
rect 4613 5593 4627 5607
rect 4553 5493 4567 5507
rect 4533 5453 4547 5467
rect 4593 5453 4607 5467
rect 4793 5633 4807 5647
rect 4773 5473 4787 5487
rect 4433 5393 4447 5407
rect 4333 5193 4347 5207
rect 4393 5193 4407 5207
rect 4313 5173 4327 5187
rect 4353 5133 4367 5147
rect 4253 5113 4267 5127
rect 4173 4973 4187 4987
rect 4213 4973 4227 4987
rect 4333 4973 4347 4987
rect 4173 4953 4187 4967
rect 4133 4893 4147 4907
rect 4293 4933 4307 4947
rect 4273 4913 4287 4927
rect 4193 4873 4207 4887
rect 3933 4693 3947 4707
rect 3973 4673 3987 4687
rect 3773 4653 3787 4667
rect 3793 4633 3807 4647
rect 3793 4553 3807 4567
rect 3753 4533 3767 4547
rect 3433 4513 3447 4527
rect 3233 4413 3247 4427
rect 3213 4293 3227 4307
rect 3093 4213 3107 4227
rect 3153 4213 3167 4227
rect 3173 4213 3187 4227
rect 3313 4433 3327 4447
rect 3273 4293 3287 4307
rect 3293 4253 3307 4267
rect 3233 4193 3247 4207
rect 3173 4173 3187 4187
rect 3293 4173 3307 4187
rect 3153 4153 3167 4167
rect 3373 4433 3387 4447
rect 3333 4253 3347 4267
rect 3413 4213 3427 4227
rect 3373 4193 3387 4207
rect 3353 4173 3367 4187
rect 3333 4153 3347 4167
rect 3233 4133 3247 4147
rect 3313 4133 3327 4147
rect 3353 4133 3367 4147
rect 3153 4013 3167 4027
rect 3113 3953 3127 3967
rect 3133 3953 3147 3967
rect 3253 3993 3267 4007
rect 3313 3993 3327 4007
rect 3313 3973 3327 3987
rect 3413 4173 3427 4187
rect 3393 4033 3407 4047
rect 3393 4013 3407 4027
rect 3193 3913 3207 3927
rect 3213 3873 3227 3887
rect 3193 3733 3207 3747
rect 3113 3693 3127 3707
rect 3093 3593 3107 3607
rect 3073 3213 3087 3227
rect 3153 3573 3167 3587
rect 3193 3533 3207 3547
rect 3153 3513 3167 3527
rect 3253 3733 3267 3747
rect 3233 3693 3247 3707
rect 3233 3613 3247 3627
rect 3293 3593 3307 3607
rect 3213 3433 3227 3447
rect 3173 3233 3187 3247
rect 3113 3213 3127 3227
rect 3093 3193 3107 3207
rect 3153 3193 3167 3207
rect 3093 3173 3107 3187
rect 3333 3953 3347 3967
rect 3633 4493 3647 4507
rect 3953 4653 3967 4667
rect 3913 4633 3927 4647
rect 3893 4593 3907 4607
rect 3833 4493 3847 4507
rect 3493 4473 3507 4487
rect 3533 4453 3547 4467
rect 3613 4453 3627 4467
rect 3653 4433 3667 4447
rect 3453 4413 3467 4427
rect 3453 4393 3467 4407
rect 3433 3853 3447 3867
rect 3373 3753 3387 3767
rect 3373 3713 3387 3727
rect 3353 3693 3367 3707
rect 3253 3393 3267 3407
rect 3313 3393 3327 3407
rect 3393 3673 3407 3687
rect 3413 3533 3427 3547
rect 3433 3493 3447 3507
rect 3393 3473 3407 3487
rect 3813 4473 3827 4487
rect 3753 4413 3767 4427
rect 3693 4373 3707 4387
rect 3493 4213 3507 4227
rect 3773 4213 3787 4227
rect 3473 4193 3487 4207
rect 3633 4193 3647 4207
rect 3613 4173 3627 4187
rect 3513 4153 3527 4167
rect 3593 4153 3607 4167
rect 3473 4053 3487 4067
rect 3513 4053 3527 4067
rect 3473 4033 3487 4047
rect 3493 4013 3507 4027
rect 3573 3993 3587 4007
rect 3473 3733 3487 3747
rect 3513 3713 3527 3727
rect 3533 3693 3547 3707
rect 3553 3653 3567 3667
rect 3553 3633 3567 3647
rect 3513 3533 3527 3547
rect 3473 3493 3487 3507
rect 3553 3513 3567 3527
rect 3493 3453 3507 3467
rect 3453 3373 3467 3387
rect 3453 3293 3467 3307
rect 3273 3233 3287 3247
rect 3313 3233 3327 3247
rect 3353 3233 3367 3247
rect 3253 3213 3267 3227
rect 3293 3213 3307 3227
rect 3293 3193 3307 3207
rect 3333 3193 3347 3207
rect 3273 3113 3287 3127
rect 3213 3093 3227 3107
rect 3233 3073 3247 3087
rect 3113 3053 3127 3067
rect 3153 3033 3167 3047
rect 3193 3033 3207 3047
rect 3093 3013 3107 3027
rect 3133 3013 3147 3027
rect 3073 2973 3087 2987
rect 3053 2953 3067 2967
rect 3033 2913 3047 2927
rect 2973 2713 2987 2727
rect 2873 2433 2887 2447
rect 2833 2333 2847 2347
rect 2933 2533 2947 2547
rect 2953 2433 2967 2447
rect 2893 2293 2907 2307
rect 2913 2253 2927 2267
rect 2793 2193 2807 2207
rect 2873 2113 2887 2127
rect 2853 2073 2867 2087
rect 2813 2053 2827 2067
rect 2693 2013 2707 2027
rect 2673 1993 2687 2007
rect 2673 1933 2687 1947
rect 2653 1813 2667 1827
rect 2233 1713 2247 1727
rect 2293 1713 2307 1727
rect 2233 1693 2247 1707
rect 2293 1693 2307 1707
rect 2253 1633 2267 1647
rect 2193 1593 2207 1607
rect 2213 1593 2227 1607
rect 2233 1573 2247 1587
rect 2133 1373 2147 1387
rect 2173 1373 2187 1387
rect 2053 1313 2067 1327
rect 2013 1233 2027 1247
rect 1953 1193 1967 1207
rect 1973 1153 1987 1167
rect 1993 1033 2007 1047
rect 1853 873 1867 887
rect 1933 873 1947 887
rect 1653 833 1667 847
rect 1633 793 1647 807
rect 1753 793 1767 807
rect 1793 773 1807 787
rect 1793 753 1807 767
rect 1773 733 1787 747
rect 1633 673 1647 687
rect 1653 673 1667 687
rect 1833 813 1847 827
rect 1813 713 1827 727
rect 1793 673 1807 687
rect 1773 653 1787 667
rect 1813 653 1827 667
rect 1653 633 1667 647
rect 1713 633 1727 647
rect 1673 613 1687 627
rect 1693 573 1707 587
rect 1553 373 1567 387
rect 1593 373 1607 387
rect 1613 373 1627 387
rect 1653 373 1667 387
rect 1453 333 1467 347
rect 1533 333 1547 347
rect 1493 313 1507 327
rect 1433 293 1447 307
rect 1373 213 1387 227
rect 1233 193 1247 207
rect 1113 173 1127 187
rect 1173 173 1187 187
rect 1293 173 1307 187
rect 1153 153 1167 167
rect 1113 133 1127 147
rect 1133 133 1147 147
rect 1593 353 1607 367
rect 1613 333 1627 347
rect 1573 313 1587 327
rect 1633 273 1647 287
rect 1453 193 1467 207
rect 1553 193 1567 207
rect 1393 173 1407 187
rect 1453 153 1467 167
rect 1273 133 1287 147
rect 1313 133 1327 147
rect 1373 133 1387 147
rect 1533 133 1547 147
rect 1753 393 1767 407
rect 1713 353 1727 367
rect 1693 313 1707 327
rect 1413 113 1427 127
rect 1553 113 1567 127
rect 1593 113 1607 127
rect 1233 93 1247 107
rect 1013 73 1027 87
rect 1733 313 1747 327
rect 1733 233 1747 247
rect 1693 133 1707 147
rect 1653 113 1667 127
rect 1753 113 1767 127
rect 1813 313 1827 327
rect 1793 273 1807 287
rect 1893 853 1907 867
rect 1913 813 1927 827
rect 1933 813 1947 827
rect 1973 813 1987 827
rect 1933 793 1947 807
rect 1973 693 1987 707
rect 1933 633 1947 647
rect 1973 633 1987 647
rect 1913 613 1927 627
rect 1953 593 1967 607
rect 1973 593 1987 607
rect 1953 533 1967 547
rect 1893 373 1907 387
rect 1973 353 1987 367
rect 1873 333 1887 347
rect 1813 133 1827 147
rect 1753 93 1767 107
rect 1773 93 1787 107
rect 1733 33 1747 47
rect 1633 13 1647 27
rect 1693 13 1707 27
rect 1933 313 1947 327
rect 1853 253 1867 267
rect 1913 253 1927 267
rect 1913 233 1927 247
rect 1933 233 1947 247
rect 2013 993 2027 1007
rect 2093 1033 2107 1047
rect 2013 893 2027 907
rect 2053 893 2067 907
rect 1893 173 1907 187
rect 1933 173 1947 187
rect 1913 133 1927 147
rect 1913 113 1927 127
rect 1873 73 1887 87
rect 1833 13 1847 27
rect 1873 13 1887 27
rect 2053 853 2067 867
rect 2033 673 2047 687
rect 2073 833 2087 847
rect 2113 773 2127 787
rect 2033 613 2047 627
rect 2053 613 2067 627
rect 2053 433 2067 447
rect 2033 413 2047 427
rect 2193 1333 2207 1347
rect 2153 1313 2167 1327
rect 2173 1293 2187 1307
rect 2153 1153 2167 1167
rect 2213 1133 2227 1147
rect 2173 873 2187 887
rect 2193 853 2207 867
rect 2153 833 2167 847
rect 2253 1113 2267 1127
rect 2493 1773 2507 1787
rect 2553 1733 2567 1747
rect 2633 1793 2647 1807
rect 2613 1773 2627 1787
rect 2653 1773 2667 1787
rect 2733 1873 2747 1887
rect 2693 1813 2707 1827
rect 2773 1813 2787 1827
rect 2713 1793 2727 1807
rect 2753 1793 2767 1807
rect 2633 1673 2647 1687
rect 2413 1633 2427 1647
rect 2453 1633 2467 1647
rect 2513 1633 2527 1647
rect 2593 1633 2607 1647
rect 2313 1593 2327 1607
rect 2373 1593 2387 1607
rect 2333 1573 2347 1587
rect 2313 1513 2327 1527
rect 2433 1593 2447 1607
rect 2493 1553 2507 1567
rect 2493 1533 2507 1547
rect 2373 1413 2387 1427
rect 2413 1413 2427 1427
rect 2313 1293 2327 1307
rect 2353 1273 2367 1287
rect 2313 1093 2327 1107
rect 2233 1033 2247 1047
rect 2273 1033 2287 1047
rect 2313 893 2327 907
rect 2233 853 2247 867
rect 2213 813 2227 827
rect 2173 733 2187 747
rect 2313 833 2327 847
rect 2333 813 2347 827
rect 2293 773 2307 787
rect 2233 673 2247 687
rect 2153 633 2167 647
rect 2193 613 2207 627
rect 2433 1293 2447 1307
rect 2553 1593 2567 1607
rect 2593 1573 2607 1587
rect 2573 1553 2587 1567
rect 2613 1553 2627 1567
rect 2573 1313 2587 1327
rect 2533 1293 2547 1307
rect 2513 1213 2527 1227
rect 2613 1173 2627 1187
rect 2393 1113 2407 1127
rect 2433 1093 2447 1107
rect 2453 1073 2467 1087
rect 2453 853 2467 867
rect 2493 853 2507 867
rect 2893 2033 2907 2047
rect 2793 1793 2807 1807
rect 2853 1793 2867 1807
rect 2773 1713 2787 1727
rect 2673 1573 2687 1587
rect 2733 1573 2747 1587
rect 2713 1553 2727 1567
rect 2673 1533 2687 1547
rect 2753 1513 2767 1527
rect 2673 1313 2687 1327
rect 2713 1313 2727 1327
rect 2773 1313 2787 1327
rect 2653 1293 2667 1307
rect 2693 1293 2707 1307
rect 2753 1293 2767 1307
rect 2733 1173 2747 1187
rect 2733 1153 2747 1167
rect 2633 1133 2647 1147
rect 2673 1133 2687 1147
rect 2613 1113 2627 1127
rect 2873 1773 2887 1787
rect 2833 1753 2847 1767
rect 2893 1633 2907 1647
rect 3013 2733 3027 2747
rect 2993 2693 3007 2707
rect 2993 2633 3007 2647
rect 3073 2813 3087 2827
rect 3013 2553 3027 2567
rect 3033 2453 3047 2467
rect 3133 2753 3147 2767
rect 3093 2733 3107 2747
rect 3113 2733 3127 2747
rect 3073 2573 3087 2587
rect 3153 2673 3167 2687
rect 3193 2993 3207 3007
rect 3253 3013 3267 3027
rect 3353 3133 3367 3147
rect 3353 3073 3367 3087
rect 3333 3033 3347 3047
rect 3393 3253 3407 3267
rect 3433 3253 3447 3267
rect 3393 3153 3407 3167
rect 3273 2893 3287 2907
rect 3233 2793 3247 2807
rect 3213 2773 3227 2787
rect 3193 2733 3207 2747
rect 3093 2513 3107 2527
rect 3053 2393 3067 2407
rect 3133 2393 3147 2407
rect 2993 2373 3007 2387
rect 2973 2253 2987 2267
rect 3033 2293 3047 2307
rect 3053 2273 3067 2287
rect 3033 2213 3047 2227
rect 2973 2193 2987 2207
rect 2953 2133 2967 2147
rect 2933 2113 2947 2127
rect 3013 2073 3027 2087
rect 2933 1833 2947 1847
rect 2993 1793 3007 1807
rect 3033 1753 3047 1767
rect 3013 1633 3027 1647
rect 2933 1613 2947 1627
rect 2973 1573 2987 1587
rect 2993 1573 3007 1587
rect 2913 1553 2927 1567
rect 2873 1533 2887 1547
rect 3073 2253 3087 2267
rect 3113 2253 3127 2267
rect 3253 2733 3267 2747
rect 3253 2593 3267 2607
rect 3273 2593 3287 2607
rect 3233 2573 3247 2587
rect 3173 2433 3187 2447
rect 3213 2373 3227 2387
rect 3153 2313 3167 2327
rect 3193 2253 3207 2267
rect 3153 2213 3167 2227
rect 3133 2073 3147 2087
rect 3153 2053 3167 2067
rect 3193 2053 3207 2067
rect 3133 2033 3147 2047
rect 3173 2013 3187 2027
rect 3433 3213 3447 3227
rect 3493 3213 3507 3227
rect 3433 3193 3447 3207
rect 3473 3193 3487 3207
rect 3613 4073 3627 4087
rect 3633 4033 3647 4047
rect 3713 4173 3727 4187
rect 3653 4013 3667 4027
rect 3653 3993 3667 4007
rect 3593 3813 3607 3827
rect 3853 4473 3867 4487
rect 3973 4573 3987 4587
rect 3953 4533 3967 4547
rect 3733 4153 3747 4167
rect 3833 4153 3847 4167
rect 3753 4073 3767 4087
rect 3733 3993 3747 4007
rect 3793 4053 3807 4067
rect 3833 3813 3847 3827
rect 3713 3733 3727 3747
rect 3673 3713 3687 3727
rect 3713 3713 3727 3727
rect 3633 3693 3647 3707
rect 3653 3693 3667 3707
rect 3773 3693 3787 3707
rect 3633 3633 3647 3647
rect 3693 3633 3707 3647
rect 3693 3613 3707 3627
rect 3673 3573 3687 3587
rect 3633 3553 3647 3567
rect 3573 3453 3587 3467
rect 3553 3253 3567 3267
rect 3613 3253 3627 3267
rect 3593 3233 3607 3247
rect 3513 3173 3527 3187
rect 3493 3153 3507 3167
rect 3413 3033 3427 3047
rect 3433 3033 3447 3047
rect 3413 2993 3427 3007
rect 3373 2973 3387 2987
rect 3373 2953 3387 2967
rect 3433 2973 3447 2987
rect 3413 2853 3427 2867
rect 3413 2753 3427 2767
rect 3393 2693 3407 2707
rect 3393 2613 3407 2627
rect 3353 2593 3367 2607
rect 3333 2573 3347 2587
rect 3293 2553 3307 2567
rect 3293 2373 3307 2387
rect 3353 2553 3367 2567
rect 3453 2833 3467 2847
rect 3573 3213 3587 3227
rect 3533 3053 3547 3067
rect 3533 3013 3547 3027
rect 3653 3513 3667 3527
rect 3813 3713 3827 3727
rect 3793 3633 3807 3647
rect 3773 3593 3787 3607
rect 3833 3593 3847 3607
rect 3793 3573 3807 3587
rect 3733 3533 3747 3547
rect 3733 3513 3747 3527
rect 3713 3493 3727 3507
rect 3653 3473 3667 3487
rect 3693 3293 3707 3307
rect 3753 3233 3767 3247
rect 3633 3213 3647 3227
rect 3653 3213 3667 3227
rect 3713 3213 3727 3227
rect 3733 3213 3747 3227
rect 3653 3113 3667 3127
rect 3633 3033 3647 3047
rect 3693 3033 3707 3047
rect 3613 3013 3627 3027
rect 3673 3013 3687 3027
rect 3573 2993 3587 3007
rect 3593 2993 3607 3007
rect 3693 2993 3707 3007
rect 3513 2793 3527 2807
rect 3633 2793 3647 2807
rect 3653 2793 3667 2807
rect 3513 2773 3527 2787
rect 3513 2753 3527 2767
rect 3473 2733 3487 2747
rect 3433 2713 3447 2727
rect 3333 2313 3347 2327
rect 3293 2293 3307 2307
rect 3273 2273 3287 2287
rect 3233 2193 3247 2207
rect 3313 2193 3327 2207
rect 3413 2313 3427 2327
rect 3353 2133 3367 2147
rect 3273 2113 3287 2127
rect 3333 2093 3347 2107
rect 3293 2053 3307 2067
rect 3273 2033 3287 2047
rect 3193 1993 3207 2007
rect 3213 1993 3227 2007
rect 3273 1993 3287 2007
rect 3133 1933 3147 1947
rect 3253 1813 3267 1827
rect 3053 1593 3067 1607
rect 3093 1593 3107 1607
rect 3053 1573 3067 1587
rect 3093 1573 3107 1587
rect 3073 1553 3087 1567
rect 3053 1533 3067 1547
rect 3093 1533 3107 1547
rect 2993 1513 3007 1527
rect 2973 1373 2987 1387
rect 2833 1333 2847 1347
rect 2873 1313 2887 1327
rect 2793 1273 2807 1287
rect 2813 1273 2827 1287
rect 2813 1113 2827 1127
rect 2993 1333 3007 1347
rect 2973 1313 2987 1327
rect 2933 1273 2947 1287
rect 2873 1213 2887 1227
rect 2913 1213 2927 1227
rect 2773 1093 2787 1107
rect 2733 1073 2747 1087
rect 2833 1073 2847 1087
rect 2553 1033 2567 1047
rect 2433 793 2447 807
rect 2513 833 2527 847
rect 2493 793 2507 807
rect 2373 773 2387 787
rect 2413 773 2427 787
rect 2473 773 2487 787
rect 2353 733 2367 747
rect 2373 733 2387 747
rect 2353 713 2367 727
rect 2333 693 2347 707
rect 2353 673 2367 687
rect 2313 613 2327 627
rect 2433 713 2447 727
rect 2413 653 2427 667
rect 2473 633 2487 647
rect 2693 873 2707 887
rect 2593 853 2607 867
rect 2633 853 2647 867
rect 2673 853 2687 867
rect 2573 833 2587 847
rect 2613 813 2627 827
rect 2613 713 2627 727
rect 2533 633 2547 647
rect 2553 633 2567 647
rect 2413 613 2427 627
rect 2453 613 2467 627
rect 2493 613 2507 627
rect 2273 493 2287 507
rect 2413 473 2427 487
rect 2353 433 2367 447
rect 2173 413 2187 427
rect 2073 373 2087 387
rect 2093 353 2107 367
rect 2133 333 2147 347
rect 2113 293 2127 307
rect 2013 133 2027 147
rect 2213 373 2227 387
rect 2233 353 2247 367
rect 2353 373 2367 387
rect 2393 373 2407 387
rect 2373 353 2387 367
rect 2273 293 2287 307
rect 2173 253 2187 267
rect 2313 153 2327 167
rect 2353 153 2367 167
rect 2493 393 2507 407
rect 2593 613 2607 627
rect 2633 613 2647 627
rect 2653 593 2667 607
rect 2653 413 2667 427
rect 2533 373 2547 387
rect 2693 813 2707 827
rect 2753 833 2767 847
rect 2793 833 2807 847
rect 2773 813 2787 827
rect 2713 773 2727 787
rect 2773 693 2787 707
rect 2733 633 2747 647
rect 2713 613 2727 627
rect 3033 1233 3047 1247
rect 3013 1193 3027 1207
rect 2993 1133 3007 1147
rect 3233 1793 3247 1807
rect 3173 1613 3187 1627
rect 3213 1613 3227 1627
rect 3133 1593 3147 1607
rect 3153 1573 3167 1587
rect 3193 1593 3207 1607
rect 3233 1593 3247 1607
rect 3313 1913 3327 1927
rect 3393 2113 3407 2127
rect 3493 2693 3507 2707
rect 3533 2653 3547 2667
rect 3553 2653 3567 2667
rect 3513 2573 3527 2587
rect 3613 2753 3627 2767
rect 3573 2613 3587 2627
rect 3673 2473 3687 2487
rect 3493 2333 3507 2347
rect 3833 3533 3847 3547
rect 3833 3493 3847 3507
rect 3813 3473 3827 3487
rect 3813 3453 3827 3467
rect 3813 3213 3827 3227
rect 3913 4413 3927 4427
rect 3873 4193 3887 4207
rect 3893 4033 3907 4047
rect 3993 4493 4007 4507
rect 4013 4453 4027 4467
rect 4153 4773 4167 4787
rect 4113 4693 4127 4707
rect 4093 4653 4107 4667
rect 4073 4613 4087 4627
rect 4133 4593 4147 4607
rect 4033 4393 4047 4407
rect 3973 4233 3987 4247
rect 3973 4193 3987 4207
rect 4013 4193 4027 4207
rect 3993 4173 4007 4187
rect 4033 4073 4047 4087
rect 4513 5413 4527 5427
rect 4573 5413 4587 5427
rect 4613 5413 4627 5427
rect 4653 5413 4667 5427
rect 4593 5313 4607 5327
rect 4533 5233 4547 5247
rect 4473 5213 4487 5227
rect 4533 5213 4547 5227
rect 4493 5173 4507 5187
rect 4533 5153 4547 5167
rect 4573 5153 4587 5167
rect 4393 5133 4407 5147
rect 4433 5133 4447 5147
rect 4473 5133 4487 5147
rect 4513 5113 4527 5127
rect 4493 5053 4507 5067
rect 4433 5013 4447 5027
rect 4413 4913 4427 4927
rect 4453 4913 4467 4927
rect 4373 4893 4387 4907
rect 4413 4893 4427 4907
rect 4213 4693 4227 4707
rect 4293 4693 4307 4707
rect 4333 4693 4347 4707
rect 4313 4673 4327 4687
rect 4213 4653 4227 4667
rect 4353 4653 4367 4667
rect 4373 4653 4387 4667
rect 4173 4493 4187 4507
rect 4253 4493 4267 4507
rect 4113 4453 4127 4467
rect 4153 4453 4167 4467
rect 4153 4393 4167 4407
rect 4113 4193 4127 4207
rect 4133 4153 4147 4167
rect 4093 4113 4107 4127
rect 4053 4013 4067 4027
rect 3913 3993 3927 4007
rect 3953 3993 3967 4007
rect 4013 3993 4027 4007
rect 3893 3973 3907 3987
rect 3893 3933 3907 3947
rect 3933 3933 3947 3947
rect 3973 3713 3987 3727
rect 4093 3973 4107 3987
rect 4053 3953 4067 3967
rect 4033 3713 4047 3727
rect 4073 3713 4087 3727
rect 4013 3673 4027 3687
rect 3933 3653 3947 3667
rect 3993 3653 4007 3667
rect 3913 3613 3927 3627
rect 3913 3573 3927 3587
rect 3953 3493 3967 3507
rect 3933 3473 3947 3487
rect 4093 3693 4107 3707
rect 4053 3673 4067 3687
rect 4093 3613 4107 3627
rect 4033 3553 4047 3567
rect 4113 3593 4127 3607
rect 4113 3553 4127 3567
rect 4133 3553 4147 3567
rect 4073 3513 4087 3527
rect 4093 3493 4107 3507
rect 4133 3493 4147 3507
rect 3893 3453 3907 3467
rect 4053 3353 4067 3367
rect 3913 3333 3927 3347
rect 3853 3253 3867 3267
rect 3853 3193 3867 3207
rect 3793 3073 3807 3087
rect 3773 3053 3787 3067
rect 3793 3013 3807 3027
rect 3813 3013 3827 3027
rect 3833 2973 3847 2987
rect 3833 2953 3847 2967
rect 3773 2773 3787 2787
rect 3733 2753 3747 2767
rect 3893 3193 3907 3207
rect 3873 3153 3887 3167
rect 3853 2853 3867 2867
rect 3713 2733 3727 2747
rect 3753 2633 3767 2647
rect 3833 2733 3847 2747
rect 3753 2613 3767 2627
rect 3793 2613 3807 2627
rect 3713 2593 3727 2607
rect 3833 2593 3847 2607
rect 4033 3233 4047 3247
rect 4013 3213 4027 3227
rect 3993 3173 4007 3187
rect 3973 3113 3987 3127
rect 3973 3093 3987 3107
rect 3953 3053 3967 3067
rect 4013 3033 4027 3047
rect 4033 3033 4047 3047
rect 3993 3013 4007 3027
rect 3933 2953 3947 2967
rect 3973 2933 3987 2947
rect 3933 2813 3947 2827
rect 3873 2773 3887 2787
rect 3913 2773 3927 2787
rect 3853 2573 3867 2587
rect 3913 2733 3927 2747
rect 3893 2713 3907 2727
rect 3933 2613 3947 2627
rect 3953 2613 3967 2627
rect 3893 2573 3907 2587
rect 3853 2533 3867 2547
rect 3873 2533 3887 2547
rect 4033 3013 4047 3027
rect 4013 2933 4027 2947
rect 3993 2833 4007 2847
rect 4013 2753 4027 2767
rect 3973 2553 3987 2567
rect 3933 2513 3947 2527
rect 3713 2333 3727 2347
rect 3953 2333 3967 2347
rect 3873 2313 3887 2327
rect 3533 2273 3547 2287
rect 3693 2273 3707 2287
rect 3733 2273 3747 2287
rect 3433 2253 3447 2267
rect 3453 2173 3467 2187
rect 3433 2153 3447 2167
rect 3413 2093 3427 2107
rect 3373 2033 3387 2047
rect 3373 1853 3387 1867
rect 3253 1553 3267 1567
rect 3133 1513 3147 1527
rect 3273 1493 3287 1507
rect 3293 1393 3307 1407
rect 3113 1353 3127 1367
rect 3093 1333 3107 1347
rect 3153 1333 3167 1347
rect 3173 1333 3187 1347
rect 3253 1333 3267 1347
rect 3133 1313 3147 1327
rect 3113 1293 3127 1307
rect 3153 1193 3167 1207
rect 3073 1153 3087 1167
rect 3053 1133 3067 1147
rect 3113 1133 3127 1147
rect 3273 1313 3287 1327
rect 3293 1273 3307 1287
rect 3253 1233 3267 1247
rect 3013 1073 3027 1087
rect 2933 1053 2947 1067
rect 2913 993 2927 1007
rect 2873 853 2887 867
rect 2913 833 2927 847
rect 2893 773 2907 787
rect 2853 733 2867 747
rect 2813 653 2827 667
rect 2833 653 2847 667
rect 2873 653 2887 667
rect 2753 593 2767 607
rect 2793 433 2807 447
rect 2673 393 2687 407
rect 3053 853 3067 867
rect 3033 833 3047 847
rect 3153 1093 3167 1107
rect 2993 813 3007 827
rect 3073 813 3087 827
rect 3173 833 3187 847
rect 3133 793 3147 807
rect 3013 713 3027 727
rect 3193 813 3207 827
rect 3033 673 3047 687
rect 3093 673 3107 687
rect 3153 673 3167 687
rect 2993 633 3007 647
rect 2893 613 2907 627
rect 2933 613 2947 627
rect 2673 353 2687 367
rect 2753 373 2767 387
rect 2693 333 2707 347
rect 2773 353 2787 367
rect 3153 653 3167 667
rect 3113 633 3127 647
rect 3093 593 3107 607
rect 3293 1113 3307 1127
rect 3333 1793 3347 1807
rect 3453 2073 3467 2087
rect 3513 2073 3527 2087
rect 3553 2073 3567 2087
rect 3493 2053 3507 2067
rect 3453 2033 3467 2047
rect 3533 2033 3547 2047
rect 3633 2253 3647 2267
rect 3613 2113 3627 2127
rect 3833 2273 3847 2287
rect 3913 2273 3927 2287
rect 3953 2273 3967 2287
rect 3773 2093 3787 2107
rect 3593 2053 3607 2067
rect 3713 2033 3727 2047
rect 3793 2073 3807 2087
rect 3773 2053 3787 2067
rect 3813 2053 3827 2067
rect 3593 2013 3607 2027
rect 3753 2013 3767 2027
rect 3573 1953 3587 1967
rect 3513 1913 3527 1927
rect 3573 1913 3587 1927
rect 3513 1833 3527 1847
rect 3513 1813 3527 1827
rect 3413 1773 3427 1787
rect 3353 1653 3367 1667
rect 3533 1773 3547 1787
rect 3493 1753 3507 1767
rect 3753 1993 3767 2007
rect 3593 1773 3607 1787
rect 3473 1633 3487 1647
rect 3333 1613 3347 1627
rect 3553 1613 3567 1627
rect 3393 1573 3407 1587
rect 3453 1573 3467 1587
rect 3373 1353 3387 1367
rect 3473 1453 3487 1467
rect 3653 1793 3667 1807
rect 3793 1813 3807 1827
rect 3633 1773 3647 1787
rect 3673 1773 3687 1787
rect 3733 1773 3747 1787
rect 3773 1773 3787 1787
rect 3813 1773 3827 1787
rect 3613 1733 3627 1747
rect 3653 1733 3667 1747
rect 3633 1613 3647 1627
rect 3573 1573 3587 1587
rect 3593 1553 3607 1567
rect 3553 1393 3567 1407
rect 3433 1353 3447 1367
rect 3393 1333 3407 1347
rect 3513 1333 3527 1347
rect 3573 1333 3587 1347
rect 3413 1313 3427 1327
rect 3533 1313 3547 1327
rect 3393 1293 3407 1307
rect 3733 1653 3747 1667
rect 3673 1613 3687 1627
rect 3773 1633 3787 1647
rect 3753 1613 3767 1627
rect 3753 1593 3767 1607
rect 3733 1573 3747 1587
rect 3773 1573 3787 1587
rect 3713 1533 3727 1547
rect 3653 1513 3667 1527
rect 3613 1433 3627 1447
rect 4333 4473 4347 4487
rect 4253 4433 4267 4447
rect 4293 4453 4307 4467
rect 4273 4413 4287 4427
rect 4193 4213 4207 4227
rect 4253 4213 4267 4227
rect 4173 3913 4187 3927
rect 4173 3693 4187 3707
rect 4153 3473 4167 3487
rect 4173 3333 4187 3347
rect 4153 3253 4167 3267
rect 4093 3233 4107 3247
rect 4153 3213 4167 3227
rect 4073 3193 4087 3207
rect 4093 3093 4107 3107
rect 4133 3073 4147 3087
rect 4073 3013 4087 3027
rect 4053 2953 4067 2967
rect 4133 2973 4147 2987
rect 4213 4193 4227 4207
rect 4273 4173 4287 4187
rect 4253 4153 4267 4167
rect 4233 4133 4247 4147
rect 4213 4013 4227 4027
rect 4253 4013 4267 4027
rect 4273 3973 4287 3987
rect 4273 3953 4287 3967
rect 4233 3893 4247 3907
rect 4213 3693 4227 3707
rect 4253 3713 4267 3727
rect 4373 4473 4387 4487
rect 4433 4693 4447 4707
rect 4473 4693 4487 4707
rect 4473 4613 4487 4627
rect 4453 4493 4467 4507
rect 4353 4453 4367 4467
rect 4393 4453 4407 4467
rect 4393 4233 4407 4247
rect 4433 4213 4447 4227
rect 4413 4193 4427 4207
rect 4333 4153 4347 4167
rect 4413 4133 4427 4147
rect 4313 4033 4327 4047
rect 4353 4013 4367 4027
rect 4313 3973 4327 3987
rect 4233 3653 4247 3667
rect 4213 3513 4227 3527
rect 4253 3513 4267 3527
rect 4233 3493 4247 3507
rect 4373 3973 4387 3987
rect 4353 3953 4367 3967
rect 4433 4073 4447 4087
rect 4433 4013 4447 4027
rect 4433 3893 4447 3907
rect 4333 3833 4347 3847
rect 4313 3613 4327 3627
rect 4253 3473 4267 3487
rect 4213 3233 4227 3247
rect 4173 2833 4187 2847
rect 4193 2833 4207 2847
rect 4113 2813 4127 2827
rect 4133 2813 4147 2827
rect 4093 2793 4107 2807
rect 4053 2753 4067 2767
rect 4233 3193 4247 3207
rect 4293 3433 4307 3447
rect 4273 3213 4287 3227
rect 4313 3033 4327 3047
rect 4273 2993 4287 3007
rect 4313 2973 4327 2987
rect 4233 2813 4247 2827
rect 4213 2793 4227 2807
rect 4213 2773 4227 2787
rect 4193 2753 4207 2767
rect 4113 2733 4127 2747
rect 4093 2693 4107 2707
rect 4073 2673 4087 2687
rect 4033 2633 4047 2647
rect 4073 2633 4087 2647
rect 3993 2513 4007 2527
rect 4033 2513 4047 2527
rect 3853 2253 3867 2267
rect 3973 2253 3987 2267
rect 3893 2173 3907 2187
rect 4033 2233 4047 2247
rect 4053 2233 4067 2247
rect 4013 2093 4027 2107
rect 3913 2073 3927 2087
rect 3973 2073 3987 2087
rect 4073 2153 4087 2167
rect 4133 2653 4147 2667
rect 4113 2613 4127 2627
rect 4153 2613 4167 2627
rect 4113 2553 4127 2567
rect 4173 2593 4187 2607
rect 4173 2553 4187 2567
rect 4173 2513 4187 2527
rect 4253 2753 4267 2767
rect 4313 2753 4327 2767
rect 4293 2653 4307 2667
rect 4273 2573 4287 2587
rect 4253 2533 4267 2547
rect 4253 2513 4267 2527
rect 4353 3733 4367 3747
rect 4393 3713 4407 3727
rect 4473 4213 4487 4227
rect 4473 4013 4487 4027
rect 4573 4993 4587 5007
rect 4533 4853 4547 4867
rect 4633 5133 4647 5147
rect 4633 4953 4647 4967
rect 4593 4873 4607 4887
rect 4553 4813 4567 4827
rect 4633 4813 4647 4827
rect 4533 4693 4547 4707
rect 4573 4693 4587 4707
rect 4613 4673 4627 4687
rect 4733 5433 4747 5447
rect 4673 5393 4687 5407
rect 4753 5413 4767 5427
rect 4713 5373 4727 5387
rect 4773 5373 4787 5387
rect 4913 5613 4927 5627
rect 4953 5513 4967 5527
rect 4873 5413 4887 5427
rect 4853 5393 4867 5407
rect 4893 5393 4907 5407
rect 4753 5353 4767 5367
rect 4833 5353 4847 5367
rect 4673 5053 4687 5067
rect 4673 4953 4687 4967
rect 4713 4953 4727 4967
rect 4893 5353 4907 5367
rect 4853 4973 4867 4987
rect 4733 4933 4747 4947
rect 5033 5653 5047 5667
rect 5053 5613 5067 5627
rect 5053 5553 5067 5567
rect 5033 5513 5047 5527
rect 4993 5433 5007 5447
rect 4973 5193 4987 5207
rect 4913 5113 4927 5127
rect 5033 5133 5047 5147
rect 5213 5913 5227 5927
rect 5133 5873 5147 5887
rect 5193 5873 5207 5887
rect 5153 5653 5167 5667
rect 5173 5633 5187 5647
rect 5213 5613 5227 5627
rect 5253 5913 5267 5927
rect 5753 5953 5767 5967
rect 5573 5933 5587 5947
rect 5713 5933 5727 5947
rect 5373 5893 5387 5907
rect 5253 5653 5267 5667
rect 5313 5653 5327 5667
rect 5233 5513 5247 5527
rect 5113 5393 5127 5407
rect 5153 5453 5167 5467
rect 5193 5453 5207 5467
rect 5233 5453 5247 5467
rect 5213 5413 5227 5427
rect 5153 5393 5167 5407
rect 5173 5393 5187 5407
rect 5133 5173 5147 5187
rect 5153 5153 5167 5167
rect 5133 5113 5147 5127
rect 5053 5093 5067 5107
rect 4953 5073 4967 5087
rect 4933 4993 4947 5007
rect 4993 4973 5007 4987
rect 4953 4953 4967 4967
rect 5033 4953 5047 4967
rect 5013 4933 5027 4947
rect 4873 4913 4887 4927
rect 4893 4913 4907 4927
rect 4933 4913 4947 4927
rect 4973 4913 4987 4927
rect 4693 4853 4707 4867
rect 4833 4853 4847 4867
rect 4673 4673 4687 4687
rect 4553 4653 4567 4667
rect 4593 4653 4607 4667
rect 4553 4633 4567 4647
rect 4653 4653 4667 4667
rect 4673 4653 4687 4667
rect 4713 4653 4727 4667
rect 4633 4613 4647 4627
rect 4553 4493 4567 4507
rect 4573 4493 4587 4507
rect 4533 4453 4547 4467
rect 4613 4473 4627 4487
rect 4653 4453 4667 4467
rect 4753 4593 4767 4607
rect 4793 4553 4807 4567
rect 4833 4533 4847 4547
rect 4773 4493 4787 4507
rect 4713 4433 4727 4447
rect 4733 4413 4747 4427
rect 4593 4373 4607 4387
rect 4593 4213 4607 4227
rect 4673 4213 4687 4227
rect 4513 4193 4527 4207
rect 4553 4193 4567 4207
rect 4773 4393 4787 4407
rect 4753 4213 4767 4227
rect 4493 3973 4507 3987
rect 4373 3653 4387 3667
rect 4393 3613 4407 3627
rect 4353 3513 4367 3527
rect 4433 3593 4447 3607
rect 4413 3493 4427 3507
rect 4413 3433 4427 3447
rect 4393 3233 4407 3247
rect 4393 3173 4407 3187
rect 4373 3153 4387 3167
rect 4473 3633 4487 3647
rect 4453 3473 4467 3487
rect 4593 4073 4607 4087
rect 4533 3993 4547 4007
rect 4733 4173 4747 4187
rect 4693 4133 4707 4147
rect 4633 4053 4647 4067
rect 4613 3993 4627 4007
rect 4653 4033 4667 4047
rect 4733 3993 4747 4007
rect 4753 3973 4767 3987
rect 4633 3933 4647 3947
rect 4533 3913 4547 3927
rect 4593 3913 4607 3927
rect 4733 3913 4747 3927
rect 4713 3853 4727 3867
rect 4573 3833 4587 3847
rect 4553 3693 4567 3707
rect 4513 3553 4527 3567
rect 4513 3493 4527 3507
rect 4493 3473 4507 3487
rect 4533 3473 4547 3487
rect 4533 3453 4547 3467
rect 4473 3313 4487 3327
rect 4473 3233 4487 3247
rect 4513 3233 4527 3247
rect 4453 3213 4467 3227
rect 4433 3193 4447 3207
rect 4433 3173 4447 3187
rect 4373 3033 4387 3047
rect 4413 3033 4427 3047
rect 4353 3013 4367 3027
rect 4393 2933 4407 2947
rect 4493 3113 4507 3127
rect 4493 3073 4507 3087
rect 4433 2773 4447 2787
rect 4353 2753 4367 2767
rect 4413 2753 4427 2767
rect 4233 2313 4247 2327
rect 4433 2733 4447 2747
rect 4393 2673 4407 2687
rect 4453 2633 4467 2647
rect 4433 2593 4447 2607
rect 4393 2533 4407 2547
rect 4173 2293 4187 2307
rect 4273 2293 4287 2307
rect 4353 2293 4367 2307
rect 4233 2253 4247 2267
rect 4333 2253 4347 2267
rect 4313 2193 4327 2207
rect 4193 2153 4207 2167
rect 4293 2133 4307 2147
rect 4173 2113 4187 2127
rect 4093 2093 4107 2107
rect 3893 2053 3907 2067
rect 3913 2013 3927 2027
rect 3853 1813 3867 1827
rect 3973 1993 3987 2007
rect 4053 2053 4067 2067
rect 4013 1893 4027 1907
rect 3933 1873 3947 1887
rect 3953 1813 3967 1827
rect 3913 1753 3927 1767
rect 3913 1653 3927 1667
rect 3873 1613 3887 1627
rect 3993 1793 4007 1807
rect 3973 1773 3987 1787
rect 3953 1753 3967 1767
rect 4073 1993 4087 2007
rect 4053 1893 4067 1907
rect 4033 1633 4047 1647
rect 3993 1613 4007 1627
rect 3933 1593 3947 1607
rect 3893 1573 3907 1587
rect 3853 1553 3867 1567
rect 3873 1353 3887 1367
rect 3593 1313 3607 1327
rect 3633 1313 3647 1327
rect 3813 1313 3827 1327
rect 3833 1313 3847 1327
rect 3913 1313 3927 1327
rect 3453 1233 3467 1247
rect 3353 1193 3367 1207
rect 3333 1153 3347 1167
rect 3293 1073 3307 1087
rect 3313 1073 3327 1087
rect 3473 1193 3487 1207
rect 3513 1193 3527 1207
rect 3573 1193 3587 1207
rect 3453 1093 3467 1107
rect 3573 1133 3587 1147
rect 3613 1133 3627 1147
rect 3553 1113 3567 1127
rect 3493 1073 3507 1087
rect 3413 853 3427 867
rect 3253 833 3267 847
rect 3293 833 3307 847
rect 3353 833 3367 847
rect 3393 833 3407 847
rect 3313 813 3327 827
rect 3273 793 3287 807
rect 3413 793 3427 807
rect 3433 773 3447 787
rect 3353 753 3367 767
rect 3353 713 3367 727
rect 3313 693 3327 707
rect 3453 653 3467 667
rect 3213 613 3227 627
rect 3293 613 3307 627
rect 3333 613 3347 627
rect 3433 613 3447 627
rect 3173 593 3187 607
rect 3533 653 3547 667
rect 3473 573 3487 587
rect 3293 553 3307 567
rect 3193 433 3207 447
rect 3173 413 3187 427
rect 3193 413 3207 427
rect 2913 373 2927 387
rect 2893 353 2907 367
rect 2953 353 2967 367
rect 3073 353 3087 367
rect 2513 313 2527 327
rect 2753 313 2767 327
rect 2793 313 2807 327
rect 2933 313 2947 327
rect 3133 373 3147 387
rect 3113 353 3127 367
rect 3173 353 3187 367
rect 3253 393 3267 407
rect 3273 333 3287 347
rect 3093 313 3107 327
rect 2933 293 2947 307
rect 2973 293 2987 307
rect 2933 273 2947 287
rect 3053 273 3067 287
rect 2833 253 2847 267
rect 2753 213 2767 227
rect 2773 213 2787 227
rect 2533 193 2547 207
rect 2633 193 2647 207
rect 2513 173 2527 187
rect 2153 133 2167 147
rect 2213 133 2227 147
rect 2373 133 2387 147
rect 2413 133 2427 147
rect 2493 133 2507 147
rect 2473 113 2487 127
rect 2593 153 2607 167
rect 2613 153 2627 167
rect 2333 93 2347 107
rect 2673 153 2687 167
rect 2873 193 2887 207
rect 2913 193 2927 207
rect 2793 153 2807 167
rect 2893 133 2907 147
rect 3153 213 3167 227
rect 3033 193 3047 207
rect 3053 193 3067 207
rect 2993 153 3007 167
rect 3173 173 3187 187
rect 3153 153 3167 167
rect 3073 133 3087 147
rect 2893 113 2907 127
rect 3713 1293 3727 1307
rect 3673 1273 3687 1287
rect 3693 1193 3707 1207
rect 3593 1073 3607 1087
rect 3713 1133 3727 1147
rect 3733 1093 3747 1107
rect 3833 1233 3847 1247
rect 3853 1233 3867 1247
rect 3813 893 3827 907
rect 4133 2073 4147 2087
rect 4333 2113 4347 2127
rect 4193 2053 4207 2067
rect 4133 2033 4147 2047
rect 4153 2033 4167 2047
rect 4313 2053 4327 2067
rect 4313 2033 4327 2047
rect 4273 2013 4287 2027
rect 4353 1873 4367 1887
rect 4413 2273 4427 2287
rect 4693 3693 4707 3707
rect 4713 3693 4727 3707
rect 4593 3613 4607 3627
rect 4813 4173 4827 4187
rect 4793 4133 4807 4147
rect 4853 4373 4867 4387
rect 4833 4013 4847 4027
rect 4853 3973 4867 3987
rect 4893 4873 4907 4887
rect 4993 4693 5007 4707
rect 4973 4673 4987 4687
rect 5033 4593 5047 4607
rect 4933 4573 4947 4587
rect 4953 4553 4967 4567
rect 4913 4473 4927 4487
rect 5013 4493 5027 4507
rect 4993 4473 5007 4487
rect 4973 4453 4987 4467
rect 4933 4413 4947 4427
rect 4893 4393 4907 4407
rect 4913 4393 4927 4407
rect 4953 4173 4967 4187
rect 4973 4173 4987 4187
rect 4953 4093 4967 4107
rect 4973 4053 4987 4067
rect 4933 3993 4947 4007
rect 4913 3873 4927 3887
rect 4973 3873 4987 3887
rect 4873 3793 4887 3807
rect 4853 3753 4867 3767
rect 4913 3733 4927 3747
rect 4773 3653 4787 3667
rect 4793 3633 4807 3647
rect 4693 3593 4707 3607
rect 4793 3553 4807 3567
rect 4573 3473 4587 3487
rect 4773 3513 4787 3527
rect 4553 3173 4567 3187
rect 4553 3053 4567 3067
rect 4513 3013 4527 3027
rect 4633 3433 4647 3447
rect 4633 3373 4647 3387
rect 4593 3233 4607 3247
rect 4753 3373 4767 3387
rect 4693 3233 4707 3247
rect 4673 3213 4687 3227
rect 4733 3213 4747 3227
rect 4653 3193 4667 3207
rect 4713 3193 4727 3207
rect 4673 3093 4687 3107
rect 4613 3033 4627 3047
rect 4573 2933 4587 2947
rect 4553 2813 4567 2827
rect 4493 2773 4507 2787
rect 4593 2773 4607 2787
rect 4573 2753 4587 2767
rect 4493 2733 4507 2747
rect 4553 2713 4567 2727
rect 4673 3013 4687 3027
rect 4653 2993 4667 3007
rect 4693 2993 4707 3007
rect 4673 2953 4687 2967
rect 4633 2833 4647 2847
rect 4613 2673 4627 2687
rect 4553 2593 4567 2607
rect 4513 2573 4527 2587
rect 4593 2553 4607 2567
rect 4493 2533 4507 2547
rect 4533 2513 4547 2527
rect 4513 2493 4527 2507
rect 4433 2253 4447 2267
rect 4633 2313 4647 2327
rect 4533 2293 4547 2307
rect 4513 2213 4527 2227
rect 4393 2193 4407 2207
rect 4513 2153 4527 2167
rect 4433 2133 4447 2147
rect 4393 2073 4407 2087
rect 4413 2053 4427 2067
rect 4493 2093 4507 2107
rect 4453 2073 4467 2087
rect 4513 2053 4527 2067
rect 4493 2033 4507 2047
rect 4393 2013 4407 2027
rect 4473 1873 4487 1887
rect 4433 1853 4447 1867
rect 4213 1813 4227 1827
rect 4373 1813 4387 1827
rect 4133 1793 4147 1807
rect 4113 1753 4127 1767
rect 4073 1573 4087 1587
rect 4073 1513 4087 1527
rect 4053 1353 4067 1367
rect 3933 1273 3947 1287
rect 3933 1233 3947 1247
rect 3893 1153 3907 1167
rect 3893 1133 3907 1147
rect 3853 1113 3867 1127
rect 4013 1333 4027 1347
rect 4033 1313 4047 1327
rect 4073 1313 4087 1327
rect 3993 1213 4007 1227
rect 4033 1193 4047 1207
rect 4073 1173 4087 1187
rect 4153 1593 4167 1607
rect 4193 1593 4207 1607
rect 4133 1393 4147 1407
rect 4153 1313 4167 1327
rect 4193 1273 4207 1287
rect 4113 1153 4127 1167
rect 4153 1113 4167 1127
rect 4193 1113 4207 1127
rect 3873 1093 3887 1107
rect 3913 993 3927 1007
rect 4193 973 4207 987
rect 3693 853 3707 867
rect 3973 853 3987 867
rect 4273 1793 4287 1807
rect 4373 1793 4387 1807
rect 4473 1793 4487 1807
rect 4253 1773 4267 1787
rect 4293 1773 4307 1787
rect 4433 1773 4447 1787
rect 4493 1773 4507 1787
rect 4393 1753 4407 1767
rect 4353 1613 4367 1627
rect 4393 1593 4407 1607
rect 4333 1553 4347 1567
rect 4293 1333 4307 1347
rect 4413 1573 4427 1587
rect 4453 1613 4467 1627
rect 4433 1553 4447 1567
rect 4373 1513 4387 1527
rect 4413 1433 4427 1447
rect 4353 1373 4367 1387
rect 4253 1313 4267 1327
rect 4313 1313 4327 1327
rect 4253 1113 4267 1127
rect 4293 1113 4307 1127
rect 4333 1113 4347 1127
rect 4273 1093 4287 1107
rect 4293 1073 4307 1087
rect 4253 1033 4267 1047
rect 3573 833 3587 847
rect 3673 833 3687 847
rect 3713 833 3727 847
rect 3813 833 3827 847
rect 3653 813 3667 827
rect 3593 793 3607 807
rect 3693 793 3707 807
rect 3793 753 3807 767
rect 3773 713 3787 727
rect 3753 673 3767 687
rect 3853 833 3867 847
rect 3893 833 3907 847
rect 3833 673 3847 687
rect 3773 633 3787 647
rect 3833 633 3847 647
rect 3613 593 3627 607
rect 3793 613 3807 627
rect 3953 813 3967 827
rect 3913 713 3927 727
rect 4073 833 4087 847
rect 4113 833 4127 847
rect 3973 693 3987 707
rect 3953 633 3967 647
rect 3853 613 3867 627
rect 3933 613 3947 627
rect 3653 573 3667 587
rect 3553 553 3567 567
rect 3513 473 3527 487
rect 3453 393 3467 407
rect 3333 373 3347 387
rect 3373 353 3387 367
rect 3393 333 3407 347
rect 3353 213 3367 227
rect 3373 193 3387 207
rect 3313 173 3327 187
rect 3353 153 3367 167
rect 3293 133 3307 147
rect 3333 133 3347 147
rect 3453 373 3467 387
rect 3453 313 3467 327
rect 4133 793 4147 807
rect 3973 613 3987 627
rect 4093 633 4107 647
rect 4053 613 4067 627
rect 4093 613 4107 627
rect 4213 833 4227 847
rect 4273 833 4287 847
rect 4233 793 4247 807
rect 4233 773 4247 787
rect 4233 713 4247 727
rect 4193 673 4207 687
rect 4213 633 4227 647
rect 4153 613 4167 627
rect 4033 453 4047 467
rect 3913 433 3927 447
rect 4173 593 4187 607
rect 4153 453 4167 467
rect 4073 413 4087 427
rect 4093 413 4107 427
rect 4133 413 4147 427
rect 3513 393 3527 407
rect 3493 273 3507 287
rect 3473 193 3487 207
rect 3433 173 3447 187
rect 3453 153 3467 167
rect 4013 373 4027 387
rect 4033 373 4047 387
rect 3533 353 3547 367
rect 3573 353 3587 367
rect 3613 353 3627 367
rect 3693 353 3707 367
rect 3733 353 3747 367
rect 3833 353 3847 367
rect 3553 333 3567 347
rect 3593 313 3607 327
rect 3613 253 3627 267
rect 3713 313 3727 327
rect 3873 293 3887 307
rect 3673 233 3687 247
rect 3813 213 3827 227
rect 3613 173 3627 187
rect 3653 153 3667 167
rect 3693 153 3707 167
rect 3773 153 3787 167
rect 3633 133 3647 147
rect 3673 133 3687 147
rect 3933 333 3947 347
rect 3933 293 3947 307
rect 3893 253 3907 267
rect 3913 253 3927 267
rect 3913 173 3927 187
rect 4053 333 4067 347
rect 4053 233 4067 247
rect 4233 613 4247 627
rect 4193 553 4207 567
rect 4253 533 4267 547
rect 4253 433 4267 447
rect 4173 393 4187 407
rect 4213 373 4227 387
rect 4113 313 4127 327
rect 4273 333 4287 347
rect 4413 1313 4427 1327
rect 4393 1273 4407 1287
rect 4433 1133 4447 1147
rect 4373 1113 4387 1127
rect 4373 1073 4387 1087
rect 4353 953 4367 967
rect 4413 933 4427 947
rect 4373 853 4387 867
rect 4333 833 4347 847
rect 4313 813 4327 827
rect 4353 813 4367 827
rect 4393 793 4407 807
rect 4373 693 4387 707
rect 4553 2273 4567 2287
rect 4633 2193 4647 2207
rect 4573 2153 4587 2167
rect 4633 2113 4647 2127
rect 4573 2093 4587 2107
rect 4633 2093 4647 2107
rect 4613 2073 4627 2087
rect 4553 2053 4567 2067
rect 4593 2053 4607 2067
rect 4633 2053 4647 2067
rect 4573 1813 4587 1827
rect 4533 1613 4547 1627
rect 4513 1553 4527 1567
rect 4553 1453 4567 1467
rect 4513 1353 4527 1367
rect 4473 1313 4487 1327
rect 4553 1313 4567 1327
rect 4533 1193 4547 1207
rect 4473 1173 4487 1187
rect 4553 1113 4567 1127
rect 4553 1093 4567 1107
rect 4473 993 4487 1007
rect 4453 873 4467 887
rect 4453 853 4467 867
rect 4453 713 4467 727
rect 4533 913 4547 927
rect 4493 853 4507 867
rect 4513 813 4527 827
rect 4433 653 4447 667
rect 4393 613 4407 627
rect 4353 593 4367 607
rect 4313 573 4327 587
rect 4453 633 4467 647
rect 4353 413 4367 427
rect 4393 413 4407 427
rect 4433 413 4447 427
rect 4313 333 4327 347
rect 4293 293 4307 307
rect 4113 253 4127 267
rect 4193 253 4207 267
rect 4093 213 4107 227
rect 3793 133 3807 147
rect 3873 133 3887 147
rect 4053 133 4067 147
rect 4153 213 4167 227
rect 4193 153 4207 167
rect 4273 153 4287 167
rect 4173 133 4187 147
rect 3693 113 3707 127
rect 3833 113 3847 127
rect 4053 113 4067 127
rect 4333 313 4347 327
rect 4353 173 4367 187
rect 4433 373 4447 387
rect 4513 693 4527 707
rect 4493 613 4507 627
rect 4473 413 4487 427
rect 4453 353 4467 367
rect 4513 353 4527 367
rect 4493 333 4507 347
rect 4453 313 4467 327
rect 4433 293 4447 307
rect 4413 173 4427 187
rect 4513 193 4527 207
rect 4453 153 4467 167
rect 4513 133 4527 147
rect 4393 113 4407 127
rect 3233 93 3247 107
rect 3473 93 3487 107
rect 2593 73 2607 87
rect 2133 33 2147 47
rect 4633 1773 4647 1787
rect 4593 1613 4607 1627
rect 4693 2753 4707 2767
rect 4733 2713 4747 2727
rect 4893 3693 4907 3707
rect 4933 3693 4947 3707
rect 5013 4393 5027 4407
rect 5133 5053 5147 5067
rect 5113 5013 5127 5027
rect 5193 5373 5207 5387
rect 5173 4953 5187 4967
rect 5073 4913 5087 4927
rect 5153 4913 5167 4927
rect 5053 4533 5067 4547
rect 5093 4673 5107 4687
rect 5133 4673 5147 4687
rect 5173 4673 5187 4687
rect 5113 4653 5127 4667
rect 5153 4573 5167 4587
rect 5073 4493 5087 4507
rect 5133 4473 5147 4487
rect 5213 5173 5227 5187
rect 5213 5113 5227 5127
rect 5273 5633 5287 5647
rect 5333 5613 5347 5627
rect 5293 5593 5307 5607
rect 5273 5573 5287 5587
rect 5293 5453 5307 5467
rect 5253 5413 5267 5427
rect 5273 5413 5287 5427
rect 5333 5413 5347 5427
rect 5313 5393 5327 5407
rect 5293 5173 5307 5187
rect 5253 5133 5267 5147
rect 5273 5113 5287 5127
rect 5293 5073 5307 5087
rect 5273 5033 5287 5047
rect 5213 4953 5227 4967
rect 5253 4953 5267 4967
rect 5253 4653 5267 4667
rect 5193 4573 5207 4587
rect 5073 4453 5087 4467
rect 5053 4433 5067 4447
rect 5093 4433 5107 4447
rect 5093 4413 5107 4427
rect 5053 4233 5067 4247
rect 5013 4033 5027 4047
rect 5093 4213 5107 4227
rect 5213 4473 5227 4487
rect 5153 4433 5167 4447
rect 5153 4393 5167 4407
rect 5133 4173 5147 4187
rect 5233 4453 5247 4467
rect 5453 5693 5467 5707
rect 5493 5913 5507 5927
rect 5473 5673 5487 5687
rect 5653 5893 5667 5907
rect 5553 5873 5567 5887
rect 5633 5873 5647 5887
rect 5673 5873 5687 5887
rect 5553 5673 5567 5687
rect 5513 5653 5527 5667
rect 5493 5613 5507 5627
rect 5433 5593 5447 5607
rect 5473 5593 5487 5607
rect 5433 5553 5447 5567
rect 5393 5473 5407 5487
rect 5413 5473 5427 5487
rect 5393 5433 5407 5447
rect 5453 5473 5467 5487
rect 5433 5433 5447 5447
rect 5533 5633 5547 5647
rect 5513 5593 5527 5607
rect 5613 5653 5627 5667
rect 5573 5633 5587 5647
rect 5613 5593 5627 5607
rect 5413 5393 5427 5407
rect 5473 5393 5487 5407
rect 5493 5393 5507 5407
rect 5393 5353 5407 5367
rect 5353 5173 5367 5187
rect 5373 5173 5387 5187
rect 5393 5153 5407 5167
rect 5433 5153 5447 5167
rect 5413 5133 5427 5147
rect 5393 5113 5407 5127
rect 5373 5093 5387 5107
rect 5353 5073 5367 5087
rect 5313 5033 5327 5047
rect 5333 4973 5347 4987
rect 5353 4913 5367 4927
rect 5373 4693 5387 4707
rect 5373 4673 5387 4687
rect 5293 4593 5307 4607
rect 5313 4593 5327 4607
rect 5293 4573 5307 4587
rect 5273 4393 5287 4407
rect 5373 4473 5387 4487
rect 5333 4453 5347 4467
rect 5373 4433 5387 4447
rect 5313 4413 5327 4427
rect 5193 4373 5207 4387
rect 5173 4333 5187 4347
rect 5173 4133 5187 4147
rect 5053 3973 5067 3987
rect 4993 3833 5007 3847
rect 5033 3713 5047 3727
rect 4993 3693 5007 3707
rect 4933 3673 4947 3687
rect 4973 3673 4987 3687
rect 4893 3653 4907 3667
rect 4853 3533 4867 3547
rect 4873 3473 4887 3487
rect 4833 3313 4847 3327
rect 4813 3273 4827 3287
rect 4853 3273 4867 3287
rect 4853 3233 4867 3247
rect 4813 3093 4827 3107
rect 4793 3053 4807 3067
rect 4833 3073 4847 3087
rect 4853 3033 4867 3047
rect 4873 3033 4887 3047
rect 4833 3013 4847 3027
rect 4773 2993 4787 3007
rect 4853 2993 4867 3007
rect 4793 2793 4807 2807
rect 4833 2753 4847 2767
rect 4813 2733 4827 2747
rect 4773 2713 4787 2727
rect 4753 2693 4767 2707
rect 4693 2673 4707 2687
rect 4673 2553 4687 2567
rect 4713 2573 4727 2587
rect 4833 2573 4847 2587
rect 4813 2293 4827 2307
rect 4753 2233 4767 2247
rect 4773 2213 4787 2227
rect 4753 2113 4767 2127
rect 4713 2093 4727 2107
rect 4693 2073 4707 2087
rect 4673 1813 4687 1827
rect 4673 1733 4687 1747
rect 4733 2053 4747 2067
rect 4793 2053 4807 2067
rect 4753 1773 4767 1787
rect 4693 1693 4707 1707
rect 4613 1593 4627 1607
rect 4653 1593 4667 1607
rect 4593 1013 4607 1027
rect 4593 953 4607 967
rect 4573 793 4587 807
rect 4553 693 4567 707
rect 4753 1653 4767 1667
rect 4953 3533 4967 3547
rect 5033 3513 5047 3527
rect 5013 3473 5027 3487
rect 5033 3473 5047 3487
rect 4973 3453 4987 3467
rect 5013 3293 5027 3307
rect 4993 3213 5007 3227
rect 5033 3193 5047 3207
rect 5153 3973 5167 3987
rect 5273 4213 5287 4227
rect 5233 4193 5247 4207
rect 5213 4153 5227 4167
rect 5233 4153 5247 4167
rect 5273 4153 5287 4167
rect 5253 4133 5267 4147
rect 5213 3993 5227 4007
rect 5233 3993 5247 4007
rect 5233 3973 5247 3987
rect 5213 3853 5227 3867
rect 5213 3813 5227 3827
rect 5193 3733 5207 3747
rect 5133 3713 5147 3727
rect 5173 3673 5187 3687
rect 5093 3653 5107 3667
rect 5073 3533 5087 3547
rect 5133 3533 5147 3547
rect 5073 3513 5087 3527
rect 5113 3513 5127 3527
rect 5093 3493 5107 3507
rect 5093 3453 5107 3467
rect 5113 3273 5127 3287
rect 5073 3253 5087 3267
rect 5133 3253 5147 3267
rect 5153 3213 5167 3227
rect 5133 3193 5147 3207
rect 4973 3113 4987 3127
rect 4993 3053 5007 3067
rect 4933 3033 4947 3047
rect 4973 3033 4987 3047
rect 4893 2993 4907 3007
rect 4893 2853 4907 2867
rect 4973 2633 4987 2647
rect 5133 3153 5147 3167
rect 5073 3053 5087 3067
rect 5033 3033 5047 3047
rect 5193 3633 5207 3647
rect 5413 4953 5427 4967
rect 5413 4853 5427 4867
rect 5473 5113 5487 5127
rect 5553 5413 5567 5427
rect 5533 5393 5547 5407
rect 5573 5373 5587 5387
rect 5533 5153 5547 5167
rect 5513 5113 5527 5127
rect 5553 5113 5567 5127
rect 5493 5053 5507 5067
rect 5553 5093 5567 5107
rect 5533 4953 5547 4967
rect 5513 4873 5527 4887
rect 5473 4693 5487 4707
rect 5513 4673 5527 4687
rect 5433 4653 5447 4667
rect 5493 4653 5507 4667
rect 5413 4613 5427 4627
rect 5393 4333 5407 4347
rect 5353 4233 5367 4247
rect 5413 4233 5427 4247
rect 5333 4213 5347 4227
rect 5313 4153 5327 4167
rect 5333 4113 5347 4127
rect 5293 4073 5307 4087
rect 5313 3973 5327 3987
rect 5333 3953 5347 3967
rect 5293 3833 5307 3847
rect 5273 3813 5287 3827
rect 5293 3793 5307 3807
rect 5273 3753 5287 3767
rect 5273 3713 5287 3727
rect 5233 3673 5247 3687
rect 5253 3653 5267 3667
rect 5313 3753 5327 3767
rect 5373 4213 5387 4227
rect 5413 4213 5427 4227
rect 5393 4193 5407 4207
rect 5533 4633 5547 4647
rect 5453 4613 5467 4627
rect 5533 4613 5547 4627
rect 5493 4473 5507 4487
rect 5633 5493 5647 5507
rect 5633 5433 5647 5447
rect 5613 5093 5627 5107
rect 5593 5073 5607 5087
rect 5633 5033 5647 5047
rect 5573 4953 5587 4967
rect 5633 4953 5647 4967
rect 5633 4933 5647 4947
rect 5573 4693 5587 4707
rect 5673 5613 5687 5627
rect 5733 5893 5747 5907
rect 5713 5593 5727 5607
rect 5713 5573 5727 5587
rect 5693 5513 5707 5527
rect 5673 5453 5687 5467
rect 5653 4713 5667 4727
rect 5633 4613 5647 4627
rect 5653 4593 5667 4607
rect 5613 4453 5627 4467
rect 5633 4433 5647 4447
rect 5533 4233 5547 4247
rect 5513 4213 5527 4227
rect 5473 4113 5487 4127
rect 5473 4093 5487 4107
rect 5433 4073 5447 4087
rect 5453 4033 5467 4047
rect 5373 3993 5387 4007
rect 5373 3953 5387 3967
rect 5433 3853 5447 3867
rect 5373 3713 5387 3727
rect 5393 3693 5407 3707
rect 5413 3673 5427 3687
rect 5453 3593 5467 3607
rect 5353 3533 5367 3547
rect 5433 3533 5447 3547
rect 5393 3513 5407 3527
rect 5353 3493 5367 3507
rect 5313 3453 5327 3467
rect 5353 3453 5367 3467
rect 5333 3433 5347 3447
rect 5333 3393 5347 3407
rect 5213 3373 5227 3387
rect 5253 3373 5267 3387
rect 5293 3373 5307 3387
rect 5313 3313 5327 3327
rect 5213 3293 5227 3307
rect 5253 3293 5267 3307
rect 5293 3233 5307 3247
rect 5273 3213 5287 3227
rect 5233 3173 5247 3187
rect 5213 3113 5227 3127
rect 5173 3073 5187 3087
rect 5013 2733 5027 2747
rect 5073 2933 5087 2947
rect 4873 2573 4887 2587
rect 4913 2573 4927 2587
rect 4933 2573 4947 2587
rect 4993 2573 5007 2587
rect 4873 2513 4887 2527
rect 4853 2273 4867 2287
rect 4893 2333 4907 2347
rect 4913 2293 4927 2307
rect 4933 2273 4947 2287
rect 4873 2253 4887 2267
rect 4873 2093 4887 2107
rect 4893 2093 4907 2107
rect 4853 2033 4867 2047
rect 4873 1833 4887 1847
rect 4893 1813 4907 1827
rect 4913 1793 4927 1807
rect 4853 1773 4867 1787
rect 4893 1753 4907 1767
rect 4793 1593 4807 1607
rect 4833 1593 4847 1607
rect 4653 1573 4667 1587
rect 4693 1573 4707 1587
rect 4773 1573 4787 1587
rect 4793 1553 4807 1567
rect 4673 1513 4687 1527
rect 4633 1453 4647 1467
rect 4673 1353 4687 1367
rect 4633 1333 4647 1347
rect 4653 1313 4667 1327
rect 4693 1313 4707 1327
rect 4773 1313 4787 1327
rect 4633 1273 4647 1287
rect 4753 1273 4767 1287
rect 4693 1233 4707 1247
rect 4713 1133 4727 1147
rect 4633 1113 4647 1127
rect 4673 1113 4687 1127
rect 4753 1113 4767 1127
rect 4693 1013 4707 1027
rect 4733 993 4747 1007
rect 4613 913 4627 927
rect 4913 1573 4927 1587
rect 4993 2293 5007 2307
rect 4973 2273 4987 2287
rect 4953 2193 4967 2207
rect 4973 2153 4987 2167
rect 4953 2093 4967 2107
rect 5033 2633 5047 2647
rect 5053 2633 5067 2647
rect 5073 2633 5087 2647
rect 5033 2573 5047 2587
rect 5033 2553 5047 2567
rect 5033 2313 5047 2327
rect 5013 2113 5027 2127
rect 5073 2553 5087 2567
rect 5153 2733 5167 2747
rect 5133 2533 5147 2547
rect 5093 2313 5107 2327
rect 5053 2293 5067 2307
rect 5073 2253 5087 2267
rect 5253 3033 5267 3047
rect 5373 3393 5387 3407
rect 5353 3153 5367 3167
rect 5373 3113 5387 3127
rect 5353 3073 5367 3087
rect 5333 3033 5347 3047
rect 5233 2733 5247 2747
rect 5273 2733 5287 2747
rect 5313 2733 5327 2747
rect 5313 2713 5327 2727
rect 5193 2593 5207 2607
rect 5253 2573 5267 2587
rect 5193 2553 5207 2567
rect 5413 3193 5427 3207
rect 5413 3033 5427 3047
rect 5413 2773 5427 2787
rect 5493 3993 5507 4007
rect 5553 3753 5567 3767
rect 5553 3733 5567 3747
rect 5533 3673 5547 3687
rect 5493 3533 5507 3547
rect 5533 3513 5547 3527
rect 5473 3493 5487 3507
rect 5513 3493 5527 3507
rect 5493 3373 5507 3387
rect 5533 3233 5547 3247
rect 5673 4233 5687 4247
rect 5613 4193 5627 4207
rect 5673 4173 5687 4187
rect 5653 4153 5667 4167
rect 5673 4093 5687 4107
rect 5713 4573 5727 4587
rect 5933 5913 5947 5927
rect 5773 5873 5787 5887
rect 5813 5873 5827 5887
rect 5753 5513 5767 5527
rect 5933 5573 5947 5587
rect 5793 5553 5807 5567
rect 5833 5433 5847 5447
rect 5813 4933 5827 4947
rect 5813 4713 5827 4727
rect 5773 4653 5787 4667
rect 5813 4633 5827 4647
rect 5753 4573 5767 4587
rect 5793 4473 5807 4487
rect 5733 4453 5747 4467
rect 5753 4433 5767 4447
rect 5733 4293 5747 4307
rect 5733 4153 5747 4167
rect 5593 4013 5607 4027
rect 5693 4013 5707 4027
rect 5673 3993 5687 4007
rect 5713 3993 5727 4007
rect 5653 3973 5667 3987
rect 5693 3973 5707 3987
rect 5693 3953 5707 3967
rect 5593 3593 5607 3607
rect 5673 3733 5687 3747
rect 5653 3673 5667 3687
rect 5673 3593 5687 3607
rect 5633 3533 5647 3547
rect 5713 3933 5727 3947
rect 5713 3713 5727 3727
rect 5773 4293 5787 4307
rect 5813 4173 5827 4187
rect 5773 4153 5787 4167
rect 5813 4153 5827 4167
rect 5753 4133 5767 4147
rect 5793 4133 5807 4147
rect 5793 4113 5807 4127
rect 5773 4013 5787 4027
rect 5793 4013 5807 4027
rect 5853 4933 5867 4947
rect 5913 4933 5927 4947
rect 5893 4653 5907 4667
rect 5853 4633 5867 4647
rect 5853 4213 5867 4227
rect 5833 3993 5847 4007
rect 5753 3973 5767 3987
rect 5793 3973 5807 3987
rect 5833 3973 5847 3987
rect 5813 3953 5827 3967
rect 5833 3933 5847 3947
rect 5773 3753 5787 3767
rect 5813 3753 5827 3767
rect 5753 3733 5767 3747
rect 5813 3733 5827 3747
rect 5793 3713 5807 3727
rect 5793 3693 5807 3707
rect 5693 3493 5707 3507
rect 5613 3393 5627 3407
rect 5593 3253 5607 3267
rect 5573 3213 5587 3227
rect 5493 3193 5507 3207
rect 5553 3173 5567 3187
rect 5453 3113 5467 3127
rect 5573 3113 5587 3127
rect 5553 3093 5567 3107
rect 5513 3013 5527 3027
rect 5613 3233 5627 3247
rect 5653 3233 5667 3247
rect 5653 3193 5667 3207
rect 5613 3113 5627 3127
rect 5693 3173 5707 3187
rect 5673 3013 5687 3027
rect 5613 2853 5627 2867
rect 5413 2633 5427 2647
rect 5393 2593 5407 2607
rect 5173 2333 5187 2347
rect 5193 2293 5207 2307
rect 5153 2273 5167 2287
rect 5093 2233 5107 2247
rect 5133 2233 5147 2247
rect 5073 2073 5087 2087
rect 4993 1813 5007 1827
rect 5033 2053 5047 2067
rect 5033 1793 5047 1807
rect 5053 1773 5067 1787
rect 5013 1753 5027 1767
rect 5033 1653 5047 1667
rect 4973 1593 4987 1607
rect 4933 1553 4947 1567
rect 4833 1533 4847 1547
rect 4873 1533 4887 1547
rect 4913 1373 4927 1387
rect 4953 1373 4967 1387
rect 4893 1313 4907 1327
rect 4953 1293 4967 1307
rect 4853 1273 4867 1287
rect 4933 1173 4947 1187
rect 4813 1113 4827 1127
rect 4993 1573 5007 1587
rect 5133 2153 5147 2167
rect 5213 2273 5227 2287
rect 5173 2253 5187 2267
rect 5193 2253 5207 2267
rect 5333 2313 5347 2327
rect 5333 2253 5347 2267
rect 5393 2253 5407 2267
rect 5173 2173 5187 2187
rect 5233 2173 5247 2187
rect 5253 2173 5267 2187
rect 5333 2173 5347 2187
rect 5373 2173 5387 2187
rect 5153 2133 5167 2147
rect 5113 2073 5127 2087
rect 5153 2073 5167 2087
rect 5233 2133 5247 2147
rect 5193 2073 5207 2087
rect 5273 2093 5287 2107
rect 5133 1793 5147 1807
rect 5153 1653 5167 1667
rect 5253 2053 5267 2067
rect 5293 2053 5307 2067
rect 5373 2153 5387 2167
rect 5353 2093 5367 2107
rect 5333 1973 5347 1987
rect 5233 1813 5247 1827
rect 5293 1793 5307 1807
rect 5233 1773 5247 1787
rect 5273 1773 5287 1787
rect 5313 1773 5327 1787
rect 5193 1693 5207 1707
rect 5213 1693 5227 1707
rect 5193 1673 5207 1687
rect 5173 1633 5187 1647
rect 5173 1573 5187 1587
rect 5253 1633 5267 1647
rect 5133 1393 5147 1407
rect 5193 1353 5207 1367
rect 5093 1333 5107 1347
rect 4993 1313 5007 1327
rect 5033 1313 5047 1327
rect 5073 1313 5087 1327
rect 5093 1313 5107 1327
rect 5133 1313 5147 1327
rect 5173 1313 5187 1327
rect 5053 1293 5067 1307
rect 5013 1233 5027 1247
rect 4933 1113 4947 1127
rect 4973 1113 4987 1127
rect 5013 1133 5027 1147
rect 4993 1093 5007 1107
rect 4833 1073 4847 1087
rect 4873 973 4887 987
rect 4673 853 4687 867
rect 4793 853 4807 867
rect 4833 853 4847 867
rect 4653 833 4667 847
rect 4733 833 4747 847
rect 4633 813 4647 827
rect 4713 813 4727 827
rect 4813 813 4827 827
rect 4613 773 4627 787
rect 4653 753 4667 767
rect 4673 673 4687 687
rect 4593 613 4607 627
rect 4633 373 4647 387
rect 4593 333 4607 347
rect 4653 333 4667 347
rect 4653 313 4667 327
rect 4573 293 4587 307
rect 4613 293 4627 307
rect 4573 233 4587 247
rect 4553 133 4567 147
rect 4593 113 4607 127
rect 4633 113 4647 127
rect 4533 13 4547 27
rect 4613 13 4627 27
rect 4773 773 4787 787
rect 4793 633 4807 647
rect 4693 553 4707 567
rect 5113 1293 5127 1307
rect 5153 1273 5167 1287
rect 5153 1193 5167 1207
rect 5153 1153 5167 1167
rect 5133 1133 5147 1147
rect 5113 1113 5127 1127
rect 5093 1053 5107 1067
rect 5073 933 5087 947
rect 4913 873 4927 887
rect 4953 833 4967 847
rect 5053 833 5067 847
rect 5093 833 5107 847
rect 4933 813 4947 827
rect 5073 813 5087 827
rect 4893 793 4907 807
rect 5033 793 5047 807
rect 5213 1333 5227 1347
rect 5233 1333 5247 1347
rect 5213 1173 5227 1187
rect 5313 1613 5327 1627
rect 5393 2053 5407 2067
rect 5553 2733 5567 2747
rect 5673 2733 5687 2747
rect 5593 2573 5607 2587
rect 5493 2553 5507 2567
rect 5513 2533 5527 2547
rect 5553 2533 5567 2547
rect 5613 2533 5627 2547
rect 5453 2513 5467 2527
rect 5433 2373 5447 2387
rect 5473 2373 5487 2387
rect 5453 2293 5467 2307
rect 5453 2193 5467 2207
rect 5353 1673 5367 1687
rect 5373 1613 5387 1627
rect 5333 1593 5347 1607
rect 5353 1593 5367 1607
rect 5333 1553 5347 1567
rect 5333 1393 5347 1407
rect 5273 1333 5287 1347
rect 5313 1333 5327 1347
rect 5293 1313 5307 1327
rect 5313 1173 5327 1187
rect 5253 1133 5267 1147
rect 5233 1113 5247 1127
rect 5273 1113 5287 1127
rect 5213 1093 5227 1107
rect 5173 1073 5187 1087
rect 5213 1073 5227 1087
rect 5153 1053 5167 1067
rect 5133 1013 5147 1027
rect 5133 833 5147 847
rect 5113 693 5127 707
rect 4853 633 4867 647
rect 5093 673 5107 687
rect 5113 673 5127 687
rect 4873 613 4887 627
rect 4873 433 4887 447
rect 4973 613 4987 627
rect 5053 433 5067 447
rect 4813 373 4827 387
rect 4753 353 4767 367
rect 4793 353 4807 367
rect 4693 333 4707 347
rect 4733 333 4747 347
rect 4813 333 4827 347
rect 4773 313 4787 327
rect 4693 233 4707 247
rect 4913 393 4927 407
rect 5013 393 5027 407
rect 4853 353 4867 367
rect 5033 353 5047 367
rect 4933 333 4947 347
rect 4893 313 4907 327
rect 5033 313 5047 327
rect 4873 293 4887 307
rect 4733 153 4747 167
rect 4713 133 4727 147
rect 4753 133 4767 147
rect 5193 893 5207 907
rect 5153 633 5167 647
rect 5213 633 5227 647
rect 5173 613 5187 627
rect 5133 593 5147 607
rect 5193 433 5207 447
rect 5113 393 5127 407
rect 5153 313 5167 327
rect 5233 273 5247 287
rect 5093 193 5107 207
rect 5133 193 5147 207
rect 4973 173 4987 187
rect 5093 173 5107 187
rect 5013 133 5027 147
rect 5293 1093 5307 1107
rect 5293 1033 5307 1047
rect 5273 613 5287 627
rect 5293 373 5307 387
rect 5273 313 5287 327
rect 5353 1333 5367 1347
rect 5353 1293 5367 1307
rect 5353 1173 5367 1187
rect 5333 1133 5347 1147
rect 5413 1553 5427 1567
rect 5533 2333 5547 2347
rect 5493 2313 5507 2327
rect 5573 2293 5587 2307
rect 5773 3533 5787 3547
rect 5813 3673 5827 3687
rect 5793 3473 5807 3487
rect 5733 3393 5747 3407
rect 5793 3253 5807 3267
rect 5733 3233 5747 3247
rect 5773 3213 5787 3227
rect 5773 3193 5787 3207
rect 5793 3033 5807 3047
rect 5773 2913 5787 2927
rect 5733 2853 5747 2867
rect 5733 2773 5747 2787
rect 5793 2733 5807 2747
rect 5773 2713 5787 2727
rect 5753 2573 5767 2587
rect 5793 2553 5807 2567
rect 5713 2293 5727 2307
rect 5773 2293 5787 2307
rect 5613 2273 5627 2287
rect 5653 2273 5667 2287
rect 5673 2273 5687 2287
rect 5713 2273 5727 2287
rect 5473 2073 5487 2087
rect 5453 2053 5467 2067
rect 5473 2053 5487 2067
rect 5513 2053 5527 2067
rect 5453 1773 5467 1787
rect 5513 1973 5527 1987
rect 5513 1793 5527 1807
rect 5513 1753 5527 1767
rect 5493 1733 5507 1747
rect 5493 1673 5507 1687
rect 5473 1613 5487 1627
rect 5453 1593 5467 1607
rect 5433 1373 5447 1387
rect 5453 1353 5467 1367
rect 5413 1333 5427 1347
rect 5493 1313 5507 1327
rect 5473 1293 5487 1307
rect 5433 1233 5447 1247
rect 5453 1193 5467 1207
rect 5393 1153 5407 1167
rect 5413 1133 5427 1147
rect 5393 1113 5407 1127
rect 5333 1093 5347 1107
rect 5353 933 5367 947
rect 5373 893 5387 907
rect 5333 753 5347 767
rect 5373 673 5387 687
rect 5333 633 5347 647
rect 5573 2233 5587 2247
rect 5633 2253 5647 2267
rect 5653 2253 5667 2267
rect 5593 2093 5607 2107
rect 5593 2073 5607 2087
rect 5573 1833 5587 1847
rect 5533 1613 5547 1627
rect 5593 1593 5607 1607
rect 5633 2033 5647 2047
rect 5673 2233 5687 2247
rect 5733 2253 5747 2267
rect 5693 2113 5707 2127
rect 5673 2093 5687 2107
rect 5713 2093 5727 2107
rect 5693 2073 5707 2087
rect 5673 2053 5687 2067
rect 5653 1853 5667 1867
rect 5653 1833 5667 1847
rect 5633 1753 5647 1767
rect 5593 1573 5607 1587
rect 5573 1553 5587 1567
rect 5533 1513 5547 1527
rect 5553 1333 5567 1347
rect 5593 1313 5607 1327
rect 5513 1293 5527 1307
rect 5613 1293 5627 1307
rect 5573 1273 5587 1287
rect 5573 1153 5587 1167
rect 5533 1113 5547 1127
rect 5513 1073 5527 1087
rect 5473 1013 5487 1027
rect 5553 1013 5567 1027
rect 5513 893 5527 907
rect 5553 833 5567 847
rect 5473 813 5487 827
rect 5493 813 5507 827
rect 5753 2113 5767 2127
rect 5893 4153 5907 4167
rect 5873 4033 5887 4047
rect 5873 3973 5887 3987
rect 5873 3673 5887 3687
rect 5853 3533 5867 3547
rect 5833 3473 5847 3487
rect 5833 3193 5847 3207
rect 5833 2913 5847 2927
rect 5833 2713 5847 2727
rect 5833 2253 5847 2267
rect 5813 2233 5827 2247
rect 5873 3493 5887 3507
rect 5873 2253 5887 2267
rect 5773 2093 5787 2107
rect 5813 2093 5827 2107
rect 5793 2073 5807 2087
rect 5733 2053 5747 2067
rect 5773 2053 5787 2067
rect 5773 2033 5787 2047
rect 5713 1873 5727 1887
rect 5713 1853 5727 1867
rect 5693 1793 5707 1807
rect 5673 1673 5687 1687
rect 5873 2233 5887 2247
rect 5853 2113 5867 2127
rect 5833 2033 5847 2047
rect 5813 1933 5827 1947
rect 5793 1873 5807 1887
rect 5773 1633 5787 1647
rect 5833 1753 5847 1767
rect 5793 1613 5807 1627
rect 5733 1573 5747 1587
rect 5733 1553 5747 1567
rect 5773 1553 5787 1567
rect 5713 1313 5727 1327
rect 5653 1293 5667 1307
rect 5633 1093 5647 1107
rect 5693 1093 5707 1107
rect 5613 993 5627 1007
rect 5573 713 5587 727
rect 5633 813 5647 827
rect 5753 1533 5767 1547
rect 5773 1313 5787 1327
rect 5773 1113 5787 1127
rect 5513 693 5527 707
rect 5613 693 5627 707
rect 5473 653 5487 667
rect 5693 713 5707 727
rect 5673 673 5687 687
rect 5453 613 5467 627
rect 5513 613 5527 627
rect 5413 413 5427 427
rect 5413 393 5427 407
rect 5413 373 5427 387
rect 5353 353 5367 367
rect 5393 353 5407 367
rect 5593 633 5607 647
rect 5613 613 5627 627
rect 5653 613 5667 627
rect 5573 593 5587 607
rect 5533 573 5547 587
rect 5533 393 5547 407
rect 5493 353 5507 367
rect 5553 333 5567 347
rect 5513 293 5527 307
rect 5453 273 5467 287
rect 5513 273 5527 287
rect 5313 213 5327 227
rect 5433 173 5447 187
rect 5473 153 5487 167
rect 5593 573 5607 587
rect 5593 313 5607 327
rect 5753 813 5767 827
rect 5713 653 5727 667
rect 5733 653 5747 667
rect 5713 613 5727 627
rect 5693 573 5707 587
rect 5673 353 5687 367
rect 5713 333 5727 347
rect 5693 313 5707 327
rect 5653 293 5667 307
rect 5653 193 5667 207
rect 5313 133 5327 147
rect 5453 133 5467 147
rect 5553 133 5567 147
rect 5613 153 5627 167
rect 5733 153 5747 167
rect 5813 1113 5827 1127
rect 5913 2093 5927 2107
rect 5913 2033 5927 2047
rect 5873 1753 5887 1767
rect 5873 1173 5887 1187
rect 5873 1113 5887 1127
rect 5873 833 5887 847
rect 5853 793 5867 807
rect 5813 613 5827 627
rect 5853 613 5867 627
rect 5773 593 5787 607
rect 5833 593 5847 607
rect 5793 573 5807 587
rect 5793 353 5807 367
rect 5833 353 5847 367
rect 5793 273 5807 287
rect 5793 213 5807 227
rect 5753 133 5767 147
rect 5213 113 5227 127
rect 5253 113 5267 127
rect 5293 113 5307 127
rect 5333 113 5347 127
rect 5493 113 5507 127
rect 5593 113 5607 127
rect 5813 173 5827 187
rect 5813 153 5827 167
rect 5853 153 5867 167
rect 5853 133 5867 147
rect 5813 113 5827 127
rect 5873 113 5887 127
rect 5793 93 5807 107
rect 5833 93 5847 107
rect 4953 73 4967 87
<< metal3 >>
rect 2327 6016 4473 6024
rect 4987 5956 5753 5964
rect 2096 5936 2173 5944
rect 227 5916 293 5924
rect 347 5916 473 5924
rect 527 5916 993 5924
rect 1176 5924 1184 5933
rect 1087 5916 1184 5924
rect 1676 5924 1684 5933
rect 2096 5927 2104 5936
rect 2187 5936 2273 5944
rect 2567 5936 2653 5944
rect 3687 5936 3833 5944
rect 3887 5936 3904 5944
rect 1587 5916 1684 5924
rect 1847 5916 1973 5924
rect 2707 5916 2833 5924
rect 2907 5916 3233 5924
rect 3327 5916 3373 5924
rect 3896 5924 3904 5936
rect 3927 5936 3993 5944
rect 4116 5936 4253 5944
rect 4116 5924 4124 5936
rect 5587 5936 5713 5944
rect 3896 5916 4124 5924
rect 4147 5916 4284 5924
rect 4276 5907 4284 5916
rect 4307 5916 4573 5924
rect 4627 5916 5213 5924
rect 5267 5916 5493 5924
rect 5947 5916 5984 5924
rect 87 5896 313 5904
rect 367 5896 693 5904
rect 847 5896 1324 5904
rect -24 5876 13 5884
rect 87 5876 113 5884
rect 207 5876 313 5884
rect 607 5876 673 5884
rect 1207 5876 1253 5884
rect 1316 5884 1324 5896
rect 1347 5896 1433 5904
rect 1487 5896 1653 5904
rect 1867 5896 2193 5904
rect 2467 5896 2673 5904
rect 2727 5896 3053 5904
rect 3227 5896 3353 5904
rect 3527 5896 3653 5904
rect 3787 5896 3833 5904
rect 4027 5896 4113 5904
rect 4327 5896 4793 5904
rect 4947 5896 5373 5904
rect 5667 5896 5733 5904
rect 1316 5876 1793 5884
rect 1907 5876 2273 5884
rect 2287 5876 2473 5884
rect 2967 5876 3033 5884
rect 3087 5876 3213 5884
rect 3707 5876 3913 5884
rect 4156 5884 4164 5893
rect 4156 5876 4433 5884
rect 4707 5876 4773 5884
rect 4787 5876 4913 5884
rect 4967 5876 5133 5884
rect 5147 5876 5193 5884
rect 5567 5876 5633 5884
rect 5687 5876 5773 5884
rect 5827 5876 5984 5884
rect 687 5856 1313 5864
rect 1527 5856 2033 5864
rect 3827 5856 4053 5864
rect 27 5836 813 5844
rect 727 5796 1333 5804
rect 1367 5796 1393 5804
rect 867 5776 1193 5784
rect 3487 5756 3773 5764
rect 4787 5756 4813 5764
rect 3427 5736 3593 5744
rect 3627 5716 4293 5724
rect 4307 5716 4493 5724
rect 1447 5696 1993 5704
rect 3047 5696 3833 5704
rect 3947 5696 5453 5704
rect 287 5676 413 5684
rect 627 5676 833 5684
rect 967 5676 1513 5684
rect 1607 5676 2393 5684
rect 2407 5676 3213 5684
rect 3227 5676 3553 5684
rect 3807 5676 4833 5684
rect 5487 5676 5553 5684
rect 247 5656 424 5664
rect 107 5636 204 5644
rect 196 5627 204 5636
rect 416 5644 424 5656
rect 567 5656 653 5664
rect 927 5656 1553 5664
rect 1567 5656 2353 5664
rect 2527 5656 2573 5664
rect 3187 5656 3513 5664
rect 3567 5656 3753 5664
rect 3787 5656 3953 5664
rect 4707 5656 4773 5664
rect 4827 5656 5033 5664
rect 5047 5656 5153 5664
rect 5267 5656 5313 5664
rect 5527 5656 5613 5664
rect 307 5636 404 5644
rect 416 5636 453 5644
rect 396 5627 404 5636
rect 796 5644 804 5653
rect 687 5636 804 5644
rect 827 5636 953 5644
rect 976 5636 1153 5644
rect 976 5624 984 5636
rect 1207 5636 1233 5644
rect 1347 5636 1593 5644
rect 1647 5636 1873 5644
rect 1887 5636 1933 5644
rect 2447 5636 2493 5644
rect 2567 5636 2853 5644
rect 3387 5636 3504 5644
rect 3496 5627 3504 5636
rect 3627 5636 3653 5644
rect 3707 5636 3813 5644
rect 3956 5636 4073 5644
rect 3956 5627 3964 5636
rect 4127 5636 4233 5644
rect 4447 5636 4533 5644
rect 4687 5636 4793 5644
rect 5187 5636 5273 5644
rect 5547 5636 5573 5644
rect 447 5616 984 5624
rect 1007 5616 1153 5624
rect 1187 5616 1313 5624
rect 1447 5616 1473 5624
rect 1587 5616 1713 5624
rect 1847 5616 1893 5624
rect 2267 5616 2333 5624
rect 2387 5616 2633 5624
rect 2767 5616 2813 5624
rect 2967 5616 3093 5624
rect 3587 5616 3593 5624
rect 3607 5616 3633 5624
rect 3687 5616 3933 5624
rect 4636 5624 4644 5633
rect 4387 5616 4644 5624
rect 4667 5616 4913 5624
rect 5067 5616 5213 5624
rect 5227 5616 5333 5624
rect 5507 5616 5673 5624
rect 687 5596 713 5604
rect 987 5596 1013 5604
rect 1027 5596 1353 5604
rect 1367 5596 1733 5604
rect 2047 5596 2133 5604
rect 2147 5596 2673 5604
rect 2687 5596 2893 5604
rect 2907 5596 3013 5604
rect 3267 5596 3273 5604
rect 3287 5596 3313 5604
rect 3367 5596 3533 5604
rect 3987 5596 4053 5604
rect 4067 5596 4173 5604
rect 4527 5596 4613 5604
rect 5307 5596 5433 5604
rect 5487 5596 5513 5604
rect 5627 5596 5713 5604
rect 127 5576 153 5584
rect 947 5576 973 5584
rect 1207 5576 1253 5584
rect 1267 5576 2293 5584
rect 3247 5576 3333 5584
rect 3627 5576 5273 5584
rect 5727 5576 5933 5584
rect 1407 5556 1553 5564
rect 1567 5556 1753 5564
rect 1767 5556 1913 5564
rect 1927 5556 5053 5564
rect 5447 5556 5793 5564
rect 2647 5536 4513 5544
rect 1967 5516 2793 5524
rect 4967 5516 5033 5524
rect 5047 5516 5233 5524
rect 5247 5516 5693 5524
rect 5707 5516 5753 5524
rect 1707 5496 2453 5504
rect 2867 5496 2973 5504
rect 3307 5496 3473 5504
rect 3487 5496 4193 5504
rect 4207 5496 4333 5504
rect 4347 5496 4473 5504
rect 4567 5496 5633 5504
rect 127 5476 593 5484
rect 607 5476 653 5484
rect 2387 5476 2533 5484
rect 2547 5476 4773 5484
rect 4796 5476 5324 5484
rect 267 5456 393 5464
rect 407 5456 433 5464
rect 567 5456 613 5464
rect 1087 5456 1273 5464
rect 1427 5456 1473 5464
rect 2427 5456 2553 5464
rect 2627 5456 2673 5464
rect 2727 5456 3613 5464
rect 4007 5456 4233 5464
rect 107 5436 193 5444
rect 207 5436 233 5444
rect 907 5436 933 5444
rect 1067 5436 1113 5444
rect 1807 5436 1993 5444
rect 2127 5436 2173 5444
rect 2347 5436 2413 5444
rect 2507 5436 2824 5444
rect 147 5416 213 5424
rect 347 5416 413 5424
rect 696 5424 704 5433
rect 2816 5427 2824 5436
rect 2847 5436 3153 5444
rect 3207 5436 3233 5444
rect 3447 5436 3553 5444
rect 3607 5436 3793 5444
rect 3807 5436 4113 5444
rect 4156 5427 4164 5456
rect 4487 5456 4533 5464
rect 4796 5464 4804 5476
rect 4607 5456 4804 5464
rect 5167 5456 5193 5464
rect 5247 5456 5293 5464
rect 5316 5464 5324 5476
rect 5407 5476 5413 5484
rect 5427 5476 5453 5484
rect 5316 5456 5673 5464
rect 4207 5436 4393 5444
rect 4747 5436 4993 5444
rect 5407 5436 5433 5444
rect 5647 5436 5833 5444
rect 587 5416 704 5424
rect 847 5416 953 5424
rect 1227 5416 1393 5424
rect 1527 5416 1813 5424
rect 1887 5416 1913 5424
rect 2107 5416 2273 5424
rect 2527 5416 2553 5424
rect 3087 5416 3413 5424
rect 3316 5407 3324 5416
rect 3727 5416 3824 5424
rect 187 5396 293 5404
rect 467 5396 853 5404
rect 867 5396 913 5404
rect 1047 5396 1293 5404
rect 1307 5396 1773 5404
rect 2107 5396 2133 5404
rect 2207 5396 2353 5404
rect 2447 5396 2493 5404
rect 2987 5396 3093 5404
rect 3247 5396 3273 5404
rect 3816 5404 3824 5416
rect 3847 5416 4104 5424
rect 3816 5396 3853 5404
rect 4096 5404 4104 5416
rect 4167 5416 4413 5424
rect 4436 5407 4444 5433
rect 4527 5416 4573 5424
rect 4627 5416 4653 5424
rect 4767 5416 4873 5424
rect 5227 5416 5253 5424
rect 5287 5416 5333 5424
rect 5347 5416 5553 5424
rect 4096 5396 4193 5404
rect 4207 5396 4273 5404
rect 4687 5396 4853 5404
rect 4907 5396 5113 5404
rect 5127 5396 5153 5404
rect 5187 5396 5313 5404
rect 5427 5396 5473 5404
rect 5507 5396 5533 5404
rect 87 5376 213 5384
rect 467 5376 513 5384
rect 1187 5376 1333 5384
rect 2327 5376 2473 5384
rect 2487 5376 2713 5384
rect 2947 5376 2973 5384
rect 2987 5376 3173 5384
rect 3567 5376 3973 5384
rect 4227 5376 4713 5384
rect 4787 5376 5193 5384
rect 5207 5376 5573 5384
rect 2267 5356 2313 5364
rect 2427 5356 2653 5364
rect 3227 5356 3733 5364
rect 3767 5356 4753 5364
rect 4847 5356 4893 5364
rect 4907 5356 5393 5364
rect 2007 5336 2613 5344
rect 1147 5316 1213 5324
rect 2707 5316 2773 5324
rect 2787 5316 4593 5324
rect 3087 5296 3573 5304
rect 3127 5276 3933 5284
rect 3547 5256 3633 5264
rect 3647 5256 3693 5264
rect 4307 5236 4533 5244
rect 687 5216 893 5224
rect 3027 5216 3653 5224
rect 4487 5216 4533 5224
rect 147 5196 173 5204
rect 187 5196 253 5204
rect 3167 5196 4333 5204
rect 4407 5196 4973 5204
rect 107 5176 193 5184
rect 647 5176 713 5184
rect 727 5176 753 5184
rect 1007 5176 1233 5184
rect 1247 5176 1613 5184
rect 1627 5176 1673 5184
rect 1687 5176 2333 5184
rect 2667 5176 2713 5184
rect 2727 5176 3013 5184
rect 3467 5176 3624 5184
rect 127 5156 153 5164
rect 387 5156 493 5164
rect 627 5156 773 5164
rect 1247 5156 1433 5164
rect 1607 5156 1633 5164
rect 1727 5156 1844 5164
rect 447 5136 473 5144
rect 787 5136 873 5144
rect 1176 5127 1184 5153
rect 1467 5136 1553 5144
rect 1836 5144 1844 5156
rect 1867 5156 1913 5164
rect 2627 5156 2693 5164
rect 2927 5156 3004 5164
rect 2996 5147 3004 5156
rect 3067 5156 3093 5164
rect 3207 5156 3273 5164
rect 3316 5156 3333 5164
rect 3316 5147 3324 5156
rect 3347 5156 3433 5164
rect 3616 5164 3624 5176
rect 3907 5176 3993 5184
rect 4127 5176 4173 5184
rect 4187 5176 4193 5184
rect 4327 5176 4493 5184
rect 5147 5176 5213 5184
rect 5307 5176 5353 5184
rect 5387 5176 5444 5184
rect 5436 5167 5444 5176
rect 3616 5156 3773 5164
rect 3787 5156 3873 5164
rect 4027 5156 4213 5164
rect 4587 5156 5153 5164
rect 5167 5156 5393 5164
rect 1836 5136 1873 5144
rect 1887 5136 1953 5144
rect 2007 5136 2053 5144
rect 2587 5136 2633 5144
rect 2867 5136 2933 5144
rect 3047 5136 3113 5144
rect 4367 5136 4393 5144
rect 4447 5136 4473 5144
rect 4536 5144 4544 5153
rect 4536 5136 4633 5144
rect 5047 5136 5144 5144
rect 5136 5127 5144 5136
rect 5267 5136 5304 5144
rect 267 5116 353 5124
rect 627 5116 733 5124
rect 907 5116 993 5124
rect 1007 5116 1113 5124
rect 1327 5116 1413 5124
rect 1847 5116 2013 5124
rect 2507 5116 2773 5124
rect 2967 5116 3133 5124
rect 4027 5116 4253 5124
rect 4527 5116 4913 5124
rect 5227 5116 5273 5124
rect 5296 5124 5304 5136
rect 5536 5144 5544 5153
rect 5427 5136 5544 5144
rect 5296 5116 5393 5124
rect 5487 5116 5513 5124
rect 5527 5116 5553 5124
rect 927 5096 1233 5104
rect 2767 5096 2873 5104
rect 2887 5096 3233 5104
rect 3847 5096 3853 5104
rect 3867 5096 4093 5104
rect 5067 5096 5373 5104
rect 5567 5096 5613 5104
rect 287 5076 393 5084
rect 467 5076 513 5084
rect 527 5076 673 5084
rect 1027 5076 1153 5084
rect 4967 5076 5293 5084
rect 5367 5076 5593 5084
rect 2407 5056 2413 5064
rect 2427 5056 4493 5064
rect 4507 5056 4673 5064
rect 5147 5056 5493 5064
rect 3567 5036 3713 5044
rect 5287 5036 5313 5044
rect 5327 5036 5633 5044
rect 4447 5016 5113 5024
rect 1487 4996 2793 5004
rect 2987 4996 3013 5004
rect 4587 4996 4933 5004
rect 447 4976 513 4984
rect 527 4976 553 4984
rect 567 4976 1073 4984
rect 1647 4976 1773 4984
rect 2607 4976 2653 4984
rect 2827 4976 2853 4984
rect 3407 4976 3693 4984
rect 4187 4976 4213 4984
rect 4347 4976 4853 4984
rect 5007 4976 5333 4984
rect 147 4956 253 4964
rect 747 4956 813 4964
rect 1007 4956 1113 4964
rect 1147 4956 1293 4964
rect 1307 4956 1333 4964
rect 1347 4956 1413 4964
rect 1856 4956 1873 4964
rect 167 4936 193 4944
rect 207 4936 213 4944
rect 367 4936 453 4944
rect 467 4936 493 4944
rect 1407 4936 1424 4944
rect 187 4916 233 4924
rect 287 4916 533 4924
rect 847 4916 973 4924
rect 1156 4924 1164 4933
rect 1416 4927 1424 4936
rect 1567 4936 1633 4944
rect 1747 4936 1773 4944
rect 1856 4944 1864 4956
rect 1887 4956 2113 4964
rect 2127 4956 2173 4964
rect 2287 4956 2393 4964
rect 2407 4956 2453 4964
rect 2467 4956 2573 4964
rect 2647 4956 2673 4964
rect 2687 4956 2733 4964
rect 2747 4956 2753 4964
rect 1807 4936 1864 4944
rect 1876 4936 1933 4944
rect 1156 4916 1253 4924
rect 1267 4916 1273 4924
rect 1447 4916 1533 4924
rect 1627 4916 1653 4924
rect 1876 4924 1884 4936
rect 2087 4936 2273 4944
rect 2756 4936 2833 4944
rect 1747 4916 1884 4924
rect 1907 4916 2053 4924
rect 2067 4916 2133 4924
rect 2227 4916 2333 4924
rect 2707 4916 2733 4924
rect 2756 4924 2764 4936
rect 2887 4936 2953 4944
rect 2967 4936 3213 4944
rect 2747 4916 2764 4924
rect 2787 4916 2813 4924
rect 2847 4916 3153 4924
rect 3256 4924 3264 4973
rect 3327 4956 3353 4964
rect 3607 4956 3633 4964
rect 3687 4956 3733 4964
rect 3747 4956 3953 4964
rect 4007 4956 4173 4964
rect 4647 4956 4673 4964
rect 4727 4956 4953 4964
rect 5047 4956 5173 4964
rect 5227 4956 5253 4964
rect 5427 4956 5533 4964
rect 5587 4956 5633 4964
rect 3427 4936 4293 4944
rect 4747 4936 5013 4944
rect 5027 4936 5633 4944
rect 5827 4936 5853 4944
rect 5867 4936 5913 4944
rect 3256 4916 3273 4924
rect 3827 4916 4273 4924
rect 4287 4916 4413 4924
rect 4467 4916 4873 4924
rect 4887 4916 4893 4924
rect 4947 4916 4973 4924
rect 5087 4916 5153 4924
rect 5167 4916 5353 4924
rect 107 4896 213 4904
rect 227 4896 293 4904
rect 547 4896 613 4904
rect 707 4896 913 4904
rect 1576 4904 1584 4913
rect 1576 4896 1693 4904
rect 2927 4896 3313 4904
rect 3647 4896 4133 4904
rect 4387 4896 4413 4904
rect 127 4876 193 4884
rect 1487 4876 1893 4884
rect 2667 4876 3373 4884
rect 3567 4876 4193 4884
rect 4607 4876 4893 4884
rect 4907 4876 5513 4884
rect 1247 4856 2253 4864
rect 2627 4856 2713 4864
rect 2727 4856 2993 4864
rect 3307 4856 4533 4864
rect 4547 4856 4693 4864
rect 4847 4856 5413 4864
rect 3107 4836 3513 4844
rect 3367 4816 4553 4824
rect 4567 4816 4633 4824
rect 2747 4796 3573 4804
rect 867 4776 1033 4784
rect 1047 4776 1813 4784
rect 1827 4776 4153 4784
rect 1087 4716 1173 4724
rect 1187 4716 2273 4724
rect 2307 4716 2433 4724
rect 3047 4716 3393 4724
rect 5667 4716 5813 4724
rect 447 4696 473 4704
rect 767 4696 804 4704
rect 107 4676 233 4684
rect 367 4676 593 4684
rect 796 4684 804 4696
rect 947 4696 1173 4704
rect 1287 4696 1453 4704
rect 1847 4696 1973 4704
rect 1987 4696 2073 4704
rect 2207 4696 2473 4704
rect 2487 4696 2644 4704
rect 2636 4687 2644 4696
rect 2667 4696 2773 4704
rect 2927 4696 2973 4704
rect 2987 4696 3553 4704
rect 3947 4696 4113 4704
rect 4227 4696 4293 4704
rect 4347 4696 4433 4704
rect 4487 4696 4533 4704
rect 4547 4696 4573 4704
rect 5007 4696 5373 4704
rect 5487 4696 5573 4704
rect 796 4676 873 4684
rect 887 4676 1093 4684
rect 1367 4676 1393 4684
rect 1507 4676 1593 4684
rect 1887 4676 1933 4684
rect 1947 4676 2313 4684
rect 2367 4676 2413 4684
rect 2467 4676 2493 4684
rect 2507 4676 2593 4684
rect 2767 4676 3093 4684
rect 3187 4676 3273 4684
rect 3587 4676 3633 4684
rect 3687 4676 3784 4684
rect 467 4656 493 4664
rect 627 4656 693 4664
rect 776 4664 784 4673
rect 747 4656 784 4664
rect 827 4656 913 4664
rect 1167 4656 1253 4664
rect 387 4636 533 4644
rect 727 4636 753 4644
rect 787 4636 893 4644
rect 1227 4636 1273 4644
rect 1316 4644 1324 4673
rect 3776 4667 3784 4676
rect 3987 4676 4313 4684
rect 4627 4676 4673 4684
rect 4987 4676 5093 4684
rect 5147 4676 5173 4684
rect 5387 4676 5513 4684
rect 1767 4656 1773 4664
rect 1787 4656 2133 4664
rect 2307 4656 2333 4664
rect 2627 4656 2833 4664
rect 2947 4656 3013 4664
rect 3127 4656 3153 4664
rect 3267 4656 3293 4664
rect 3967 4656 4093 4664
rect 4227 4656 4353 4664
rect 4387 4656 4553 4664
rect 4607 4656 4653 4664
rect 4687 4656 4713 4664
rect 5127 4656 5253 4664
rect 5447 4656 5493 4664
rect 5787 4656 5893 4664
rect 1316 4636 1353 4644
rect 1627 4636 1733 4644
rect 2127 4636 2353 4644
rect 2847 4636 2873 4644
rect 2907 4636 2953 4644
rect 3287 4636 3313 4644
rect 3447 4636 3473 4644
rect 3807 4636 3913 4644
rect 4567 4636 5533 4644
rect 5827 4636 5853 4644
rect 587 4616 993 4624
rect 1487 4616 1693 4624
rect 1727 4616 1833 4624
rect 2067 4616 2173 4624
rect 2327 4616 2713 4624
rect 2827 4616 2973 4624
rect 3667 4616 4073 4624
rect 4487 4616 4633 4624
rect 5427 4616 5453 4624
rect 5547 4616 5633 4624
rect 3067 4596 3133 4604
rect 3147 4596 3893 4604
rect 4147 4596 4753 4604
rect 4767 4596 5033 4604
rect 5047 4596 5293 4604
rect 5307 4596 5313 4604
rect 5327 4596 5653 4604
rect 1647 4576 1673 4584
rect 2667 4576 3613 4584
rect 3627 4576 3973 4584
rect 4947 4576 5153 4584
rect 5207 4576 5293 4584
rect 5727 4576 5753 4584
rect 1667 4556 1913 4564
rect 2587 4556 2693 4564
rect 3207 4556 3453 4564
rect 3467 4556 3793 4564
rect 4807 4556 4953 4564
rect 1367 4536 2013 4544
rect 2387 4536 2553 4544
rect 3767 4536 3953 4544
rect 4847 4536 5053 4544
rect 1047 4516 1573 4524
rect 2347 4516 2413 4524
rect 2427 4516 2913 4524
rect 3227 4516 3433 4524
rect 67 4496 353 4504
rect 467 4496 493 4504
rect 2267 4496 2573 4504
rect 2587 4496 2653 4504
rect 2747 4496 3113 4504
rect 3267 4496 3633 4504
rect 3847 4496 3993 4504
rect 4187 4496 4253 4504
rect 4467 4496 4553 4504
rect 4587 4496 4773 4504
rect 5027 4496 5073 4504
rect 76 4476 193 4484
rect 76 4444 84 4476
rect 287 4476 553 4484
rect 727 4476 853 4484
rect 1547 4476 1613 4484
rect 1747 4476 1793 4484
rect 2127 4476 2473 4484
rect 3027 4476 3073 4484
rect 3307 4476 3493 4484
rect 3827 4476 3853 4484
rect 4347 4476 4373 4484
rect 4627 4476 4913 4484
rect 4927 4476 4993 4484
rect 5147 4476 5213 4484
rect 5387 4476 5493 4484
rect 107 4456 213 4464
rect 256 4464 264 4473
rect 256 4456 324 4464
rect 76 4436 193 4444
rect 247 4436 293 4444
rect 316 4444 324 4456
rect 627 4456 744 4464
rect 736 4447 744 4456
rect 907 4456 1073 4464
rect 1147 4456 1264 4464
rect 1256 4447 1264 4456
rect 1407 4456 1484 4464
rect 316 4436 353 4444
rect 427 4436 473 4444
rect 487 4436 693 4444
rect 927 4436 1153 4444
rect 1347 4436 1373 4444
rect 1427 4436 1453 4444
rect 1476 4444 1484 4456
rect 1587 4456 1633 4464
rect 1827 4456 1973 4464
rect 2547 4456 2593 4464
rect 2607 4456 2953 4464
rect 3136 4464 3144 4473
rect 3007 4456 3144 4464
rect 3547 4456 3613 4464
rect 4027 4456 4113 4464
rect 4167 4456 4293 4464
rect 4367 4456 4393 4464
rect 4547 4456 4653 4464
rect 4987 4456 5073 4464
rect 5247 4456 5333 4464
rect 5627 4456 5733 4464
rect 1476 4436 1513 4444
rect 1867 4436 1993 4444
rect 3327 4436 3373 4444
rect 3667 4436 4253 4444
rect 4727 4436 5053 4444
rect 5107 4436 5153 4444
rect 5167 4436 5373 4444
rect 5387 4436 5633 4444
rect 5796 4444 5804 4473
rect 5767 4436 5804 4444
rect 207 4416 273 4424
rect 547 4416 693 4424
rect 876 4424 884 4433
rect 707 4416 884 4424
rect 1376 4424 1384 4433
rect 1376 4416 1393 4424
rect 1556 4424 1564 4433
rect 1547 4416 1564 4424
rect 2007 4416 2493 4424
rect 2507 4416 2513 4424
rect 2687 4416 2813 4424
rect 2827 4416 2933 4424
rect 3247 4416 3453 4424
rect 3767 4416 3913 4424
rect 3927 4416 4273 4424
rect 4747 4416 4933 4424
rect 5107 4416 5313 4424
rect 227 4396 293 4404
rect 787 4396 1113 4404
rect 1947 4396 2853 4404
rect 2867 4396 3453 4404
rect 4047 4396 4153 4404
rect 4787 4396 4893 4404
rect 4927 4396 5013 4404
rect 5167 4396 5273 4404
rect 3707 4376 4593 4384
rect 4867 4376 5193 4384
rect 127 4356 293 4364
rect 1307 4336 1373 4344
rect 5187 4336 5393 4344
rect 387 4316 593 4324
rect 607 4316 713 4324
rect 727 4316 1053 4324
rect 1067 4316 1293 4324
rect 1907 4316 2713 4324
rect 3227 4296 3273 4304
rect 5747 4296 5773 4304
rect 527 4276 733 4284
rect -24 4256 13 4264
rect 667 4256 873 4264
rect 3307 4256 3333 4264
rect -24 4236 2473 4244
rect -24 4216 -16 4236
rect 3987 4236 4393 4244
rect 4407 4236 5053 4244
rect 5367 4236 5413 4244
rect 5547 4236 5673 4244
rect 107 4216 133 4224
rect 147 4216 253 4224
rect 307 4216 393 4224
rect 507 4216 653 4224
rect 667 4216 833 4224
rect 847 4216 1013 4224
rect 1627 4216 1764 4224
rect 1756 4207 1764 4216
rect 1787 4216 1904 4224
rect 1896 4207 1904 4216
rect 2487 4216 2633 4224
rect 2647 4216 2653 4224
rect 2887 4216 2993 4224
rect 3107 4216 3153 4224
rect 3187 4216 3413 4224
rect 3507 4216 3773 4224
rect 4207 4216 4253 4224
rect 4447 4216 4473 4224
rect 4487 4216 4593 4224
rect 4616 4216 4673 4224
rect 147 4196 173 4204
rect 247 4196 253 4204
rect 267 4196 373 4204
rect 387 4196 493 4204
rect 547 4196 613 4204
rect 627 4196 633 4204
rect 687 4196 713 4204
rect 867 4196 933 4204
rect 947 4196 1024 4204
rect 207 4176 233 4184
rect 407 4176 473 4184
rect 1016 4184 1024 4196
rect 1047 4196 1153 4204
rect 1327 4196 1453 4204
rect 1507 4196 1733 4204
rect 2367 4196 2384 4204
rect 1016 4176 1173 4184
rect 1187 4176 1333 4184
rect 1427 4176 1493 4184
rect 1587 4176 1873 4184
rect 2376 4184 2384 4196
rect 2447 4196 2493 4204
rect 2707 4196 2753 4204
rect 2987 4196 3233 4204
rect 3387 4196 3473 4204
rect 3887 4196 3973 4204
rect 4027 4196 4113 4204
rect 4427 4196 4513 4204
rect 4616 4204 4624 4216
rect 4687 4216 4753 4224
rect 5107 4216 5273 4224
rect 5347 4216 5373 4224
rect 5427 4216 5513 4224
rect 5527 4216 5853 4224
rect 4567 4196 4624 4204
rect 5407 4196 5613 4204
rect 2376 4176 2393 4184
rect 2796 4184 2804 4193
rect 2796 4176 3173 4184
rect 3307 4176 3353 4184
rect 3427 4176 3613 4184
rect 3636 4184 3644 4193
rect 3636 4176 3713 4184
rect 4216 4184 4224 4193
rect 4007 4176 4224 4184
rect 4287 4176 4733 4184
rect 4827 4176 4953 4184
rect 4987 4176 5133 4184
rect 5236 4167 5244 4193
rect 5687 4176 5813 4184
rect 127 4156 293 4164
rect 387 4156 773 4164
rect 827 4156 1033 4164
rect 1207 4156 1633 4164
rect 1647 4156 1713 4164
rect 1867 4156 1953 4164
rect 1967 4156 2033 4164
rect 2047 4156 2053 4164
rect 2287 4156 2373 4164
rect 2567 4156 2613 4164
rect 2787 4156 2933 4164
rect 3167 4156 3333 4164
rect 3527 4156 3593 4164
rect 3747 4156 3833 4164
rect 4147 4156 4253 4164
rect 4347 4156 5213 4164
rect 5287 4156 5313 4164
rect 5667 4156 5733 4164
rect 5747 4156 5773 4164
rect 5827 4156 5893 4164
rect 447 4136 493 4144
rect 987 4136 1113 4144
rect 1407 4136 1473 4144
rect 2607 4136 2793 4144
rect 3027 4136 3233 4144
rect 3327 4136 3353 4144
rect 4247 4136 4413 4144
rect 4707 4136 4793 4144
rect 5187 4136 5253 4144
rect 5767 4136 5793 4144
rect 287 4116 313 4124
rect 327 4116 413 4124
rect 427 4116 533 4124
rect 1327 4116 1513 4124
rect 1527 4116 1593 4124
rect 2607 4116 2693 4124
rect 2707 4116 2853 4124
rect 4107 4116 5333 4124
rect 5347 4116 5473 4124
rect 5487 4116 5793 4124
rect 4967 4096 5473 4104
rect 5487 4096 5673 4104
rect 1067 4076 1433 4084
rect 1507 4076 2153 4084
rect 2807 4076 3053 4084
rect 3067 4076 3613 4084
rect 3627 4076 3753 4084
rect 4047 4076 4433 4084
rect 4607 4076 5293 4084
rect 5307 4076 5433 4084
rect 2027 4056 2193 4064
rect 3487 4056 3513 4064
rect 3527 4056 3793 4064
rect 4647 4056 4973 4064
rect 2867 4036 2993 4044
rect 3407 4036 3473 4044
rect 3487 4036 3633 4044
rect 3907 4036 4313 4044
rect 4667 4036 5013 4044
rect 5027 4036 5453 4044
rect 5716 4036 5873 4044
rect 207 4016 213 4024
rect 227 4016 553 4024
rect 1167 4016 1333 4024
rect 1347 4016 1633 4024
rect 1767 4016 1993 4024
rect 2447 4016 2493 4024
rect 2527 4016 2553 4024
rect 2907 4016 3153 4024
rect 3407 4016 3493 4024
rect 3667 4016 4053 4024
rect 4067 4016 4213 4024
rect 4267 4016 4353 4024
rect 4447 4016 4473 4024
rect 4736 4016 4833 4024
rect 4736 4007 4744 4016
rect 5607 4016 5693 4024
rect 5716 4007 5724 4036
rect 156 3996 413 4004
rect 156 3984 164 3996
rect 487 3996 533 4004
rect 547 3996 573 4004
rect 627 3996 713 4004
rect 1027 3996 1053 4004
rect 1227 3996 1293 4004
rect 1307 3996 1453 4004
rect 1496 3996 1533 4004
rect 87 3976 164 3984
rect 187 3976 233 3984
rect 327 3976 433 3984
rect 456 3984 464 3993
rect 456 3976 593 3984
rect 907 3976 913 3984
rect 927 3976 953 3984
rect 1007 3976 1033 3984
rect 1047 3976 1113 3984
rect 1367 3976 1433 3984
rect 1496 3984 1504 3996
rect 1547 3996 1553 4004
rect 1627 3996 1693 4004
rect 1747 3996 1853 4004
rect 2007 3996 2053 4004
rect 2287 3996 2433 4004
rect 2456 3996 2773 4004
rect 1447 3976 1504 3984
rect 1527 3976 1593 3984
rect 1907 3976 1993 3984
rect 2147 3976 2253 3984
rect 2307 3976 2353 3984
rect 2456 3984 2464 3996
rect 2987 3996 3033 4004
rect 3267 3996 3313 4004
rect 3587 3996 3653 4004
rect 3667 3996 3733 4004
rect 3927 3996 3944 4004
rect 2436 3976 2464 3984
rect 627 3956 653 3964
rect 1187 3956 1333 3964
rect 1347 3956 1393 3964
rect 1887 3956 1973 3964
rect 1987 3956 2033 3964
rect 2047 3956 2153 3964
rect 2436 3964 2444 3976
rect 2507 3976 2533 3984
rect 2727 3976 2833 3984
rect 3327 3976 3893 3984
rect 3936 3984 3944 3996
rect 3967 3996 4013 4004
rect 4547 3996 4613 4004
rect 5247 3996 5373 4004
rect 5507 3996 5673 4004
rect 3907 3976 3924 3984
rect 3936 3976 4093 3984
rect 2427 3956 2444 3964
rect 2476 3964 2484 3973
rect 2476 3956 2573 3964
rect 2607 3956 2633 3964
rect 2667 3956 2733 3964
rect 3127 3956 3133 3964
rect 3147 3956 3333 3964
rect 3916 3964 3924 3976
rect 4287 3976 4313 3984
rect 4387 3976 4493 3984
rect 4767 3976 4853 3984
rect 4936 3984 4944 3993
rect 4867 3976 4944 3984
rect 5067 3976 5153 3984
rect 5216 3984 5224 3993
rect 5216 3976 5233 3984
rect 5327 3976 5653 3984
rect 5676 3976 5693 3984
rect 3916 3956 4053 3964
rect 4287 3956 4353 3964
rect 5347 3956 5373 3964
rect 167 3936 233 3944
rect 307 3936 433 3944
rect 1687 3936 1973 3944
rect 2456 3944 2464 3953
rect 2456 3936 2473 3944
rect 2487 3936 2513 3944
rect 3907 3936 3933 3944
rect 3947 3936 4633 3944
rect 5676 3944 5684 3976
rect 5756 3964 5764 3973
rect 5707 3956 5764 3964
rect 5676 3936 5713 3944
rect 5776 3944 5784 4013
rect 5796 3987 5804 4013
rect 5816 3996 5833 4004
rect 5816 3967 5824 3996
rect 5847 3976 5873 3984
rect 5776 3936 5833 3944
rect 1727 3916 2213 3924
rect 2227 3916 3193 3924
rect 4187 3916 4533 3924
rect 4607 3916 4733 3924
rect 27 3896 1433 3904
rect 1447 3896 1933 3904
rect 4247 3896 4433 3904
rect 1747 3876 1793 3884
rect 2707 3876 2873 3884
rect 2887 3876 3213 3884
rect 4927 3876 4973 3884
rect 27 3856 693 3864
rect 707 3856 1233 3864
rect 3447 3856 4713 3864
rect 5227 3856 5433 3864
rect 1907 3836 2853 3844
rect 2867 3836 4333 3844
rect 4587 3836 4993 3844
rect 5007 3836 5293 3844
rect 1567 3816 2313 3824
rect 3607 3816 3833 3824
rect 5227 3816 5273 3824
rect 467 3796 2673 3804
rect 4887 3796 5293 3804
rect 887 3776 1113 3784
rect 1647 3776 1873 3784
rect 1887 3776 2613 3784
rect 927 3756 1013 3764
rect 1967 3756 2033 3764
rect 2187 3756 2253 3764
rect 2267 3756 2373 3764
rect 2707 3756 2773 3764
rect 2787 3756 3373 3764
rect 4867 3756 5273 3764
rect 5327 3756 5553 3764
rect 5567 3756 5773 3764
rect 5827 3756 5844 3764
rect 327 3736 353 3744
rect 407 3736 413 3744
rect 427 3736 513 3744
rect 887 3736 953 3744
rect 1087 3736 1153 3744
rect 1407 3736 1553 3744
rect 1847 3736 1933 3744
rect 2027 3736 2053 3744
rect 2216 3736 2293 3744
rect 2216 3727 2224 3736
rect 2527 3736 2553 3744
rect 2567 3736 2653 3744
rect 2847 3736 2893 3744
rect 3207 3736 3253 3744
rect 3267 3736 3473 3744
rect 3656 3736 3713 3744
rect 147 3716 253 3724
rect 287 3716 373 3724
rect 787 3716 933 3724
rect 1107 3716 1293 3724
rect 1427 3716 1513 3724
rect 1687 3716 1793 3724
rect 1827 3716 1873 3724
rect 1967 3716 2073 3724
rect 2276 3716 2353 3724
rect 487 3696 513 3704
rect 87 3676 413 3684
rect 536 3684 544 3713
rect 2276 3707 2284 3716
rect 2387 3716 2493 3724
rect 2507 3716 2753 3724
rect 3387 3716 3513 3724
rect 3656 3707 3664 3736
rect 4256 3736 4353 3744
rect 4256 3727 4264 3736
rect 4927 3736 5193 3744
rect 5207 3736 5553 3744
rect 5687 3736 5753 3744
rect 5767 3736 5813 3744
rect 3727 3716 3813 3724
rect 3827 3716 3973 3724
rect 4047 3716 4073 3724
rect 4156 3716 4253 3724
rect 607 3696 673 3704
rect 687 3696 793 3704
rect 1047 3696 1213 3704
rect 1227 3696 1573 3704
rect 2127 3696 2233 3704
rect 2307 3696 2533 3704
rect 2547 3696 2793 3704
rect 2807 3696 3013 3704
rect 3067 3696 3113 3704
rect 3247 3696 3353 3704
rect 3547 3696 3633 3704
rect 3676 3704 3684 3713
rect 3676 3696 3773 3704
rect 4156 3704 4164 3716
rect 4276 3716 4393 3724
rect 4107 3696 4164 3704
rect 4187 3696 4213 3704
rect 4276 3704 4284 3716
rect 4936 3716 5033 3724
rect 4936 3707 4944 3716
rect 5047 3716 5133 3724
rect 5287 3716 5373 3724
rect 5727 3716 5793 3724
rect 4227 3696 4284 3704
rect 4567 3696 4693 3704
rect 4727 3696 4893 3704
rect 5007 3696 5393 3704
rect 5836 3704 5844 3756
rect 5807 3696 5844 3704
rect 536 3676 653 3684
rect 767 3676 813 3684
rect 947 3676 1373 3684
rect 1587 3676 1653 3684
rect 1667 3676 1773 3684
rect 2387 3676 2553 3684
rect 2647 3676 2693 3684
rect 3407 3676 4013 3684
rect 4027 3676 4053 3684
rect 4947 3676 4973 3684
rect 5187 3676 5233 3684
rect 5427 3676 5533 3684
rect 5547 3676 5653 3684
rect 5827 3676 5873 3684
rect 507 3656 553 3664
rect 627 3656 653 3664
rect 847 3656 1193 3664
rect 1216 3656 1853 3664
rect 727 3636 1073 3644
rect 1216 3644 1224 3656
rect 1867 3656 1953 3664
rect 1967 3656 3053 3664
rect 3567 3656 3933 3664
rect 4007 3656 4233 3664
rect 4247 3656 4373 3664
rect 4787 3656 4893 3664
rect 5107 3656 5253 3664
rect 1087 3636 1224 3644
rect 1747 3636 1853 3644
rect 2727 3636 3553 3644
rect 3647 3636 3693 3644
rect 3707 3636 3793 3644
rect 4487 3636 4793 3644
rect 4807 3636 5193 3644
rect 1667 3616 3233 3624
rect 3707 3616 3913 3624
rect 4107 3616 4313 3624
rect 4407 3616 4593 3624
rect 107 3596 233 3604
rect 247 3596 313 3604
rect 2807 3596 2873 3604
rect 2927 3596 3053 3604
rect 3107 3596 3293 3604
rect 3307 3596 3773 3604
rect 3847 3596 4113 3604
rect 4447 3596 4693 3604
rect 4707 3596 5453 3604
rect 5467 3596 5593 3604
rect 5607 3596 5673 3604
rect 227 3576 253 3584
rect 587 3576 853 3584
rect 867 3576 953 3584
rect 1207 3576 1493 3584
rect 1507 3576 1553 3584
rect 3167 3576 3673 3584
rect 3687 3576 3793 3584
rect 3807 3576 3913 3584
rect 687 3556 1053 3564
rect 1067 3556 1593 3564
rect 1947 3556 1973 3564
rect 2527 3556 2573 3564
rect 2587 3556 2733 3564
rect 3647 3556 4033 3564
rect 4047 3556 4113 3564
rect 4127 3556 4133 3564
rect 4527 3556 4793 3564
rect 187 3536 313 3544
rect 627 3536 784 3544
rect 776 3527 784 3536
rect 1467 3536 1673 3544
rect 1687 3536 1753 3544
rect 1767 3536 2013 3544
rect 2116 3536 2193 3544
rect 107 3516 353 3524
rect 227 3496 253 3504
rect 387 3496 493 3504
rect 636 3504 644 3513
rect 627 3496 644 3504
rect 767 3496 793 3504
rect 876 3487 884 3533
rect 1167 3516 1213 3524
rect 1707 3516 1813 3524
rect 2116 3524 2124 3536
rect 2207 3536 2213 3544
rect 2227 3536 2273 3544
rect 2507 3536 2533 3544
rect 2587 3536 2653 3544
rect 2987 3536 3193 3544
rect 3427 3536 3513 3544
rect 3747 3536 3833 3544
rect 4776 3536 4853 3544
rect 4776 3527 4784 3536
rect 4867 3536 4953 3544
rect 5087 3536 5133 3544
rect 5367 3536 5433 3544
rect 5507 3536 5633 3544
rect 5787 3536 5853 3544
rect 1887 3516 2124 3524
rect 2407 3516 2433 3524
rect 2447 3516 2633 3524
rect 2787 3516 2913 3524
rect 3567 3516 3644 3524
rect 967 3496 1033 3504
rect 1287 3496 1393 3504
rect 1747 3496 1793 3504
rect 1847 3496 1993 3504
rect 2087 3496 2113 3504
rect 2347 3496 2373 3504
rect 2407 3496 2473 3504
rect 2487 3496 2513 3504
rect 2767 3496 2833 3504
rect 3156 3504 3164 3513
rect 2867 3496 3164 3504
rect 3447 3496 3473 3504
rect 3636 3504 3644 3516
rect 3667 3516 3733 3524
rect 4087 3516 4213 3524
rect 4096 3507 4104 3516
rect 4267 3516 4353 3524
rect 5047 3516 5073 3524
rect 5407 3516 5533 3524
rect 3636 3496 3713 3504
rect 3727 3496 3833 3504
rect 3847 3496 3953 3504
rect 4147 3496 4233 3504
rect 4427 3496 4513 3504
rect 5116 3504 5124 3513
rect 5107 3496 5124 3504
rect 5367 3496 5473 3504
rect 5527 3496 5693 3504
rect 5707 3496 5873 3504
rect 787 3476 813 3484
rect 1787 3476 2093 3484
rect 2287 3476 2353 3484
rect 2547 3476 2953 3484
rect 2967 3476 3033 3484
rect 3407 3476 3653 3484
rect 3827 3476 3933 3484
rect 4167 3476 4253 3484
rect 4467 3476 4493 3484
rect 4547 3476 4573 3484
rect 4887 3476 5013 3484
rect 5027 3476 5033 3484
rect 5807 3476 5833 3484
rect 767 3456 973 3464
rect 2147 3456 2293 3464
rect 2307 3456 2313 3464
rect 3507 3456 3573 3464
rect 3827 3456 3893 3464
rect 4547 3456 4973 3464
rect 4987 3456 5093 3464
rect 5327 3456 5353 3464
rect 367 3436 453 3444
rect 467 3436 473 3444
rect 1247 3436 1373 3444
rect 1387 3436 3213 3444
rect 4307 3436 4413 3444
rect 4647 3436 5333 3444
rect 1927 3416 2233 3424
rect 207 3396 1413 3404
rect 1427 3396 1893 3404
rect 3267 3396 3313 3404
rect 5347 3396 5373 3404
rect 5627 3396 5733 3404
rect 2167 3376 2233 3384
rect 3467 3376 4633 3384
rect 4767 3376 5213 3384
rect 5267 3376 5293 3384
rect 5307 3376 5493 3384
rect 2407 3356 2613 3364
rect 2787 3356 4053 3364
rect 1207 3336 1253 3344
rect 1267 3336 1353 3344
rect 1367 3336 1513 3344
rect 1527 3336 1693 3344
rect 2307 3336 2773 3344
rect 3927 3336 4173 3344
rect 347 3316 4473 3324
rect 4847 3316 5313 3324
rect 267 3296 953 3304
rect 967 3296 973 3304
rect 2707 3296 3453 3304
rect 3467 3296 3693 3304
rect 5027 3296 5213 3304
rect 5227 3296 5253 3304
rect 587 3276 693 3284
rect 1887 3276 1913 3284
rect 1927 3276 1933 3284
rect 2007 3276 2113 3284
rect 2127 3276 2133 3284
rect 2147 3276 2153 3284
rect 2547 3276 2653 3284
rect 2747 3276 2913 3284
rect 2927 3276 4813 3284
rect 4867 3276 5113 3284
rect 247 3256 493 3264
rect 576 3256 593 3264
rect -24 3236 224 3244
rect 216 3227 224 3236
rect 427 3236 453 3244
rect 576 3244 584 3256
rect 607 3256 813 3264
rect 827 3256 893 3264
rect 2047 3256 2093 3264
rect 2247 3256 2333 3264
rect 2356 3256 2373 3264
rect 2356 3247 2364 3256
rect 2507 3256 2593 3264
rect 2827 3256 3393 3264
rect 3567 3256 3613 3264
rect 3867 3256 4153 3264
rect 5087 3256 5133 3264
rect 5607 3256 5793 3264
rect 496 3236 584 3244
rect 496 3224 504 3236
rect 607 3236 613 3244
rect 627 3236 633 3244
rect 1007 3236 1093 3244
rect 1247 3236 1453 3244
rect 1507 3236 1733 3244
rect 1927 3236 2013 3244
rect 2527 3236 2693 3244
rect 2767 3236 2873 3244
rect 3187 3236 3273 3244
rect 3327 3236 3353 3244
rect 3436 3244 3444 3253
rect 3436 3236 3593 3244
rect 3767 3236 4033 3244
rect 4107 3236 4213 3244
rect 4407 3236 4473 3244
rect 4527 3236 4593 3244
rect 4607 3236 4684 3244
rect 4676 3227 4684 3236
rect 4707 3236 4853 3244
rect 5307 3236 5533 3244
rect 5547 3236 5613 3244
rect 5667 3236 5733 3244
rect 487 3216 504 3224
rect 527 3216 673 3224
rect 687 3216 733 3224
rect 847 3216 873 3224
rect 1807 3216 1853 3224
rect 1867 3216 1973 3224
rect 2567 3216 2613 3224
rect 2687 3216 2753 3224
rect 2867 3216 2893 3224
rect 2947 3216 2993 3224
rect 3087 3216 3113 3224
rect 3267 3216 3293 3224
rect 3447 3216 3493 3224
rect 3587 3216 3633 3224
rect 3667 3216 3713 3224
rect 3747 3216 3813 3224
rect 4027 3216 4153 3224
rect 4287 3216 4453 3224
rect 4747 3216 4993 3224
rect 5167 3216 5273 3224
rect 5587 3216 5773 3224
rect 447 3196 673 3204
rect 727 3196 793 3204
rect 1107 3196 1273 3204
rect 1767 3196 1813 3204
rect 1987 3196 2293 3204
rect 2427 3196 2673 3204
rect 2727 3196 2893 3204
rect 3047 3196 3093 3204
rect 3167 3196 3293 3204
rect 3347 3196 3433 3204
rect 3447 3196 3473 3204
rect 3867 3196 3893 3204
rect 3907 3196 4073 3204
rect 4247 3196 4433 3204
rect 4667 3196 4713 3204
rect 5047 3196 5124 3204
rect 627 3176 773 3184
rect 787 3176 813 3184
rect 1027 3176 1033 3184
rect 1047 3176 1153 3184
rect 1167 3176 1233 3184
rect 1327 3176 1433 3184
rect 2487 3176 2973 3184
rect 3107 3176 3513 3184
rect 4007 3176 4393 3184
rect 4447 3176 4553 3184
rect 5116 3184 5124 3196
rect 5147 3196 5413 3204
rect 5507 3196 5653 3204
rect 5787 3196 5833 3204
rect 5116 3176 5233 3184
rect 5567 3176 5693 3184
rect 127 3156 233 3164
rect 307 3156 393 3164
rect 627 3156 753 3164
rect 3407 3156 3493 3164
rect 3887 3156 4373 3164
rect 5147 3156 5353 3164
rect 87 3136 213 3144
rect 307 3136 853 3144
rect 2387 3136 2433 3144
rect 2807 3136 3353 3144
rect 147 3116 253 3124
rect 267 3116 313 3124
rect 2407 3116 2433 3124
rect 3287 3116 3653 3124
rect 3987 3116 4493 3124
rect 4507 3116 4973 3124
rect 5227 3116 5373 3124
rect 5387 3116 5453 3124
rect 5587 3116 5613 3124
rect 567 3096 693 3104
rect 1067 3096 1833 3104
rect 3227 3096 3973 3104
rect 4107 3096 4673 3104
rect 4827 3096 5553 3104
rect 67 3076 93 3084
rect 227 3076 413 3084
rect 1127 3076 1353 3084
rect 1767 3076 2093 3084
rect 2267 3076 2333 3084
rect 3247 3076 3344 3084
rect 107 3056 153 3064
rect 327 3056 513 3064
rect 527 3056 1093 3064
rect 1307 3056 1313 3064
rect 1327 3056 1393 3064
rect 1607 3056 1893 3064
rect 2067 3056 2133 3064
rect 2147 3056 2793 3064
rect 2887 3056 2933 3064
rect 3027 3056 3113 3064
rect 3336 3064 3344 3076
rect 3367 3076 3793 3084
rect 3807 3076 4133 3084
rect 4147 3076 4493 3084
rect 4847 3076 5173 3084
rect 5187 3076 5353 3084
rect 3336 3056 3533 3064
rect 3547 3056 3773 3064
rect 3967 3056 4553 3064
rect 4807 3056 4993 3064
rect 5007 3056 5073 3064
rect 76 3036 273 3044
rect 76 3027 84 3036
rect 567 3036 753 3044
rect 1087 3036 1113 3044
rect 1127 3036 1133 3044
rect 1207 3036 1253 3044
rect 1907 3036 1953 3044
rect 2107 3036 2133 3044
rect 2207 3036 2233 3044
rect 2247 3036 2304 3044
rect 127 3016 153 3024
rect 167 3016 373 3024
rect 387 3016 473 3024
rect 787 3016 873 3024
rect 1387 3016 1413 3024
rect 1467 3016 1553 3024
rect 1967 3016 2013 3024
rect 2127 3016 2213 3024
rect 2296 3024 2304 3036
rect 2327 3036 2513 3044
rect 2887 3036 3124 3044
rect 2296 3016 2393 3024
rect 2507 3016 2593 3024
rect 2607 3016 2673 3024
rect 2727 3016 2833 3024
rect 2987 3016 3093 3024
rect 3116 3024 3124 3036
rect 3167 3036 3193 3044
rect 3347 3036 3413 3044
rect 3447 3036 3633 3044
rect 3707 3036 4013 3044
rect 4047 3036 4313 3044
rect 4387 3036 4404 3044
rect 3116 3016 3133 3024
rect 3547 3016 3613 3024
rect 3687 3016 3793 3024
rect 3827 3016 3993 3024
rect 4047 3016 4073 3024
rect 4087 3016 4353 3024
rect 4396 3024 4404 3036
rect 4427 3036 4613 3044
rect 4627 3036 4853 3044
rect 4887 3036 4933 3044
rect 4987 3036 5033 3044
rect 5267 3036 5333 3044
rect 5347 3036 5413 3044
rect 5716 3036 5793 3044
rect 4376 3016 4513 3024
rect 447 2996 573 3004
rect 587 2996 633 3004
rect 747 2996 893 3004
rect 907 2996 933 3004
rect 1167 2996 1193 3004
rect 1427 2996 1573 3004
rect 1587 2996 1633 3004
rect 1947 2996 1993 3004
rect 2007 2996 2253 3004
rect 2647 2996 2693 3004
rect 2767 2996 2993 3004
rect 3007 2996 3193 3004
rect 547 2976 853 2984
rect 867 2976 1533 2984
rect 1547 2976 1973 2984
rect 3256 2984 3264 3013
rect 3427 2996 3573 3004
rect 3607 2996 3693 3004
rect 4376 3004 4384 3016
rect 4687 3016 4833 3024
rect 5527 3016 5673 3024
rect 5716 3024 5724 3036
rect 5687 3016 5724 3024
rect 4287 2996 4384 3004
rect 4436 2996 4653 3004
rect 3087 2976 3264 2984
rect 3387 2976 3433 2984
rect 3847 2976 4133 2984
rect 4436 2984 4444 2996
rect 4707 2996 4773 3004
rect 4867 2996 4893 3004
rect 4327 2976 4444 2984
rect 547 2956 613 2964
rect 867 2956 913 2964
rect 1887 2956 2153 2964
rect 2307 2956 2353 2964
rect 2367 2956 2753 2964
rect 3067 2956 3373 2964
rect 3847 2956 3933 2964
rect 4067 2956 4673 2964
rect 2367 2936 2453 2944
rect 3987 2936 4013 2944
rect 4027 2936 4393 2944
rect 4587 2936 5073 2944
rect 2967 2916 3033 2924
rect 5787 2916 5833 2924
rect 1867 2896 3273 2904
rect 2047 2856 3413 2864
rect 3867 2856 4893 2864
rect 5627 2856 5733 2864
rect 3467 2836 3993 2844
rect 4007 2836 4173 2844
rect 4207 2836 4633 2844
rect 1167 2816 1213 2824
rect 1707 2816 2033 2824
rect 2447 2816 2953 2824
rect 3087 2816 3933 2824
rect 3947 2816 4113 2824
rect 4147 2816 4233 2824
rect 4247 2816 4553 2824
rect 1827 2796 1864 2804
rect 1347 2776 1373 2784
rect 1467 2776 1553 2784
rect 1767 2776 1793 2784
rect 1816 2776 1833 2784
rect 67 2756 113 2764
rect 127 2756 353 2764
rect 527 2756 613 2764
rect 787 2756 873 2764
rect 1147 2756 1233 2764
rect 1407 2756 1653 2764
rect 1676 2747 1684 2773
rect 1816 2764 1824 2776
rect 1807 2756 1824 2764
rect 1856 2764 1864 2796
rect 1976 2796 2073 2804
rect 1956 2767 1964 2793
rect 1976 2787 1984 2796
rect 2407 2796 2493 2804
rect 2516 2796 2573 2804
rect 2067 2776 2133 2784
rect 2187 2776 2253 2784
rect 2516 2784 2524 2796
rect 2596 2796 2733 2804
rect 2276 2776 2524 2784
rect 1856 2756 1913 2764
rect 2027 2756 2093 2764
rect 2276 2764 2284 2776
rect 2596 2784 2604 2796
rect 3247 2796 3513 2804
rect 3527 2796 3633 2804
rect 3647 2796 3653 2804
rect 4107 2796 4213 2804
rect 4227 2796 4793 2804
rect 2547 2776 2604 2784
rect 2667 2776 2733 2784
rect 2747 2776 2773 2784
rect 2987 2776 3213 2784
rect 3527 2776 3764 2784
rect 2116 2756 2284 2764
rect 107 2736 233 2744
rect 367 2736 413 2744
rect 427 2736 593 2744
rect 687 2736 753 2744
rect 1267 2736 1493 2744
rect 1727 2736 1773 2744
rect 1887 2736 1933 2744
rect 2116 2744 2124 2756
rect 2307 2756 2413 2764
rect 2567 2756 2793 2764
rect 2976 2756 3133 2764
rect 2087 2736 2124 2744
rect 2347 2736 2513 2744
rect 2916 2744 2924 2753
rect 2747 2736 2924 2744
rect 2976 2727 2984 2756
rect 3427 2756 3513 2764
rect 3627 2756 3733 2764
rect 3756 2764 3764 2776
rect 3787 2776 3873 2784
rect 3887 2776 3913 2784
rect 3996 2776 4213 2784
rect 3996 2764 4004 2776
rect 4507 2776 4593 2784
rect 5427 2776 5733 2784
rect 3756 2756 4004 2764
rect 4027 2756 4053 2764
rect 4207 2756 4253 2764
rect 4327 2756 4353 2764
rect 4436 2764 4444 2773
rect 4436 2756 4573 2764
rect 4707 2756 4833 2764
rect 3027 2736 3093 2744
rect 3127 2736 3193 2744
rect 3207 2736 3253 2744
rect 3487 2736 3713 2744
rect 3847 2736 3913 2744
rect 4416 2744 4424 2753
rect 4127 2736 4424 2744
rect 4447 2736 4493 2744
rect 4827 2736 5013 2744
rect 5167 2736 5233 2744
rect 5247 2736 5273 2744
rect 5327 2736 5553 2744
rect 5687 2736 5793 2744
rect 167 2716 273 2724
rect 287 2716 313 2724
rect 567 2716 693 2724
rect 1007 2716 1213 2724
rect 1227 2716 1293 2724
rect 1447 2716 1713 2724
rect 1767 2716 1853 2724
rect 2007 2716 2233 2724
rect 2527 2716 2613 2724
rect 3447 2716 3893 2724
rect 4567 2716 4733 2724
rect 4747 2716 4773 2724
rect 4787 2716 5313 2724
rect 5787 2716 5833 2724
rect 387 2696 453 2704
rect 467 2696 573 2704
rect 587 2696 973 2704
rect 1807 2696 2013 2704
rect 2287 2696 2673 2704
rect 2727 2696 2993 2704
rect 3407 2696 3493 2704
rect 4107 2696 4753 2704
rect 587 2676 653 2684
rect 907 2676 1013 2684
rect 1027 2676 1333 2684
rect 1547 2676 1813 2684
rect 2847 2676 3153 2684
rect 3167 2676 4073 2684
rect 4407 2676 4613 2684
rect 4627 2676 4693 2684
rect 3547 2656 3553 2664
rect 3567 2656 4133 2664
rect 4147 2656 4293 2664
rect 3007 2636 3753 2644
rect 4047 2636 4073 2644
rect 4087 2636 4453 2644
rect 4987 2636 5033 2644
rect 5067 2636 5073 2644
rect 5087 2636 5413 2644
rect 487 2616 733 2624
rect 807 2616 833 2624
rect 847 2616 1173 2624
rect 1187 2616 1433 2624
rect 3407 2616 3573 2624
rect 3587 2616 3753 2624
rect 3767 2616 3793 2624
rect 3807 2616 3933 2624
rect 3947 2616 3953 2624
rect 3967 2616 4113 2624
rect 4127 2616 4153 2624
rect 507 2596 713 2604
rect 1847 2596 3253 2604
rect 3287 2596 3353 2604
rect 3727 2596 3833 2604
rect 3847 2596 4173 2604
rect 4447 2596 4553 2604
rect 5207 2596 5393 2604
rect 247 2576 433 2584
rect 527 2576 693 2584
rect 927 2576 1093 2584
rect 1707 2576 2133 2584
rect 2727 2576 2793 2584
rect 2827 2576 2853 2584
rect 3087 2576 3233 2584
rect 3347 2576 3513 2584
rect 3867 2576 3893 2584
rect 4527 2576 4713 2584
rect 4847 2576 4873 2584
rect 4927 2576 4933 2584
rect 4947 2576 4993 2584
rect 5047 2576 5253 2584
rect 5267 2576 5593 2584
rect 5607 2576 5753 2584
rect 496 2556 593 2564
rect 496 2547 504 2556
rect 667 2556 973 2564
rect 1287 2556 1473 2564
rect 1507 2556 1533 2564
rect 1767 2556 1813 2564
rect 1887 2556 1913 2564
rect 2267 2556 2393 2564
rect 2467 2556 3013 2564
rect 3307 2556 3353 2564
rect 3987 2556 4113 2564
rect 4276 2564 4284 2573
rect 4187 2556 4593 2564
rect 4687 2556 5033 2564
rect 5087 2556 5193 2564
rect 5507 2556 5793 2564
rect 347 2536 453 2544
rect 747 2536 1253 2544
rect 1307 2536 1393 2544
rect 2007 2536 2153 2544
rect 2267 2536 2293 2544
rect 2307 2536 2373 2544
rect 2396 2536 2533 2544
rect 227 2516 313 2524
rect 327 2516 473 2524
rect 487 2516 553 2524
rect 687 2516 693 2524
rect 707 2516 893 2524
rect 907 2516 993 2524
rect 1367 2516 1413 2524
rect 1427 2516 1713 2524
rect 1727 2516 1753 2524
rect 1787 2516 1853 2524
rect 1927 2516 2013 2524
rect 2067 2516 2113 2524
rect 2247 2516 2273 2524
rect 2396 2524 2404 2536
rect 2547 2536 2733 2544
rect 2747 2536 2833 2544
rect 2947 2536 3853 2544
rect 3887 2536 4253 2544
rect 4407 2536 4493 2544
rect 5147 2536 5513 2544
rect 5567 2536 5613 2544
rect 2287 2516 2404 2524
rect 2487 2516 3093 2524
rect 3947 2516 3993 2524
rect 4047 2516 4173 2524
rect 4267 2516 4533 2524
rect 4887 2516 5453 2524
rect 327 2496 933 2504
rect 947 2496 4513 2504
rect 107 2476 753 2484
rect 1007 2476 1113 2484
rect 1127 2476 1353 2484
rect 1367 2476 1453 2484
rect 1467 2476 1673 2484
rect 2167 2476 2193 2484
rect 2647 2476 3673 2484
rect 207 2456 253 2464
rect 967 2456 1413 2464
rect 2247 2456 2813 2464
rect 2827 2456 3033 2464
rect 2087 2436 2413 2444
rect 2427 2436 2573 2444
rect 2767 2436 2873 2444
rect 2967 2436 3173 2444
rect 1227 2416 1373 2424
rect 1387 2416 1433 2424
rect 1447 2416 1513 2424
rect 1527 2416 1793 2424
rect 1807 2416 1973 2424
rect 2047 2396 2393 2404
rect 3067 2396 3133 2404
rect 1587 2376 2993 2384
rect 3227 2376 3293 2384
rect 5447 2376 5473 2384
rect 127 2356 173 2364
rect 2367 2356 2633 2364
rect 707 2336 1133 2344
rect 1507 2336 2833 2344
rect 3316 2336 3493 2344
rect 387 2316 453 2324
rect 627 2316 893 2324
rect 927 2316 1533 2324
rect 1747 2316 2313 2324
rect 2327 2316 2333 2324
rect 2587 2316 3153 2324
rect 3316 2324 3324 2336
rect 3507 2336 3713 2344
rect 3967 2336 4893 2344
rect 5187 2336 5533 2344
rect 3167 2316 3324 2324
rect 3347 2316 3413 2324
rect 3887 2316 4233 2324
rect 4647 2316 5033 2324
rect 5107 2316 5324 2324
rect 287 2296 493 2304
rect 747 2296 1033 2304
rect 1147 2296 1173 2304
rect 1687 2296 1733 2304
rect 2387 2296 2453 2304
rect 2467 2296 2493 2304
rect 2907 2296 2924 2304
rect 147 2276 233 2284
rect 247 2276 333 2284
rect 347 2276 373 2284
rect 767 2276 793 2284
rect 847 2276 913 2284
rect 1056 2276 1093 2284
rect 547 2256 593 2264
rect 636 2244 644 2273
rect 667 2256 733 2264
rect 827 2256 853 2264
rect 567 2236 953 2244
rect 1056 2244 1064 2276
rect 1247 2276 1433 2284
rect 1547 2276 1753 2284
rect 2047 2276 2193 2284
rect 2207 2276 2353 2284
rect 2367 2276 2413 2284
rect 2547 2276 2673 2284
rect 1087 2256 1313 2264
rect 1936 2264 1944 2273
rect 1527 2256 2024 2264
rect 1056 2236 1993 2244
rect 2016 2244 2024 2256
rect 2107 2256 2253 2264
rect 2267 2256 2273 2264
rect 2327 2256 2513 2264
rect 2016 2236 2173 2244
rect 407 2216 773 2224
rect 1027 2216 1153 2224
rect 1207 2216 1453 2224
rect 1807 2216 1853 2224
rect 1867 2216 2533 2224
rect 2716 2224 2724 2273
rect 2916 2267 2924 2296
rect 3047 2296 3293 2304
rect 3307 2296 4173 2304
rect 4187 2296 4273 2304
rect 4367 2296 4533 2304
rect 4827 2296 4913 2304
rect 5007 2296 5053 2304
rect 5136 2296 5193 2304
rect 3067 2276 3273 2284
rect 3707 2276 3733 2284
rect 3847 2276 3913 2284
rect 3927 2276 3953 2284
rect 4427 2276 4553 2284
rect 4867 2276 4933 2284
rect 5136 2284 5144 2296
rect 5316 2304 5324 2316
rect 5347 2316 5493 2324
rect 5316 2296 5453 2304
rect 5467 2296 5573 2304
rect 5727 2296 5773 2304
rect 4987 2276 5144 2284
rect 5167 2276 5213 2284
rect 5627 2276 5653 2284
rect 5687 2276 5713 2284
rect 2987 2256 3073 2264
rect 3127 2256 3193 2264
rect 3207 2256 3433 2264
rect 3536 2264 3544 2273
rect 3447 2256 3544 2264
rect 3647 2256 3853 2264
rect 3867 2256 3973 2264
rect 4247 2256 4333 2264
rect 4447 2256 4873 2264
rect 5087 2256 5173 2264
rect 5207 2256 5333 2264
rect 5407 2256 5633 2264
rect 5647 2256 5653 2264
rect 5747 2256 5833 2264
rect 5976 2264 5984 2284
rect 5887 2256 5984 2264
rect 2787 2236 4033 2244
rect 4067 2236 4753 2244
rect 5107 2236 5133 2244
rect 5587 2236 5673 2244
rect 5827 2236 5873 2244
rect 2716 2216 2773 2224
rect 3047 2216 3153 2224
rect 3167 2216 4424 2224
rect 367 2196 573 2204
rect 1327 2196 2133 2204
rect 2147 2196 2793 2204
rect 2807 2196 2973 2204
rect 3247 2196 3313 2204
rect 4327 2196 4393 2204
rect 4416 2204 4424 2216
rect 4527 2216 4773 2224
rect 4416 2196 4633 2204
rect 4967 2196 5453 2204
rect 447 2176 993 2184
rect 2007 2176 3453 2184
rect 3907 2176 5173 2184
rect 5187 2176 5233 2184
rect 5267 2176 5333 2184
rect 5347 2176 5373 2184
rect 1727 2156 2013 2164
rect 2507 2156 2553 2164
rect 3447 2156 4073 2164
rect 4207 2156 4513 2164
rect 4527 2156 4573 2164
rect 4587 2156 4973 2164
rect 5147 2156 5373 2164
rect 1187 2136 1313 2144
rect 1647 2136 1773 2144
rect 1927 2136 2053 2144
rect 2707 2136 2953 2144
rect 3367 2136 4293 2144
rect 4307 2136 4433 2144
rect 5167 2136 5233 2144
rect 247 2116 293 2124
rect 307 2116 433 2124
rect 727 2116 833 2124
rect 1007 2116 2233 2124
rect 2267 2116 2873 2124
rect 2947 2116 3273 2124
rect 3287 2116 3393 2124
rect 3627 2116 4173 2124
rect 4347 2116 4633 2124
rect 4767 2116 5013 2124
rect 5027 2116 5693 2124
rect 5767 2116 5853 2124
rect 267 2096 313 2104
rect 327 2096 393 2104
rect 467 2096 493 2104
rect 607 2096 664 2104
rect 387 2076 573 2084
rect 656 2084 664 2096
rect 687 2096 713 2104
rect 907 2096 1113 2104
rect 1767 2096 1973 2104
rect 2167 2096 2273 2104
rect 3347 2096 3413 2104
rect 4027 2096 4093 2104
rect 4507 2096 4573 2104
rect 4647 2096 4713 2104
rect 4887 2096 4893 2104
rect 4907 2096 4953 2104
rect 5287 2096 5353 2104
rect 5607 2096 5673 2104
rect 5727 2096 5773 2104
rect 5827 2096 5913 2104
rect 656 2076 744 2084
rect 127 2056 224 2064
rect 216 2047 224 2056
rect 467 2056 513 2064
rect 616 2064 624 2073
rect 736 2067 744 2076
rect 887 2076 1133 2084
rect 1207 2076 1253 2084
rect 1427 2076 1513 2084
rect 1527 2076 1653 2084
rect 1827 2076 2173 2084
rect 616 2056 693 2064
rect 927 2056 973 2064
rect 1027 2056 1413 2064
rect 1507 2056 1553 2064
rect 1816 2064 1824 2073
rect 1956 2067 1964 2076
rect 2187 2076 2193 2084
rect 2567 2076 2593 2084
rect 2647 2076 2853 2084
rect 3027 2076 3133 2084
rect 3147 2076 3453 2084
rect 3527 2076 3553 2084
rect 3776 2067 3784 2093
rect 3807 2076 3913 2084
rect 3987 2076 4133 2084
rect 4407 2076 4453 2084
rect 4627 2076 4693 2084
rect 5087 2076 5113 2084
rect 5167 2076 5193 2084
rect 5487 2076 5593 2084
rect 5707 2076 5793 2084
rect 1647 2056 1824 2064
rect 2307 2056 2653 2064
rect 2827 2056 3153 2064
rect 3207 2056 3293 2064
rect 3507 2056 3593 2064
rect 3827 2056 3893 2064
rect 4067 2056 4193 2064
rect 4327 2056 4413 2064
rect 4527 2056 4553 2064
rect 4607 2056 4633 2064
rect 4747 2056 4793 2064
rect 5047 2056 5253 2064
rect 5307 2056 5393 2064
rect 5467 2056 5473 2064
rect 5487 2056 5513 2064
rect 5687 2056 5733 2064
rect 5756 2056 5773 2064
rect 687 2036 853 2044
rect 1307 2036 1393 2044
rect 1727 2036 1833 2044
rect 1876 2044 1884 2053
rect 1867 2036 1884 2044
rect 2447 2036 2533 2044
rect 2607 2036 2633 2044
rect 2907 2036 3133 2044
rect 3147 2036 3273 2044
rect 3287 2036 3373 2044
rect 3467 2036 3533 2044
rect 3547 2036 3713 2044
rect 4147 2036 4153 2044
rect 4167 2036 4313 2044
rect 4507 2036 4853 2044
rect 5756 2044 5764 2056
rect 5647 2036 5764 2044
rect 5787 2036 5833 2044
rect 5927 2036 5984 2044
rect 107 2016 373 2024
rect 907 2016 1253 2024
rect 1567 2016 1593 2024
rect 2287 2016 2393 2024
rect 2647 2016 2693 2024
rect 3187 2016 3593 2024
rect 3607 2016 3753 2024
rect 3927 2016 4273 2024
rect 4287 2016 4393 2024
rect 947 1996 993 2004
rect 1587 1996 1633 2004
rect 1647 1996 1673 2004
rect 2687 1996 3193 2004
rect 3227 1996 3273 2004
rect 3767 1996 3973 2004
rect 3987 1996 4073 2004
rect 87 1976 293 1984
rect 1587 1976 1613 1984
rect 5347 1976 5513 1984
rect 1387 1956 2173 1964
rect 2187 1956 2453 1964
rect 2467 1956 3573 1964
rect 1187 1936 1713 1944
rect 2067 1936 2573 1944
rect 2587 1936 2673 1944
rect 3147 1936 5813 1944
rect 3327 1916 3513 1924
rect 3527 1916 3573 1924
rect 4027 1896 4053 1904
rect 2547 1876 2733 1884
rect 3947 1876 4353 1884
rect 4367 1876 4473 1884
rect 5727 1876 5793 1884
rect 467 1856 553 1864
rect 2127 1856 3373 1864
rect 4447 1856 5653 1864
rect 5667 1856 5713 1864
rect 487 1836 613 1844
rect 907 1836 933 1844
rect 1167 1836 1633 1844
rect 1787 1836 2033 1844
rect 2087 1836 2113 1844
rect 2487 1836 2933 1844
rect 3527 1836 4873 1844
rect 5587 1836 5653 1844
rect 507 1816 533 1824
rect 707 1816 793 1824
rect 807 1816 853 1824
rect 867 1816 993 1824
rect 1007 1816 1293 1824
rect 1327 1816 1473 1824
rect 1867 1816 1904 1824
rect 487 1796 573 1804
rect 827 1796 893 1804
rect 907 1796 1033 1804
rect 1507 1796 1593 1804
rect 1896 1804 1904 1816
rect 2127 1816 2213 1824
rect 2627 1816 2653 1824
rect 2707 1816 2773 1824
rect 3267 1816 3513 1824
rect 3807 1816 3853 1824
rect 3867 1816 3953 1824
rect 4227 1816 4373 1824
rect 4587 1816 4673 1824
rect 4907 1816 4924 1824
rect 4916 1807 4924 1816
rect 5007 1816 5233 1824
rect 1896 1796 1973 1804
rect 2167 1796 2633 1804
rect 2647 1796 2684 1804
rect 547 1776 633 1784
rect 1127 1776 1173 1784
rect 1256 1784 1264 1793
rect 1256 1776 1353 1784
rect 1527 1776 1573 1784
rect 1587 1776 1773 1784
rect 1876 1784 1884 1793
rect 1787 1776 2493 1784
rect 2627 1776 2653 1784
rect 2676 1784 2684 1796
rect 2727 1796 2753 1804
rect 2807 1796 2853 1804
rect 2867 1796 2993 1804
rect 3247 1796 3333 1804
rect 3667 1796 3993 1804
rect 4147 1796 4273 1804
rect 4387 1796 4473 1804
rect 5047 1796 5133 1804
rect 5216 1796 5293 1804
rect 2676 1776 2873 1784
rect 3427 1776 3533 1784
rect 3607 1776 3633 1784
rect 3687 1776 3733 1784
rect 3787 1776 3813 1784
rect 3987 1776 4253 1784
rect 4307 1776 4433 1784
rect 4507 1776 4633 1784
rect 4656 1776 4753 1784
rect 216 1764 224 1773
rect 216 1756 313 1764
rect 327 1756 433 1764
rect 507 1756 673 1764
rect 767 1756 813 1764
rect 847 1756 1013 1764
rect 1027 1756 1153 1764
rect 1247 1756 1453 1764
rect 1707 1756 1773 1764
rect 1947 1756 1993 1764
rect 2007 1756 2833 1764
rect 2847 1756 3033 1764
rect 3507 1756 3913 1764
rect 3967 1756 4113 1764
rect 4656 1764 4664 1776
rect 4767 1776 4853 1784
rect 5216 1784 5224 1796
rect 5527 1796 5693 1804
rect 5067 1776 5224 1784
rect 5247 1776 5273 1784
rect 5327 1776 5453 1784
rect 4407 1756 4664 1764
rect 4907 1756 5013 1764
rect 5527 1756 5633 1764
rect 5847 1756 5873 1764
rect 607 1736 873 1744
rect 1787 1736 2553 1744
rect 3627 1736 3653 1744
rect 4687 1736 5493 1744
rect 1447 1716 1753 1724
rect 1767 1716 1833 1724
rect 2027 1716 2233 1724
rect 2307 1716 2773 1724
rect 1367 1696 2133 1704
rect 2247 1696 2293 1704
rect 4707 1696 5193 1704
rect 5207 1696 5213 1704
rect 1227 1676 1353 1684
rect 1907 1676 2633 1684
rect 5207 1676 5353 1684
rect 5507 1676 5673 1684
rect 407 1656 653 1664
rect 667 1656 1273 1664
rect 3367 1656 3733 1664
rect 3927 1656 4753 1664
rect 4767 1656 5033 1664
rect 5047 1656 5153 1664
rect 367 1636 613 1644
rect 627 1636 733 1644
rect 767 1636 913 1644
rect 927 1636 1453 1644
rect 1647 1636 1733 1644
rect 1827 1636 1913 1644
rect 1927 1636 1973 1644
rect 2267 1636 2413 1644
rect 2467 1636 2513 1644
rect 2607 1636 2893 1644
rect 2907 1636 3013 1644
rect 3027 1636 3473 1644
rect 3787 1636 4033 1644
rect 5187 1636 5253 1644
rect 5787 1636 5824 1644
rect 387 1616 433 1624
rect 647 1616 713 1624
rect 827 1616 933 1624
rect 1007 1616 1113 1624
rect 1287 1616 1473 1624
rect 1587 1616 1853 1624
rect 1867 1616 1873 1624
rect 1887 1616 1913 1624
rect 2107 1616 2933 1624
rect 2947 1616 3173 1624
rect 3187 1616 3213 1624
rect 3347 1616 3553 1624
rect 3567 1616 3633 1624
rect 3647 1616 3673 1624
rect 3767 1616 3873 1624
rect 4007 1616 4353 1624
rect 4467 1616 4533 1624
rect 4607 1616 5313 1624
rect 5387 1616 5473 1624
rect 5547 1616 5793 1624
rect 147 1596 193 1604
rect 207 1596 353 1604
rect 427 1596 533 1604
rect 547 1596 833 1604
rect 907 1596 993 1604
rect 1047 1596 1484 1604
rect 47 1576 73 1584
rect 127 1576 273 1584
rect 387 1576 473 1584
rect 787 1576 873 1584
rect 927 1576 1173 1584
rect 1407 1576 1433 1584
rect 1476 1584 1484 1596
rect 1507 1596 1533 1604
rect 1687 1596 1853 1604
rect 1967 1596 2133 1604
rect 2147 1596 2193 1604
rect 2227 1596 2313 1604
rect 2387 1596 2433 1604
rect 2567 1596 3053 1604
rect 3067 1596 3093 1604
rect 3147 1596 3193 1604
rect 3247 1596 3753 1604
rect 3947 1596 4153 1604
rect 4207 1596 4393 1604
rect 4627 1596 4653 1604
rect 4847 1596 4973 1604
rect 5367 1596 5453 1604
rect 5607 1596 5744 1604
rect 1476 1576 1513 1584
rect 1567 1576 1593 1584
rect 1627 1576 1653 1584
rect 1707 1576 1793 1584
rect 1947 1576 1973 1584
rect 2247 1576 2333 1584
rect 2436 1584 2444 1593
rect 2436 1576 2593 1584
rect 2607 1576 2673 1584
rect 2747 1576 2973 1584
rect 3007 1576 3053 1584
rect 3107 1576 3153 1584
rect 3407 1576 3453 1584
rect 3747 1576 3764 1584
rect 267 1556 353 1564
rect 367 1556 493 1564
rect 607 1556 753 1564
rect 1327 1556 1893 1564
rect 2107 1556 2133 1564
rect 2507 1556 2573 1564
rect 2627 1556 2713 1564
rect 2927 1556 3073 1564
rect 3087 1556 3253 1564
rect 3576 1564 3584 1573
rect 3576 1556 3593 1564
rect 3756 1564 3764 1576
rect 3787 1576 3893 1584
rect 3907 1576 4073 1584
rect 4427 1576 4653 1584
rect 4707 1576 4773 1584
rect 4796 1567 4804 1593
rect 4927 1576 4993 1584
rect 5007 1576 5173 1584
rect 5336 1584 5344 1593
rect 5736 1587 5744 1596
rect 5336 1576 5593 1584
rect 5616 1576 5733 1584
rect 3756 1556 3853 1564
rect 4347 1556 4433 1564
rect 4447 1556 4513 1564
rect 4947 1556 5333 1564
rect 5347 1556 5413 1564
rect 5616 1564 5624 1576
rect 5587 1556 5624 1564
rect 5747 1556 5773 1564
rect 127 1536 173 1544
rect 727 1536 1253 1544
rect 1267 1536 1313 1544
rect 1867 1536 2493 1544
rect 2687 1536 2873 1544
rect 3067 1536 3093 1544
rect 3727 1536 4833 1544
rect 4847 1536 4873 1544
rect 5816 1544 5824 1636
rect 5767 1536 5824 1544
rect 187 1516 513 1524
rect 527 1516 793 1524
rect 1427 1516 1573 1524
rect 1587 1516 1733 1524
rect 2327 1516 2753 1524
rect 3007 1516 3133 1524
rect 3667 1516 4073 1524
rect 4387 1516 4673 1524
rect 4687 1516 5533 1524
rect 1427 1496 1713 1504
rect 1867 1496 3273 1504
rect 2107 1456 3473 1464
rect 3487 1456 4553 1464
rect 4567 1456 4633 1464
rect 3627 1436 4413 1444
rect 2387 1416 2413 1424
rect 1107 1396 1613 1404
rect 3307 1396 3553 1404
rect 3567 1396 4133 1404
rect 5147 1396 5333 1404
rect 1507 1376 1953 1384
rect 2027 1376 2053 1384
rect 2147 1376 2173 1384
rect 2987 1376 4353 1384
rect 4927 1376 4953 1384
rect 4967 1376 5433 1384
rect 347 1356 3113 1364
rect 3387 1356 3433 1364
rect 3447 1356 3873 1364
rect 3887 1356 4053 1364
rect 4527 1356 4673 1364
rect 5207 1356 5453 1364
rect -24 1336 13 1344
rect 27 1336 333 1344
rect 767 1336 953 1344
rect 1227 1336 1253 1344
rect 1447 1336 1504 1344
rect 47 1316 93 1324
rect 167 1316 193 1324
rect 207 1316 344 1324
rect 336 1304 344 1316
rect 367 1316 433 1324
rect 827 1316 913 1324
rect 336 1296 573 1304
rect 976 1304 984 1333
rect 1496 1327 1504 1336
rect 2047 1336 2193 1344
rect 2207 1336 2833 1344
rect 2847 1336 2993 1344
rect 3107 1336 3153 1344
rect 3187 1336 3253 1344
rect 3407 1336 3424 1344
rect 3416 1327 3424 1336
rect 3527 1336 3573 1344
rect 4027 1336 4293 1344
rect 4307 1336 4633 1344
rect 5107 1336 5213 1344
rect 5247 1336 5273 1344
rect 5327 1336 5353 1344
rect 5427 1336 5553 1344
rect 1147 1316 1193 1324
rect 1247 1316 1353 1324
rect 1667 1316 1753 1324
rect 2067 1316 2153 1324
rect 2587 1316 2673 1324
rect 2727 1316 2773 1324
rect 2887 1316 2973 1324
rect 3147 1316 3273 1324
rect 3547 1316 3593 1324
rect 3647 1316 3813 1324
rect 3827 1316 3833 1324
rect 3927 1316 4033 1324
rect 4087 1316 4153 1324
rect 4267 1316 4313 1324
rect 4427 1316 4473 1324
rect 4567 1316 4653 1324
rect 4707 1316 4773 1324
rect 4907 1316 4993 1324
rect 5047 1316 5073 1324
rect 5107 1316 5133 1324
rect 5187 1316 5293 1324
rect 5507 1316 5593 1324
rect 5727 1316 5773 1324
rect 947 1296 984 1304
rect 1067 1296 1233 1304
rect 1947 1296 1993 1304
rect 2187 1296 2313 1304
rect 2447 1296 2533 1304
rect 2667 1296 2693 1304
rect 2767 1296 3113 1304
rect 3407 1296 3713 1304
rect 4967 1296 5053 1304
rect 5127 1296 5353 1304
rect 5487 1296 5513 1304
rect 5627 1296 5653 1304
rect 867 1276 973 1284
rect 1447 1276 1573 1284
rect 2367 1276 2793 1284
rect 2827 1276 2933 1284
rect 3307 1276 3673 1284
rect 3687 1276 3933 1284
rect 4207 1276 4393 1284
rect 4647 1276 4753 1284
rect 4767 1276 4853 1284
rect 5167 1276 5573 1284
rect 387 1256 613 1264
rect 707 1256 1033 1264
rect 1047 1256 1113 1264
rect 1127 1256 1173 1264
rect 1187 1256 1873 1264
rect 2027 1236 3033 1244
rect 3047 1236 3253 1244
rect 3467 1236 3833 1244
rect 3847 1236 3853 1244
rect 3947 1236 4693 1244
rect 5027 1236 5433 1244
rect 2527 1216 2873 1224
rect 2927 1216 3993 1224
rect 1967 1196 3013 1204
rect 3167 1196 3353 1204
rect 3367 1196 3473 1204
rect 3527 1196 3573 1204
rect 3587 1196 3693 1204
rect 4047 1196 4533 1204
rect 5167 1196 5453 1204
rect 647 1176 1053 1184
rect 2627 1176 2733 1184
rect 4087 1176 4473 1184
rect 4487 1176 4933 1184
rect 5227 1176 5313 1184
rect 5367 1176 5873 1184
rect 587 1156 593 1164
rect 607 1156 933 1164
rect 1647 1156 1973 1164
rect 1987 1156 2153 1164
rect 2747 1156 3073 1164
rect 3347 1156 3893 1164
rect 4127 1156 5153 1164
rect 5407 1156 5573 1164
rect 87 1136 173 1144
rect 727 1136 753 1144
rect 1627 1136 1713 1144
rect 1727 1136 1853 1144
rect 2227 1136 2633 1144
rect 2687 1136 2993 1144
rect 3007 1136 3053 1144
rect 3067 1136 3113 1144
rect 3127 1136 3573 1144
rect 3627 1136 3713 1144
rect 3907 1136 4433 1144
rect 4727 1136 5013 1144
rect 5147 1136 5253 1144
rect 5347 1136 5413 1144
rect 127 1116 153 1124
rect 427 1116 653 1124
rect 907 1116 1133 1124
rect 1347 1116 1453 1124
rect 1467 1116 1593 1124
rect 1607 1116 1673 1124
rect 1687 1116 1873 1124
rect 1887 1116 2253 1124
rect 2267 1116 2393 1124
rect 2407 1116 2613 1124
rect 2827 1116 3293 1124
rect 3567 1116 3853 1124
rect 4167 1116 4193 1124
rect 4267 1116 4293 1124
rect 4347 1116 4373 1124
rect 4567 1116 4633 1124
rect 4767 1116 4813 1124
rect 4947 1116 4973 1124
rect 4987 1116 5113 1124
rect 5247 1116 5273 1124
rect 5407 1116 5533 1124
rect 5547 1116 5644 1124
rect 67 1096 93 1104
rect 147 1096 253 1104
rect 407 1096 513 1104
rect 687 1096 733 1104
rect 1087 1096 1113 1104
rect 1307 1096 1393 1104
rect 1567 1096 1813 1104
rect 2327 1096 2433 1104
rect 2787 1096 3153 1104
rect 3167 1096 3453 1104
rect 3747 1096 3873 1104
rect 3887 1096 4273 1104
rect 4676 1104 4684 1113
rect 5636 1107 5644 1116
rect 5696 1116 5773 1124
rect 5696 1107 5704 1116
rect 5827 1116 5873 1124
rect 4567 1096 4684 1104
rect 5007 1096 5213 1104
rect 5307 1096 5333 1104
rect 107 1076 233 1084
rect 247 1076 353 1084
rect 367 1076 493 1084
rect 787 1076 1273 1084
rect 1447 1076 1453 1084
rect 1467 1076 1533 1084
rect 2467 1076 2733 1084
rect 2747 1076 2833 1084
rect 3027 1076 3293 1084
rect 3327 1076 3493 1084
rect 3507 1076 3593 1084
rect 4307 1076 4373 1084
rect 4847 1076 5173 1084
rect 5227 1076 5513 1084
rect 1027 1056 1433 1064
rect 1867 1056 2933 1064
rect 5107 1056 5153 1064
rect 1107 1036 1993 1044
rect 2007 1036 2093 1044
rect 2247 1036 2273 1044
rect 2287 1036 2553 1044
rect 4267 1036 5293 1044
rect 307 1016 833 1024
rect 1147 1016 1153 1024
rect 1167 1016 4593 1024
rect 4707 1016 5133 1024
rect 5487 1016 5553 1024
rect 2027 996 2913 1004
rect 3927 996 4473 1004
rect 4487 996 4733 1004
rect 4747 996 5613 1004
rect 4207 976 4873 984
rect 4367 956 4593 964
rect 4427 936 5073 944
rect 5087 936 5353 944
rect 4547 916 4613 924
rect 547 896 973 904
rect 987 896 2013 904
rect 2067 896 2313 904
rect 3827 896 5193 904
rect 5207 896 5373 904
rect 5387 896 5513 904
rect 287 876 1093 884
rect 1207 876 1493 884
rect 1867 876 1933 884
rect 2187 876 2693 884
rect 4467 876 4913 884
rect 407 856 473 864
rect 527 856 553 864
rect 847 856 1013 864
rect 1027 856 1133 864
rect 1267 856 1293 864
rect 1307 856 1893 864
rect 1907 856 2053 864
rect 2207 856 2233 864
rect 2247 856 2453 864
rect 2507 856 2593 864
rect 2647 856 2673 864
rect 2756 856 2873 864
rect 2756 847 2764 856
rect 3067 856 3413 864
rect 3707 856 3724 864
rect 3716 847 3724 856
rect 3987 856 4364 864
rect 327 836 453 844
rect 647 836 804 844
rect 47 816 73 824
rect 107 816 173 824
rect 367 816 553 824
rect 607 816 653 824
rect 747 816 773 824
rect 796 824 804 836
rect 887 836 993 844
rect 1087 836 1113 844
rect 1207 836 1253 844
rect 1287 836 1373 844
rect 1567 836 1653 844
rect 2087 836 2153 844
rect 2167 836 2313 844
rect 2527 836 2573 844
rect 2807 836 2913 844
rect 2927 836 3033 844
rect 3187 836 3253 844
rect 3276 836 3293 844
rect 796 816 853 824
rect 1407 816 1573 824
rect 1847 816 1913 824
rect 1927 816 1933 824
rect 1987 816 2213 824
rect 2347 816 2613 824
rect 2707 816 2773 824
rect 2787 816 2993 824
rect 3087 816 3193 824
rect 3276 824 3284 836
rect 3367 836 3393 844
rect 3587 836 3673 844
rect 3827 836 3853 844
rect 3867 836 3893 844
rect 4127 836 4213 844
rect 4287 836 4333 844
rect 4356 844 4364 856
rect 4387 856 4453 864
rect 4687 856 4784 864
rect 4496 844 4504 853
rect 4356 836 4504 844
rect 4667 836 4733 844
rect 4776 844 4784 856
rect 4807 856 4833 864
rect 4776 836 4953 844
rect 5107 836 5133 844
rect 5567 836 5873 844
rect 3207 816 3284 824
rect 3327 816 3653 824
rect 4076 824 4084 833
rect 3967 816 4084 824
rect 4327 816 4353 824
rect 4527 816 4633 824
rect 4647 816 4713 824
rect 4827 816 4924 824
rect 127 796 593 804
rect 1447 796 1633 804
rect 1647 796 1753 804
rect 1947 796 2433 804
rect 2447 796 2493 804
rect 3147 796 3273 804
rect 3427 796 3593 804
rect 3707 796 4133 804
rect 4147 796 4233 804
rect 4407 796 4573 804
rect 4587 796 4893 804
rect 4916 804 4924 816
rect 5056 824 5064 833
rect 4947 816 5064 824
rect 5087 816 5473 824
rect 5507 816 5633 824
rect 5767 816 5864 824
rect 5856 807 5864 816
rect 4916 796 5033 804
rect 1247 776 1453 784
rect 1807 776 2113 784
rect 2307 776 2373 784
rect 2427 776 2473 784
rect 2487 776 2713 784
rect 2907 776 3433 784
rect 4247 776 4613 784
rect 4627 776 4773 784
rect 1047 756 1313 764
rect 1327 756 1793 764
rect 3367 756 3793 764
rect 4667 756 5333 764
rect 867 736 1353 744
rect 1787 736 2173 744
rect 2187 736 2353 744
rect 2387 736 2853 744
rect 827 716 953 724
rect 1287 716 1813 724
rect 2367 716 2433 724
rect 2447 716 2613 724
rect 3027 716 3353 724
rect 3787 716 3913 724
rect 4247 716 4453 724
rect 5587 716 5693 724
rect 667 696 1973 704
rect 2347 696 2773 704
rect 3327 696 3973 704
rect 4387 696 4513 704
rect 4567 696 5113 704
rect 5527 696 5613 704
rect 247 676 373 684
rect 387 676 613 684
rect 807 676 873 684
rect 1007 676 1153 684
rect 1167 676 1633 684
rect 1667 676 1793 684
rect 2047 676 2233 684
rect 2247 676 2353 684
rect 3047 676 3093 684
rect 3107 676 3153 684
rect 3767 676 3833 684
rect 4207 676 4673 684
rect 5107 676 5113 684
rect 5127 676 5373 684
rect 5387 676 5673 684
rect 827 656 1013 664
rect 1167 656 1213 664
rect 1487 656 1773 664
rect 1827 656 2413 664
rect 2827 656 2833 664
rect 2847 656 2873 664
rect 3167 656 3453 664
rect 3467 656 3524 664
rect 216 636 313 644
rect 216 627 224 636
rect 327 636 413 644
rect 507 636 524 644
rect 227 616 233 624
rect 496 584 504 613
rect 516 607 524 636
rect 627 636 833 644
rect 847 636 853 644
rect 927 636 993 644
rect 1016 636 1033 644
rect 547 616 733 624
rect 1016 624 1024 636
rect 1267 636 1653 644
rect 1727 636 1933 644
rect 1987 636 2064 644
rect 2056 627 2064 636
rect 2167 636 2324 644
rect 2316 627 2324 636
rect 2487 636 2533 644
rect 2567 636 2733 644
rect 3007 636 3113 644
rect 3516 644 3524 656
rect 3547 656 4433 664
rect 5487 656 5713 664
rect 5727 656 5733 664
rect 3516 636 3773 644
rect 3847 636 3953 644
rect 3967 636 4093 644
rect 4107 636 4204 644
rect 907 616 1024 624
rect 1427 616 1673 624
rect 1927 616 2033 624
rect 2076 616 2193 624
rect 767 596 813 604
rect 827 596 873 604
rect 1147 596 1273 604
rect 1407 596 1553 604
rect 1967 596 1973 604
rect 2076 604 2084 616
rect 2427 616 2453 624
rect 2507 616 2593 624
rect 2647 616 2713 624
rect 2907 616 2933 624
rect 3227 616 3293 624
rect 3347 616 3433 624
rect 3807 616 3853 624
rect 3876 616 3933 624
rect 1987 596 2084 604
rect 2667 596 2753 604
rect 3107 596 3173 604
rect 3876 604 3884 616
rect 3987 616 4053 624
rect 4107 616 4153 624
rect 4196 624 4204 636
rect 4227 636 4453 644
rect 4807 636 4853 644
rect 5167 636 5213 644
rect 5347 636 5593 644
rect 4196 616 4233 624
rect 4407 616 4493 624
rect 4607 616 4873 624
rect 4987 616 5173 624
rect 5287 616 5453 624
rect 5527 616 5613 624
rect 5667 616 5713 624
rect 5827 616 5853 624
rect 3627 596 3884 604
rect 4187 596 4353 604
rect 4367 596 5133 604
rect 5147 596 5573 604
rect 5787 596 5833 604
rect 496 576 1693 584
rect 3487 576 3653 584
rect 3667 576 4313 584
rect 5547 576 5593 584
rect 5707 576 5793 584
rect 267 556 333 564
rect 347 556 533 564
rect 3307 556 3553 564
rect 4207 556 4693 564
rect 1967 536 4253 544
rect 1067 496 2273 504
rect 2427 476 3513 484
rect 4047 456 4153 464
rect 2067 436 2353 444
rect 2807 436 3193 444
rect 3927 436 4253 444
rect 4887 436 5053 444
rect 5067 436 5193 444
rect 747 416 793 424
rect 2047 416 2173 424
rect 2667 416 3173 424
rect 3207 416 4073 424
rect 4087 416 4093 424
rect 4147 416 4353 424
rect 4407 416 4433 424
rect 4447 416 4473 424
rect 4487 416 5413 424
rect 87 396 413 404
rect 807 396 833 404
rect 1547 396 1753 404
rect 2196 396 2493 404
rect 947 376 973 384
rect 1027 376 1093 384
rect 1567 376 1593 384
rect 1627 376 1653 384
rect 1907 376 2073 384
rect 2196 384 2204 396
rect 2687 396 3253 404
rect 3267 396 3453 404
rect 3527 396 4173 404
rect 4927 396 5013 404
rect 5027 396 5113 404
rect 5427 396 5533 404
rect 2087 376 2204 384
rect 2227 376 2353 384
rect 2407 376 2533 384
rect 2767 376 2913 384
rect 2927 376 3124 384
rect 47 356 73 364
rect 227 356 344 364
rect 116 327 124 353
rect 147 336 173 344
rect 336 344 344 356
rect 367 356 453 364
rect 716 364 724 373
rect 3116 367 3124 376
rect 3147 376 3333 384
rect 3467 376 4013 384
rect 4027 376 4033 384
rect 4227 376 4433 384
rect 4447 376 4633 384
rect 4647 376 4813 384
rect 5307 376 5413 384
rect 607 356 833 364
rect 676 347 684 356
rect 1267 356 1433 364
rect 1447 356 1473 364
rect 1527 356 1593 364
rect 1607 356 1713 364
rect 1987 356 2093 364
rect 2107 356 2233 364
rect 2387 356 2673 364
rect 2687 356 2773 364
rect 2907 356 2953 364
rect 2967 356 3073 364
rect 3187 356 3373 364
rect 3387 356 3533 364
rect 3587 356 3613 364
rect 3747 356 3833 364
rect 4467 356 4513 364
rect 4676 356 4753 364
rect 336 336 473 344
rect 907 336 1053 344
rect 1147 336 1444 344
rect 527 316 933 324
rect 947 316 1073 324
rect 1347 316 1393 324
rect 1436 324 1444 336
rect 1467 336 1533 344
rect 1627 336 1873 344
rect 2147 336 2693 344
rect 2707 336 2804 344
rect 2796 327 2804 336
rect 3287 336 3393 344
rect 3696 344 3704 353
rect 3567 336 3704 344
rect 3947 336 4053 344
rect 4287 336 4313 344
rect 4507 336 4593 344
rect 4676 344 4684 356
rect 4807 356 4853 364
rect 5047 356 5353 364
rect 5407 356 5493 364
rect 5507 356 5673 364
rect 5807 356 5833 364
rect 4667 336 4684 344
rect 4707 336 4733 344
rect 4827 336 4933 344
rect 5567 336 5713 344
rect 1436 316 1493 324
rect 1507 316 1573 324
rect 1707 316 1733 324
rect 1827 316 1933 324
rect 2527 316 2753 324
rect 2947 316 3093 324
rect 3467 316 3593 324
rect 3727 316 4113 324
rect 4347 316 4453 324
rect 4467 316 4653 324
rect 4787 316 4893 324
rect 4907 316 5033 324
rect 5167 316 5273 324
rect 5607 316 5693 324
rect 107 296 1093 304
rect 1107 296 1273 304
rect 1447 296 2113 304
rect 2287 296 2933 304
rect 2987 296 3873 304
rect 3887 296 3933 304
rect 4307 296 4433 304
rect 4587 296 4613 304
rect 4887 296 5513 304
rect 5527 296 5653 304
rect 1647 276 1793 284
rect 1807 276 2933 284
rect 2947 276 3053 284
rect 3507 276 5233 284
rect 5467 276 5513 284
rect 5527 276 5793 284
rect 1867 256 1913 264
rect 1927 256 2173 264
rect 2847 256 3613 264
rect 3627 256 3893 264
rect 3907 256 3913 264
rect 4127 256 4193 264
rect 107 236 293 244
rect 307 236 353 244
rect 407 236 573 244
rect 587 236 813 244
rect 827 236 1033 244
rect 1747 236 1913 244
rect 1947 236 3673 244
rect 4067 236 4573 244
rect 4587 236 4693 244
rect 347 216 493 224
rect 507 216 793 224
rect 867 216 973 224
rect 987 216 1073 224
rect 1387 216 2753 224
rect 2787 216 3153 224
rect 3367 216 3813 224
rect 4107 216 4153 224
rect 5327 216 5793 224
rect 467 196 833 204
rect 847 196 1233 204
rect 1256 196 1453 204
rect 927 176 1113 184
rect 1256 184 1264 196
rect 1567 196 2533 204
rect 2547 196 2633 204
rect 2647 196 2873 204
rect 2927 196 3033 204
rect 3067 196 3373 204
rect 3387 196 3473 204
rect 3636 196 4513 204
rect 1187 176 1264 184
rect 1407 176 1884 184
rect 547 156 633 164
rect 687 156 944 164
rect 136 144 144 153
rect 136 136 213 144
rect 227 136 313 144
rect 387 136 453 144
rect 527 136 573 144
rect 707 136 773 144
rect 936 144 944 156
rect 967 156 1144 164
rect 1136 147 1144 156
rect 1167 156 1284 164
rect 1276 147 1284 156
rect 936 136 1113 144
rect 667 116 713 124
rect 867 116 913 124
rect 927 116 953 124
rect 1296 124 1304 173
rect 1876 164 1884 176
rect 1907 176 1933 184
rect 2296 176 2513 184
rect 2296 164 2304 176
rect 2527 176 3173 184
rect 3187 176 3313 184
rect 3447 176 3613 184
rect 1467 156 1564 164
rect 1876 156 2304 164
rect 1327 136 1373 144
rect 1007 116 1413 124
rect 1536 124 1544 133
rect 1556 127 1564 156
rect 2367 156 2593 164
rect 2687 156 2793 164
rect 2807 156 2993 164
rect 3167 156 3344 164
rect 1707 136 1813 144
rect 1927 136 1944 144
rect 1427 116 1544 124
rect 1607 116 1653 124
rect 1767 116 1913 124
rect 1936 124 1944 136
rect 2027 136 2153 144
rect 2316 144 2324 153
rect 2227 136 2324 144
rect 2387 136 2413 144
rect 2616 144 2624 153
rect 3336 147 3344 156
rect 3367 156 3453 164
rect 3636 147 3644 196
rect 5107 196 5133 204
rect 5147 196 5653 204
rect 3927 176 4353 184
rect 4367 176 4413 184
rect 4987 176 5093 184
rect 5136 176 5433 184
rect 3667 156 3693 164
rect 3716 156 3773 164
rect 2507 136 2893 144
rect 3087 136 3293 144
rect 3716 144 3724 156
rect 4207 156 4273 164
rect 4287 156 4453 164
rect 5136 164 5144 176
rect 5796 176 5813 184
rect 4747 156 5144 164
rect 5487 156 5613 164
rect 5796 164 5804 176
rect 5747 156 5804 164
rect 5827 156 5853 164
rect 3687 136 3724 144
rect 3807 136 3873 144
rect 4067 136 4173 144
rect 4527 136 4553 144
rect 4567 136 4713 144
rect 5027 136 5313 144
rect 5467 136 5553 144
rect 5767 136 5853 144
rect 1936 116 2473 124
rect 2907 116 3693 124
rect 3847 116 4053 124
rect 4407 116 4593 124
rect 4756 124 4764 133
rect 4647 116 4764 124
rect 5227 116 5253 124
rect 5267 116 5293 124
rect 5347 116 5493 124
rect 5507 116 5593 124
rect 5827 116 5873 124
rect 1247 96 1753 104
rect 1787 96 2333 104
rect 3247 96 3473 104
rect 5807 96 5833 104
rect 1027 76 1873 84
rect 2607 76 4953 84
rect 1747 36 2133 44
rect 1647 16 1693 24
rect 1847 16 1873 24
rect 4547 16 4613 24
use INVX1  _863_
timestamp 0
transform 1 0 5130 0 1 5050
box -6 -8 66 248
use NAND2X1  _864_
timestamp 0
transform -1 0 4970 0 -1 6010
box -6 -8 86 248
use OAI21X1  _865_
timestamp 0
transform 1 0 5370 0 1 5050
box -6 -8 106 248
use NOR2X1  _866_
timestamp 0
transform -1 0 5490 0 -1 5530
box -6 -8 86 248
use INVX1  _867_
timestamp 0
transform 1 0 5290 0 -1 5530
box -6 -8 66 248
use NAND2X1  _868_
timestamp 0
transform -1 0 4470 0 -1 5050
box -6 -8 86 248
use INVX2  _869_
timestamp 0
transform -1 0 5270 0 -1 3610
box -6 -8 66 248
use NAND2X1  _870_
timestamp 0
transform 1 0 5530 0 -1 5530
box -6 -8 86 248
use OAI21X1  _871_
timestamp 0
transform -1 0 5190 0 -1 5050
box -6 -8 106 248
use AOI21X1  _872_
timestamp 0
transform 1 0 5530 0 1 5050
box -6 -8 106 248
use NOR2X1  _873_
timestamp 0
transform 1 0 5750 0 1 2650
box -6 -8 86 248
use INVX2  _874_
timestamp 0
transform 1 0 5810 0 -1 5530
box -6 -8 66 248
use INVX1  _875_
timestamp 0
transform -1 0 5510 0 -1 3130
box -6 -8 66 248
use NOR2X1  _876_
timestamp 0
transform 1 0 5330 0 -1 3130
box -6 -8 86 248
use AOI22X1  _877_
timestamp 0
transform -1 0 5310 0 1 4090
box -6 -8 126 248
use OAI21X1  _878_
timestamp 0
transform -1 0 5330 0 1 5050
box -6 -8 106 248
use INVX1  _879_
timestamp 0
transform 1 0 5190 0 -1 5530
box -6 -8 66 248
use NAND2X1  _880_
timestamp 0
transform -1 0 5210 0 1 5530
box -6 -8 86 248
use OAI21X1  _881_
timestamp 0
transform -1 0 5350 0 1 5530
box -6 -8 106 248
use INVX1  _882_
timestamp 0
transform 1 0 3390 0 -1 6010
box -6 -8 66 248
use NAND2X1  _883_
timestamp 0
transform 1 0 3790 0 1 5530
box -6 -8 86 248
use OAI21X1  _884_
timestamp 0
transform 1 0 3630 0 1 5530
box -6 -8 106 248
use AOI21X1  _885_
timestamp 0
transform 1 0 5410 0 1 5530
box -6 -8 106 248
use AOI22X1  _886_
timestamp 0
transform 1 0 5450 0 1 4570
box -6 -8 126 248
use OAI21X1  _887_
timestamp 0
transform -1 0 5650 0 1 5530
box -6 -8 106 248
use INVX1  _888_
timestamp 0
transform 1 0 5330 0 1 730
box -6 -8 66 248
use NAND2X1  _889_
timestamp 0
transform -1 0 4930 0 1 1210
box -6 -8 86 248
use OAI21X1  _890_
timestamp 0
transform -1 0 5070 0 1 1210
box -6 -8 106 248
use INVX1  _891_
timestamp 0
transform 1 0 5810 0 1 250
box -6 -8 66 248
use INVX1  _892_
timestamp 0
transform -1 0 4870 0 -1 1210
box -6 -8 66 248
use OAI22X1  _893_
timestamp 0
transform 1 0 5150 0 -1 1210
box -6 -8 126 248
use AOI21X1  _894_
timestamp 0
transform 1 0 5410 0 1 1210
box -6 -8 106 248
use AOI22X1  _895_
timestamp 0
transform -1 0 5650 0 1 2170
box -6 -8 126 248
use OAI21X1  _896_
timestamp 0
transform -1 0 5810 0 -1 2170
box -6 -8 106 248
use INVX1  _897_
timestamp 0
transform 1 0 5490 0 -1 2170
box -6 -8 66 248
use INVX1  _898_
timestamp 0
transform -1 0 5010 0 -1 730
box -6 -8 66 248
use NAND2X1  _899_
timestamp 0
transform 1 0 5270 0 1 1210
box -6 -8 86 248
use OAI21X1  _900_
timestamp 0
transform 1 0 5110 0 1 1210
box -6 -8 106 248
use INVX1  _901_
timestamp 0
transform -1 0 5670 0 -1 1210
box -6 -8 66 248
use INVX1  _902_
timestamp 0
transform 1 0 5850 0 1 730
box -6 -8 66 248
use OAI22X1  _903_
timestamp 0
transform 1 0 5450 0 -1 1210
box -6 -8 126 248
use AOI21X1  _904_
timestamp 0
transform 1 0 5550 0 1 1210
box -6 -8 106 248
use AOI22X1  _905_
timestamp 0
transform 1 0 5710 0 -1 1690
box -6 -8 126 248
use OAI21X1  _906_
timestamp 0
transform 1 0 5690 0 1 2170
box -6 -8 106 248
use INVX1  _907_
timestamp 0
transform 1 0 1890 0 -1 5530
box -6 -8 66 248
use NAND2X1  _908_
timestamp 0
transform -1 0 1370 0 -1 6010
box -6 -8 86 248
use OAI21X1  _909_
timestamp 0
transform 1 0 1910 0 1 5530
box -6 -8 106 248
use INVX1  _910_
timestamp 0
transform 1 0 1670 0 -1 6010
box -6 -8 66 248
use INVX1  _911_
timestamp 0
transform 1 0 2830 0 1 5530
box -6 -8 66 248
use OAI22X1  _912_
timestamp 0
transform -1 0 2550 0 -1 5530
box -6 -8 126 248
use AOI21X1  _913_
timestamp 0
transform 1 0 2770 0 -1 5530
box -6 -8 106 248
use AOI22X1  _914_
timestamp 0
transform -1 0 4470 0 -1 4570
box -6 -8 126 248
use OAI21X1  _915_
timestamp 0
transform 1 0 4310 0 1 5050
box -6 -8 106 248
use INVX1  _916_
timestamp 0
transform 1 0 1270 0 -1 5530
box -6 -8 66 248
use NAND2X1  _917_
timestamp 0
transform -1 0 1550 0 -1 5530
box -6 -8 86 248
use OAI21X1  _918_
timestamp 0
transform 1 0 1750 0 -1 5530
box -6 -8 106 248
use INVX1  _919_
timestamp 0
transform 1 0 1170 0 -1 6010
box -6 -8 66 248
use INVX1  _920_
timestamp 0
transform -1 0 2230 0 -1 5530
box -6 -8 66 248
use OAI22X1  _921_
timestamp 0
transform -1 0 2390 0 -1 5530
box -6 -8 126 248
use AOI21X1  _922_
timestamp 0
transform -1 0 2710 0 -1 5530
box -6 -8 106 248
use AOI22X1  _923_
timestamp 0
transform -1 0 4650 0 1 4570
box -6 -8 126 248
use OAI21X1  _924_
timestamp 0
transform 1 0 4550 0 -1 5530
box -6 -8 106 248
use INVX1  _925_
timestamp 0
transform -1 0 5650 0 -1 2650
box -6 -8 66 248
use INVX1  _926_
timestamp 0
transform -1 0 4410 0 1 1690
box -6 -8 66 248
use INVX8  _927_
timestamp 0
transform 1 0 1070 0 -1 2650
box -6 -8 126 248
use INVX1  _928_
timestamp 0
transform -1 0 3050 0 1 3130
box -6 -8 66 248
use NAND2X1  _929_
timestamp 0
transform -1 0 3010 0 -1 3130
box -6 -8 86 248
use OAI21X1  _930_
timestamp 0
transform -1 0 3170 0 -1 3130
box -6 -8 106 248
use INVX1  _931_
timestamp 0
transform 1 0 4070 0 1 3130
box -6 -8 66 248
use NAND2X1  _932_
timestamp 0
transform -1 0 4050 0 -1 2650
box -6 -8 86 248
use OAI21X1  _933_
timestamp 0
transform -1 0 4130 0 1 2650
box -6 -8 106 248
use MUX2X1  _934_
timestamp 0
transform 1 0 3070 0 1 2650
box -6 -8 126 248
use INVX1  _935_
timestamp 0
transform 1 0 1270 0 -1 3130
box -6 -8 66 248
use NAND2X1  _936_
timestamp 0
transform -1 0 1170 0 1 2650
box -6 -8 86 248
use OAI21X1  _937_
timestamp 0
transform -1 0 1310 0 1 2650
box -6 -8 106 248
use INVX1  _938_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 66 248
use NAND2X1  _939_
timestamp 0
transform 1 0 1990 0 1 3130
box -6 -8 86 248
use OAI21X1  _940_
timestamp 0
transform 1 0 1850 0 1 3130
box -6 -8 106 248
use MUX2X1  _941_
timestamp 0
transform 1 0 1510 0 -1 2650
box -6 -8 126 248
use MUX2X1  _942_
timestamp 0
transform -1 0 3110 0 1 2170
box -6 -8 126 248
use NOR2X1  _943_
timestamp 0
transform -1 0 4350 0 1 2170
box -6 -8 86 248
use NAND2X1  _944_
timestamp 0
transform -1 0 4230 0 1 2170
box -6 -8 86 248
use INVX1  _945_
timestamp 0
transform -1 0 4590 0 1 2170
box -6 -8 66 248
use INVX4  _946_
timestamp 0
transform 1 0 1830 0 1 1690
box -6 -8 86 248
use NAND2X1  _947_
timestamp 0
transform -1 0 2330 0 -1 2650
box -6 -8 86 248
use OAI21X1  _948_
timestamp 0
transform 1 0 2330 0 1 4090
box -6 -8 106 248
use INVX2  _949_
timestamp 0
transform -1 0 1090 0 1 4570
box -6 -8 66 248
use OAI21X1  _950_
timestamp 0
transform 1 0 4390 0 1 2170
box -6 -8 106 248
use OAI21X1  _951_
timestamp 0
transform -1 0 5550 0 -1 2650
box -6 -8 106 248
use INVX8  _952_
timestamp 0
transform -1 0 5610 0 -1 5050
box -6 -8 126 248
use NAND2X1  _953_
timestamp 0
transform 1 0 5570 0 -1 1690
box -6 -8 86 248
use NOR2X1  _954_
timestamp 0
transform -1 0 4170 0 -1 2650
box -6 -8 86 248
use NAND2X1  _955_
timestamp 0
transform 1 0 3490 0 -1 2650
box -6 -8 86 248
use INVX2  _956_
timestamp 0
transform 1 0 3510 0 -1 730
box -6 -8 66 248
use MUX2X1  _957_
timestamp 0
transform -1 0 3110 0 -1 2650
box -6 -8 126 248
use MUX2X1  _958_
timestamp 0
transform -1 0 3930 0 -1 2650
box -6 -8 126 248
use MUX2X1  _959_
timestamp 0
transform 1 0 2830 0 -1 2650
box -6 -8 126 248
use MUX2X1  _960_
timestamp 0
transform -1 0 1230 0 -1 3130
box -6 -8 126 248
use MUX2X1  _961_
timestamp 0
transform -1 0 2230 0 -1 3130
box -6 -8 126 248
use MUX2X1  _962_
timestamp 0
transform 1 0 1430 0 1 2170
box -6 -8 126 248
use MUX2X1  _963_
timestamp 0
transform -1 0 2950 0 1 2170
box -6 -8 126 248
use INVX1  _964_
timestamp 0
transform 1 0 4110 0 1 1690
box -6 -8 66 248
use INVX8  _965_
timestamp 0
transform 1 0 1670 0 -1 4090
box -6 -8 126 248
use INVX1  _966_
timestamp 0
transform -1 0 2510 0 -1 3610
box -6 -8 66 248
use NAND2X1  _967_
timestamp 0
transform 1 0 2310 0 -1 3610
box -6 -8 86 248
use OAI21X1  _968_
timestamp 0
transform -1 0 2430 0 1 3130
box -6 -8 106 248
use INVX1  _969_
timestamp 0
transform -1 0 4290 0 -1 2650
box -6 -8 66 248
use NAND2X1  _970_
timestamp 0
transform 1 0 3590 0 1 2650
box -6 -8 86 248
use OAI21X1  _971_
timestamp 0
transform -1 0 3810 0 1 2650
box -6 -8 106 248
use MUX2X1  _972_
timestamp 0
transform 1 0 2910 0 1 2650
box -6 -8 126 248
use INVX1  _973_
timestamp 0
transform 1 0 1110 0 -1 3610
box -6 -8 66 248
use NAND2X1  _974_
timestamp 0
transform -1 0 1030 0 1 3130
box -6 -8 86 248
use OAI21X1  _975_
timestamp 0
transform -1 0 1170 0 1 3130
box -6 -8 106 248
use INVX1  _976_
timestamp 0
transform -1 0 2050 0 1 4090
box -6 -8 66 248
use NAND2X1  _977_
timestamp 0
transform 1 0 1470 0 1 3130
box -6 -8 86 248
use OAI21X1  _978_
timestamp 0
transform -1 0 1810 0 1 3130
box -6 -8 106 248
use MUX2X1  _979_
timestamp 0
transform 1 0 1790 0 -1 2650
box -6 -8 126 248
use MUX2X1  _980_
timestamp 0
transform 1 0 3170 0 -1 2650
box -6 -8 126 248
use NAND3X1  _981_
timestamp 0
transform 1 0 3270 0 1 2170
box -6 -8 106 248
use MUX2X1  _982_
timestamp 0
transform -1 0 2490 0 -1 2650
box -6 -8 126 248
use MUX2X1  _983_
timestamp 0
transform -1 0 3750 0 -1 2650
box -6 -8 126 248
use MUX2X1  _984_
timestamp 0
transform 1 0 2530 0 -1 2650
box -6 -8 126 248
use MUX2X1  _985_
timestamp 0
transform 1 0 890 0 -1 2650
box -6 -8 126 248
use MUX2X1  _986_
timestamp 0
transform -1 0 1790 0 -1 3130
box -6 -8 126 248
use MUX2X1  _987_
timestamp 0
transform 1 0 1630 0 -1 2170
box -6 -8 126 248
use MUX2X1  _988_
timestamp 0
transform -1 0 2650 0 1 1690
box -6 -8 126 248
use OAI21X1  _989_
timestamp 0
transform -1 0 3550 0 1 1690
box -6 -8 106 248
use AOI21X1  _990_
timestamp 0
transform 1 0 4270 0 -1 2170
box -6 -8 106 248
use INVX1  _991_
timestamp 0
transform 1 0 4710 0 -1 2170
box -6 -8 66 248
use NAND3X1  _992_
timestamp 0
transform 1 0 4410 0 -1 2170
box -6 -8 106 248
use AND2X2  _993_
timestamp 0
transform 1 0 4810 0 -1 2170
box -6 -8 106 248
use OAI21X1  _994_
timestamp 0
transform 1 0 4850 0 1 1690
box -6 -8 106 248
use OR2X2  _995_
timestamp 0
transform 1 0 4950 0 -1 2170
box -6 -8 106 248
use AOI21X1  _996_
timestamp 0
transform 1 0 4990 0 1 1690
box -6 -8 106 248
use OAI21X1  _997_
timestamp 0
transform 1 0 5270 0 1 1690
box -6 -8 106 248
use NAND2X1  _998_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 86 248
use INVX1  _999_
timestamp 0
transform -1 0 4050 0 -1 1690
box -6 -8 66 248
use NAND2X1  _1000_
timestamp 0
transform 1 0 4130 0 1 1210
box -6 -8 86 248
use OAI21X1  _1001_
timestamp 0
transform -1 0 3690 0 1 1690
box -6 -8 106 248
use NAND2X1  _1002_
timestamp 0
transform 1 0 3750 0 1 1690
box -6 -8 86 248
use OAI21X1  _1003_
timestamp 0
transform -1 0 3970 0 -1 2170
box -6 -8 106 248
use MUX2X1  _1004_
timestamp 0
transform 1 0 3710 0 -1 2170
box -6 -8 126 248
use NAND2X1  _1005_
timestamp 0
transform 1 0 3710 0 1 2170
box -6 -8 86 248
use INVX1  _1006_
timestamp 0
transform 1 0 2530 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1007_
timestamp 0
transform 1 0 2410 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1008_
timestamp 0
transform 1 0 2250 0 -1 1210
box -6 -8 106 248
use INVX1  _1009_
timestamp 0
transform -1 0 3530 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1010_
timestamp 0
transform -1 0 3310 0 1 1210
box -6 -8 86 248
use OAI21X1  _1011_
timestamp 0
transform 1 0 3070 0 1 1210
box -6 -8 106 248
use MUX2X1  _1012_
timestamp 0
transform 1 0 2210 0 1 1690
box -6 -8 126 248
use NAND2X1  _1013_
timestamp 0
transform 1 0 3370 0 -1 3130
box -6 -8 86 248
use AND2X2  _1014_
timestamp 0
transform 1 0 3490 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1015_
timestamp 0
transform -1 0 3910 0 1 3130
box -6 -8 86 248
use INVX1  _1016_
timestamp 0
transform -1 0 3570 0 -1 3130
box -6 -8 66 248
use OAI21X1  _1017_
timestamp 0
transform 1 0 3530 0 1 3130
box -6 -8 106 248
use OAI21X1  _1018_
timestamp 0
transform 1 0 4210 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1019_
timestamp 0
transform 1 0 4350 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1020_
timestamp 0
transform 1 0 5050 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1021_
timestamp 0
transform 1 0 4070 0 -1 3610
box -6 -8 86 248
use INVX1  _1022_
timestamp 0
transform 1 0 4390 0 1 1210
box -6 -8 66 248
use NAND2X1  _1023_
timestamp 0
transform -1 0 3570 0 1 1210
box -6 -8 86 248
use OAI21X1  _1024_
timestamp 0
transform -1 0 3650 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1025_
timestamp 0
transform -1 0 4090 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1026_
timestamp 0
transform 1 0 4130 0 -1 2170
box -6 -8 106 248
use MUX2X1  _1027_
timestamp 0
transform 1 0 3530 0 -1 2170
box -6 -8 126 248
use INVX1  _1028_
timestamp 0
transform 1 0 2870 0 -1 730
box -6 -8 66 248
use NAND2X1  _1029_
timestamp 0
transform -1 0 1590 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1030_
timestamp 0
transform -1 0 1890 0 -1 1210
box -6 -8 106 248
use INVX1  _1031_
timestamp 0
transform -1 0 3190 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1032_
timestamp 0
transform -1 0 2610 0 1 1210
box -6 -8 86 248
use OAI21X1  _1033_
timestamp 0
transform -1 0 2750 0 1 1210
box -6 -8 106 248
use MUX2X1  _1034_
timestamp 0
transform 1 0 1950 0 -1 2170
box -6 -8 126 248
use MUX2X1  _1035_
timestamp 0
transform -1 0 3550 0 1 2170
box -6 -8 126 248
use OAI21X1  _1036_
timestamp 0
transform 1 0 4050 0 1 3610
box -6 -8 106 248
use INVX1  _1037_
timestamp 0
transform -1 0 3850 0 -1 3610
box -6 -8 66 248
use NAND3X1  _1038_
timestamp 0
transform 1 0 3910 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1039_
timestamp 0
transform 1 0 4350 0 1 3610
box -6 -8 106 248
use INVX1  _1040_
timestamp 0
transform 1 0 4470 0 -1 4090
box -6 -8 66 248
use NAND3X1  _1041_
timestamp 0
transform 1 0 4210 0 1 3610
box -6 -8 106 248
use NAND3X1  _1042_
timestamp 0
transform 1 0 4330 0 -1 4090
box -6 -8 106 248
use INVX1  _1043_
timestamp 0
transform -1 0 3910 0 1 4090
box -6 -8 66 248
use INVX1  _1044_
timestamp 0
transform -1 0 4150 0 1 4090
box -6 -8 66 248
use OAI21X1  _1045_
timestamp 0
transform -1 0 4050 0 1 4090
box -6 -8 106 248
use AOI21X1  _1046_
timestamp 0
transform 1 0 4210 0 1 4090
box -6 -8 106 248
use OAI21X1  _1047_
timestamp 0
transform 1 0 4910 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1048_
timestamp 0
transform 1 0 4290 0 1 4570
box -6 -8 86 248
use AOI21X1  _1049_
timestamp 0
transform -1 0 4290 0 -1 4090
box -6 -8 106 248
use INVX1  _1050_
timestamp 0
transform 1 0 3650 0 1 4570
box -6 -8 66 248
use INVX1  _1051_
timestamp 0
transform 1 0 750 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1052_
timestamp 0
transform -1 0 1330 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1053_
timestamp 0
transform -1 0 1470 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1054_
timestamp 0
transform 1 0 1950 0 1 1690
box -6 -8 86 248
use OAI21X1  _1055_
timestamp 0
transform 1 0 1810 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1056_
timestamp 0
transform -1 0 2390 0 1 2170
box -6 -8 86 248
use INVX1  _1057_
timestamp 0
transform 1 0 2410 0 -1 2170
box -6 -8 66 248
use NAND2X1  _1058_
timestamp 0
transform 1 0 2690 0 1 1690
box -6 -8 86 248
use INVX1  _1059_
timestamp 0
transform 1 0 2870 0 -1 2170
box -6 -8 66 248
use NAND2X1  _1060_
timestamp 0
transform -1 0 3190 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1061_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 86 248
use AOI21X1  _1062_
timestamp 0
transform 1 0 2670 0 1 2170
box -6 -8 106 248
use OAI21X1  _1063_
timestamp 0
transform -1 0 3750 0 -1 3610
box -6 -8 106 248
use OR2X2  _1064_
timestamp 0
transform 1 0 3910 0 1 3610
box -6 -8 106 248
use AOI21X1  _1065_
timestamp 0
transform -1 0 3450 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1066_
timestamp 0
transform 1 0 3490 0 1 3610
box -6 -8 106 248
use NAND3X1  _1067_
timestamp 0
transform 1 0 3770 0 1 3610
box -6 -8 106 248
use INVX1  _1068_
timestamp 0
transform -1 0 3530 0 1 4090
box -6 -8 66 248
use AOI21X1  _1069_
timestamp 0
transform -1 0 3730 0 1 3610
box -6 -8 106 248
use NOR2X1  _1070_
timestamp 0
transform 1 0 3710 0 1 4090
box -6 -8 86 248
use NOR2X1  _1071_
timestamp 0
transform 1 0 3770 0 1 4570
box -6 -8 86 248
use INVX1  _1072_
timestamp 0
transform 1 0 3990 0 -1 4570
box -6 -8 66 248
use OAI21X1  _1073_
timestamp 0
transform 1 0 4090 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1074_
timestamp 0
transform 1 0 3910 0 1 4570
box -6 -8 106 248
use NAND2X1  _1075_
timestamp 0
transform -1 0 4490 0 1 4570
box -6 -8 86 248
use OAI21X1  _1076_
timestamp 0
transform -1 0 3670 0 1 4090
box -6 -8 106 248
use INVX1  _1077_
timestamp 0
transform 1 0 3190 0 1 4090
box -6 -8 66 248
use NAND2X1  _1078_
timestamp 0
transform 1 0 2730 0 1 3610
box -6 -8 86 248
use INVX1  _1079_
timestamp 0
transform 1 0 50 0 -1 730
box -6 -8 66 248
use NAND2X1  _1080_
timestamp 0
transform -1 0 850 0 1 1210
box -6 -8 86 248
use OAI21X1  _1081_
timestamp 0
transform -1 0 990 0 1 1210
box -6 -8 106 248
use NAND2X1  _1082_
timestamp 0
transform 1 0 1390 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1083_
timestamp 0
transform 1 0 950 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1084_
timestamp 0
transform -1 0 2590 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1085_
timestamp 0
transform -1 0 3330 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1086_
timestamp 0
transform 1 0 2630 0 -1 2170
box -6 -8 86 248
use AOI21X1  _1087_
timestamp 0
transform 1 0 2250 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1088_
timestamp 0
transform -1 0 2550 0 1 3610
box -6 -8 106 248
use INVX1  _1089_
timestamp 0
transform -1 0 2170 0 -1 4090
box -6 -8 66 248
use INVX1  _1090_
timestamp 0
transform -1 0 2390 0 1 3610
box -6 -8 66 248
use OAI21X1  _1091_
timestamp 0
transform 1 0 2230 0 -1 4090
box -6 -8 106 248
use AOI21X1  _1092_
timestamp 0
transform 1 0 2530 0 -1 4090
box -6 -8 106 248
use INVX1  _1093_
timestamp 0
transform 1 0 2850 0 1 4090
box -6 -8 66 248
use NAND3X1  _1094_
timestamp 0
transform -1 0 2490 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1095_
timestamp 0
transform 1 0 2950 0 1 4090
box -6 -8 86 248
use OR2X2  _1096_
timestamp 0
transform 1 0 3470 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1097_
timestamp 0
transform -1 0 3290 0 -1 4570
box -6 -8 86 248
use AOI21X1  _1098_
timestamp 0
transform 1 0 3610 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1099_
timestamp 0
transform -1 0 4630 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1100_
timestamp 0
transform -1 0 2810 0 1 4090
box -6 -8 106 248
use NAND3X1  _1101_
timestamp 0
transform -1 0 2690 0 1 3610
box -6 -8 106 248
use NAND2X1  _1102_
timestamp 0
transform -1 0 410 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1103_
timestamp 0
transform -1 0 550 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1104_
timestamp 0
transform -1 0 910 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1105_
timestamp 0
transform -1 0 1210 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1106_
timestamp 0
transform -1 0 1430 0 1 2650
box -6 -8 86 248
use OAI21X1  _1107_
timestamp 0
transform -1 0 1730 0 1 2650
box -6 -8 106 248
use INVX1  _1108_
timestamp 0
transform -1 0 1770 0 -1 3610
box -6 -8 66 248
use NAND3X1  _1109_
timestamp 0
transform 1 0 1770 0 1 3610
box -6 -8 106 248
use INVX1  _1110_
timestamp 0
transform 1 0 1970 0 -1 3610
box -6 -8 66 248
use AOI21X1  _1111_
timestamp 0
transform 1 0 1630 0 1 3610
box -6 -8 106 248
use OAI21X1  _1112_
timestamp 0
transform 1 0 1810 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1113_
timestamp 0
transform -1 0 2290 0 1 3610
box -6 -8 106 248
use NAND2X1  _1114_
timestamp 0
transform 1 0 2050 0 1 3610
box -6 -8 86 248
use NAND3X1  _1115_
timestamp 0
transform 1 0 1910 0 1 3610
box -6 -8 106 248
use AND2X2  _1116_
timestamp 0
transform -1 0 1750 0 -1 4570
box -6 -8 106 248
use INVX1  _1117_
timestamp 0
transform 1 0 1770 0 -1 5050
box -6 -8 66 248
use OR2X2  _1118_
timestamp 0
transform 1 0 2150 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1119_
timestamp 0
transform -1 0 2110 0 -1 5050
box -6 -8 86 248
use NAND2X1  _1120_
timestamp 0
transform 1 0 2290 0 -1 5050
box -6 -8 86 248
use AOI22X1  _1121_
timestamp 0
transform -1 0 2430 0 1 5530
box -6 -8 126 248
use OAI21X1  _1122_
timestamp 0
transform 1 0 1870 0 -1 5050
box -6 -8 106 248
use NOR2X1  _1123_
timestamp 0
transform 1 0 1290 0 -1 4090
box -6 -8 86 248
use INVX1  _1124_
timestamp 0
transform 1 0 1590 0 1 4090
box -6 -8 66 248
use NOR2X1  _1125_
timestamp 0
transform -1 0 990 0 1 2170
box -6 -8 86 248
use INVX1  _1126_
timestamp 0
transform -1 0 470 0 1 1210
box -6 -8 66 248
use NOR2X1  _1127_
timestamp 0
transform -1 0 630 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1128_
timestamp 0
transform 1 0 610 0 1 2170
box -6 -8 106 248
use OAI21X1  _1129_
timestamp 0
transform -1 0 1130 0 1 2170
box -6 -8 106 248
use NAND3X1  _1130_
timestamp 0
transform 1 0 1710 0 1 4090
box -6 -8 106 248
use INVX1  _1131_
timestamp 0
transform 1 0 1410 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1132_
timestamp 0
transform -1 0 1630 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1133_
timestamp 0
transform 1 0 1850 0 1 4090
box -6 -8 106 248
use NAND3X1  _1134_
timestamp 0
transform -1 0 1590 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1135_
timestamp 0
transform 1 0 1430 0 1 4090
box -6 -8 106 248
use NAND3X1  _1136_
timestamp 0
transform 1 0 1350 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1137_
timestamp 0
transform 1 0 1650 0 -1 5050
box -6 -8 86 248
use INVX1  _1138_
timestamp 0
transform 1 0 1690 0 1 5050
box -6 -8 66 248
use AND2X2  _1139_
timestamp 0
transform 1 0 1930 0 1 5050
box -6 -8 106 248
use OAI21X1  _1140_
timestamp 0
transform -1 0 1890 0 1 5050
box -6 -8 106 248
use OAI22X1  _1141_
timestamp 0
transform -1 0 2130 0 -1 5530
box -6 -8 126 248
use NOR3X1  _1142_
timestamp 0
transform -1 0 1250 0 -1 4090
box -6 -8 186 248
use INVX1  _1143_
timestamp 0
transform -1 0 1070 0 1 4090
box -6 -8 66 248
use AOI21X1  _1144_
timestamp 0
transform 1 0 690 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1145_
timestamp 0
transform 1 0 1730 0 1 2170
box -6 -8 86 248
use OAI21X1  _1146_
timestamp 0
transform 1 0 770 0 1 2170
box -6 -8 106 248
use INVX1  _1147_
timestamp 0
transform 1 0 910 0 1 4090
box -6 -8 66 248
use NAND3X1  _1148_
timestamp 0
transform -1 0 1210 0 1 4090
box -6 -8 106 248
use OAI21X1  _1149_
timestamp 0
transform -1 0 1030 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1150_
timestamp 0
transform 1 0 1110 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1151_
timestamp 0
transform -1 0 1310 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1152_
timestamp 0
transform 1 0 870 0 1 4570
box -6 -8 106 248
use AND2X2  _1153_
timestamp 0
transform -1 0 1230 0 1 4570
box -6 -8 106 248
use NAND3X1  _1154_
timestamp 0
transform -1 0 1610 0 -1 5050
box -6 -8 106 248
use INVX1  _1155_
timestamp 0
transform -1 0 1630 0 1 4570
box -6 -8 66 248
use AOI21X1  _1156_
timestamp 0
transform -1 0 1370 0 1 4570
box -6 -8 106 248
use AOI21X1  _1157_
timestamp 0
transform -1 0 1510 0 1 4570
box -6 -8 106 248
use OAI21X1  _1158_
timestamp 0
transform -1 0 1470 0 -1 5050
box -6 -8 106 248
use AND2X2  _1159_
timestamp 0
transform -1 0 1310 0 -1 5050
box -6 -8 106 248
use NOR2X1  _1160_
timestamp 0
transform 1 0 1290 0 1 5050
box -6 -8 86 248
use OAI21X1  _1161_
timestamp 0
transform 1 0 1410 0 1 5050
box -6 -8 106 248
use NAND2X1  _1162_
timestamp 0
transform -1 0 1630 0 1 5050
box -6 -8 86 248
use OAI21X1  _1163_
timestamp 0
transform -1 0 1710 0 -1 5530
box -6 -8 106 248
use AOI21X1  _1164_
timestamp 0
transform -1 0 810 0 1 4570
box -6 -8 106 248
use NOR2X1  _1165_
timestamp 0
transform 1 0 870 0 1 5050
box -6 -8 86 248
use NAND3X1  _1166_
timestamp 0
transform -1 0 1370 0 1 4090
box -6 -8 106 248
use NOR2X1  _1167_
timestamp 0
transform 1 0 310 0 -1 2170
box -6 -8 86 248
use AOI21X1  _1168_
timestamp 0
transform -1 0 430 0 1 2170
box -6 -8 106 248
use NAND3X1  _1169_
timestamp 0
transform 1 0 630 0 1 4090
box -6 -8 106 248
use INVX1  _1170_
timestamp 0
transform -1 0 390 0 1 4570
box -6 -8 66 248
use AOI21X1  _1171_
timestamp 0
transform -1 0 1070 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1172_
timestamp 0
transform 1 0 570 0 1 4570
box -6 -8 106 248
use INVX1  _1173_
timestamp 0
transform 1 0 450 0 -1 4570
box -6 -8 66 248
use NAND2X1  _1174_
timestamp 0
transform -1 0 650 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1175_
timestamp 0
transform 1 0 690 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1176_
timestamp 0
transform -1 0 910 0 -1 4570
box -6 -8 106 248
use AND2X2  _1177_
timestamp 0
transform 1 0 930 0 -1 5050
box -6 -8 106 248
use OR2X2  _1178_
timestamp 0
transform 1 0 990 0 1 5050
box -6 -8 106 248
use AOI21X1  _1179_
timestamp 0
transform 1 0 1130 0 1 5050
box -6 -8 106 248
use AOI22X1  _1180_
timestamp 0
transform -1 0 1210 0 -1 5530
box -6 -8 126 248
use NAND2X1  _1181_
timestamp 0
transform 1 0 670 0 -1 6010
box -6 -8 86 248
use NAND2X1  _1182_
timestamp 0
transform 1 0 790 0 -1 5050
box -6 -8 86 248
use AND2X2  _1183_
timestamp 0
transform -1 0 750 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1184_
timestamp 0
transform -1 0 1170 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1185_
timestamp 0
transform 1 0 370 0 -1 5050
box -6 -8 86 248
use NAND3X1  _1186_
timestamp 0
transform -1 0 870 0 1 4090
box -6 -8 106 248
use INVX1  _1187_
timestamp 0
transform -1 0 910 0 1 2650
box -6 -8 66 248
use INVX1  _1188_
timestamp 0
transform -1 0 130 0 1 2170
box -6 -8 66 248
use OAI21X1  _1189_
timestamp 0
transform -1 0 810 0 1 2650
box -6 -8 106 248
use NAND3X1  _1190_
timestamp 0
transform -1 0 430 0 1 4090
box -6 -8 106 248
use INVX1  _1191_
timestamp 0
transform -1 0 130 0 1 4090
box -6 -8 66 248
use OAI21X1  _1192_
timestamp 0
transform -1 0 410 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1193_
timestamp 0
transform -1 0 130 0 1 4570
box -6 -8 86 248
use NAND3X1  _1194_
timestamp 0
transform -1 0 290 0 1 4570
box -6 -8 106 248
use INVX1  _1195_
timestamp 0
transform -1 0 210 0 -1 4090
box -6 -8 66 248
use NAND3X1  _1196_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 106 248
use NAND2X1  _1197_
timestamp 0
transform -1 0 130 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1198_
timestamp 0
transform -1 0 270 0 -1 4570
box -6 -8 106 248
use AND2X2  _1199_
timestamp 0
transform 1 0 70 0 -1 5050
box -6 -8 106 248
use OR2X2  _1200_
timestamp 0
transform -1 0 290 0 1 5050
box -6 -8 106 248
use INVX1  _1201_
timestamp 0
transform -1 0 110 0 -1 6010
box -6 -8 66 248
use INVX1  _1202_
timestamp 0
transform 1 0 350 0 1 5050
box -6 -8 66 248
use AOI21X1  _1203_
timestamp 0
transform -1 0 550 0 1 5050
box -6 -8 106 248
use INVX1  _1204_
timestamp 0
transform 1 0 390 0 -1 5530
box -6 -8 66 248
use NAND2X1  _1205_
timestamp 0
transform -1 0 250 0 -1 6010
box -6 -8 86 248
use OAI21X1  _1206_
timestamp 0
transform 1 0 290 0 -1 6010
box -6 -8 106 248
use INVX1  _1207_
timestamp 0
transform -1 0 1430 0 -1 5530
box -6 -8 66 248
use INVX1  _1208_
timestamp 0
transform -1 0 130 0 1 5530
box -6 -8 66 248
use OR2X2  _1209_
timestamp 0
transform -1 0 570 0 1 2170
box -6 -8 106 248
use AOI21X1  _1210_
timestamp 0
transform -1 0 290 0 1 2170
box -6 -8 106 248
use OAI21X1  _1211_
timestamp 0
transform 1 0 470 0 1 4090
box -6 -8 106 248
use NAND2X1  _1212_
timestamp 0
transform 1 0 350 0 1 3610
box -6 -8 86 248
use OR2X2  _1213_
timestamp 0
transform 1 0 70 0 1 3610
box -6 -8 106 248
use NAND3X1  _1214_
timestamp 0
transform -1 0 310 0 1 3610
box -6 -8 106 248
use INVX1  _1215_
timestamp 0
transform -1 0 410 0 -1 3130
box -6 -8 66 248
use AND2X2  _1216_
timestamp 0
transform 1 0 210 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1217_
timestamp 0
transform -1 0 130 0 1 3130
box -6 -8 86 248
use OAI21X1  _1218_
timestamp 0
transform 1 0 50 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1219_
timestamp 0
transform -1 0 150 0 1 5050
box -6 -8 86 248
use NOR3X1  _1220_
timestamp 0
transform 1 0 170 0 1 5530
box -6 -8 186 248
use AOI22X1  _1221_
timestamp 0
transform 1 0 230 0 -1 5530
box -6 -8 126 248
use OAI21X1  _1222_
timestamp 0
transform 1 0 390 0 1 5530
box -6 -8 106 248
use OAI21X1  _1223_
timestamp 0
transform -1 0 1230 0 1 5530
box -6 -8 106 248
use OAI21X1  _1224_
timestamp 0
transform -1 0 850 0 -1 2650
box -6 -8 106 248
use OR2X2  _1225_
timestamp 0
transform 1 0 250 0 -1 4090
box -6 -8 106 248
use INVX1  _1226_
timestamp 0
transform -1 0 110 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1227_
timestamp 0
transform 1 0 410 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1228_
timestamp 0
transform 1 0 750 0 1 3610
box -6 -8 86 248
use INVX1  _1229_
timestamp 0
transform -1 0 630 0 1 3130
box -6 -8 66 248
use OAI21X1  _1230_
timestamp 0
transform -1 0 530 0 1 3130
box -6 -8 106 248
use NOR2X1  _1231_
timestamp 0
transform -1 0 650 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1232_
timestamp 0
transform -1 0 790 0 -1 3610
box -6 -8 106 248
use INVX1  _1233_
timestamp 0
transform -1 0 250 0 -1 2650
box -6 -8 66 248
use NOR2X1  _1234_
timestamp 0
transform 1 0 830 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1235_
timestamp 0
transform 1 0 630 0 1 3610
box -6 -8 86 248
use OAI21X1  _1236_
timestamp 0
transform -1 0 570 0 1 3610
box -6 -8 106 248
use AND2X2  _1237_
timestamp 0
transform -1 0 530 0 1 4570
box -6 -8 106 248
use OAI21X1  _1238_
timestamp 0
transform -1 0 170 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1239_
timestamp 0
transform 1 0 210 0 -1 5050
box -6 -8 106 248
use AOI21X1  _1240_
timestamp 0
transform 1 0 490 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1241_
timestamp 0
transform -1 0 610 0 -1 5530
box -6 -8 106 248
use INVX1  _1242_
timestamp 0
transform 1 0 530 0 1 5530
box -6 -8 66 248
use NOR2X1  _1243_
timestamp 0
transform 1 0 650 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1244_
timestamp 0
transform 1 0 650 0 1 5530
box -6 -8 86 248
use NAND2X1  _1245_
timestamp 0
transform -1 0 850 0 1 5530
box -6 -8 86 248
use AOI22X1  _1246_
timestamp 0
transform -1 0 1630 0 1 5530
box -6 -8 126 248
use INVX1  _1247_
timestamp 0
transform 1 0 310 0 1 1690
box -6 -8 66 248
use NAND2X1  _1248_
timestamp 0
transform -1 0 270 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1249_
timestamp 0
transform -1 0 150 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1250_
timestamp 0
transform -1 0 270 0 -1 2170
box -6 -8 86 248
use INVX1  _1251_
timestamp 0
transform 1 0 430 0 -1 2170
box -6 -8 66 248
use OAI21X1  _1252_
timestamp 0
transform -1 0 1070 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1253_
timestamp 0
transform -1 0 750 0 1 3130
box -6 -8 86 248
use OAI21X1  _1254_
timestamp 0
transform 1 0 790 0 1 3130
box -6 -8 106 248
use NAND2X1  _1255_
timestamp 0
transform -1 0 970 0 1 3610
box -6 -8 86 248
use AOI21X1  _1256_
timestamp 0
transform 1 0 590 0 1 5050
box -6 -8 106 248
use NAND3X1  _1257_
timestamp 0
transform 1 0 730 0 1 5050
box -6 -8 106 248
use NAND2X1  _1258_
timestamp 0
transform -1 0 870 0 -1 5530
box -6 -8 86 248
use OAI22X1  _1259_
timestamp 0
transform -1 0 1030 0 -1 5530
box -6 -8 126 248
use INVX1  _1260_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 66 248
use INVX1  _1261_
timestamp 0
transform 1 0 4290 0 1 2650
box -6 -8 66 248
use NAND2X1  _1262_
timestamp 0
transform -1 0 2550 0 1 3130
box -6 -8 86 248
use OAI21X1  _1263_
timestamp 0
transform -1 0 3790 0 1 3130
box -6 -8 106 248
use NOR2X1  _1264_
timestamp 0
transform 1 0 4930 0 -1 4090
box -6 -8 86 248
use AND2X2  _1265_
timestamp 0
transform 1 0 4630 0 1 4090
box -6 -8 106 248
use OR2X2  _1266_
timestamp 0
transform 1 0 4790 0 1 4090
box -6 -8 106 248
use NAND2X1  _1267_
timestamp 0
transform 1 0 5310 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1268_
timestamp 0
transform 1 0 5170 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1269_
timestamp 0
transform 1 0 5590 0 -1 4570
box -6 -8 86 248
use INVX2  _1270_
timestamp 0
transform -1 0 2170 0 1 3130
box -6 -8 66 248
use OAI21X1  _1271_
timestamp 0
transform -1 0 3710 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1272_
timestamp 0
transform -1 0 3350 0 1 3130
box -6 -8 106 248
use OAI21X1  _1273_
timestamp 0
transform -1 0 3970 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1274_
timestamp 0
transform 1 0 4030 0 -1 4090
box -6 -8 106 248
use OR2X2  _1275_
timestamp 0
transform 1 0 5470 0 1 4090
box -6 -8 106 248
use NAND2X1  _1276_
timestamp 0
transform -1 0 5430 0 1 4090
box -6 -8 86 248
use NAND2X1  _1277_
timestamp 0
transform 1 0 5630 0 1 4090
box -6 -8 86 248
use NOR2X1  _1278_
timestamp 0
transform -1 0 5830 0 1 4090
box -6 -8 86 248
use NAND2X1  _1279_
timestamp 0
transform 1 0 5790 0 -1 730
box -6 -8 86 248
use NAND2X1  _1280_
timestamp 0
transform 1 0 5830 0 -1 250
box -6 -8 86 248
use OAI21X1  _1281_
timestamp 0
transform -1 0 5810 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1282_
timestamp 0
transform -1 0 5350 0 -1 4090
box -6 -8 86 248
use INVX1  _1283_
timestamp 0
transform 1 0 5850 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1284_
timestamp 0
transform 1 0 5770 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1285_
timestamp 0
transform -1 0 4150 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1286_
timestamp 0
transform 1 0 4630 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1287_
timestamp 0
transform -1 0 4870 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1288_
timestamp 0
transform 1 0 5630 0 1 3130
box -6 -8 86 248
use OR2X2  _1289_
timestamp 0
transform 1 0 5550 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1290_
timestamp 0
transform 1 0 5750 0 1 3130
box -6 -8 86 248
use INVX1  _1291_
timestamp 0
transform -1 0 5590 0 -1 6010
box -6 -8 66 248
use NOR2X1  _1292_
timestamp 0
transform 1 0 5850 0 1 4570
box -6 -8 86 248
use NAND2X1  _1293_
timestamp 0
transform 1 0 5630 0 -1 6010
box -6 -8 86 248
use NAND2X1  _1294_
timestamp 0
transform 1 0 5770 0 1 3610
box -6 -8 86 248
use OAI21X1  _1295_
timestamp 0
transform -1 0 5730 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1296_
timestamp 0
transform 1 0 5630 0 1 3610
box -6 -8 86 248
use INVX1  _1297_
timestamp 0
transform 1 0 5530 0 1 3610
box -6 -8 66 248
use INVX1  _1298_
timestamp 0
transform 1 0 4850 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1299_
timestamp 0
transform -1 0 3970 0 1 2650
box -6 -8 106 248
use NAND2X1  _1300_
timestamp 0
transform -1 0 3990 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1301_
timestamp 0
transform -1 0 4430 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1302_
timestamp 0
transform 1 0 4490 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1303_
timestamp 0
transform 1 0 5070 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1304_
timestamp 0
transform -1 0 5030 0 -1 3610
box -6 -8 86 248
use INVX1  _1305_
timestamp 0
transform 1 0 5010 0 1 3610
box -6 -8 66 248
use OAI21X1  _1306_
timestamp 0
transform 1 0 5110 0 1 3610
box -6 -8 106 248
use INVX1  _1307_
timestamp 0
transform 1 0 5250 0 1 3610
box -6 -8 66 248
use NAND3X1  _1308_
timestamp 0
transform 1 0 5370 0 1 3610
box -6 -8 106 248
use NAND2X1  _1309_
timestamp 0
transform -1 0 5230 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1310_
timestamp 0
transform -1 0 5010 0 1 4570
box -6 -8 86 248
use OAI21X1  _1311_
timestamp 0
transform -1 0 5170 0 1 4570
box -6 -8 106 248
use NAND2X1  _1312_
timestamp 0
transform 1 0 4270 0 -1 5050
box -6 -8 86 248
use NOR2X1  _1313_
timestamp 0
transform 1 0 3210 0 -1 4090
box -6 -8 86 248
use NAND3X1  _1314_
timestamp 0
transform 1 0 3210 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1315_
timestamp 0
transform -1 0 3190 0 1 3130
box -6 -8 106 248
use NOR2X1  _1316_
timestamp 0
transform 1 0 3090 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1317_
timestamp 0
transform 1 0 2670 0 -1 4570
box -6 -8 86 248
use INVX1  _1318_
timestamp 0
transform 1 0 2570 0 -1 4570
box -6 -8 66 248
use OAI21X1  _1319_
timestamp 0
transform -1 0 3030 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1320_
timestamp 0
transform -1 0 4950 0 1 3610
box -6 -8 106 248
use AOI21X1  _1321_
timestamp 0
transform 1 0 2830 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1322_
timestamp 0
transform -1 0 2790 0 -1 5050
box -6 -8 86 248
use INVX1  _1323_
timestamp 0
transform 1 0 2970 0 -1 5050
box -6 -8 66 248
use OAI21X1  _1324_
timestamp 0
transform -1 0 2650 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1325_
timestamp 0
transform 1 0 3350 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1326_
timestamp 0
transform 1 0 3030 0 -1 6010
box -6 -8 86 248
use OAI21X1  _1327_
timestamp 0
transform -1 0 2690 0 1 5050
box -6 -8 106 248
use OAI21X1  _1328_
timestamp 0
transform -1 0 3550 0 1 2650
box -6 -8 106 248
use INVX1  _1329_
timestamp 0
transform -1 0 3410 0 1 2650
box -6 -8 66 248
use OAI21X1  _1330_
timestamp 0
transform 1 0 2570 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1331_
timestamp 0
transform 1 0 2590 0 1 4090
box -6 -8 86 248
use NOR2X1  _1332_
timestamp 0
transform -1 0 2390 0 -1 4570
box -6 -8 86 248
use AND2X2  _1333_
timestamp 0
transform -1 0 2130 0 1 4570
box -6 -8 106 248
use INVX1  _1334_
timestamp 0
transform 1 0 2170 0 1 4570
box -6 -8 66 248
use INVX1  _1335_
timestamp 0
transform -1 0 1970 0 1 4570
box -6 -8 66 248
use OAI21X1  _1336_
timestamp 0
transform -1 0 2390 0 1 4570
box -6 -8 106 248
use NAND2X1  _1337_
timestamp 0
transform 1 0 2430 0 1 4570
box -6 -8 86 248
use INVX1  _1338_
timestamp 0
transform 1 0 2470 0 1 5050
box -6 -8 66 248
use NOR2X1  _1339_
timestamp 0
transform 1 0 2530 0 -1 6010
box -6 -8 86 248
use NAND2X1  _1340_
timestamp 0
transform 1 0 2470 0 1 5530
box -6 -8 86 248
use NAND2X1  _1341_
timestamp 0
transform -1 0 2490 0 -1 6010
box -6 -8 86 248
use OAI21X1  _1342_
timestamp 0
transform 1 0 2650 0 -1 6010
box -6 -8 106 248
use NOR2X1  _1343_
timestamp 0
transform 1 0 2730 0 1 5050
box -6 -8 86 248
use OAI21X1  _1344_
timestamp 0
transform 1 0 2570 0 1 4570
box -6 -8 106 248
use AOI21X1  _1345_
timestamp 0
transform 1 0 3210 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1346_
timestamp 0
transform -1 0 3490 0 1 3130
box -6 -8 106 248
use NOR2X1  _1347_
timestamp 0
transform 1 0 3610 0 -1 4090
box -6 -8 86 248
use AND2X2  _1348_
timestamp 0
transform 1 0 3730 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1349_
timestamp 0
transform 1 0 3470 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1350_
timestamp 0
transform 1 0 3330 0 -1 4090
box -6 -8 86 248
use INVX1  _1351_
timestamp 0
transform -1 0 3130 0 1 4090
box -6 -8 66 248
use OAI21X1  _1352_
timestamp 0
transform -1 0 3410 0 1 4090
box -6 -8 106 248
use NAND2X1  _1353_
timestamp 0
transform 1 0 3330 0 -1 4570
box -6 -8 86 248
use AND2X2  _1354_
timestamp 0
transform 1 0 4510 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1355_
timestamp 0
transform 1 0 4670 0 -1 5050
box -6 -8 106 248
use OAI22X1  _1356_
timestamp 0
transform -1 0 5050 0 -1 5050
box -6 -8 126 248
use OAI21X1  _1357_
timestamp 0
transform -1 0 3350 0 1 4570
box -6 -8 106 248
use NAND3X1  _1358_
timestamp 0
transform 1 0 3770 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1359_
timestamp 0
transform 1 0 4390 0 1 2650
box -6 -8 106 248
use NAND2X1  _1360_
timestamp 0
transform -1 0 4610 0 1 2650
box -6 -8 86 248
use INVX1  _1361_
timestamp 0
transform 1 0 4250 0 -1 4570
box -6 -8 66 248
use NAND2X1  _1362_
timestamp 0
transform 1 0 3870 0 -1 4570
box -6 -8 86 248
use INVX1  _1363_
timestamp 0
transform -1 0 3070 0 1 4570
box -6 -8 66 248
use NOR2X1  _1364_
timestamp 0
transform -1 0 3830 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1365_
timestamp 0
transform -1 0 3470 0 1 4570
box -6 -8 86 248
use INVX1  _1366_
timestamp 0
transform -1 0 3470 0 1 5050
box -6 -8 66 248
use OR2X2  _1367_
timestamp 0
transform 1 0 3310 0 1 5530
box -6 -8 106 248
use AOI21X1  _1368_
timestamp 0
transform -1 0 3270 0 1 5530
box -6 -8 106 248
use AOI22X1  _1369_
timestamp 0
transform -1 0 3590 0 1 5530
box -6 -8 126 248
use NAND2X1  _1370_
timestamp 0
transform 1 0 4770 0 -1 6010
box -6 -8 86 248
use NAND2X1  _1371_
timestamp 0
transform 1 0 4170 0 1 2650
box -6 -8 86 248
use NAND2X1  _1372_
timestamp 0
transform -1 0 4290 0 -1 3130
box -6 -8 86 248
use INVX1  _1373_
timestamp 0
transform -1 0 4030 0 1 5050
box -6 -8 66 248
use NAND2X1  _1374_
timestamp 0
transform 1 0 3850 0 1 5050
box -6 -8 86 248
use INVX1  _1375_
timestamp 0
transform 1 0 4090 0 1 5050
box -6 -8 66 248
use NAND2X1  _1376_
timestamp 0
transform 1 0 4190 0 1 5050
box -6 -8 86 248
use NAND2X1  _1377_
timestamp 0
transform -1 0 4010 0 1 5530
box -6 -8 86 248
use INVX1  _1378_
timestamp 0
transform -1 0 3810 0 -1 6010
box -6 -8 66 248
use OAI21X1  _1379_
timestamp 0
transform -1 0 3210 0 1 4570
box -6 -8 106 248
use OR2X2  _1380_
timestamp 0
transform -1 0 3350 0 1 5050
box -6 -8 106 248
use INVX1  _1381_
timestamp 0
transform -1 0 3190 0 1 5050
box -6 -8 66 248
use AOI21X1  _1382_
timestamp 0
transform -1 0 3170 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1383_
timestamp 0
transform -1 0 2950 0 1 5050
box -6 -8 86 248
use OAI21X1  _1384_
timestamp 0
transform 1 0 2990 0 1 5050
box -6 -8 106 248
use NOR2X1  _1385_
timestamp 0
transform 1 0 3850 0 -1 6010
box -6 -8 86 248
use INVX1  _1386_
timestamp 0
transform 1 0 3990 0 -1 6010
box -6 -8 66 248
use OAI21X1  _1387_
timestamp 0
transform 1 0 4090 0 -1 6010
box -6 -8 106 248
use OAI21X1  _1388_
timestamp 0
transform 1 0 4250 0 -1 6010
box -6 -8 106 248
use NAND2X1  _1389_
timestamp 0
transform -1 0 4830 0 1 5530
box -6 -8 86 248
use INVX1  _1390_
timestamp 0
transform 1 0 3490 0 -1 6010
box -6 -8 66 248
use AOI21X1  _1391_
timestamp 0
transform -1 0 3710 0 -1 6010
box -6 -8 106 248
use INVX1  _1392_
timestamp 0
transform -1 0 2970 0 -1 5530
box -6 -8 66 248
use NAND2X1  _1393_
timestamp 0
transform -1 0 3230 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1394_
timestamp 0
transform -1 0 3110 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1395_
timestamp 0
transform 1 0 3270 0 -1 5530
box -6 -8 86 248
use AND2X2  _1396_
timestamp 0
transform 1 0 4310 0 1 5530
box -6 -8 106 248
use OAI21X1  _1397_
timestamp 0
transform 1 0 4470 0 1 5530
box -6 -8 106 248
use OAI21X1  _1398_
timestamp 0
transform 1 0 4610 0 1 5530
box -6 -8 106 248
use OAI21X1  _1399_
timestamp 0
transform -1 0 3490 0 -1 5530
box -6 -8 106 248
use OR2X2  _1400_
timestamp 0
transform 1 0 4170 0 1 5530
box -6 -8 106 248
use INVX1  _1401_
timestamp 0
transform -1 0 4110 0 1 5530
box -6 -8 66 248
use AOI21X1  _1402_
timestamp 0
transform 1 0 3930 0 -1 5530
box -6 -8 106 248
use INVX1  _1403_
timestamp 0
transform -1 0 3570 0 1 5050
box -6 -8 66 248
use NAND2X1  _1404_
timestamp 0
transform -1 0 3750 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1405_
timestamp 0
transform -1 0 3630 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1406_
timestamp 0
transform -1 0 3870 0 -1 5530
box -6 -8 86 248
use AND2X2  _1407_
timestamp 0
transform 1 0 4230 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1408_
timestamp 0
transform 1 0 4390 0 -1 5530
box -6 -8 106 248
use OAI22X1  _1409_
timestamp 0
transform -1 0 4570 0 1 5050
box -6 -8 126 248
use NAND2X1  _1410_
timestamp 0
transform -1 0 4910 0 -1 5530
box -6 -8 86 248
use OAI21X1  _1411_
timestamp 0
transform -1 0 4190 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1412_
timestamp 0
transform 1 0 4690 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1413_
timestamp 0
transform -1 0 4990 0 1 2170
box -6 -8 106 248
use NOR2X1  _1414_
timestamp 0
transform 1 0 4750 0 1 2170
box -6 -8 86 248
use NAND2X1  _1415_
timestamp 0
transform 1 0 850 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1416_
timestamp 0
transform 1 0 710 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1417_
timestamp 0
transform -1 0 130 0 1 1210
box -6 -8 86 248
use OAI21X1  _1418_
timestamp 0
transform -1 0 150 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1419_
timestamp 0
transform 1 0 5450 0 -1 1690
box -6 -8 86 248
use AND2X2  _1420_
timestamp 0
transform -1 0 5390 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1421_
timestamp 0
transform -1 0 530 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1422_
timestamp 0
transform 1 0 310 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1423_
timestamp 0
transform -1 0 130 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1424_
timestamp 0
transform -1 0 150 0 1 2650
box -6 -8 106 248
use NOR2X1  _1425_
timestamp 0
transform 1 0 4930 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1426_
timestamp 0
transform 1 0 1530 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1427_
timestamp 0
transform 1 0 1390 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1428_
timestamp 0
transform -1 0 1430 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1429_
timestamp 0
transform 1 0 1210 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1430_
timestamp 0
transform 1 0 4010 0 1 2170
box -6 -8 86 248
use NAND2X1  _1431_
timestamp 0
transform -1 0 2290 0 1 3130
box -6 -8 86 248
use OAI21X1  _1432_
timestamp 0
transform 1 0 2270 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1433_
timestamp 0
transform -1 0 1930 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1434_
timestamp 0
transform -1 0 2070 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1435_
timestamp 0
transform -1 0 2790 0 1 3130
box -6 -8 86 248
use OAI21X1  _1436_
timestamp 0
transform -1 0 2950 0 1 3130
box -6 -8 106 248
use NAND2X1  _1437_
timestamp 0
transform 1 0 2850 0 1 3610
box -6 -8 86 248
use OAI21X1  _1438_
timestamp 0
transform 1 0 2730 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1439_
timestamp 0
transform -1 0 4730 0 1 2650
box -6 -8 86 248
use OAI21X1  _1440_
timestamp 0
transform 1 0 4770 0 1 2650
box -6 -8 106 248
use NAND2X1  _1441_
timestamp 0
transform -1 0 4430 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1442_
timestamp 0
transform -1 0 4570 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1443_
timestamp 0
transform -1 0 290 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1444_
timestamp 0
transform 1 0 70 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1445_
timestamp 0
transform -1 0 550 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1446_
timestamp 0
transform 1 0 330 0 -1 1210
box -6 -8 106 248
use INVX1  _1447_
timestamp 0
transform 1 0 1230 0 1 730
box -6 -8 66 248
use NAND2X1  _1448_
timestamp 0
transform 1 0 1090 0 1 730
box -6 -8 86 248
use OAI21X1  _1449_
timestamp 0
transform -1 0 1190 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1450_
timestamp 0
transform 1 0 970 0 1 730
box -6 -8 86 248
use OAI21X1  _1451_
timestamp 0
transform 1 0 810 0 1 730
box -6 -8 106 248
use NAND2X1  _1452_
timestamp 0
transform -1 0 2090 0 1 1210
box -6 -8 86 248
use OAI21X1  _1453_
timestamp 0
transform -1 0 2230 0 1 1210
box -6 -8 106 248
use NAND2X1  _1454_
timestamp 0
transform 1 0 2950 0 1 1210
box -6 -8 86 248
use OAI21X1  _1455_
timestamp 0
transform 1 0 2810 0 1 1210
box -6 -8 106 248
use NAND2X1  _1456_
timestamp 0
transform -1 0 3490 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1457_
timestamp 0
transform 1 0 3350 0 1 1210
box -6 -8 106 248
use NAND2X1  _1458_
timestamp 0
transform 1 0 4010 0 1 1210
box -6 -8 86 248
use OAI21X1  _1459_
timestamp 0
transform 1 0 3850 0 1 1210
box -6 -8 106 248
use NAND2X1  _1460_
timestamp 0
transform 1 0 4630 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1461_
timestamp 0
transform 1 0 4350 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1462_
timestamp 0
transform 1 0 4630 0 1 1210
box -6 -8 86 248
use OAI21X1  _1463_
timestamp 0
transform 1 0 4490 0 1 1210
box -6 -8 106 248
use NAND2X1  _1464_
timestamp 0
transform 1 0 4510 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1465_
timestamp 0
transform 1 0 4450 0 1 1690
box -6 -8 106 248
use NAND2X1  _1466_
timestamp 0
transform -1 0 4350 0 1 1210
box -6 -8 86 248
use OAI21X1  _1467_
timestamp 0
transform -1 0 4310 0 1 1690
box -6 -8 106 248
use NAND2X1  _1468_
timestamp 0
transform -1 0 2790 0 1 4570
box -6 -8 86 248
use OAI21X1  _1469_
timestamp 0
transform -1 0 3610 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1470_
timestamp 0
transform -1 0 1450 0 1 3610
box -6 -8 86 248
use OAI21X1  _1471_
timestamp 0
transform -1 0 1590 0 1 3610
box -6 -8 106 248
use NAND2X1  _1472_
timestamp 0
transform -1 0 3610 0 1 4570
box -6 -8 86 248
use OAI21X1  _1473_
timestamp 0
transform -1 0 4230 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1474_
timestamp 0
transform -1 0 2870 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1475_
timestamp 0
transform -1 0 2950 0 1 4570
box -6 -8 106 248
use NAND2X1  _1476_
timestamp 0
transform -1 0 2750 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1477_
timestamp 0
transform -1 0 2910 0 -1 4090
box -6 -8 106 248
use INVX1  _1478_
timestamp 0
transform -1 0 4630 0 1 3130
box -6 -8 66 248
use NOR2X1  _1479_
timestamp 0
transform -1 0 4030 0 1 3130
box -6 -8 86 248
use AOI21X1  _1480_
timestamp 0
transform -1 0 4530 0 1 3130
box -6 -8 106 248
use NAND2X1  _1481_
timestamp 0
transform 1 0 2470 0 1 4090
box -6 -8 86 248
use OAI21X1  _1482_
timestamp 0
transform -1 0 2530 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1483_
timestamp 0
transform 1 0 1950 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1484_
timestamp 0
transform -1 0 1890 0 -1 4570
box -6 -8 106 248
use INVX1  _1485_
timestamp 0
transform 1 0 5050 0 -1 4090
box -6 -8 66 248
use INVX1  _1486_
timestamp 0
transform 1 0 4830 0 1 3130
box -6 -8 66 248
use OAI21X1  _1487_
timestamp 0
transform 1 0 5230 0 1 3130
box -6 -8 106 248
use OAI21X1  _1488_
timestamp 0
transform 1 0 5090 0 1 3130
box -6 -8 106 248
use OAI21X1  _1489_
timestamp 0
transform -1 0 5050 0 1 3130
box -6 -8 106 248
use OAI21X1  _1490_
timestamp 0
transform 1 0 4670 0 1 3130
box -6 -8 106 248
use NAND2X1  _1491_
timestamp 0
transform -1 0 4450 0 1 4090
box -6 -8 86 248
use OAI21X1  _1492_
timestamp 0
transform -1 0 4590 0 1 4090
box -6 -8 106 248
use NAND2X1  _1493_
timestamp 0
transform -1 0 5390 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1494_
timestamp 0
transform -1 0 5550 0 -1 3610
box -6 -8 106 248
use INVX1  _1495_
timestamp 0
transform 1 0 2170 0 -1 6010
box -6 -8 66 248
use NAND2X1  _1496_
timestamp 0
transform -1 0 870 0 -1 6010
box -6 -8 86 248
use OAI21X1  _1497_
timestamp 0
transform -1 0 1890 0 -1 6010
box -6 -8 106 248
use NAND2X1  _1498_
timestamp 0
transform -1 0 5110 0 1 2170
box -6 -8 86 248
use AOI21X1  _1499_
timestamp 0
transform 1 0 4550 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1500_
timestamp 0
transform -1 0 3090 0 -1 1690
box -6 -8 86 248
use MUX2X1  _1501_
timestamp 0
transform -1 0 690 0 -1 2650
box -6 -8 126 248
use MUX2X1  _1502_
timestamp 0
transform -1 0 1270 0 1 1690
box -6 -8 126 248
use OAI22X1  _1503_
timestamp 0
transform -1 0 2270 0 1 2170
box -6 -8 126 248
use AOI21X1  _1504_
timestamp 0
transform -1 0 2170 0 1 1690
box -6 -8 106 248
use NAND3X1  _1505_
timestamp 0
transform 1 0 3150 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1506_
timestamp 0
transform 1 0 2810 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1507_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 86 248
use NAND3X1  _1508_
timestamp 0
transform 1 0 2670 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1509_
timestamp 0
transform 1 0 2770 0 1 2650
box -6 -8 86 248
use NAND3X1  _1510_
timestamp 0
transform 1 0 2510 0 1 2650
box -6 -8 106 248
use NAND2X1  _1511_
timestamp 0
transform -1 0 2050 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1512_
timestamp 0
transform -1 0 2150 0 -1 3610
box -6 -8 86 248
use NAND3X1  _1513_
timestamp 0
transform -1 0 2010 0 1 2650
box -6 -8 106 248
use NAND2X1  _1514_
timestamp 0
transform -1 0 1570 0 1 2650
box -6 -8 86 248
use NAND3X1  _1515_
timestamp 0
transform 1 0 1770 0 1 2650
box -6 -8 106 248
use NAND2X1  _1516_
timestamp 0
transform 1 0 2390 0 1 2650
box -6 -8 86 248
use NAND2X1  _1517_
timestamp 0
transform 1 0 2650 0 1 2650
box -6 -8 86 248
use NAND3X1  _1518_
timestamp 0
transform -1 0 2330 0 1 2650
box -6 -8 106 248
use NAND2X1  _1519_
timestamp 0
transform 1 0 1970 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1520_
timestamp 0
transform 1 0 1670 0 -1 2650
box -6 -8 86 248
use NAND3X1  _1521_
timestamp 0
transform -1 0 2190 0 -1 2650
box -6 -8 106 248
use AOI22X1  _1522_
timestamp 0
transform 1 0 2070 0 1 2650
box -6 -8 126 248
use INVX1  _1523_
timestamp 0
transform 1 0 3210 0 1 1690
box -6 -8 66 248
use OAI21X1  _1524_
timestamp 0
transform -1 0 3410 0 1 1690
box -6 -8 106 248
use AOI21X1  _1525_
timestamp 0
transform 1 0 3850 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1526_
timestamp 0
transform -1 0 3790 0 -1 1690
box -6 -8 106 248
use INVX1  _1527_
timestamp 0
transform 1 0 4890 0 -1 1690
box -6 -8 66 248
use OR2X2  _1528_
timestamp 0
transform 1 0 5010 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1529_
timestamp 0
transform -1 0 5170 0 -1 2170
box -6 -8 86 248
use INVX1  _1530_
timestamp 0
transform 1 0 5370 0 -1 2170
box -6 -8 66 248
use OAI21X1  _1531_
timestamp 0
transform 1 0 5150 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1532_
timestamp 0
transform -1 0 5310 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1533_
timestamp 0
transform 1 0 3850 0 1 2170
box -6 -8 106 248
use OAI21X1  _1534_
timestamp 0
transform -1 0 5250 0 1 2170
box -6 -8 106 248
use INVX1  _1535_
timestamp 0
transform -1 0 5750 0 -1 730
box -6 -8 66 248
use INVX2  _1536_
timestamp 0
transform 1 0 5150 0 1 1690
box -6 -8 66 248
use OAI21X1  _1537_
timestamp 0
transform 1 0 4750 0 -1 1690
box -6 -8 106 248
use INVX1  _1538_
timestamp 0
transform 1 0 4830 0 -1 250
box -6 -8 66 248
use NAND3X1  _1539_
timestamp 0
transform -1 0 2950 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1540_
timestamp 0
transform 1 0 590 0 1 2650
box -6 -8 86 248
use OAI21X1  _1541_
timestamp 0
transform 1 0 450 0 1 2650
box -6 -8 106 248
use NAND2X1  _1542_
timestamp 0
transform -1 0 1590 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1543_
timestamp 0
transform -1 0 1670 0 1 1690
box -6 -8 106 248
use OAI22X1  _1544_
timestamp 0
transform -1 0 2110 0 1 2170
box -6 -8 126 248
use INVX1  _1545_
timestamp 0
transform -1 0 1830 0 -1 1690
box -6 -8 66 248
use OAI21X1  _1546_
timestamp 0
transform 1 0 1630 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1547_
timestamp 0
transform 1 0 2550 0 -1 1690
box -6 -8 106 248
use INVX1  _1548_
timestamp 0
transform -1 0 2370 0 -1 1690
box -6 -8 66 248
use NAND2X1  _1549_
timestamp 0
transform -1 0 370 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1550_
timestamp 0
transform -1 0 530 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1551_
timestamp 0
transform 1 0 1370 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1552_
timestamp 0
transform 1 0 1230 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1553_
timestamp 0
transform 1 0 1890 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1554_
timestamp 0
transform -1 0 2270 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1555_
timestamp 0
transform 1 0 2710 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1556_
timestamp 0
transform 1 0 5010 0 1 250
box -6 -8 86 248
use NOR2X1  _1557_
timestamp 0
transform 1 0 5130 0 1 250
box -6 -8 86 248
use INVX1  _1558_
timestamp 0
transform 1 0 5270 0 1 250
box -6 -8 66 248
use NAND2X1  _1559_
timestamp 0
transform 1 0 5370 0 1 250
box -6 -8 86 248
use AOI21X1  _1560_
timestamp 0
transform 1 0 5490 0 1 250
box -6 -8 106 248
use OAI21X1  _1561_
timestamp 0
transform 1 0 5650 0 1 250
box -6 -8 106 248
use AOI22X1  _1562_
timestamp 0
transform -1 0 5650 0 -1 730
box -6 -8 126 248
use NAND3X1  _1563_
timestamp 0
transform -1 0 2130 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1564_
timestamp 0
transform -1 0 510 0 1 1690
box -6 -8 86 248
use OAI21X1  _1565_
timestamp 0
transform -1 0 650 0 1 1690
box -6 -8 106 248
use NAND2X1  _1566_
timestamp 0
transform -1 0 810 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1567_
timestamp 0
transform -1 0 950 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1568_
timestamp 0
transform -1 0 1070 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1569_
timestamp 0
transform -1 0 1590 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1570_
timestamp 0
transform 1 0 2990 0 -1 1210
box -6 -8 106 248
use NOR2X1  _1571_
timestamp 0
transform -1 0 2490 0 -1 1690
box -6 -8 86 248
use INVX1  _1572_
timestamp 0
transform -1 0 3070 0 1 730
box -6 -8 66 248
use OAI21X1  _1573_
timestamp 0
transform 1 0 2850 0 1 730
box -6 -8 106 248
use NAND3X1  _1574_
timestamp 0
transform 1 0 3390 0 1 730
box -6 -8 106 248
use INVX1  _1575_
timestamp 0
transform -1 0 3610 0 1 730
box -6 -8 66 248
use AOI21X1  _1576_
timestamp 0
transform 1 0 3250 0 1 730
box -6 -8 106 248
use OAI21X1  _1577_
timestamp 0
transform 1 0 3650 0 1 730
box -6 -8 106 248
use NAND2X1  _1578_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 86 248
use OAI21X1  _1579_
timestamp 0
transform -1 0 4910 0 -1 730
box -6 -8 106 248
use AND2X2  _1580_
timestamp 0
transform 1 0 4870 0 1 250
box -6 -8 106 248
use AOI21X1  _1581_
timestamp 0
transform 1 0 4430 0 1 250
box -6 -8 106 248
use OAI21X1  _1582_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 106 248
use AOI22X1  _1583_
timestamp 0
transform -1 0 4770 0 -1 1210
box -6 -8 126 248
use AOI21X1  _1584_
timestamp 0
transform -1 0 4810 0 1 250
box -6 -8 106 248
use INVX1  _1585_
timestamp 0
transform 1 0 4710 0 -1 730
box -6 -8 66 248
use NOR2X1  _1586_
timestamp 0
transform -1 0 790 0 1 1690
box -6 -8 86 248
use AOI21X1  _1587_
timestamp 0
transform 1 0 990 0 1 1690
box -6 -8 106 248
use NAND2X1  _1588_
timestamp 0
transform 1 0 1730 0 1 1210
box -6 -8 86 248
use OAI21X1  _1589_
timestamp 0
transform 1 0 1590 0 1 1210
box -6 -8 106 248
use INVX1  _1590_
timestamp 0
transform 1 0 2150 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1591_
timestamp 0
transform -1 0 3210 0 1 730
box -6 -8 106 248
use NOR2X1  _1592_
timestamp 0
transform 1 0 2990 0 -1 730
box -6 -8 86 248
use INVX1  _1593_
timestamp 0
transform 1 0 3790 0 1 730
box -6 -8 66 248
use NAND2X1  _1594_
timestamp 0
transform 1 0 3130 0 -1 730
box -6 -8 86 248
use NAND3X1  _1595_
timestamp 0
transform 1 0 3750 0 -1 730
box -6 -8 106 248
use INVX1  _1596_
timestamp 0
transform -1 0 3470 0 -1 730
box -6 -8 66 248
use OAI21X1  _1597_
timestamp 0
transform -1 0 3370 0 -1 730
box -6 -8 106 248
use AND2X2  _1598_
timestamp 0
transform 1 0 4450 0 1 730
box -6 -8 106 248
use AOI21X1  _1599_
timestamp 0
transform 1 0 4750 0 1 730
box -6 -8 106 248
use NAND3X1  _1600_
timestamp 0
transform 1 0 4610 0 1 730
box -6 -8 106 248
use OAI21X1  _1601_
timestamp 0
transform 1 0 4890 0 1 730
box -6 -8 106 248
use OAI21X1  _1602_
timestamp 0
transform 1 0 5030 0 1 730
box -6 -8 106 248
use OAI21X1  _1603_
timestamp 0
transform -1 0 5550 0 1 730
box -6 -8 106 248
use NAND3X1  _1604_
timestamp 0
transform -1 0 2810 0 1 730
box -6 -8 106 248
use AOI21X1  _1605_
timestamp 0
transform 1 0 850 0 1 1690
box -6 -8 106 248
use NAND2X1  _1606_
timestamp 0
transform -1 0 1430 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1607_
timestamp 0
transform 1 0 1430 0 1 1210
box -6 -8 106 248
use NAND3X1  _1608_
timestamp 0
transform 1 0 2590 0 -1 730
box -6 -8 106 248
use NOR3X1  _1609_
timestamp 0
transform 1 0 1930 0 -1 1210
box -6 -8 186 248
use INVX1  _1610_
timestamp 0
transform 1 0 2170 0 1 730
box -6 -8 66 248
use OAI21X1  _1611_
timestamp 0
transform 1 0 2290 0 -1 730
box -6 -8 106 248
use NAND3X1  _1612_
timestamp 0
transform 1 0 2730 0 -1 730
box -6 -8 106 248
use NAND3X1  _1613_
timestamp 0
transform 1 0 2430 0 1 730
box -6 -8 106 248
use OAI21X1  _1614_
timestamp 0
transform 1 0 2290 0 1 730
box -6 -8 106 248
use NAND3X1  _1615_
timestamp 0
transform 1 0 2570 0 1 730
box -6 -8 106 248
use NAND2X1  _1616_
timestamp 0
transform -1 0 4090 0 1 250
box -6 -8 86 248
use NAND2X1  _1617_
timestamp 0
transform -1 0 4130 0 -1 730
box -6 -8 86 248
use OAI21X1  _1618_
timestamp 0
transform 1 0 4170 0 -1 730
box -6 -8 106 248
use AOI21X1  _1619_
timestamp 0
transform 1 0 4550 0 -1 250
box -6 -8 106 248
use OAI21X1  _1620_
timestamp 0
transform 1 0 4690 0 -1 250
box -6 -8 106 248
use AOI22X1  _1621_
timestamp 0
transform -1 0 5530 0 -1 250
box -6 -8 126 248
use INVX1  _1622_
timestamp 0
transform 1 0 4030 0 -1 250
box -6 -8 66 248
use AND2X2  _1623_
timestamp 0
transform -1 0 3710 0 -1 730
box -6 -8 106 248
use NAND3X1  _1624_
timestamp 0
transform -1 0 3990 0 -1 730
box -6 -8 106 248
use INVX1  _1625_
timestamp 0
transform -1 0 4250 0 1 730
box -6 -8 66 248
use AOI21X1  _1626_
timestamp 0
transform 1 0 3890 0 1 730
box -6 -8 106 248
use AOI21X1  _1627_
timestamp 0
transform -1 0 4130 0 1 730
box -6 -8 106 248
use OAI21X1  _1628_
timestamp 0
transform -1 0 4250 0 1 250
box -6 -8 106 248
use AOI21X1  _1629_
timestamp 0
transform 1 0 4130 0 -1 250
box -6 -8 106 248
use NAND2X1  _1630_
timestamp 0
transform -1 0 2230 0 -1 730
box -6 -8 86 248
use NOR2X1  _1631_
timestamp 0
transform -1 0 670 0 -1 1690
box -6 -8 86 248
use AOI21X1  _1632_
timestamp 0
transform -1 0 1310 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1633_
timestamp 0
transform 1 0 2050 0 1 250
box -6 -8 106 248
use INVX1  _1634_
timestamp 0
transform 1 0 2030 0 -1 730
box -6 -8 66 248
use OAI21X1  _1635_
timestamp 0
transform 1 0 2430 0 -1 730
box -6 -8 106 248
use NAND2X1  _1636_
timestamp 0
transform 1 0 2350 0 1 250
box -6 -8 86 248
use AOI21X1  _1637_
timestamp 0
transform 1 0 2770 0 1 250
box -6 -8 106 248
use NAND3X1  _1638_
timestamp 0
transform 1 0 2190 0 1 250
box -6 -8 106 248
use NAND2X1  _1639_
timestamp 0
transform 1 0 2490 0 1 250
box -6 -8 86 248
use AOI21X1  _1640_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 106 248
use NOR2X1  _1641_
timestamp 0
transform 1 0 3890 0 -1 250
box -6 -8 86 248
use NOR2X1  _1642_
timestamp 0
transform 1 0 4410 0 -1 250
box -6 -8 86 248
use NAND2X1  _1643_
timestamp 0
transform -1 0 4350 0 -1 250
box -6 -8 86 248
use OAI21X1  _1644_
timestamp 0
transform -1 0 4410 0 1 730
box -6 -8 106 248
use OAI21X1  _1645_
timestamp 0
transform 1 0 3570 0 -1 1210
box -6 -8 106 248
use INVX1  _1646_
timestamp 0
transform 1 0 3710 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1647_
timestamp 0
transform -1 0 4350 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1648_
timestamp 0
transform -1 0 5410 0 -1 1210
box -6 -8 106 248
use INVX1  _1649_
timestamp 0
transform 1 0 4750 0 1 1210
box -6 -8 66 248
use NAND3X1  _1650_
timestamp 0
transform 1 0 3070 0 1 250
box -6 -8 106 248
use AOI21X1  _1651_
timestamp 0
transform -1 0 3850 0 -1 250
box -6 -8 106 248
use AND2X2  _1652_
timestamp 0
transform 1 0 3210 0 1 250
box -6 -8 106 248
use NAND3X1  _1653_
timestamp 0
transform -1 0 2730 0 1 250
box -6 -8 106 248
use NAND3X1  _1654_
timestamp 0
transform 1 0 3350 0 1 250
box -6 -8 106 248
use OAI21X1  _1655_
timestamp 0
transform 1 0 3610 0 -1 250
box -6 -8 106 248
use NAND3X1  _1656_
timestamp 0
transform 1 0 2030 0 1 730
box -6 -8 106 248
use INVX1  _1657_
timestamp 0
transform 1 0 1110 0 -1 1690
box -6 -8 66 248
use INVX1  _1658_
timestamp 0
transform 1 0 1330 0 1 1210
box -6 -8 66 248
use OAI21X1  _1659_
timestamp 0
transform 1 0 1170 0 1 1210
box -6 -8 106 248
use INVX1  _1660_
timestamp 0
transform -1 0 1170 0 -1 730
box -6 -8 66 248
use NAND3X1  _1661_
timestamp 0
transform -1 0 1850 0 1 730
box -6 -8 106 248
use INVX1  _1662_
timestamp 0
transform 1 0 1630 0 1 730
box -6 -8 66 248
use AOI21X1  _1663_
timestamp 0
transform 1 0 1330 0 1 730
box -6 -8 106 248
use OAI21X1  _1664_
timestamp 0
transform -1 0 1590 0 1 730
box -6 -8 106 248
use OAI21X1  _1665_
timestamp 0
transform -1 0 1990 0 -1 730
box -6 -8 106 248
use NAND2X1  _1666_
timestamp 0
transform 1 0 1650 0 -1 730
box -6 -8 86 248
use NAND3X1  _1667_
timestamp 0
transform -1 0 1470 0 -1 730
box -6 -8 106 248
use AND2X2  _1668_
timestamp 0
transform 1 0 1510 0 -1 730
box -6 -8 106 248
use AND2X2  _1669_
timestamp 0
transform 1 0 2610 0 -1 250
box -6 -8 106 248
use OAI21X1  _1670_
timestamp 0
transform 1 0 2870 0 -1 250
box -6 -8 106 248
use OR2X2  _1671_
timestamp 0
transform 1 0 3010 0 -1 250
box -6 -8 106 248
use AOI22X1  _1672_
timestamp 0
transform -1 0 3950 0 -1 1210
box -6 -8 126 248
use INVX1  _1673_
timestamp 0
transform 1 0 1330 0 1 250
box -6 -8 66 248
use NOR2X1  _1674_
timestamp 0
transform 1 0 2750 0 -1 250
box -6 -8 86 248
use NOR2X1  _1675_
timestamp 0
transform 1 0 990 0 -1 730
box -6 -8 86 248
use OAI21X1  _1676_
timestamp 0
transform -1 0 1130 0 1 1210
box -6 -8 106 248
use INVX1  _1677_
timestamp 0
transform 1 0 570 0 1 250
box -6 -8 66 248
use OAI21X1  _1678_
timestamp 0
transform -1 0 910 0 1 250
box -6 -8 106 248
use NOR2X1  _1679_
timestamp 0
transform 1 0 1770 0 -1 730
box -6 -8 86 248
use NAND3X1  _1680_
timestamp 0
transform -1 0 1310 0 -1 730
box -6 -8 106 248
use NAND3X1  _1681_
timestamp 0
transform 1 0 790 0 -1 250
box -6 -8 106 248
use NAND3X1  _1682_
timestamp 0
transform 1 0 930 0 -1 250
box -6 -8 106 248
use AOI21X1  _1683_
timestamp 0
transform 1 0 470 0 -1 250
box -6 -8 106 248
use OAI21X1  _1684_
timestamp 0
transform -1 0 930 0 -1 730
box -6 -8 106 248
use NOR2X1  _1685_
timestamp 0
transform 1 0 670 0 1 250
box -6 -8 86 248
use OAI21X1  _1686_
timestamp 0
transform 1 0 630 0 -1 250
box -6 -8 106 248
use AND2X2  _1687_
timestamp 0
transform -1 0 1470 0 -1 250
box -6 -8 106 248
use AND2X2  _1688_
timestamp 0
transform 1 0 3150 0 -1 250
box -6 -8 106 248
use OAI21X1  _1689_
timestamp 0
transform 1 0 3310 0 -1 250
box -6 -8 106 248
use OAI21X1  _1690_
timestamp 0
transform 1 0 3450 0 -1 250
box -6 -8 106 248
use OAI21X1  _1691_
timestamp 0
transform 1 0 5170 0 1 730
box -6 -8 106 248
use OAI21X1  _1692_
timestamp 0
transform -1 0 710 0 -1 1210
box -6 -8 106 248
use INVX1  _1693_
timestamp 0
transform -1 0 250 0 -1 250
box -6 -8 66 248
use OAI21X1  _1694_
timestamp 0
transform -1 0 410 0 -1 250
box -6 -8 106 248
use OR2X2  _1695_
timestamp 0
transform 1 0 290 0 1 250
box -6 -8 106 248
use NAND2X1  _1696_
timestamp 0
transform 1 0 710 0 -1 730
box -6 -8 86 248
use AOI21X1  _1697_
timestamp 0
transform -1 0 270 0 -1 730
box -6 -8 106 248
use INVX1  _1698_
timestamp 0
transform 1 0 190 0 1 250
box -6 -8 66 248
use NAND3X1  _1699_
timestamp 0
transform 1 0 430 0 1 250
box -6 -8 106 248
use NOR2X1  _1700_
timestamp 0
transform -1 0 150 0 -1 250
box -6 -8 86 248
use OAI21X1  _1701_
timestamp 0
transform -1 0 150 0 1 250
box -6 -8 106 248
use NAND2X1  _1702_
timestamp 0
transform -1 0 1030 0 1 250
box -6 -8 86 248
use AOI21X1  _1703_
timestamp 0
transform 1 0 1090 0 -1 250
box -6 -8 106 248
use AOI21X1  _1704_
timestamp 0
transform -1 0 1330 0 -1 250
box -6 -8 106 248
use NAND3X1  _1705_
timestamp 0
transform -1 0 2550 0 -1 250
box -6 -8 106 248
use AOI21X1  _1706_
timestamp 0
transform -1 0 1930 0 -1 250
box -6 -8 106 248
use AND2X2  _1707_
timestamp 0
transform 1 0 1070 0 1 250
box -6 -8 106 248
use OAI21X1  _1708_
timestamp 0
transform -1 0 3610 0 1 250
box -6 -8 106 248
use NOR3X1  _1709_
timestamp 0
transform -1 0 3970 0 1 250
box -6 -8 186 248
use AOI21X1  _1710_
timestamp 0
transform -1 0 3750 0 1 250
box -6 -8 106 248
use NAND3X1  _1711_
timestamp 0
transform 1 0 1530 0 -1 250
box -6 -8 106 248
use OAI21X1  _1712_
timestamp 0
transform 1 0 1670 0 -1 250
box -6 -8 106 248
use OAI21X1  _1713_
timestamp 0
transform 1 0 1570 0 1 250
box -6 -8 106 248
use OR2X2  _1714_
timestamp 0
transform 1 0 1890 0 1 250
box -6 -8 106 248
use AOI22X1  _1715_
timestamp 0
transform -1 0 4430 0 -1 730
box -6 -8 126 248
use NAND2X1  _1716_
timestamp 0
transform 1 0 5290 0 -1 250
box -6 -8 86 248
use INVX1  _1717_
timestamp 0
transform -1 0 1290 0 1 250
box -6 -8 66 248
use OAI21X1  _1718_
timestamp 0
transform 1 0 310 0 -1 730
box -6 -8 106 248
use NAND2X1  _1719_
timestamp 0
transform -1 0 530 0 1 730
box -6 -8 86 248
use OR2X2  _1720_
timestamp 0
transform -1 0 390 0 1 730
box -6 -8 106 248
use NAND2X1  _1721_
timestamp 0
transform -1 0 530 0 -1 730
box -6 -8 86 248
use INVX1  _1722_
timestamp 0
transform 1 0 1990 0 -1 250
box -6 -8 66 248
use NOR3X1  _1723_
timestamp 0
transform 1 0 2090 0 -1 250
box -6 -8 186 248
use AOI21X1  _1724_
timestamp 0
transform -1 0 1530 0 1 250
box -6 -8 106 248
use OAI21X1  _1725_
timestamp 0
transform 1 0 1730 0 1 250
box -6 -8 106 248
use OAI21X1  _1726_
timestamp 0
transform 1 0 2310 0 -1 250
box -6 -8 106 248
use NAND2X1  _1727_
timestamp 0
transform -1 0 5010 0 -1 250
box -6 -8 86 248
use DFFPOSX1  _1728_
timestamp 0
transform -1 0 5890 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1729_
timestamp 0
transform 1 0 5370 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1730_
timestamp 0
transform -1 0 4690 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1731_
timestamp 0
transform -1 0 4890 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1732_
timestamp 0
transform 1 0 4010 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1733_
timestamp 0
transform -1 0 4870 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1734_
timestamp 0
transform 1 0 2550 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1735_
timestamp 0
transform 1 0 2010 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1736_
timestamp 0
transform 1 0 1370 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1737_
timestamp 0
transform 1 0 870 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1738_
timestamp 0
transform 1 0 390 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1739_
timestamp 0
transform 1 0 1230 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1740_
timestamp 0
transform 1 0 1630 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1741_
timestamp 0
transform 1 0 850 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1742_
timestamp 0
transform 1 0 4890 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1743_
timestamp 0
transform -1 0 5810 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1744_
timestamp 0
transform -1 0 5590 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1745_
timestamp 0
transform 1 0 5170 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1746_
timestamp 0
transform 1 0 3610 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1747_
timestamp 0
transform 1 0 2750 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1748_
timestamp 0
transform -1 0 5430 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1749_
timestamp 0
transform 1 0 3110 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1750_
timestamp 0
transform 1 0 4490 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1751_
timestamp 0
transform 1 0 4830 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1752_
timestamp 0
transform 1 0 4830 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _1753_
timestamp 0
transform 1 0 4910 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _1754_
timestamp 0
transform -1 0 650 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1755_
timestamp 0
transform 1 0 10 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1756_
timestamp 0
transform 1 0 10 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1757_
timestamp 0
transform 1 0 150 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1758_
timestamp 0
transform -1 0 1410 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1759_
timestamp 0
transform -1 0 1330 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1760_
timestamp 0
transform -1 0 2610 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1761_
timestamp 0
transform -1 0 2290 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1762_
timestamp 0
transform 1 0 3070 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1763_
timestamp 0
transform 1 0 2830 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1764_
timestamp 0
transform -1 0 5110 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1765_
timestamp 0
transform -1 0 4810 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1766_
timestamp 0
transform -1 0 250 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1767_
timestamp 0
transform -1 0 710 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1768_
timestamp 0
transform 1 0 810 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1769_
timestamp 0
transform 1 0 530 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1770_
timestamp 0
transform 1 0 2230 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1771_
timestamp 0
transform -1 0 2950 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1772_
timestamp 0
transform -1 0 3810 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1773_
timestamp 0
transform -1 0 3430 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1774_
timestamp 0
transform -1 0 4290 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _1775_
timestamp 0
transform 1 0 3950 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1776_
timestamp 0
transform 1 0 4550 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1777_
timestamp 0
transform -1 0 4070 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1778_
timestamp 0
transform -1 0 3810 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _1779_
timestamp 0
transform 1 0 1430 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1780_
timestamp 0
transform -1 0 4090 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1781_
timestamp 0
transform 1 0 2890 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1782_
timestamp 0
transform 1 0 2910 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1783_
timestamp 0
transform -1 0 4370 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1784_
timestamp 0
transform 1 0 2030 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1785_
timestamp 0
transform 1 0 1630 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1786_
timestamp 0
transform 1 0 5330 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1787_
timestamp 0
transform 1 0 4570 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1788_
timestamp 0
transform 1 0 4530 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1789_
timestamp 0
transform 1 0 5550 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1790_
timestamp 0
transform 1 0 130 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1791_
timestamp 0
transform 1 0 5470 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1792_
timestamp 0
transform -1 0 5890 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1793_
timestamp 0
transform -1 0 5890 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1794_
timestamp 0
transform -1 0 5350 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1795_
timestamp 0
transform -1 0 5410 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1796_
timestamp 0
transform -1 0 5170 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1797_
timestamp 0
transform 1 0 1890 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _1798_
timestamp 0
transform 1 0 5250 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1799_
timestamp 0
transform 1 0 5250 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1800_
timestamp 0
transform -1 0 5110 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1801_
timestamp 0
transform 1 0 5550 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1802_
timestamp 0
transform 1 0 5530 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1803_
timestamp 0
transform -1 0 5910 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1804_
timestamp 0
transform 1 0 4350 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1805_
timestamp 0
transform -1 0 5250 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1806_
timestamp 0
transform 1 0 4430 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1807_
timestamp 0
transform 1 0 5010 0 -1 250
box -6 -8 246 248
use BUFX2  _1808_
timestamp 0
transform -1 0 5110 0 -1 6010
box -6 -8 86 248
use BUFX2  _1809_
timestamp 0
transform -1 0 5470 0 -1 6010
box -6 -8 86 248
use BUFX2  _1810_
timestamp 0
transform 1 0 2270 0 -1 6010
box -6 -8 86 248
use BUFX2  _1811_
timestamp 0
transform 1 0 4410 0 -1 6010
box -6 -8 86 248
use BUFX2  _1812_
timestamp 0
transform 1 0 5750 0 -1 6010
box -6 -8 86 248
use BUFX2  _1813_
timestamp 0
transform 1 0 5670 0 -1 5530
box -6 -8 86 248
use BUFX2  _1814_
timestamp 0
transform 1 0 5850 0 -1 2170
box -6 -8 86 248
use BUFX2  _1815_
timestamp 0
transform 1 0 5830 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 3350 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform -1 0 1030 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 1830 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform -1 0 1070 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 3290 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform -1 0 3310 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 1730 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 4810 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 4830 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 5590 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform -1 0 5470 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 5450 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 2130 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform -1 0 1330 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform 1 0 2710 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 2970 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 1170 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 5070 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert26
timestamp 0
transform -1 0 4930 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert27
timestamp 0
transform 1 0 2410 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert28
timestamp 0
transform -1 0 2410 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert29
timestamp 0
transform -1 0 4690 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert30
timestamp 0
transform -1 0 1930 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert31
timestamp 0
transform -1 0 1950 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert32
timestamp 0
transform 1 0 3150 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert33
timestamp 0
transform 1 0 2830 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert34
timestamp 0
transform 1 0 4630 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert35
timestamp 0
transform -1 0 4810 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert36
timestamp 0
transform 1 0 5210 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert37
timestamp 0
transform 1 0 5150 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert38
timestamp 0
transform 1 0 5270 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert39
timestamp 0
transform -1 0 1410 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert40
timestamp 0
transform 1 0 2430 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert41
timestamp 0
transform 1 0 3590 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert42
timestamp 0
transform -1 0 1390 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert43
timestamp 0
transform 1 0 2550 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert44
timestamp 0
transform -1 0 1530 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert45
timestamp 0
transform 1 0 1610 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert46
timestamp 0
transform -1 0 1790 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert47
timestamp 0
transform 1 0 3390 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert48
timestamp 0
transform -1 0 1670 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert49
timestamp 0
transform 1 0 3350 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert50
timestamp 0
transform -1 0 2470 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert51
timestamp 0
transform 1 0 3230 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert52
timestamp 0
transform 1 0 2630 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert53
timestamp 0
transform -1 0 1990 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert54
timestamp 0
transform -1 0 630 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert55
timestamp 0
transform 1 0 3110 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert56
timestamp 0
transform -1 0 670 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert57
timestamp 0
transform -1 0 1090 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert58
timestamp 0
transform -1 0 3070 0 1 3610
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform -1 0 5870 0 1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform 1 0 670 0 -1 4090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform -1 0 5870 0 1 1690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert15
timestamp 0
transform -1 0 370 0 1 1210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert16
timestamp 0
transform -1 0 2270 0 1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert17
timestamp 0
transform -1 0 3170 0 1 1690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert18
timestamp 0
transform -1 0 5890 0 1 1210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert19
timestamp 0
transform -1 0 5850 0 -1 5050
box -6 -8 206 248
use FILL  FILL87150x64950
timestamp 0
transform -1 0 5830 0 -1 4570
box -6 -8 26 248
use FILL  FILL87450x21750
timestamp 0
transform -1 0 5850 0 -1 1690
box -6 -8 26 248
use FILL  FILL87450x39750
timestamp 0
transform 1 0 5830 0 1 2650
box -6 -8 26 248
use FILL  FILL87450x46950
timestamp 0
transform 1 0 5830 0 1 3130
box -6 -8 26 248
use FILL  FILL87450x61350
timestamp 0
transform 1 0 5830 0 1 4090
box -6 -8 26 248
use FILL  FILL87450x64950
timestamp 0
transform -1 0 5850 0 -1 4570
box -6 -8 26 248
use FILL  FILL87450x86550
timestamp 0
transform -1 0 5850 0 -1 6010
box -6 -8 26 248
use FILL  FILL87750x21750
timestamp 0
transform -1 0 5870 0 -1 1690
box -6 -8 26 248
use FILL  FILL87750x39750
timestamp 0
transform 1 0 5850 0 1 2650
box -6 -8 26 248
use FILL  FILL87750x46950
timestamp 0
transform 1 0 5850 0 1 3130
box -6 -8 26 248
use FILL  FILL87750x54150
timestamp 0
transform 1 0 5850 0 1 3610
box -6 -8 26 248
use FILL  FILL87750x61350
timestamp 0
transform 1 0 5850 0 1 4090
box -6 -8 26 248
use FILL  FILL87750x64950
timestamp 0
transform -1 0 5870 0 -1 4570
box -6 -8 26 248
use FILL  FILL87750x72150
timestamp 0
transform -1 0 5870 0 -1 5050
box -6 -8 26 248
use FILL  FILL87750x86550
timestamp 0
transform -1 0 5870 0 -1 6010
box -6 -8 26 248
use FILL  FILL88050x3750
timestamp 0
transform 1 0 5870 0 1 250
box -6 -8 26 248
use FILL  FILL88050x7350
timestamp 0
transform -1 0 5890 0 -1 730
box -6 -8 26 248
use FILL  FILL88050x21750
timestamp 0
transform -1 0 5890 0 -1 1690
box -6 -8 26 248
use FILL  FILL88050x25350
timestamp 0
transform 1 0 5870 0 1 1690
box -6 -8 26 248
use FILL  FILL88050x39750
timestamp 0
transform 1 0 5870 0 1 2650
box -6 -8 26 248
use FILL  FILL88050x46950
timestamp 0
transform 1 0 5870 0 1 3130
box -6 -8 26 248
use FILL  FILL88050x54150
timestamp 0
transform 1 0 5870 0 1 3610
box -6 -8 26 248
use FILL  FILL88050x57750
timestamp 0
transform -1 0 5890 0 -1 4090
box -6 -8 26 248
use FILL  FILL88050x61350
timestamp 0
transform 1 0 5870 0 1 4090
box -6 -8 26 248
use FILL  FILL88050x64950
timestamp 0
transform -1 0 5890 0 -1 4570
box -6 -8 26 248
use FILL  FILL88050x72150
timestamp 0
transform -1 0 5890 0 -1 5050
box -6 -8 26 248
use FILL  FILL88050x75750
timestamp 0
transform 1 0 5870 0 1 5050
box -6 -8 26 248
use FILL  FILL88050x79350
timestamp 0
transform -1 0 5890 0 -1 5530
box -6 -8 26 248
use FILL  FILL88050x86550
timestamp 0
transform -1 0 5890 0 -1 6010
box -6 -8 26 248
use FILL  FILL88350x3750
timestamp 0
transform 1 0 5890 0 1 250
box -6 -8 26 248
use FILL  FILL88350x7350
timestamp 0
transform -1 0 5910 0 -1 730
box -6 -8 26 248
use FILL  FILL88350x18150
timestamp 0
transform 1 0 5890 0 1 1210
box -6 -8 26 248
use FILL  FILL88350x21750
timestamp 0
transform -1 0 5910 0 -1 1690
box -6 -8 26 248
use FILL  FILL88350x25350
timestamp 0
transform 1 0 5890 0 1 1690
box -6 -8 26 248
use FILL  FILL88350x36150
timestamp 0
transform -1 0 5910 0 -1 2650
box -6 -8 26 248
use FILL  FILL88350x39750
timestamp 0
transform 1 0 5890 0 1 2650
box -6 -8 26 248
use FILL  FILL88350x43350
timestamp 0
transform -1 0 5910 0 -1 3130
box -6 -8 26 248
use FILL  FILL88350x46950
timestamp 0
transform 1 0 5890 0 1 3130
box -6 -8 26 248
use FILL  FILL88350x54150
timestamp 0
transform 1 0 5890 0 1 3610
box -6 -8 26 248
use FILL  FILL88350x57750
timestamp 0
transform -1 0 5910 0 -1 4090
box -6 -8 26 248
use FILL  FILL88350x61350
timestamp 0
transform 1 0 5890 0 1 4090
box -6 -8 26 248
use FILL  FILL88350x64950
timestamp 0
transform -1 0 5910 0 -1 4570
box -6 -8 26 248
use FILL  FILL88350x72150
timestamp 0
transform -1 0 5910 0 -1 5050
box -6 -8 26 248
use FILL  FILL88350x75750
timestamp 0
transform 1 0 5890 0 1 5050
box -6 -8 26 248
use FILL  FILL88350x79350
timestamp 0
transform -1 0 5910 0 -1 5530
box -6 -8 26 248
use FILL  FILL88350x82950
timestamp 0
transform 1 0 5890 0 1 5530
box -6 -8 26 248
use FILL  FILL88350x86550
timestamp 0
transform -1 0 5910 0 -1 6010
box -6 -8 26 248
use FILL  FILL88650x150
timestamp 0
transform -1 0 5930 0 -1 250
box -6 -8 26 248
use FILL  FILL88650x3750
timestamp 0
transform 1 0 5910 0 1 250
box -6 -8 26 248
use FILL  FILL88650x7350
timestamp 0
transform -1 0 5930 0 -1 730
box -6 -8 26 248
use FILL  FILL88650x10950
timestamp 0
transform 1 0 5910 0 1 730
box -6 -8 26 248
use FILL  FILL88650x14550
timestamp 0
transform -1 0 5930 0 -1 1210
box -6 -8 26 248
use FILL  FILL88650x18150
timestamp 0
transform 1 0 5910 0 1 1210
box -6 -8 26 248
use FILL  FILL88650x21750
timestamp 0
transform -1 0 5930 0 -1 1690
box -6 -8 26 248
use FILL  FILL88650x25350
timestamp 0
transform 1 0 5910 0 1 1690
box -6 -8 26 248
use FILL  FILL88650x32550
timestamp 0
transform 1 0 5910 0 1 2170
box -6 -8 26 248
use FILL  FILL88650x36150
timestamp 0
transform -1 0 5930 0 -1 2650
box -6 -8 26 248
use FILL  FILL88650x39750
timestamp 0
transform 1 0 5910 0 1 2650
box -6 -8 26 248
use FILL  FILL88650x43350
timestamp 0
transform -1 0 5930 0 -1 3130
box -6 -8 26 248
use FILL  FILL88650x46950
timestamp 0
transform 1 0 5910 0 1 3130
box -6 -8 26 248
use FILL  FILL88650x50550
timestamp 0
transform -1 0 5930 0 -1 3610
box -6 -8 26 248
use FILL  FILL88650x54150
timestamp 0
transform 1 0 5910 0 1 3610
box -6 -8 26 248
use FILL  FILL88650x57750
timestamp 0
transform -1 0 5930 0 -1 4090
box -6 -8 26 248
use FILL  FILL88650x61350
timestamp 0
transform 1 0 5910 0 1 4090
box -6 -8 26 248
use FILL  FILL88650x64950
timestamp 0
transform -1 0 5930 0 -1 4570
box -6 -8 26 248
use FILL  FILL88650x72150
timestamp 0
transform -1 0 5930 0 -1 5050
box -6 -8 26 248
use FILL  FILL88650x75750
timestamp 0
transform 1 0 5910 0 1 5050
box -6 -8 26 248
use FILL  FILL88650x79350
timestamp 0
transform -1 0 5930 0 -1 5530
box -6 -8 26 248
use FILL  FILL88650x82950
timestamp 0
transform 1 0 5910 0 1 5530
box -6 -8 26 248
use FILL  FILL88650x86550
timestamp 0
transform -1 0 5930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__863_
timestamp 0
transform 1 0 5070 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__864_
timestamp 0
transform -1 0 4870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__865_
timestamp 0
transform 1 0 5330 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__866_
timestamp 0
transform -1 0 5370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__867_
timestamp 0
transform 1 0 5250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__868_
timestamp 0
transform -1 0 4370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__869_
timestamp 0
transform -1 0 5170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__870_
timestamp 0
transform 1 0 5490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__871_
timestamp 0
transform -1 0 5070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__872_
timestamp 0
transform 1 0 5470 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__873_
timestamp 0
transform 1 0 5710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__874_
timestamp 0
transform 1 0 5750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__875_
timestamp 0
transform -1 0 5430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__876_
timestamp 0
transform 1 0 5290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__877_
timestamp 0
transform -1 0 5150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__878_
timestamp 0
transform -1 0 5210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__879_
timestamp 0
transform 1 0 5150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__880_
timestamp 0
transform -1 0 5090 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__881_
timestamp 0
transform -1 0 5230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__882_
timestamp 0
transform 1 0 3350 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__883_
timestamp 0
transform 1 0 3730 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__884_
timestamp 0
transform 1 0 3590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__885_
timestamp 0
transform 1 0 5350 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__886_
timestamp 0
transform 1 0 5410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__887_
timestamp 0
transform -1 0 5530 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__888_
timestamp 0
transform 1 0 5270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__889_
timestamp 0
transform -1 0 4830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__890_
timestamp 0
transform -1 0 4950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__891_
timestamp 0
transform 1 0 5750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__892_
timestamp 0
transform -1 0 4790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__893_
timestamp 0
transform 1 0 5110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__894_
timestamp 0
transform 1 0 5350 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__895_
timestamp 0
transform -1 0 5510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__896_
timestamp 0
transform -1 0 5690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__897_
timestamp 0
transform 1 0 5430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__898_
timestamp 0
transform -1 0 4930 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__899_
timestamp 0
transform 1 0 5210 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__900_
timestamp 0
transform 1 0 5070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__901_
timestamp 0
transform -1 0 5590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__902_
timestamp 0
transform 1 0 5790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__903_
timestamp 0
transform 1 0 5410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__904_
timestamp 0
transform 1 0 5510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__905_
timestamp 0
transform 1 0 5650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__906_
timestamp 0
transform 1 0 5650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__907_
timestamp 0
transform 1 0 1850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__908_
timestamp 0
transform -1 0 1250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__909_
timestamp 0
transform 1 0 1870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__910_
timestamp 0
transform 1 0 1610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__911_
timestamp 0
transform 1 0 2790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__912_
timestamp 0
transform -1 0 2410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__913_
timestamp 0
transform 1 0 2710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__914_
timestamp 0
transform -1 0 4330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__915_
timestamp 0
transform 1 0 4270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__916_
timestamp 0
transform 1 0 1210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__917_
timestamp 0
transform -1 0 1450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__918_
timestamp 0
transform 1 0 1710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__919_
timestamp 0
transform 1 0 1110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__920_
timestamp 0
transform -1 0 2150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__921_
timestamp 0
transform -1 0 2250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__922_
timestamp 0
transform -1 0 2570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__923_
timestamp 0
transform -1 0 4510 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__924_
timestamp 0
transform 1 0 4490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__925_
timestamp 0
transform -1 0 5570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__926_
timestamp 0
transform -1 0 4330 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__927_
timestamp 0
transform 1 0 1010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__928_
timestamp 0
transform -1 0 2970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__929_
timestamp 0
transform -1 0 2910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__930_
timestamp 0
transform -1 0 3030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__931_
timestamp 0
transform 1 0 4030 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__932_
timestamp 0
transform -1 0 3950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__933_
timestamp 0
transform -1 0 3990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__934_
timestamp 0
transform 1 0 3030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__935_
timestamp 0
transform 1 0 1230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__936_
timestamp 0
transform -1 0 1050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__937_
timestamp 0
transform -1 0 1190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__938_
timestamp 0
transform 1 0 2150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__939_
timestamp 0
transform 1 0 1950 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__940_
timestamp 0
transform 1 0 1810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__941_
timestamp 0
transform 1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__942_
timestamp 0
transform -1 0 2970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__943_
timestamp 0
transform -1 0 4250 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__944_
timestamp 0
transform -1 0 4110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__945_
timestamp 0
transform -1 0 4510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__946_
timestamp 0
transform 1 0 1790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__947_
timestamp 0
transform -1 0 2210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__948_
timestamp 0
transform 1 0 2290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__949_
timestamp 0
transform -1 0 990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__950_
timestamp 0
transform 1 0 4350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__951_
timestamp 0
transform -1 0 5430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__952_
timestamp 0
transform -1 0 5450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__953_
timestamp 0
transform 1 0 5530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__954_
timestamp 0
transform -1 0 4070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__955_
timestamp 0
transform 1 0 3430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__956_
timestamp 0
transform 1 0 3470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__957_
timestamp 0
transform -1 0 2970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__958_
timestamp 0
transform -1 0 3770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__959_
timestamp 0
transform 1 0 2790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__960_
timestamp 0
transform -1 0 1090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__961_
timestamp 0
transform -1 0 2070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__962_
timestamp 0
transform 1 0 1390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__963_
timestamp 0
transform -1 0 2790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__964_
timestamp 0
transform 1 0 4070 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__965_
timestamp 0
transform 1 0 1630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__966_
timestamp 0
transform -1 0 2410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__967_
timestamp 0
transform 1 0 2270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__968_
timestamp 0
transform -1 0 2310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__969_
timestamp 0
transform -1 0 4190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__970_
timestamp 0
transform 1 0 3550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__971_
timestamp 0
transform -1 0 3690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__972_
timestamp 0
transform 1 0 2850 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__973_
timestamp 0
transform 1 0 1070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__974_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__975_
timestamp 0
transform -1 0 1050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__976_
timestamp 0
transform -1 0 1970 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__977_
timestamp 0
transform 1 0 1410 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__978_
timestamp 0
transform -1 0 1690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__979_
timestamp 0
transform 1 0 1750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__980_
timestamp 0
transform 1 0 3110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__981_
timestamp 0
transform 1 0 3230 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__982_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__983_
timestamp 0
transform -1 0 3590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__984_
timestamp 0
transform 1 0 2490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__985_
timestamp 0
transform 1 0 850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__986_
timestamp 0
transform -1 0 1630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__987_
timestamp 0
transform 1 0 1590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__988_
timestamp 0
transform -1 0 2490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__989_
timestamp 0
transform -1 0 3430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__990_
timestamp 0
transform 1 0 4230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__991_
timestamp 0
transform 1 0 4650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__992_
timestamp 0
transform 1 0 4370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__993_
timestamp 0
transform 1 0 4770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__994_
timestamp 0
transform 1 0 4790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__995_
timestamp 0
transform 1 0 4910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__996_
timestamp 0
transform 1 0 4950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__997_
timestamp 0
transform 1 0 5210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__998_
timestamp 0
transform 1 0 4450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__999_
timestamp 0
transform -1 0 3970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1000_
timestamp 0
transform 1 0 4090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 3570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1002_
timestamp 0
transform 1 0 3690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1003_
timestamp 0
transform -1 0 3850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1004_
timestamp 0
transform 1 0 3650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1005_
timestamp 0
transform 1 0 3670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1006_
timestamp 0
transform 1 0 2490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 2350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1008_
timestamp 0
transform 1 0 2210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1009_
timestamp 0
transform -1 0 3450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 3190 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1011_
timestamp 0
transform 1 0 3030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1012_
timestamp 0
transform 1 0 2170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 3310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1014_
timestamp 0
transform 1 0 3450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 3810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1016_
timestamp 0
transform -1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1017_
timestamp 0
transform 1 0 3490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1018_
timestamp 0
transform 1 0 4150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1019_
timestamp 0
transform 1 0 4310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1020_
timestamp 0
transform 1 0 5010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1021_
timestamp 0
transform 1 0 4010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1022_
timestamp 0
transform 1 0 4350 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 3470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1024_
timestamp 0
transform -1 0 3510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1025_
timestamp 0
transform -1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1026_
timestamp 0
transform 1 0 4090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1028_
timestamp 0
transform 1 0 2830 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1029_
timestamp 0
transform -1 0 1490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 1750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 3110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1032_
timestamp 0
transform -1 0 2490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1033_
timestamp 0
transform -1 0 2630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 1910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1035_
timestamp 0
transform -1 0 3390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1036_
timestamp 0
transform 1 0 4010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1037_
timestamp 0
transform -1 0 3770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1038_
timestamp 0
transform 1 0 3850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 4310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 4430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 4150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 4290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 3810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1044_
timestamp 0
transform -1 0 4070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1045_
timestamp 0
transform -1 0 3930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1046_
timestamp 0
transform 1 0 4150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 4870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1048_
timestamp 0
transform 1 0 4250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 4150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 3610 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1051_
timestamp 0
transform 1 0 710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 1210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1053_
timestamp 0
transform -1 0 1350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 1910 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1055_
timestamp 0
transform 1 0 1750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 2290 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 2350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1058_
timestamp 0
transform 1 0 2650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1059_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 3070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1061_
timestamp 0
transform 1 0 2710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 2630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1063_
timestamp 0
transform -1 0 3610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 3870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 3330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 3430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1067_
timestamp 0
transform 1 0 3730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1068_
timestamp 0
transform -1 0 3430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1069_
timestamp 0
transform -1 0 3610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 3670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1071_
timestamp 0
transform 1 0 3710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1072_
timestamp 0
transform 1 0 3950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 4050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1074_
timestamp 0
transform 1 0 3850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1075_
timestamp 0
transform -1 0 4390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 3550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 3130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 2690 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 10 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1080_
timestamp 0
transform -1 0 730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1081_
timestamp 0
transform -1 0 870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 1330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1083_
timestamp 0
transform 1 0 910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1084_
timestamp 0
transform -1 0 2490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 3210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1086_
timestamp 0
transform 1 0 2590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1087_
timestamp 0
transform 1 0 2210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 2410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1089_
timestamp 0
transform -1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 2310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 2170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 2490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1093_
timestamp 0
transform 1 0 2810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1094_
timestamp 0
transform -1 0 2350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 2910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1096_
timestamp 0
transform 1 0 3410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1097_
timestamp 0
transform -1 0 3190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1098_
timestamp 0
transform 1 0 3570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 4490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1100_
timestamp 0
transform -1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 2570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1102_
timestamp 0
transform -1 0 290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1103_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 1070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1106_
timestamp 0
transform -1 0 1330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 1590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1108_
timestamp 0
transform -1 0 1690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1109_
timestamp 0
transform 1 0 1730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1110_
timestamp 0
transform 1 0 1910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 1590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1112_
timestamp 0
transform 1 0 1770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1113_
timestamp 0
transform -1 0 2150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1114_
timestamp 0
transform 1 0 2010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 1870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1116_
timestamp 0
transform -1 0 1610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1117_
timestamp 0
transform 1 0 1730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 2110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1119_
timestamp 0
transform -1 0 1990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1120_
timestamp 0
transform 1 0 2250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 2270 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1122_
timestamp 0
transform 1 0 1830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 1250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 1530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1125_
timestamp 0
transform -1 0 890 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1126_
timestamp 0
transform -1 0 390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1129_
timestamp 0
transform -1 0 1010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 1650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1131_
timestamp 0
transform 1 0 1370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1132_
timestamp 0
transform -1 0 1490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1133_
timestamp 0
transform 1 0 1810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1134_
timestamp 0
transform -1 0 1470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 1370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1136_
timestamp 0
transform 1 0 1310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1137_
timestamp 0
transform 1 0 1610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1138_
timestamp 0
transform 1 0 1630 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 1890 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1140_
timestamp 0
transform -1 0 1770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1141_
timestamp 0
transform -1 0 1970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 1050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 990 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1144_
timestamp 0
transform 1 0 630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1145_
timestamp 0
transform 1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 710 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1147_
timestamp 0
transform 1 0 870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1148_
timestamp 0
transform -1 0 1090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1149_
timestamp 0
transform -1 0 890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 1070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1151_
timestamp 0
transform -1 0 1210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1152_
timestamp 0
transform 1 0 810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1153_
timestamp 0
transform -1 0 1110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1154_
timestamp 0
transform -1 0 1490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1155_
timestamp 0
transform -1 0 1530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1156_
timestamp 0
transform -1 0 1250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 1390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 1330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 1190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1160_
timestamp 0
transform 1 0 1230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1161_
timestamp 0
transform 1 0 1370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 1530 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 1570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1164_
timestamp 0
transform -1 0 690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1165_
timestamp 0
transform 1 0 830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1166_
timestamp 0
transform -1 0 1230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1167_
timestamp 0
transform 1 0 270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1168_
timestamp 0
transform -1 0 310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1170_
timestamp 0
transform -1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1171_
timestamp 0
transform -1 0 930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1174_
timestamp 0
transform -1 0 530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1176_
timestamp 0
transform -1 0 790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1177_
timestamp 0
transform 1 0 870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1178_
timestamp 0
transform 1 0 950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1179_
timestamp 0
transform 1 0 1090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1180_
timestamp 0
transform -1 0 1050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1182_
timestamp 0
transform 1 0 750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1183_
timestamp 0
transform -1 0 610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1184_
timestamp 0
transform -1 0 1050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1185_
timestamp 0
transform 1 0 310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1186_
timestamp 0
transform -1 0 750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1188_
timestamp 0
transform -1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1191_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1192_
timestamp 0
transform -1 0 290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1194_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1195_
timestamp 0
transform -1 0 130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1197_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1198_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1199_
timestamp 0
transform 1 0 10 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1200_
timestamp 0
transform -1 0 170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1201_
timestamp 0
transform -1 0 30 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1204_
timestamp 0
transform 1 0 350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1205_
timestamp 0
transform -1 0 130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 1350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 30 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1212_
timestamp 0
transform 1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 10 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1215_
timestamp 0
transform -1 0 330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1216_
timestamp 0
transform 1 0 150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1217_
timestamp 0
transform -1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1218_
timestamp 0
transform 1 0 10 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1219_
timestamp 0
transform -1 0 30 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 130 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 350 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1223_
timestamp 0
transform -1 0 1110 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1224_
timestamp 0
transform -1 0 710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1226_
timestamp 0
transform -1 0 30 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1230_
timestamp 0
transform -1 0 390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1231_
timestamp 0
transform -1 0 550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1234_
timestamp 0
transform 1 0 790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1235_
timestamp 0
transform 1 0 570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1236_
timestamp 0
transform -1 0 450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1237_
timestamp 0
transform -1 0 410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1238_
timestamp 0
transform -1 0 30 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1239_
timestamp 0
transform 1 0 170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1241_
timestamp 0
transform -1 0 470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1243_
timestamp 0
transform 1 0 610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1245_
timestamp 0
transform -1 0 750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1246_
timestamp 0
transform -1 0 1490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1247_
timestamp 0
transform 1 0 250 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1248_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1250_
timestamp 0
transform -1 0 170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1254_
timestamp 0
transform 1 0 750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1255_
timestamp 0
transform -1 0 850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1256_
timestamp 0
transform 1 0 550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1258_
timestamp 0
transform -1 0 750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1259_
timestamp 0
transform -1 0 890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1260_
timestamp 0
transform 1 0 4770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1261_
timestamp 0
transform 1 0 4250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1262_
timestamp 0
transform -1 0 2450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 3650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1264_
timestamp 0
transform 1 0 4890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1265_
timestamp 0
transform 1 0 4590 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 4730 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 5270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1268_
timestamp 0
transform 1 0 5130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1269_
timestamp 0
transform 1 0 5530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1270_
timestamp 0
transform -1 0 2090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1271_
timestamp 0
transform -1 0 3590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1272_
timestamp 0
transform -1 0 3210 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1273_
timestamp 0
transform -1 0 3850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1274_
timestamp 0
transform 1 0 3970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1275_
timestamp 0
transform 1 0 5430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 5330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 5570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1278_
timestamp 0
transform -1 0 5730 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1279_
timestamp 0
transform 1 0 5750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 5770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 5690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 5250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 5790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 5730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1286_
timestamp 0
transform 1 0 4590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 4750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1288_
timestamp 0
transform 1 0 5570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1289_
timestamp 0
transform 1 0 5510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 5710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1291_
timestamp 0
transform -1 0 5490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1292_
timestamp 0
transform 1 0 5810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 5590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1294_
timestamp 0
transform 1 0 5710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1295_
timestamp 0
transform -1 0 5610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 5590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 5470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1298_
timestamp 0
transform 1 0 4810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1299_
timestamp 0
transform -1 0 3830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 3890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1301_
timestamp 0
transform -1 0 4310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1302_
timestamp 0
transform 1 0 4430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1303_
timestamp 0
transform 1 0 5030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1304_
timestamp 0
transform -1 0 4930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1305_
timestamp 0
transform 1 0 4950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1307_
timestamp 0
transform 1 0 5210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 5310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1309_
timestamp 0
transform -1 0 5130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1310_
timestamp 0
transform -1 0 4910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1311_
timestamp 0
transform -1 0 5030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1312_
timestamp 0
transform 1 0 4230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 3150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1314_
timestamp 0
transform 1 0 3170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1315_
timestamp 0
transform -1 0 3070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 3030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 2630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 2530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1319_
timestamp 0
transform -1 0 2890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 4830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1321_
timestamp 0
transform 1 0 2790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 2670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 2930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1324_
timestamp 0
transform -1 0 2510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 3310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 2990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1327_
timestamp 0
transform -1 0 2550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1328_
timestamp 0
transform -1 0 3430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 3330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 2510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 2550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1332_
timestamp 0
transform -1 0 2290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1333_
timestamp 0
transform -1 0 1990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1334_
timestamp 0
transform 1 0 2130 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1335_
timestamp 0
transform -1 0 1890 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1336_
timestamp 0
transform -1 0 2250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1337_
timestamp 0
transform 1 0 2390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 2410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1339_
timestamp 0
transform 1 0 2490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1340_
timestamp 0
transform 1 0 2430 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 2370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 2610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 2690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1344_
timestamp 0
transform 1 0 2510 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 3170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1346_
timestamp 0
transform -1 0 3370 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 3550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1348_
timestamp 0
transform 1 0 3690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1350_
timestamp 0
transform 1 0 3290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1351_
timestamp 0
transform -1 0 3050 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 3270 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1353_
timestamp 0
transform 1 0 3290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1354_
timestamp 0
transform 1 0 4470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 4610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1356_
timestamp 0
transform -1 0 4910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 3230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 3710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 4350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1360_
timestamp 0
transform -1 0 4510 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1361_
timestamp 0
transform 1 0 4190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1362_
timestamp 0
transform 1 0 3830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1363_
timestamp 0
transform -1 0 2970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 3730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 3370 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 3370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1367_
timestamp 0
transform 1 0 3270 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 3150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1369_
timestamp 0
transform -1 0 3430 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1370_
timestamp 0
transform 1 0 4730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1371_
timestamp 0
transform 1 0 4130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 4170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 3950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1374_
timestamp 0
transform 1 0 3810 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1375_
timestamp 0
transform 1 0 4030 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 4150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 3890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 3730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 3090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1380_
timestamp 0
transform -1 0 3210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1381_
timestamp 0
transform -1 0 3110 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 3050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 2830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1384_
timestamp 0
transform 1 0 2950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1385_
timestamp 0
transform 1 0 3810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1386_
timestamp 0
transform 1 0 3930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 4050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 4190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1389_
timestamp 0
transform -1 0 4730 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1390_
timestamp 0
transform 1 0 3450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1391_
timestamp 0
transform -1 0 3570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1392_
timestamp 0
transform -1 0 2890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1393_
timestamp 0
transform -1 0 3130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 2990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1395_
timestamp 0
transform 1 0 3230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1396_
timestamp 0
transform 1 0 4270 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1397_
timestamp 0
transform 1 0 4410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 4570 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1399_
timestamp 0
transform -1 0 3370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1400_
timestamp 0
transform 1 0 4110 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 4030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1402_
timestamp 0
transform 1 0 3870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 3490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 3650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 3510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 3770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 4190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 4330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1409_
timestamp 0
transform -1 0 4430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 4810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1411_
timestamp 0
transform -1 0 4050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 4650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1413_
timestamp 0
transform -1 0 4850 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 4710 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1415_
timestamp 0
transform 1 0 810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1417_
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1419_
timestamp 0
transform 1 0 5390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1420_
timestamp 0
transform -1 0 5270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1423_
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1424_
timestamp 0
transform -1 0 30 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 4870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 1490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1427_
timestamp 0
transform 1 0 1330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1428_
timestamp 0
transform -1 0 1330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 1170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 3950 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 2190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 2230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 1810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1434_
timestamp 0
transform -1 0 1950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1435_
timestamp 0
transform -1 0 2690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1436_
timestamp 0
transform -1 0 2810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 2810 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1438_
timestamp 0
transform 1 0 2670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1439_
timestamp 0
transform -1 0 4630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1440_
timestamp 0
transform 1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 4310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1442_
timestamp 0
transform -1 0 4450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1443_
timestamp 0
transform -1 0 190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 10 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1445_
timestamp 0
transform -1 0 450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1446_
timestamp 0
transform 1 0 290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1447_
timestamp 0
transform 1 0 1170 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 1050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1449_
timestamp 0
transform -1 0 1070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1450_
timestamp 0
transform 1 0 910 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1451_
timestamp 0
transform 1 0 770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1452_
timestamp 0
transform -1 0 1970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1453_
timestamp 0
transform -1 0 2110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1454_
timestamp 0
transform 1 0 2910 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1455_
timestamp 0
transform 1 0 2750 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1456_
timestamp 0
transform -1 0 3390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1457_
timestamp 0
transform 1 0 3310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1458_
timestamp 0
transform 1 0 3950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1459_
timestamp 0
transform 1 0 3810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 4590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 4290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1462_
timestamp 0
transform 1 0 4590 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1463_
timestamp 0
transform 1 0 4450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1464_
timestamp 0
transform 1 0 4450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 4410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1466_
timestamp 0
transform -1 0 4230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1467_
timestamp 0
transform -1 0 4190 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1468_
timestamp 0
transform -1 0 2690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1469_
timestamp 0
transform -1 0 3470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1470_
timestamp 0
transform -1 0 1350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1471_
timestamp 0
transform -1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1472_
timestamp 0
transform -1 0 3490 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1473_
timestamp 0
transform -1 0 4110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1474_
timestamp 0
transform -1 0 2770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1475_
timestamp 0
transform -1 0 2810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1476_
timestamp 0
transform -1 0 2650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1477_
timestamp 0
transform -1 0 2770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1478_
timestamp 0
transform -1 0 4550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1479_
timestamp 0
transform -1 0 3930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1480_
timestamp 0
transform -1 0 4390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 2430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1482_
timestamp 0
transform -1 0 2410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1483_
timestamp 0
transform 1 0 1890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 1770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1485_
timestamp 0
transform 1 0 5010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1486_
timestamp 0
transform 1 0 4770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1487_
timestamp 0
transform 1 0 5190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 5050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1489_
timestamp 0
transform -1 0 4910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1490_
timestamp 0
transform 1 0 4630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 4330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1492_
timestamp 0
transform -1 0 4470 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1493_
timestamp 0
transform -1 0 5290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1494_
timestamp 0
transform -1 0 5410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1495_
timestamp 0
transform 1 0 2130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1496_
timestamp 0
transform -1 0 770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1497_
timestamp 0
transform -1 0 1750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1498_
timestamp 0
transform -1 0 5010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1499_
timestamp 0
transform 1 0 4510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1500_
timestamp 0
transform -1 0 2970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1501_
timestamp 0
transform -1 0 550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1502_
timestamp 0
transform -1 0 1110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1503_
timestamp 0
transform -1 0 2130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1504_
timestamp 0
transform -1 0 2050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1505_
timestamp 0
transform 1 0 3090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1506_
timestamp 0
transform 1 0 2770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1507_
timestamp 0
transform -1 0 2570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1508_
timestamp 0
transform 1 0 2610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1509_
timestamp 0
transform 1 0 2730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1510_
timestamp 0
transform 1 0 2470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1511_
timestamp 0
transform -1 0 1930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1512_
timestamp 0
transform -1 0 2050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1513_
timestamp 0
transform -1 0 1890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1514_
timestamp 0
transform -1 0 1450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1515_
timestamp 0
transform 1 0 1730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1516_
timestamp 0
transform 1 0 2330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1517_
timestamp 0
transform 1 0 2610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1518_
timestamp 0
transform -1 0 2210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1519_
timestamp 0
transform 1 0 1910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1520_
timestamp 0
transform 1 0 1630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1521_
timestamp 0
transform -1 0 2070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1522_
timestamp 0
transform 1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 3170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1524_
timestamp 0
transform -1 0 3290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1525_
timestamp 0
transform 1 0 3790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1526_
timestamp 0
transform -1 0 3670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 4850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 4950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1529_
timestamp 0
transform -1 0 5070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 5310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 5110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1532_
timestamp 0
transform -1 0 5190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1533_
timestamp 0
transform 1 0 3790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 5130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 5670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1536_
timestamp 0
transform 1 0 5090 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1537_
timestamp 0
transform 1 0 4710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1538_
timestamp 0
transform 1 0 4790 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1539_
timestamp 0
transform -1 0 2810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1540_
timestamp 0
transform 1 0 550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1541_
timestamp 0
transform 1 0 390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1542_
timestamp 0
transform -1 0 1490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1543_
timestamp 0
transform -1 0 1550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1544_
timestamp 0
transform -1 0 1950 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1545_
timestamp 0
transform -1 0 1750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 1590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1547_
timestamp 0
transform 1 0 2490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1548_
timestamp 0
transform -1 0 2290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1549_
timestamp 0
transform -1 0 270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1550_
timestamp 0
transform -1 0 390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1551_
timestamp 0
transform 1 0 1330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1552_
timestamp 0
transform 1 0 1190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1553_
timestamp 0
transform 1 0 1830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1554_
timestamp 0
transform -1 0 2150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1555_
timestamp 0
transform 1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1556_
timestamp 0
transform 1 0 4970 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1557_
timestamp 0
transform 1 0 5090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1558_
timestamp 0
transform 1 0 5210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1559_
timestamp 0
transform 1 0 5330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1560_
timestamp 0
transform 1 0 5450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1561_
timestamp 0
transform 1 0 5590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1562_
timestamp 0
transform -1 0 5510 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 2010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1564_
timestamp 0
transform -1 0 390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1565_
timestamp 0
transform -1 0 530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1566_
timestamp 0
transform -1 0 690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1567_
timestamp 0
transform -1 0 830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1568_
timestamp 0
transform -1 0 970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 1450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1570_
timestamp 0
transform 1 0 2950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1571_
timestamp 0
transform -1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1572_
timestamp 0
transform -1 0 2970 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1573_
timestamp 0
transform 1 0 2810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1574_
timestamp 0
transform 1 0 3350 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1575_
timestamp 0
transform -1 0 3510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1576_
timestamp 0
transform 1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1577_
timestamp 0
transform 1 0 3610 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1578_
timestamp 0
transform 1 0 4250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1579_
timestamp 0
transform -1 0 4790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1581_
timestamp 0
transform 1 0 4390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1582_
timestamp 0
transform -1 0 4550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 4610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1584_
timestamp 0
transform -1 0 4690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1585_
timestamp 0
transform 1 0 4670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1586_
timestamp 0
transform -1 0 670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1587_
timestamp 0
transform 1 0 950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1588_
timestamp 0
transform 1 0 1690 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1589_
timestamp 0
transform 1 0 1530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1590_
timestamp 0
transform 1 0 2110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1591_
timestamp 0
transform -1 0 3090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1592_
timestamp 0
transform 1 0 2930 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1593_
timestamp 0
transform 1 0 3750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1594_
timestamp 0
transform 1 0 3070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1595_
timestamp 0
transform 1 0 3710 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1596_
timestamp 0
transform -1 0 3390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1597_
timestamp 0
transform -1 0 3230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1598_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1599_
timestamp 0
transform 1 0 4710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1600_
timestamp 0
transform 1 0 4550 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1601_
timestamp 0
transform 1 0 4850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1602_
timestamp 0
transform 1 0 4990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1603_
timestamp 0
transform -1 0 5410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1604_
timestamp 0
transform -1 0 2690 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1606_
timestamp 0
transform -1 0 1330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1607_
timestamp 0
transform 1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1608_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1609_
timestamp 0
transform 1 0 1890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1610_
timestamp 0
transform 1 0 2130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1611_
timestamp 0
transform 1 0 2230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1612_
timestamp 0
transform 1 0 2690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1613_
timestamp 0
transform 1 0 2390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1614_
timestamp 0
transform 1 0 2230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1615_
timestamp 0
transform 1 0 2530 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1616_
timestamp 0
transform -1 0 3990 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1617_
timestamp 0
transform -1 0 4010 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1618_
timestamp 0
transform 1 0 4130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1619_
timestamp 0
transform 1 0 4490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1620_
timestamp 0
transform 1 0 4650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1621_
timestamp 0
transform -1 0 5390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1622_
timestamp 0
transform 1 0 3970 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1623_
timestamp 0
transform -1 0 3590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1624_
timestamp 0
transform -1 0 3870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1625_
timestamp 0
transform -1 0 4150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1626_
timestamp 0
transform 1 0 3850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1627_
timestamp 0
transform -1 0 4010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1628_
timestamp 0
transform -1 0 4110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1629_
timestamp 0
transform 1 0 4090 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1630_
timestamp 0
transform -1 0 2110 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1631_
timestamp 0
transform -1 0 570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1632_
timestamp 0
transform -1 0 1190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1633_
timestamp 0
transform 1 0 1990 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1634_
timestamp 0
transform 1 0 1990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1635_
timestamp 0
transform 1 0 2390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1636_
timestamp 0
transform 1 0 2290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1637_
timestamp 0
transform 1 0 2730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1638_
timestamp 0
transform 1 0 2150 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1639_
timestamp 0
transform 1 0 2430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1641_
timestamp 0
transform 1 0 3850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1642_
timestamp 0
transform 1 0 4350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1643_
timestamp 0
transform -1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1644_
timestamp 0
transform -1 0 4270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1645_
timestamp 0
transform 1 0 3530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1646_
timestamp 0
transform 1 0 3670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1647_
timestamp 0
transform -1 0 4210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1648_
timestamp 0
transform -1 0 5290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1649_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1650_
timestamp 0
transform 1 0 3010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1651_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1652_
timestamp 0
transform 1 0 3170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1653_
timestamp 0
transform -1 0 2590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1654_
timestamp 0
transform 1 0 3310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1655_
timestamp 0
transform 1 0 3550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1656_
timestamp 0
transform 1 0 1990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1657_
timestamp 0
transform 1 0 1070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 1270 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1659_
timestamp 0
transform 1 0 1130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1660_
timestamp 0
transform -1 0 1090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1661_
timestamp 0
transform -1 0 1710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1662_
timestamp 0
transform 1 0 1590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1663_
timestamp 0
transform 1 0 1290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1664_
timestamp 0
transform -1 0 1450 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1665_
timestamp 0
transform -1 0 1870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1666_
timestamp 0
transform 1 0 1610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1667_
timestamp 0
transform -1 0 1330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1668_
timestamp 0
transform 1 0 1470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1669_
timestamp 0
transform 1 0 2550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1670_
timestamp 0
transform 1 0 2830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1671_
timestamp 0
transform 1 0 2970 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1672_
timestamp 0
transform -1 0 3790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1673_
timestamp 0
transform 1 0 1290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1674_
timestamp 0
transform 1 0 2710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1675_
timestamp 0
transform 1 0 930 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1676_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1677_
timestamp 0
transform 1 0 530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1678_
timestamp 0
transform -1 0 770 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1679_
timestamp 0
transform 1 0 1730 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1680_
timestamp 0
transform -1 0 1190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1681_
timestamp 0
transform 1 0 730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1682_
timestamp 0
transform 1 0 890 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1683_
timestamp 0
transform 1 0 410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1684_
timestamp 0
transform -1 0 810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1685_
timestamp 0
transform 1 0 630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1686_
timestamp 0
transform 1 0 570 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1687_
timestamp 0
transform -1 0 1350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1688_
timestamp 0
transform 1 0 3110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1689_
timestamp 0
transform 1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1690_
timestamp 0
transform 1 0 3410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1691_
timestamp 0
transform 1 0 5130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1692_
timestamp 0
transform -1 0 570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1693_
timestamp 0
transform -1 0 170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1694_
timestamp 0
transform -1 0 270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1695_
timestamp 0
transform 1 0 250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1696_
timestamp 0
transform 1 0 670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1698_
timestamp 0
transform 1 0 150 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1699_
timestamp 0
transform 1 0 390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1700_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1701_
timestamp 0
transform -1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1702_
timestamp 0
transform -1 0 930 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1703_
timestamp 0
transform 1 0 1030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1704_
timestamp 0
transform -1 0 1210 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1705_
timestamp 0
transform -1 0 2430 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1706_
timestamp 0
transform -1 0 1790 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1707_
timestamp 0
transform 1 0 1030 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1708_
timestamp 0
transform -1 0 3470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1709_
timestamp 0
transform -1 0 3770 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1710_
timestamp 0
transform -1 0 3630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1711_
timestamp 0
transform 1 0 1470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1712_
timestamp 0
transform 1 0 1630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1713_
timestamp 0
transform 1 0 1530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1714_
timestamp 0
transform 1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1715_
timestamp 0
transform -1 0 4290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1716_
timestamp 0
transform 1 0 5250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1717_
timestamp 0
transform -1 0 1190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1718_
timestamp 0
transform 1 0 270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1719_
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1721_
timestamp 0
transform -1 0 430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1722_
timestamp 0
transform 1 0 1930 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 2050 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1724_
timestamp 0
transform -1 0 1410 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1725_
timestamp 0
transform 1 0 1670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1726_
timestamp 0
transform 1 0 2270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1727_
timestamp 0
transform -1 0 4910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1808_
timestamp 0
transform -1 0 4990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1809_
timestamp 0
transform -1 0 5370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1810_
timestamp 0
transform 1 0 2230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1811_
timestamp 0
transform 1 0 4350 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1812_
timestamp 0
transform 1 0 5710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 5610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1814_
timestamp 0
transform 1 0 5810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 5790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 3290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform -1 0 930 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 1790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform -1 0 950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform 1 0 3250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform -1 0 3210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 1610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 4770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 4710 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 5550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform -1 0 5370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 5390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 2070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform -1 0 1230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform 1 0 2650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform 1 0 2930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 1130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 5010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform -1 0 4830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform 1 0 2370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform -1 0 2290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert29
timestamp 0
transform -1 0 4590 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert30
timestamp 0
transform -1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform -1 0 1830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert32
timestamp 0
transform 1 0 3110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert33
timestamp 0
transform 1 0 2770 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert34
timestamp 0
transform 1 0 4590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert35
timestamp 0
transform -1 0 4710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert36
timestamp 0
transform 1 0 5150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert37
timestamp 0
transform 1 0 5110 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert38
timestamp 0
transform 1 0 5230 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert39
timestamp 0
transform -1 0 1290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert40
timestamp 0
transform 1 0 2390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert41
timestamp 0
transform 1 0 3550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert42
timestamp 0
transform -1 0 1270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert43
timestamp 0
transform 1 0 2510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert44
timestamp 0
transform -1 0 1430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert45
timestamp 0
transform 1 0 1550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert46
timestamp 0
transform -1 0 1690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert47
timestamp 0
transform 1 0 3330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert48
timestamp 0
transform -1 0 1570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert49
timestamp 0
transform 1 0 3310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert50
timestamp 0
transform -1 0 2350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert51
timestamp 0
transform 1 0 3190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert52
timestamp 0
transform 1 0 2590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert53
timestamp 0
transform -1 0 1870 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert54
timestamp 0
transform -1 0 530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert55
timestamp 0
transform 1 0 3070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert56
timestamp 0
transform -1 0 550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert57
timestamp 0
transform -1 0 990 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert58
timestamp 0
transform -1 0 2950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert12
timestamp 0
transform -1 0 5650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert13
timestamp 0
transform 1 0 630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert14
timestamp 0
transform -1 0 5630 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert15
timestamp 0
transform -1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert16
timestamp 0
transform -1 0 2050 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert17
timestamp 0
transform -1 0 2930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert18
timestamp 0
transform -1 0 5670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert19
timestamp 0
transform -1 0 5630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__863_
timestamp 0
transform 1 0 5090 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__864_
timestamp 0
transform -1 0 4890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__865_
timestamp 0
transform 1 0 5350 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__866_
timestamp 0
transform -1 0 5390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__867_
timestamp 0
transform 1 0 5270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__868_
timestamp 0
transform -1 0 4390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__869_
timestamp 0
transform -1 0 5190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__870_
timestamp 0
transform 1 0 5510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__871_
timestamp 0
transform -1 0 5090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__872_
timestamp 0
transform 1 0 5490 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__873_
timestamp 0
transform 1 0 5730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__874_
timestamp 0
transform 1 0 5770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__875_
timestamp 0
transform -1 0 5450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__876_
timestamp 0
transform 1 0 5310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__877_
timestamp 0
transform -1 0 5170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__878_
timestamp 0
transform -1 0 5230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__879_
timestamp 0
transform 1 0 5170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__880_
timestamp 0
transform -1 0 5110 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__881_
timestamp 0
transform -1 0 5250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__882_
timestamp 0
transform 1 0 3370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__883_
timestamp 0
transform 1 0 3750 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__884_
timestamp 0
transform 1 0 3610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__885_
timestamp 0
transform 1 0 5370 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__886_
timestamp 0
transform 1 0 5430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__887_
timestamp 0
transform -1 0 5550 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__888_
timestamp 0
transform 1 0 5290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__889_
timestamp 0
transform -1 0 4850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__890_
timestamp 0
transform -1 0 4970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__891_
timestamp 0
transform 1 0 5770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__892_
timestamp 0
transform -1 0 4810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__893_
timestamp 0
transform 1 0 5130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__894_
timestamp 0
transform 1 0 5370 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__895_
timestamp 0
transform -1 0 5530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__896_
timestamp 0
transform -1 0 5710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__897_
timestamp 0
transform 1 0 5450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__898_
timestamp 0
transform -1 0 4950 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__899_
timestamp 0
transform 1 0 5230 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__900_
timestamp 0
transform 1 0 5090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__901_
timestamp 0
transform -1 0 5610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__902_
timestamp 0
transform 1 0 5810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__903_
timestamp 0
transform 1 0 5430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__904_
timestamp 0
transform 1 0 5530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__905_
timestamp 0
transform 1 0 5670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__906_
timestamp 0
transform 1 0 5670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__907_
timestamp 0
transform 1 0 1870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__908_
timestamp 0
transform -1 0 1270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__909_
timestamp 0
transform 1 0 1890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__910_
timestamp 0
transform 1 0 1630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__911_
timestamp 0
transform 1 0 2810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__912_
timestamp 0
transform -1 0 2430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__913_
timestamp 0
transform 1 0 2730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__914_
timestamp 0
transform -1 0 4350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__915_
timestamp 0
transform 1 0 4290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__916_
timestamp 0
transform 1 0 1230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__917_
timestamp 0
transform -1 0 1470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__918_
timestamp 0
transform 1 0 1730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__919_
timestamp 0
transform 1 0 1130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__920_
timestamp 0
transform -1 0 2170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__921_
timestamp 0
transform -1 0 2270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__922_
timestamp 0
transform -1 0 2590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__923_
timestamp 0
transform -1 0 4530 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__924_
timestamp 0
transform 1 0 4510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__925_
timestamp 0
transform -1 0 5590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__926_
timestamp 0
transform -1 0 4350 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__927_
timestamp 0
transform 1 0 1030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__928_
timestamp 0
transform -1 0 2990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__929_
timestamp 0
transform -1 0 2930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__930_
timestamp 0
transform -1 0 3050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__931_
timestamp 0
transform 1 0 4050 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__932_
timestamp 0
transform -1 0 3970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__933_
timestamp 0
transform -1 0 4010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__934_
timestamp 0
transform 1 0 3050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__935_
timestamp 0
transform 1 0 1250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__936_
timestamp 0
transform -1 0 1070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__937_
timestamp 0
transform -1 0 1210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__938_
timestamp 0
transform 1 0 2170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__939_
timestamp 0
transform 1 0 1970 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__940_
timestamp 0
transform 1 0 1830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__941_
timestamp 0
transform 1 0 1470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__942_
timestamp 0
transform -1 0 2990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__943_
timestamp 0
transform -1 0 4270 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__944_
timestamp 0
transform -1 0 4130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__945_
timestamp 0
transform -1 0 4530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__946_
timestamp 0
transform 1 0 1810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__947_
timestamp 0
transform -1 0 2230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__948_
timestamp 0
transform 1 0 2310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__949_
timestamp 0
transform -1 0 1010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__950_
timestamp 0
transform 1 0 4370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__951_
timestamp 0
transform -1 0 5450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__952_
timestamp 0
transform -1 0 5470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__953_
timestamp 0
transform 1 0 5550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__954_
timestamp 0
transform -1 0 4090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__955_
timestamp 0
transform 1 0 3450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__956_
timestamp 0
transform 1 0 3490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__957_
timestamp 0
transform -1 0 2990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__958_
timestamp 0
transform -1 0 3790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__959_
timestamp 0
transform 1 0 2810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__960_
timestamp 0
transform -1 0 1110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__961_
timestamp 0
transform -1 0 2090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__962_
timestamp 0
transform 1 0 1410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__963_
timestamp 0
transform -1 0 2810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__964_
timestamp 0
transform 1 0 4090 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__965_
timestamp 0
transform 1 0 1650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__966_
timestamp 0
transform -1 0 2430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__967_
timestamp 0
transform 1 0 2290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__968_
timestamp 0
transform -1 0 2330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__969_
timestamp 0
transform -1 0 4210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__970_
timestamp 0
transform 1 0 3570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__971_
timestamp 0
transform -1 0 3710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__972_
timestamp 0
transform 1 0 2870 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__973_
timestamp 0
transform 1 0 1090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__974_
timestamp 0
transform -1 0 930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__975_
timestamp 0
transform -1 0 1070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__976_
timestamp 0
transform -1 0 1990 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__977_
timestamp 0
transform 1 0 1430 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__978_
timestamp 0
transform -1 0 1710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__979_
timestamp 0
transform 1 0 1770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__980_
timestamp 0
transform 1 0 3130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__981_
timestamp 0
transform 1 0 3250 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__982_
timestamp 0
transform -1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__983_
timestamp 0
transform -1 0 3610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__984_
timestamp 0
transform 1 0 2510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__985_
timestamp 0
transform 1 0 870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__986_
timestamp 0
transform -1 0 1650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__987_
timestamp 0
transform 1 0 1610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__988_
timestamp 0
transform -1 0 2510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__989_
timestamp 0
transform -1 0 3450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__990_
timestamp 0
transform 1 0 4250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__991_
timestamp 0
transform 1 0 4670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__992_
timestamp 0
transform 1 0 4390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__993_
timestamp 0
transform 1 0 4790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__994_
timestamp 0
transform 1 0 4810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__995_
timestamp 0
transform 1 0 4930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__996_
timestamp 0
transform 1 0 4970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__997_
timestamp 0
transform 1 0 5230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__998_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__999_
timestamp 0
transform -1 0 3990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1000_
timestamp 0
transform 1 0 4110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 3590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1002_
timestamp 0
transform 1 0 3710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1003_
timestamp 0
transform -1 0 3870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1004_
timestamp 0
transform 1 0 3670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1005_
timestamp 0
transform 1 0 3690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1006_
timestamp 0
transform 1 0 2510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1007_
timestamp 0
transform 1 0 2370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1008_
timestamp 0
transform 1 0 2230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1009_
timestamp 0
transform -1 0 3470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 3210 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1011_
timestamp 0
transform 1 0 3050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1012_
timestamp 0
transform 1 0 2190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 3330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1014_
timestamp 0
transform 1 0 3470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 3830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1016_
timestamp 0
transform -1 0 3490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1017_
timestamp 0
transform 1 0 3510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1018_
timestamp 0
transform 1 0 4170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1019_
timestamp 0
transform 1 0 4330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1020_
timestamp 0
transform 1 0 5030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1021_
timestamp 0
transform 1 0 4030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1022_
timestamp 0
transform 1 0 4370 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 3490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1024_
timestamp 0
transform -1 0 3530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1025_
timestamp 0
transform -1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1026_
timestamp 0
transform 1 0 4110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 3490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1028_
timestamp 0
transform 1 0 2850 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1029_
timestamp 0
transform -1 0 1510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 1770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 3130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1032_
timestamp 0
transform -1 0 2510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1033_
timestamp 0
transform -1 0 2650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 1930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1035_
timestamp 0
transform -1 0 3410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1036_
timestamp 0
transform 1 0 4030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1037_
timestamp 0
transform -1 0 3790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1038_
timestamp 0
transform 1 0 3870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 4450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 4170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 4310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 3830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1044_
timestamp 0
transform -1 0 4090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1045_
timestamp 0
transform -1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1046_
timestamp 0
transform 1 0 4170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1048_
timestamp 0
transform 1 0 4270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 4170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 3630 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1051_
timestamp 0
transform 1 0 730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 1230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1053_
timestamp 0
transform -1 0 1370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 1930 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1055_
timestamp 0
transform 1 0 1770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 2310 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 2370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1058_
timestamp 0
transform 1 0 2670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1059_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 3090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1061_
timestamp 0
transform 1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 2650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1063_
timestamp 0
transform -1 0 3630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 3890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1065_
timestamp 0
transform -1 0 3350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 3450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1067_
timestamp 0
transform 1 0 3750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1068_
timestamp 0
transform -1 0 3450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1069_
timestamp 0
transform -1 0 3630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 3690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1071_
timestamp 0
transform 1 0 3730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1072_
timestamp 0
transform 1 0 3970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 4070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1074_
timestamp 0
transform 1 0 3870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1075_
timestamp 0
transform -1 0 4410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 3570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1077_
timestamp 0
transform 1 0 3150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 2710 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1080_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1081_
timestamp 0
transform -1 0 890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 1350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1083_
timestamp 0
transform 1 0 930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1084_
timestamp 0
transform -1 0 2510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 3230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1086_
timestamp 0
transform 1 0 2610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1087_
timestamp 0
transform 1 0 2230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 2430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1089_
timestamp 0
transform -1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 2330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 2190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 2510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1093_
timestamp 0
transform 1 0 2830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1094_
timestamp 0
transform -1 0 2370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 2930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1096_
timestamp 0
transform 1 0 3430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1097_
timestamp 0
transform -1 0 3210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1098_
timestamp 0
transform 1 0 3590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 4510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1100_
timestamp 0
transform -1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 2590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1102_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1103_
timestamp 0
transform -1 0 450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1104_
timestamp 0
transform -1 0 830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 1090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1106_
timestamp 0
transform -1 0 1350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1108_
timestamp 0
transform -1 0 1710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1109_
timestamp 0
transform 1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1110_
timestamp 0
transform 1 0 1930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 1610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1112_
timestamp 0
transform 1 0 1790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1113_
timestamp 0
transform -1 0 2170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1114_
timestamp 0
transform 1 0 2030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 1890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1116_
timestamp 0
transform -1 0 1630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1117_
timestamp 0
transform 1 0 1750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 2130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1119_
timestamp 0
transform -1 0 2010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1120_
timestamp 0
transform 1 0 2270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 2290 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1122_
timestamp 0
transform 1 0 1850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 1270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 1550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1125_
timestamp 0
transform -1 0 910 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1126_
timestamp 0
transform -1 0 410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1129_
timestamp 0
transform -1 0 1030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 1670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1131_
timestamp 0
transform 1 0 1390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1132_
timestamp 0
transform -1 0 1510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1133_
timestamp 0
transform 1 0 1830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1134_
timestamp 0
transform -1 0 1490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 1390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1136_
timestamp 0
transform 1 0 1330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1137_
timestamp 0
transform 1 0 1630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1138_
timestamp 0
transform 1 0 1650 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1139_
timestamp 0
transform 1 0 1910 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1140_
timestamp 0
transform -1 0 1790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1141_
timestamp 0
transform -1 0 1990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 1070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1143_
timestamp 0
transform -1 0 1010 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1144_
timestamp 0
transform 1 0 650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1145_
timestamp 0
transform 1 0 1710 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1147_
timestamp 0
transform 1 0 890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1148_
timestamp 0
transform -1 0 1110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1149_
timestamp 0
transform -1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 1090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1151_
timestamp 0
transform -1 0 1230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1152_
timestamp 0
transform 1 0 830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1153_
timestamp 0
transform -1 0 1130 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1154_
timestamp 0
transform -1 0 1510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1155_
timestamp 0
transform -1 0 1550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1156_
timestamp 0
transform -1 0 1270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 1410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 1350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 1210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1160_
timestamp 0
transform 1 0 1250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1161_
timestamp 0
transform 1 0 1390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 1550 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 1590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1164_
timestamp 0
transform -1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1165_
timestamp 0
transform 1 0 850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1166_
timestamp 0
transform -1 0 1250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1167_
timestamp 0
transform 1 0 290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1168_
timestamp 0
transform -1 0 330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1170_
timestamp 0
transform -1 0 330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1171_
timestamp 0
transform -1 0 950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1174_
timestamp 0
transform -1 0 550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1176_
timestamp 0
transform -1 0 810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1177_
timestamp 0
transform 1 0 890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1178_
timestamp 0
transform 1 0 970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1179_
timestamp 0
transform 1 0 1110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1180_
timestamp 0
transform -1 0 1070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1182_
timestamp 0
transform 1 0 770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1183_
timestamp 0
transform -1 0 630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1184_
timestamp 0
transform -1 0 1070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1185_
timestamp 0
transform 1 0 330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1186_
timestamp 0
transform -1 0 770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1188_
timestamp 0
transform -1 0 50 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1191_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1192_
timestamp 0
transform -1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1193_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1194_
timestamp 0
transform -1 0 170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1195_
timestamp 0
transform -1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1197_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1198_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1199_
timestamp 0
transform 1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1200_
timestamp 0
transform -1 0 190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1201_
timestamp 0
transform -1 0 50 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1204_
timestamp 0
transform 1 0 370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1205_
timestamp 0
transform -1 0 150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 1370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 50 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1212_
timestamp 0
transform 1 0 330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1215_
timestamp 0
transform -1 0 350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1216_
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1217_
timestamp 0
transform -1 0 50 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1218_
timestamp 0
transform 1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1219_
timestamp 0
transform -1 0 50 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 150 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 370 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1223_
timestamp 0
transform -1 0 1130 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1224_
timestamp 0
transform -1 0 730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1226_
timestamp 0
transform -1 0 50 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1228_
timestamp 0
transform 1 0 730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1230_
timestamp 0
transform -1 0 410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1231_
timestamp 0
transform -1 0 570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1234_
timestamp 0
transform 1 0 810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1235_
timestamp 0
transform 1 0 590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1236_
timestamp 0
transform -1 0 470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1237_
timestamp 0
transform -1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1238_
timestamp 0
transform -1 0 50 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1239_
timestamp 0
transform 1 0 190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1240_
timestamp 0
transform 1 0 470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1241_
timestamp 0
transform -1 0 490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1243_
timestamp 0
transform 1 0 630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1245_
timestamp 0
transform -1 0 770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1246_
timestamp 0
transform -1 0 1510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1247_
timestamp 0
transform 1 0 270 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1248_
timestamp 0
transform -1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 50 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1250_
timestamp 0
transform -1 0 190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1254_
timestamp 0
transform 1 0 770 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1255_
timestamp 0
transform -1 0 870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1256_
timestamp 0
transform 1 0 570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1258_
timestamp 0
transform -1 0 770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1259_
timestamp 0
transform -1 0 910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1260_
timestamp 0
transform 1 0 4790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1261_
timestamp 0
transform 1 0 4270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1262_
timestamp 0
transform -1 0 2470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 3670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1264_
timestamp 0
transform 1 0 4910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1265_
timestamp 0
transform 1 0 4610 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 4750 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 5290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1268_
timestamp 0
transform 1 0 5150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1269_
timestamp 0
transform 1 0 5550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1270_
timestamp 0
transform -1 0 2110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1271_
timestamp 0
transform -1 0 3610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1272_
timestamp 0
transform -1 0 3230 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1273_
timestamp 0
transform -1 0 3870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1274_
timestamp 0
transform 1 0 3990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1275_
timestamp 0
transform 1 0 5450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 5350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 5590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1278_
timestamp 0
transform -1 0 5750 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1279_
timestamp 0
transform 1 0 5770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 5790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 5710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1282_
timestamp 0
transform -1 0 5270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 5810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 5750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 4030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1286_
timestamp 0
transform 1 0 4610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 4770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1288_
timestamp 0
transform 1 0 5590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1289_
timestamp 0
transform 1 0 5530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1290_
timestamp 0
transform 1 0 5730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1291_
timestamp 0
transform -1 0 5510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1292_
timestamp 0
transform 1 0 5830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 5610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1294_
timestamp 0
transform 1 0 5730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1295_
timestamp 0
transform -1 0 5630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 5610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 5490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1298_
timestamp 0
transform 1 0 4830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1299_
timestamp 0
transform -1 0 3850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 3910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1301_
timestamp 0
transform -1 0 4330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1302_
timestamp 0
transform 1 0 4450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1303_
timestamp 0
transform 1 0 5050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1304_
timestamp 0
transform -1 0 4950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1305_
timestamp 0
transform 1 0 4970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 5090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1307_
timestamp 0
transform 1 0 5230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 5330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1309_
timestamp 0
transform -1 0 5150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1310_
timestamp 0
transform -1 0 4930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1311_
timestamp 0
transform -1 0 5050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1312_
timestamp 0
transform 1 0 4250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 3170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1314_
timestamp 0
transform 1 0 3190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1315_
timestamp 0
transform -1 0 3090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 2650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 2550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1319_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 4850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1321_
timestamp 0
transform 1 0 2810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 2690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 2950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1324_
timestamp 0
transform -1 0 2530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1325_
timestamp 0
transform 1 0 3330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 3010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1327_
timestamp 0
transform -1 0 2570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1328_
timestamp 0
transform -1 0 3450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 3350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 2530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 2570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1332_
timestamp 0
transform -1 0 2310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1333_
timestamp 0
transform -1 0 2010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1334_
timestamp 0
transform 1 0 2150 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1335_
timestamp 0
transform -1 0 1910 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1336_
timestamp 0
transform -1 0 2270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1337_
timestamp 0
transform 1 0 2410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 2430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1339_
timestamp 0
transform 1 0 2510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1340_
timestamp 0
transform 1 0 2450 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1341_
timestamp 0
transform -1 0 2390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 2630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 2710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1344_
timestamp 0
transform 1 0 2530 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 3190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1346_
timestamp 0
transform -1 0 3390 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 3570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1348_
timestamp 0
transform 1 0 3710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 3430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1350_
timestamp 0
transform 1 0 3310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1351_
timestamp 0
transform -1 0 3070 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 3290 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1353_
timestamp 0
transform 1 0 3310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1354_
timestamp 0
transform 1 0 4490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 4630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1356_
timestamp 0
transform -1 0 4930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 3250 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 4370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1360_
timestamp 0
transform -1 0 4530 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1361_
timestamp 0
transform 1 0 4210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1362_
timestamp 0
transform 1 0 3850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1363_
timestamp 0
transform -1 0 2990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1364_
timestamp 0
transform -1 0 3750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 3390 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 3390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1367_
timestamp 0
transform 1 0 3290 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 3170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1369_
timestamp 0
transform -1 0 3450 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1370_
timestamp 0
transform 1 0 4750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1371_
timestamp 0
transform 1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 4190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 3970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1374_
timestamp 0
transform 1 0 3830 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1375_
timestamp 0
transform 1 0 4050 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 4170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 3910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 3750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 3110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1380_
timestamp 0
transform -1 0 3230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1381_
timestamp 0
transform -1 0 3130 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 3070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 2850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1384_
timestamp 0
transform 1 0 2970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1385_
timestamp 0
transform 1 0 3830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1386_
timestamp 0
transform 1 0 3950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1387_
timestamp 0
transform 1 0 4070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 4210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1389_
timestamp 0
transform -1 0 4750 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1390_
timestamp 0
transform 1 0 3470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1391_
timestamp 0
transform -1 0 3590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1392_
timestamp 0
transform -1 0 2910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1393_
timestamp 0
transform -1 0 3150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 3010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1395_
timestamp 0
transform 1 0 3250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1396_
timestamp 0
transform 1 0 4290 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1397_
timestamp 0
transform 1 0 4430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 4590 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1399_
timestamp 0
transform -1 0 3390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1400_
timestamp 0
transform 1 0 4130 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 4050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1402_
timestamp 0
transform 1 0 3890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 3510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 3670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 3530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1406_
timestamp 0
transform -1 0 3790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 4210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 4350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1409_
timestamp 0
transform -1 0 4450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 4830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1411_
timestamp 0
transform -1 0 4070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 4670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1413_
timestamp 0
transform -1 0 4870 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 4730 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1415_
timestamp 0
transform 1 0 830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1417_
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1419_
timestamp 0
transform 1 0 5410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1420_
timestamp 0
transform -1 0 5290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1423_
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1424_
timestamp 0
transform -1 0 50 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 4890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 1510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1427_
timestamp 0
transform 1 0 1350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1428_
timestamp 0
transform -1 0 1350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 1190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1430_
timestamp 0
transform 1 0 3970 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 2210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 2250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 1830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1434_
timestamp 0
transform -1 0 1970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1435_
timestamp 0
transform -1 0 2710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1436_
timestamp 0
transform -1 0 2830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 2830 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1438_
timestamp 0
transform 1 0 2690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1439_
timestamp 0
transform -1 0 4650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1440_
timestamp 0
transform 1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1441_
timestamp 0
transform -1 0 4330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1442_
timestamp 0
transform -1 0 4470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1443_
timestamp 0
transform -1 0 210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1445_
timestamp 0
transform -1 0 470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1446_
timestamp 0
transform 1 0 310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1447_
timestamp 0
transform 1 0 1190 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 1070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1449_
timestamp 0
transform -1 0 1090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1450_
timestamp 0
transform 1 0 930 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1451_
timestamp 0
transform 1 0 790 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1452_
timestamp 0
transform -1 0 1990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1453_
timestamp 0
transform -1 0 2130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1454_
timestamp 0
transform 1 0 2930 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1455_
timestamp 0
transform 1 0 2770 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1456_
timestamp 0
transform -1 0 3410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1457_
timestamp 0
transform 1 0 3330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1458_
timestamp 0
transform 1 0 3970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1459_
timestamp 0
transform 1 0 3830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 4610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1461_
timestamp 0
transform 1 0 4310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1462_
timestamp 0
transform 1 0 4610 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1463_
timestamp 0
transform 1 0 4470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1464_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 4430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1466_
timestamp 0
transform -1 0 4250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1467_
timestamp 0
transform -1 0 4210 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1468_
timestamp 0
transform -1 0 2710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1469_
timestamp 0
transform -1 0 3490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1470_
timestamp 0
transform -1 0 1370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1471_
timestamp 0
transform -1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1472_
timestamp 0
transform -1 0 3510 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1473_
timestamp 0
transform -1 0 4130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1474_
timestamp 0
transform -1 0 2790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1475_
timestamp 0
transform -1 0 2830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1476_
timestamp 0
transform -1 0 2670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1477_
timestamp 0
transform -1 0 2790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1478_
timestamp 0
transform -1 0 4570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1479_
timestamp 0
transform -1 0 3950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1480_
timestamp 0
transform -1 0 4410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 2450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1482_
timestamp 0
transform -1 0 2430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1483_
timestamp 0
transform 1 0 1910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 1790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1485_
timestamp 0
transform 1 0 5030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1486_
timestamp 0
transform 1 0 4790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1487_
timestamp 0
transform 1 0 5210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1488_
timestamp 0
transform 1 0 5070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1489_
timestamp 0
transform -1 0 4930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1490_
timestamp 0
transform 1 0 4650 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 4350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1492_
timestamp 0
transform -1 0 4490 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1493_
timestamp 0
transform -1 0 5310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1494_
timestamp 0
transform -1 0 5430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1495_
timestamp 0
transform 1 0 2150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1496_
timestamp 0
transform -1 0 790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1497_
timestamp 0
transform -1 0 1770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1498_
timestamp 0
transform -1 0 5030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1499_
timestamp 0
transform 1 0 4530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1500_
timestamp 0
transform -1 0 2990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1501_
timestamp 0
transform -1 0 570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1502_
timestamp 0
transform -1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1503_
timestamp 0
transform -1 0 2150 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1504_
timestamp 0
transform -1 0 2070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1505_
timestamp 0
transform 1 0 3110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1506_
timestamp 0
transform 1 0 2790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1507_
timestamp 0
transform -1 0 2590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1508_
timestamp 0
transform 1 0 2630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1509_
timestamp 0
transform 1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1510_
timestamp 0
transform 1 0 2490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1511_
timestamp 0
transform -1 0 1950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1512_
timestamp 0
transform -1 0 2070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1513_
timestamp 0
transform -1 0 1910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1514_
timestamp 0
transform -1 0 1470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1515_
timestamp 0
transform 1 0 1750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1516_
timestamp 0
transform 1 0 2350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1517_
timestamp 0
transform 1 0 2630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1518_
timestamp 0
transform -1 0 2230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1519_
timestamp 0
transform 1 0 1930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1520_
timestamp 0
transform 1 0 1650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1521_
timestamp 0
transform -1 0 2090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1522_
timestamp 0
transform 1 0 2030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1523_
timestamp 0
transform 1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1524_
timestamp 0
transform -1 0 3310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1525_
timestamp 0
transform 1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1526_
timestamp 0
transform -1 0 3690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 4870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 4970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1529_
timestamp 0
transform -1 0 5090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 5330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 5130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1532_
timestamp 0
transform -1 0 5210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1533_
timestamp 0
transform 1 0 3810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1534_
timestamp 0
transform -1 0 5150 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 5690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1536_
timestamp 0
transform 1 0 5110 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1537_
timestamp 0
transform 1 0 4730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1538_
timestamp 0
transform 1 0 4810 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1539_
timestamp 0
transform -1 0 2830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1540_
timestamp 0
transform 1 0 570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1541_
timestamp 0
transform 1 0 410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1542_
timestamp 0
transform -1 0 1510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1543_
timestamp 0
transform -1 0 1570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1544_
timestamp 0
transform -1 0 1970 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1545_
timestamp 0
transform -1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1546_
timestamp 0
transform 1 0 1610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1547_
timestamp 0
transform 1 0 2510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1548_
timestamp 0
transform -1 0 2310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1549_
timestamp 0
transform -1 0 290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1550_
timestamp 0
transform -1 0 410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1551_
timestamp 0
transform 1 0 1350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1552_
timestamp 0
transform 1 0 1210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1553_
timestamp 0
transform 1 0 1850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1554_
timestamp 0
transform -1 0 2170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1555_
timestamp 0
transform 1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1556_
timestamp 0
transform 1 0 4990 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1557_
timestamp 0
transform 1 0 5110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1558_
timestamp 0
transform 1 0 5230 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1559_
timestamp 0
transform 1 0 5350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1560_
timestamp 0
transform 1 0 5470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1561_
timestamp 0
transform 1 0 5610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1562_
timestamp 0
transform -1 0 5530 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 2030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1564_
timestamp 0
transform -1 0 410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1565_
timestamp 0
transform -1 0 550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1566_
timestamp 0
transform -1 0 710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1567_
timestamp 0
transform -1 0 850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1568_
timestamp 0
transform -1 0 990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1569_
timestamp 0
transform -1 0 1470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1570_
timestamp 0
transform 1 0 2970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1571_
timestamp 0
transform -1 0 2410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1572_
timestamp 0
transform -1 0 2990 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1573_
timestamp 0
transform 1 0 2830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1574_
timestamp 0
transform 1 0 3370 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1575_
timestamp 0
transform -1 0 3530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1576_
timestamp 0
transform 1 0 3230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1577_
timestamp 0
transform 1 0 3630 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1578_
timestamp 0
transform 1 0 4270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1579_
timestamp 0
transform -1 0 4810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 4830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1581_
timestamp 0
transform 1 0 4410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1582_
timestamp 0
transform -1 0 4570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 4630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1584_
timestamp 0
transform -1 0 4710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1585_
timestamp 0
transform 1 0 4690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1586_
timestamp 0
transform -1 0 690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1587_
timestamp 0
transform 1 0 970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1588_
timestamp 0
transform 1 0 1710 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1589_
timestamp 0
transform 1 0 1550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1590_
timestamp 0
transform 1 0 2130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1591_
timestamp 0
transform -1 0 3110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1592_
timestamp 0
transform 1 0 2950 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1593_
timestamp 0
transform 1 0 3770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1594_
timestamp 0
transform 1 0 3090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1595_
timestamp 0
transform 1 0 3730 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1596_
timestamp 0
transform -1 0 3410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1597_
timestamp 0
transform -1 0 3250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1598_
timestamp 0
transform 1 0 4430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1599_
timestamp 0
transform 1 0 4730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1600_
timestamp 0
transform 1 0 4570 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1601_
timestamp 0
transform 1 0 4870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1602_
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1603_
timestamp 0
transform -1 0 5430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1604_
timestamp 0
transform -1 0 2710 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1606_
timestamp 0
transform -1 0 1350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1607_
timestamp 0
transform 1 0 1410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1608_
timestamp 0
transform 1 0 2550 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1609_
timestamp 0
transform 1 0 1910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1610_
timestamp 0
transform 1 0 2150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1611_
timestamp 0
transform 1 0 2250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1612_
timestamp 0
transform 1 0 2710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1613_
timestamp 0
transform 1 0 2410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1614_
timestamp 0
transform 1 0 2250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1615_
timestamp 0
transform 1 0 2550 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1616_
timestamp 0
transform -1 0 4010 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1617_
timestamp 0
transform -1 0 4030 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1618_
timestamp 0
transform 1 0 4150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1619_
timestamp 0
transform 1 0 4510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1620_
timestamp 0
transform 1 0 4670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1621_
timestamp 0
transform -1 0 5410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1622_
timestamp 0
transform 1 0 3990 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1623_
timestamp 0
transform -1 0 3610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1624_
timestamp 0
transform -1 0 3890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1625_
timestamp 0
transform -1 0 4170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1626_
timestamp 0
transform 1 0 3870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1627_
timestamp 0
transform -1 0 4030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1628_
timestamp 0
transform -1 0 4130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1629_
timestamp 0
transform 1 0 4110 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1630_
timestamp 0
transform -1 0 2130 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1631_
timestamp 0
transform -1 0 590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1632_
timestamp 0
transform -1 0 1210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1633_
timestamp 0
transform 1 0 2010 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1634_
timestamp 0
transform 1 0 2010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1635_
timestamp 0
transform 1 0 2410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1636_
timestamp 0
transform 1 0 2310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1637_
timestamp 0
transform 1 0 2750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1638_
timestamp 0
transform 1 0 2170 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1639_
timestamp 0
transform 1 0 2450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 2890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1641_
timestamp 0
transform 1 0 3870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1642_
timestamp 0
transform 1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1643_
timestamp 0
transform -1 0 4270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1644_
timestamp 0
transform -1 0 4290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1645_
timestamp 0
transform 1 0 3550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1646_
timestamp 0
transform 1 0 3690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1647_
timestamp 0
transform -1 0 4230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1648_
timestamp 0
transform -1 0 5310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1649_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1650_
timestamp 0
transform 1 0 3030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1651_
timestamp 0
transform -1 0 3750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1652_
timestamp 0
transform 1 0 3190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1653_
timestamp 0
transform -1 0 2610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1654_
timestamp 0
transform 1 0 3330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1655_
timestamp 0
transform 1 0 3570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1656_
timestamp 0
transform 1 0 2010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1657_
timestamp 0
transform 1 0 1090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1658_
timestamp 0
transform 1 0 1290 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1659_
timestamp 0
transform 1 0 1150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1660_
timestamp 0
transform -1 0 1110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1661_
timestamp 0
transform -1 0 1730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1662_
timestamp 0
transform 1 0 1610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1663_
timestamp 0
transform 1 0 1310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1664_
timestamp 0
transform -1 0 1470 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1665_
timestamp 0
transform -1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1666_
timestamp 0
transform 1 0 1630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1667_
timestamp 0
transform -1 0 1350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1668_
timestamp 0
transform 1 0 1490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1669_
timestamp 0
transform 1 0 2570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1670_
timestamp 0
transform 1 0 2850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1671_
timestamp 0
transform 1 0 2990 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1672_
timestamp 0
transform -1 0 3810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1673_
timestamp 0
transform 1 0 1310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1674_
timestamp 0
transform 1 0 2730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1675_
timestamp 0
transform 1 0 950 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1676_
timestamp 0
transform -1 0 1030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1677_
timestamp 0
transform 1 0 550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1678_
timestamp 0
transform -1 0 790 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1679_
timestamp 0
transform 1 0 1750 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1680_
timestamp 0
transform -1 0 1210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1681_
timestamp 0
transform 1 0 750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1682_
timestamp 0
transform 1 0 910 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1683_
timestamp 0
transform 1 0 430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1684_
timestamp 0
transform -1 0 830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1685_
timestamp 0
transform 1 0 650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1686_
timestamp 0
transform 1 0 590 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1687_
timestamp 0
transform -1 0 1370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1688_
timestamp 0
transform 1 0 3130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1689_
timestamp 0
transform 1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1690_
timestamp 0
transform 1 0 3430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1691_
timestamp 0
transform 1 0 5150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1692_
timestamp 0
transform -1 0 590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1693_
timestamp 0
transform -1 0 190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1694_
timestamp 0
transform -1 0 290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1695_
timestamp 0
transform 1 0 270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1696_
timestamp 0
transform 1 0 690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1697_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1698_
timestamp 0
transform 1 0 170 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1699_
timestamp 0
transform 1 0 410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1700_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1701_
timestamp 0
transform -1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1702_
timestamp 0
transform -1 0 950 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1703_
timestamp 0
transform 1 0 1050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1704_
timestamp 0
transform -1 0 1230 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1705_
timestamp 0
transform -1 0 2450 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1706_
timestamp 0
transform -1 0 1810 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1707_
timestamp 0
transform 1 0 1050 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1708_
timestamp 0
transform -1 0 3490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1709_
timestamp 0
transform -1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1710_
timestamp 0
transform -1 0 3650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1711_
timestamp 0
transform 1 0 1490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1712_
timestamp 0
transform 1 0 1650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1713_
timestamp 0
transform 1 0 1550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1714_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1715_
timestamp 0
transform -1 0 4310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1716_
timestamp 0
transform 1 0 5270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1717_
timestamp 0
transform -1 0 1210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1718_
timestamp 0
transform 1 0 290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1719_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1721_
timestamp 0
transform -1 0 450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1722_
timestamp 0
transform 1 0 1950 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 2070 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1724_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1725_
timestamp 0
transform 1 0 1690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1726_
timestamp 0
transform 1 0 2290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1727_
timestamp 0
transform -1 0 4930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1808_
timestamp 0
transform -1 0 5010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1809_
timestamp 0
transform -1 0 5390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1810_
timestamp 0
transform 1 0 2250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1811_
timestamp 0
transform 1 0 4370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1812_
timestamp 0
transform 1 0 5730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__1813_
timestamp 0
transform 1 0 5630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1814_
timestamp 0
transform 1 0 5830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 5810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 3310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform -1 0 950 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 1810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform -1 0 970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform 1 0 3270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform -1 0 3230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 1630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 4790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 4730 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 5570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform -1 0 5390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 5410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 2090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform -1 0 1250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform 1 0 2670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform 1 0 2950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 5030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform -1 0 4850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform 1 0 2390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform -1 0 2310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert29
timestamp 0
transform -1 0 4610 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert30
timestamp 0
transform -1 0 1850 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert31
timestamp 0
transform -1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert32
timestamp 0
transform 1 0 3130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert33
timestamp 0
transform 1 0 2790 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert34
timestamp 0
transform 1 0 4610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert35
timestamp 0
transform -1 0 4730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert36
timestamp 0
transform 1 0 5170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert37
timestamp 0
transform 1 0 5130 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert38
timestamp 0
transform 1 0 5250 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert39
timestamp 0
transform -1 0 1310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert40
timestamp 0
transform 1 0 2410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert41
timestamp 0
transform 1 0 3570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert42
timestamp 0
transform -1 0 1290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert43
timestamp 0
transform 1 0 2530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert44
timestamp 0
transform -1 0 1450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert45
timestamp 0
transform 1 0 1570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert46
timestamp 0
transform -1 0 1710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert47
timestamp 0
transform 1 0 3350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert48
timestamp 0
transform -1 0 1590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert49
timestamp 0
transform 1 0 3330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert50
timestamp 0
transform -1 0 2370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert51
timestamp 0
transform 1 0 3210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert52
timestamp 0
transform 1 0 2610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert53
timestamp 0
transform -1 0 1890 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert54
timestamp 0
transform -1 0 550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert55
timestamp 0
transform 1 0 3090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert56
timestamp 0
transform -1 0 570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert57
timestamp 0
transform -1 0 1010 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert58
timestamp 0
transform -1 0 2970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert12
timestamp 0
transform -1 0 5670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert13
timestamp 0
transform 1 0 650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert14
timestamp 0
transform -1 0 5650 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert15
timestamp 0
transform -1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert16
timestamp 0
transform -1 0 2070 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert17
timestamp 0
transform -1 0 2950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert18
timestamp 0
transform -1 0 5690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert19
timestamp 0
transform -1 0 5650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__863_
timestamp 0
transform 1 0 5110 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__866_
timestamp 0
transform -1 0 5410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__869_
timestamp 0
transform -1 0 5210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__872_
timestamp 0
transform 1 0 5510 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__874_
timestamp 0
transform 1 0 5790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__877_
timestamp 0
transform -1 0 5190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__880_
timestamp 0
transform -1 0 5130 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__883_
timestamp 0
transform 1 0 3770 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__885_
timestamp 0
transform 1 0 5390 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__888_
timestamp 0
transform 1 0 5310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__891_
timestamp 0
transform 1 0 5790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__894_
timestamp 0
transform 1 0 5390 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__897_
timestamp 0
transform 1 0 5470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__899_
timestamp 0
transform 1 0 5250 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__902_
timestamp 0
transform 1 0 5830 0 1 730
box -6 -8 26 248
use FILL  FILL_2__905_
timestamp 0
transform 1 0 5690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__908_
timestamp 0
transform -1 0 1290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__910_
timestamp 0
transform 1 0 1650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__913_
timestamp 0
transform 1 0 2750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__916_
timestamp 0
transform 1 0 1250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__919_
timestamp 0
transform 1 0 1150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__922_
timestamp 0
transform -1 0 2610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__924_
timestamp 0
transform 1 0 4530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__927_
timestamp 0
transform 1 0 1050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__930_
timestamp 0
transform -1 0 3070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__933_
timestamp 0
transform -1 0 4030 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__936_
timestamp 0
transform -1 0 1090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__938_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__941_
timestamp 0
transform 1 0 1490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__944_
timestamp 0
transform -1 0 4150 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__947_
timestamp 0
transform -1 0 2250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__949_
timestamp 0
transform -1 0 1030 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__952_
timestamp 0
transform -1 0 5490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__955_
timestamp 0
transform 1 0 3470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__958_
timestamp 0
transform -1 0 3810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__961_
timestamp 0
transform -1 0 2110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__963_
timestamp 0
transform -1 0 2830 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__966_
timestamp 0
transform -1 0 2450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__969_
timestamp 0
transform -1 0 4230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__972_
timestamp 0
transform 1 0 2890 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__974_
timestamp 0
transform -1 0 950 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__977_
timestamp 0
transform 1 0 1450 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__980_
timestamp 0
transform 1 0 3150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__983_
timestamp 0
transform -1 0 3630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__986_
timestamp 0
transform -1 0 1670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__988_
timestamp 0
transform -1 0 2530 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__991_
timestamp 0
transform 1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__994_
timestamp 0
transform 1 0 4830 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__997_
timestamp 0
transform 1 0 5250 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1002_
timestamp 0
transform 1 0 3730 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1004_
timestamp 0
transform 1 0 3690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1007_
timestamp 0
transform 1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 3230 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 3350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1016_
timestamp 0
transform -1 0 3510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1018_
timestamp 0
transform 1 0 4190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1021_
timestamp 0
transform 1 0 4050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1024_
timestamp 0
transform -1 0 3550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 3510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1030_
timestamp 0
transform -1 0 1790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1032_
timestamp 0
transform -1 0 2530 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1035_
timestamp 0
transform -1 0 3430 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1038_
timestamp 0
transform 1 0 3890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1041_
timestamp 0
transform 1 0 4190 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 3850 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1046_
timestamp 0
transform 1 0 4190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1049_
timestamp 0
transform -1 0 4190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1052_
timestamp 0
transform -1 0 1250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1055_
timestamp 0
transform 1 0 1790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1057_
timestamp 0
transform 1 0 2390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1060_
timestamp 0
transform -1 0 3110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1063_
timestamp 0
transform -1 0 3650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1066_
timestamp 0
transform 1 0 3470 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1068_
timestamp 0
transform -1 0 3470 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1071_
timestamp 0
transform 1 0 3750 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1074_
timestamp 0
transform 1 0 3890 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1077_
timestamp 0
transform 1 0 3170 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1080_
timestamp 0
transform -1 0 770 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 1370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1085_
timestamp 0
transform -1 0 3250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1088_
timestamp 0
transform -1 0 2450 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1091_
timestamp 0
transform 1 0 2210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1094_
timestamp 0
transform -1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1096_
timestamp 0
transform 1 0 3450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1099_
timestamp 0
transform -1 0 4530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1102_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1105_
timestamp 0
transform -1 0 1110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1110_
timestamp 0
transform 1 0 1950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1113_
timestamp 0
transform -1 0 2190 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1116_
timestamp 0
transform -1 0 1650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1119_
timestamp 0
transform -1 0 2030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 2310 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1124_
timestamp 0
transform 1 0 1570 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1127_
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1130_
timestamp 0
transform 1 0 1690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1132_
timestamp 0
transform -1 0 1530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 1410 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1138_
timestamp 0
transform 1 0 1670 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1141_
timestamp 0
transform -1 0 2010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1144_
timestamp 0
transform 1 0 670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 750 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1149_
timestamp 0
transform -1 0 930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1152_
timestamp 0
transform 1 0 850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1155_
timestamp 0
transform -1 0 1570 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1158_
timestamp 0
transform -1 0 1370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1160_
timestamp 0
transform 1 0 1270 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1163_
timestamp 0
transform -1 0 1610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1166_
timestamp 0
transform -1 0 1270 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1169_
timestamp 0
transform 1 0 610 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1171_
timestamp 0
transform -1 0 970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1174_
timestamp 0
transform -1 0 570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1177_
timestamp 0
transform 1 0 910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1180_
timestamp 0
transform -1 0 1090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1183_
timestamp 0
transform -1 0 650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1185_
timestamp 0
transform 1 0 350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1188_
timestamp 0
transform -1 0 70 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1191_
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1194_
timestamp 0
transform -1 0 190 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1196_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1199_
timestamp 0
transform 1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 330 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1205_
timestamp 0
transform -1 0 170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1208_
timestamp 0
transform -1 0 70 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1216_
timestamp 0
transform 1 0 190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1219_
timestamp 0
transform -1 0 70 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1221_
timestamp 0
transform 1 0 210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1224_
timestamp 0
transform -1 0 750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1227_
timestamp 0
transform 1 0 390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1230_
timestamp 0
transform -1 0 430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1233_
timestamp 0
transform -1 0 190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1235_
timestamp 0
transform 1 0 610 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1238_
timestamp 0
transform -1 0 70 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1241_
timestamp 0
transform -1 0 510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 630 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1247_
timestamp 0
transform 1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1249_
timestamp 0
transform -1 0 70 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1252_
timestamp 0
transform -1 0 970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1255_
timestamp 0
transform -1 0 890 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1258_
timestamp 0
transform -1 0 790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1260_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1263_
timestamp 0
transform -1 0 3690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1266_
timestamp 0
transform 1 0 4770 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1269_
timestamp 0
transform 1 0 5570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1272_
timestamp 0
transform -1 0 3250 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1274_
timestamp 0
transform 1 0 4010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 5610 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1280_
timestamp 0
transform 1 0 5810 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1283_
timestamp 0
transform 1 0 5830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 4050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1288_
timestamp 0
transform 1 0 5610 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1291_
timestamp 0
transform -1 0 5530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1294_
timestamp 0
transform 1 0 5750 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1297_
timestamp 0
transform 1 0 5510 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1299_
timestamp 0
transform -1 0 3870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1302_
timestamp 0
transform 1 0 4470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1305_
timestamp 0
transform 1 0 4990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1308_
timestamp 0
transform 1 0 5350 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1311_
timestamp 0
transform -1 0 5070 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1313_
timestamp 0
transform 1 0 3190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 3070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1319_
timestamp 0
transform -1 0 2930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1322_
timestamp 0
transform -1 0 2710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1324_
timestamp 0
transform -1 0 2550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1327_
timestamp 0
transform -1 0 2590 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 2550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1333_
timestamp 0
transform -1 0 2030 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1336_
timestamp 0
transform -1 0 2290 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 2450 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1341_
timestamp 0
transform -1 0 2410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1344_
timestamp 0
transform 1 0 2550 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 3590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1349_
timestamp 0
transform 1 0 3450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1352_
timestamp 0
transform -1 0 3310 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1355_
timestamp 0
transform 1 0 4650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1358_
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1361_
timestamp 0
transform 1 0 4230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1363_
timestamp 0
transform -1 0 3010 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1366_
timestamp 0
transform -1 0 3410 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1369_
timestamp 0
transform -1 0 3470 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1372_
timestamp 0
transform -1 0 4210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1375_
timestamp 0
transform 1 0 4070 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1377_
timestamp 0
transform -1 0 3930 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1380_
timestamp 0
transform -1 0 3250 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 2870 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1386_
timestamp 0
transform 1 0 3970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 4230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1391_
timestamp 0
transform -1 0 3610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1394_
timestamp 0
transform -1 0 3030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1397_
timestamp 0
transform 1 0 4450 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1400_
timestamp 0
transform 1 0 4150 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1402_
timestamp 0
transform 1 0 3910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1405_
timestamp 0
transform -1 0 3550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 4370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1411_
timestamp 0
transform -1 0 4090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1413_
timestamp 0
transform -1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1416_
timestamp 0
transform 1 0 690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1419_
timestamp 0
transform 1 0 5430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1425_
timestamp 0
transform 1 0 4910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1427_
timestamp 0
transform 1 0 1370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1430_
timestamp 0
transform 1 0 3990 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 1850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1436_
timestamp 0
transform -1 0 2850 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1438_
timestamp 0
transform 1 0 2710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1441_
timestamp 0
transform -1 0 4350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1444_
timestamp 0
transform 1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1447_
timestamp 0
transform 1 0 1210 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1450_
timestamp 0
transform 1 0 950 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1452_
timestamp 0
transform -1 0 2010 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1455_
timestamp 0
transform 1 0 2790 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1458_
timestamp 0
transform 1 0 3990 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1461_
timestamp 0
transform 1 0 4330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1464_
timestamp 0
transform 1 0 4490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1466_
timestamp 0
transform -1 0 4270 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1469_
timestamp 0
transform -1 0 3510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1472_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1475_
timestamp 0
transform -1 0 2850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1477_
timestamp 0
transform -1 0 2810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1480_
timestamp 0
transform -1 0 4430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1483_
timestamp 0
transform 1 0 1930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1486_
timestamp 0
transform 1 0 4810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1489_
timestamp 0
transform -1 0 4950 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1491_
timestamp 0
transform -1 0 4370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1494_
timestamp 0
transform -1 0 5450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1497_
timestamp 0
transform -1 0 1790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1500_
timestamp 0
transform -1 0 3010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1502_
timestamp 0
transform -1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1505_
timestamp 0
transform 1 0 3130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1508_
timestamp 0
transform 1 0 2650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1511_
timestamp 0
transform -1 0 1970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1514_
timestamp 0
transform -1 0 1490 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1516_
timestamp 0
transform 1 0 2370 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1519_
timestamp 0
transform 1 0 1950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1522_
timestamp 0
transform 1 0 2050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1525_
timestamp 0
transform 1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1528_
timestamp 0
transform 1 0 4990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 5350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1533_
timestamp 0
transform 1 0 3830 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1536_
timestamp 0
transform 1 0 5130 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1539_
timestamp 0
transform -1 0 2850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1541_
timestamp 0
transform 1 0 430 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1544_
timestamp 0
transform -1 0 1990 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1547_
timestamp 0
transform 1 0 2530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1550_
timestamp 0
transform -1 0 430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1553_
timestamp 0
transform 1 0 1870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1555_
timestamp 0
transform 1 0 2690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1558_
timestamp 0
transform 1 0 5250 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1561_
timestamp 0
transform 1 0 5630 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1564_
timestamp 0
transform -1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1566_
timestamp 0
transform -1 0 730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1569_
timestamp 0
transform -1 0 1490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1572_
timestamp 0
transform -1 0 3010 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1575_
timestamp 0
transform -1 0 3550 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1578_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1580_
timestamp 0
transform 1 0 4850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1583_
timestamp 0
transform -1 0 4650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1586_
timestamp 0
transform -1 0 710 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1589_
timestamp 0
transform 1 0 1570 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1592_
timestamp 0
transform 1 0 2970 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1594_
timestamp 0
transform 1 0 3110 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1597_
timestamp 0
transform -1 0 3270 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1600_
timestamp 0
transform 1 0 4590 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1603_
timestamp 0
transform -1 0 5450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1605_
timestamp 0
transform 1 0 830 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1608_
timestamp 0
transform 1 0 2570 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1611_
timestamp 0
transform 1 0 2270 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1614_
timestamp 0
transform 1 0 2270 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1617_
timestamp 0
transform -1 0 4050 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1619_
timestamp 0
transform 1 0 4530 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1622_
timestamp 0
transform 1 0 4010 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1625_
timestamp 0
transform -1 0 4190 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1628_
timestamp 0
transform -1 0 4150 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1630_
timestamp 0
transform -1 0 2150 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1633_
timestamp 0
transform 1 0 2030 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1636_
timestamp 0
transform 1 0 2330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1639_
timestamp 0
transform 1 0 2470 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1642_
timestamp 0
transform 1 0 4390 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1644_
timestamp 0
transform -1 0 4310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1647_
timestamp 0
transform -1 0 4250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1650_
timestamp 0
transform 1 0 3050 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1653_
timestamp 0
transform -1 0 2630 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1655_
timestamp 0
transform 1 0 3590 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1658_
timestamp 0
transform 1 0 1310 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1661_
timestamp 0
transform -1 0 1750 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1664_
timestamp 0
transform -1 0 1490 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1667_
timestamp 0
transform -1 0 1370 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1669_
timestamp 0
transform 1 0 2590 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1672_
timestamp 0
transform -1 0 3830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1675_
timestamp 0
transform 1 0 970 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1678_
timestamp 0
transform -1 0 810 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1681_
timestamp 0
transform 1 0 770 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1683_
timestamp 0
transform 1 0 450 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1686_
timestamp 0
transform 1 0 610 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1689_
timestamp 0
transform 1 0 3290 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1692_
timestamp 0
transform -1 0 610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1694_
timestamp 0
transform -1 0 310 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1697_
timestamp 0
transform -1 0 170 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1700_
timestamp 0
transform -1 0 70 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1703_
timestamp 0
transform 1 0 1070 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1706_
timestamp 0
transform -1 0 1830 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1708_
timestamp 0
transform -1 0 3510 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1711_
timestamp 0
transform 1 0 1510 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1714_
timestamp 0
transform 1 0 1870 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1717_
timestamp 0
transform -1 0 1230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1719_
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1722_
timestamp 0
transform 1 0 1970 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1725_
timestamp 0
transform 1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1808_
timestamp 0
transform -1 0 5030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1811_
timestamp 0
transform 1 0 4390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__1813_
timestamp 0
transform 1 0 5650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform 1 0 3330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform -1 0 990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform -1 0 1650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 4750 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform 1 0 5430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 2110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform 1 0 2690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform 1 0 5050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert28
timestamp 0
transform -1 0 2330 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert31
timestamp 0
transform -1 0 1870 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert33
timestamp 0
transform 1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert36
timestamp 0
transform 1 0 5190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert39
timestamp 0
transform -1 0 1330 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert42
timestamp 0
transform -1 0 1310 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert45
timestamp 0
transform 1 0 1590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert47
timestamp 0
transform 1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert50
timestamp 0
transform -1 0 2390 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert53
timestamp 0
transform -1 0 1910 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert56
timestamp 0
transform -1 0 590 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert58
timestamp 0
transform -1 0 2990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert14
timestamp 0
transform -1 0 5670 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert17
timestamp 0
transform -1 0 2970 0 1 1690
box -6 -8 26 248
<< labels >>
flabel metal1 s 5942 2 6002 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 4256 -16 4264 7 FreeSans 16 0 0 0 Ain[1]
port 2 nsew
flabel metal3 s -24 4216 -16 4224 7 FreeSans 16 0 0 0 Ain[0]
port 3 nsew
flabel metal2 s 5417 6057 5423 6063 3 FreeSans 16 90 0 0 Aout[1]
port 4 nsew
flabel metal2 s 5057 6057 5063 6063 3 FreeSans 16 90 0 0 Aout[0]
port 5 nsew
flabel metal3 s -24 5876 -16 5884 7 FreeSans 16 0 0 0 ISin
port 6 nsew
flabel metal2 s 4477 6057 4483 6063 3 FreeSans 16 90 0 0 ISout
port 7 nsew
flabel metal3 s -24 3236 -16 3244 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal2 s 1877 -23 1883 -17 7 FreeSans 16 270 0 0 Stg[2]
port 9 nsew
flabel metal2 s 1737 -23 1743 -17 7 FreeSans 16 270 0 0 Stg[1]
port 10 nsew
flabel metal2 s 1697 -23 1703 -17 7 FreeSans 16 270 0 0 Stg[0]
port 11 nsew
flabel metal2 s 4437 6057 4443 6063 3 FreeSans 16 90 0 0 Vld
port 12 nsew
flabel metal2 s 4657 -23 4663 -17 7 FreeSans 16 270 0 0 Xin[1]
port 13 nsew
flabel metal2 s 4617 -23 4623 -17 7 FreeSans 16 270 0 0 Xin[0]
port 14 nsew
flabel metal3 s 5976 5916 5984 5924 3 FreeSans 16 0 0 0 Xout[1]
port 15 nsew
flabel metal3 s 5976 5876 5984 5884 3 FreeSans 16 0 0 0 Xout[0]
port 16 nsew
flabel metal2 s 2037 -23 2043 -17 7 FreeSans 16 270 0 0 Yin[1]
port 17 nsew
flabel metal2 s 1997 -23 2003 -17 7 FreeSans 16 270 0 0 Yin[0]
port 18 nsew
flabel metal3 s 5976 2276 5984 2284 3 FreeSans 16 0 0 0 Yout[1]
port 19 nsew
flabel metal3 s 5976 2036 5984 2044 3 FreeSans 16 0 0 0 Yout[0]
port 20 nsew
flabel metal3 s -24 1336 -16 1344 7 FreeSans 16 0 0 0 clk
port 21 nsew
<< properties >>
string FIXED_BBOX -40 -40 5980 6060
<< end >>
