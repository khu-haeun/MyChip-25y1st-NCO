magic
tech scmos
magscale 1 30
timestamp 1761282813
<< checkpaint >>
rect 9150 9150 180850 180850
use IOFILLER18  IOFILLER18_0
timestamp 1569536352
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1569536352
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1569536352
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1569536352
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1569536352
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1569536352
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1569536352
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1569536352
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1569536352
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1569536352
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1569536352
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1569536352
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1569536352
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1569536352
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1569536352
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1569536352
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1569536352
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1569536352
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1569536352
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1569536352
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1569536352
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1569536352
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1569536352
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1569536352
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50$1  IOFILLER50_0
timestamp 1569536352
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_1
timestamp 1569536352
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_2
timestamp 1569536352
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_3
timestamp 1569536352
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_4
timestamp 1569536352
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_5
timestamp 1569536352
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_6
timestamp 1569536352
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50$1  IOFILLER50_7
timestamp 1569536352
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PVDD$1  PAD_1_VDD
timestamp 1569536352
transform 0 1 18900 -1 0 141500
box 0 -9150 12000 25300
use PIC$1  PAD_2_CLK
timestamp 1569536352
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC$1  PAD_3_En
timestamp 1569536352
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC$1  PAD_4_FCW0
timestamp 1569536352
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC$1  PAD_5_FCW1
timestamp 1569536352
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC$1  PAD_6_FCW2
timestamp 1569536352
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PIC$1  PAD_7_FCW3
timestamp 1569536352
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PIC$1  PAD_8_FCW4
timestamp 1569536352
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_9_FCW5
timestamp 1569536352
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_10_FCW6
timestamp 1569536352
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_11_FCW7
timestamp 1569536352
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_12_FCW8
timestamp 1569536352
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_13_FCW9
timestamp 1569536352
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_14_FCW10
timestamp 1569536352
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC$1  PAD_15_FCW11
timestamp 1569536352
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC$1  PAD_16_FCW12
timestamp 1569536352
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC$1  PAD_17_FCW13
timestamp 1569536352
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC$1  PAD_18_FCW14
timestamp 1569536352
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC$1  PAD_19_FCW15
timestamp 1569536352
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use PIC$1  PAD_20_FCW16
timestamp 1569536352
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PIC$1  PAD_21_FCW17
timestamp 1569536352
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC$1  PAD_22_FCW18
timestamp 1569536352
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC$1  PAD_23_FCW19
timestamp 1569536352
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use POB8$1  PAD_24_Aout0
timestamp 1569536352
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB8$1  PAD_25_Aout1
timestamp 1569536352
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8$1  PAD_26_ISout
timestamp 1569536352
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8$1  PAD_27_Vld
timestamp 1569536352
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PVSS$1  PAD_28_VSS
timestamp 1569536352
transform 1 0 48500 0 -1 171100
box 0 -9150 12000 25300
use PCORNER$1  PCORNER_0
timestamp 1569536352
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER$1  PCORNER_1
timestamp 1569536352
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER$1  PCORNER_2
timestamp 1569536352
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER$1  PCORNER_3
timestamp 1569536352
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use phase_accumulator_Core_F  phase_accumulator_Core_F_0
timestamp 1569536352
transform 1 0 56700 0 1 59105
box -930 -365 77430 72950
use phase_accumulator_Pin_Route_F  phase_accumulator_Pin_Route_F_0
timestamp 1569536352
transform 1 0 0 0 1 0
box 44100 44100 145900 145900
<< end >>
