magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -604 -84 1287 876
<< ndiffusion >>
rect -484 36 1167 296
<< psubstratepdiff >>
rect -484 496 1167 756
<< metal1 >>
rect -484 496 1167 756
rect -484 36 1167 296
use CONT$3  CONT$3_0
array 0 44 36 0 5 36
timestamp 1569543463
transform 1 0 -460 0 1 76
box -6 -6 6 6
use CONT$3  CONT$3_1
array 0 44 36 0 5 36
timestamp 1569543463
transform 1 0 -460 0 1 536
box -6 -6 6 6
<< end >>
