magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -120 -120 5180 5180
<< metal1 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5030
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal2 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5031
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal3 >>
rect 0 2260 1560 5060
rect 2260 4220 3820 5060
rect 4220 4552 4552 5060
rect 4680 5012 5012 5060
tri 5012 5012 5060 5060 sw
rect 4680 4817 5060 5012
tri 4680 4680 4817 4817 ne
rect 4817 4680 5060 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5060 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5060 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5060 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5060 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5060 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5060 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5060 1560
use VIA1$5  VIA1$5_0
timestamp 1569543463
transform 1 0 4744 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_1
timestamp 1569543463
transform 1 0 4872 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_2
timestamp 1569543463
transform 1 0 4808 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_3
timestamp 1569543463
transform 1 0 4680 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_4
timestamp 1569543463
transform 1 0 4680 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_5
timestamp 1569543463
transform 1 0 4744 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_6
timestamp 1569543463
transform 1 0 4744 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_7
timestamp 1569543463
transform 1 0 4872 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_8
timestamp 1569543463
transform 1 0 4680 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_9
timestamp 1569543463
transform 1 0 4808 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_10
timestamp 1569543463
transform 1 0 4872 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_11
timestamp 1569543463
transform 1 0 4680 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_12
timestamp 1569543463
transform 1 0 4808 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_13
timestamp 1569543463
transform 1 0 4744 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_14
timestamp 1569543463
transform 1 0 4680 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_15
timestamp 1569543463
transform 1 0 4808 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_16
timestamp 1569543463
transform 1 0 4808 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_17
timestamp 1569543463
transform 1 0 4872 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_18
timestamp 1569543463
transform 1 0 4744 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_19
timestamp 1569543463
transform 1 0 4872 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_20
timestamp 1569543463
transform 1 0 4552 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_21
timestamp 1569543463
transform 1 0 4488 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_22
timestamp 1569543463
transform 1 0 4616 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_23
timestamp 1569543463
transform 1 0 4552 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_24
timestamp 1569543463
transform 1 0 4616 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_25
timestamp 1569543463
transform 1 0 4488 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_26
timestamp 1569543463
transform 1 0 4424 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_27
timestamp 1569543463
transform 1 0 4616 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_28
timestamp 1569543463
transform 1 0 4552 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_29
timestamp 1569543463
transform 1 0 4488 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_30
timestamp 1569543463
transform 1 0 4424 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_31
timestamp 1569543463
transform 1 0 4424 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_32
timestamp 1569543463
transform 1 0 4552 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_33
timestamp 1569543463
transform 1 0 4616 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_34
timestamp 1569543463
transform 1 0 4424 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_35
timestamp 1569543463
transform 1 0 4424 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_36
timestamp 1569543463
transform 1 0 4552 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_37
timestamp 1569543463
transform 1 0 4488 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_38
timestamp 1569543463
transform 1 0 4488 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_39
timestamp 1569543463
transform 1 0 4616 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_40
timestamp 1569543463
transform 1 0 4616 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_41
timestamp 1569543463
transform 1 0 4424 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_42
timestamp 1569543463
transform 1 0 4424 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_43
timestamp 1569543463
transform 1 0 4552 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_44
timestamp 1569543463
transform 1 0 4488 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_45
timestamp 1569543463
transform 1 0 4488 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_46
timestamp 1569543463
transform 1 0 4552 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_47
timestamp 1569543463
transform 1 0 4424 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_48
timestamp 1569543463
transform 1 0 4552 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_49
timestamp 1569543463
transform 1 0 4616 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_50
timestamp 1569543463
transform 1 0 4552 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_51
timestamp 1569543463
transform 1 0 4616 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_52
timestamp 1569543463
transform 1 0 4616 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_53
timestamp 1569543463
transform 1 0 4488 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_54
timestamp 1569543463
transform 1 0 4488 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_55
timestamp 1569543463
transform 1 0 4424 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_56
timestamp 1569543463
transform 1 0 4872 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_57
timestamp 1569543463
transform 1 0 4680 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_58
timestamp 1569543463
transform 1 0 4808 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_59
timestamp 1569543463
transform 1 0 4872 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_60
timestamp 1569543463
transform 1 0 4808 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_61
timestamp 1569543463
transform 1 0 4744 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_62
timestamp 1569543463
transform 1 0 4744 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_63
timestamp 1569543463
transform 1 0 4808 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_64
timestamp 1569543463
transform 1 0 4680 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_65
timestamp 1569543463
transform 1 0 4872 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_66
timestamp 1569543463
transform 1 0 4808 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_67
timestamp 1569543463
transform 1 0 4744 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_68
timestamp 1569543463
transform 1 0 4872 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_69
timestamp 1569543463
transform 1 0 4680 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_70
timestamp 1569543463
transform 1 0 4680 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_71
timestamp 1569543463
transform 1 0 4744 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_72
timestamp 1569543463
transform 1 0 4232 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_73
timestamp 1569543463
transform 1 0 4168 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_74
timestamp 1569543463
transform 1 0 4168 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_75
timestamp 1569543463
transform 1 0 4296 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_76
timestamp 1569543463
transform 1 0 4296 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_77
timestamp 1569543463
transform 1 0 4296 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_78
timestamp 1569543463
transform 1 0 4232 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_79
timestamp 1569543463
transform 1 0 4104 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_80
timestamp 1569543463
transform 1 0 4168 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_81
timestamp 1569543463
transform 1 0 4168 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_82
timestamp 1569543463
transform 1 0 4232 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_83
timestamp 1569543463
transform 1 0 4104 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_84
timestamp 1569543463
transform 1 0 4104 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_85
timestamp 1569543463
transform 1 0 4104 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_86
timestamp 1569543463
transform 1 0 4232 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_87
timestamp 1569543463
transform 1 0 4232 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_88
timestamp 1569543463
transform 1 0 4104 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_89
timestamp 1569543463
transform 1 0 4296 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_90
timestamp 1569543463
transform 1 0 4296 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_91
timestamp 1569543463
transform 1 0 4168 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_92
timestamp 1569543463
transform 1 0 3784 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_93
timestamp 1569543463
transform 1 0 3848 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_94
timestamp 1569543463
transform 1 0 3912 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_95
timestamp 1569543463
transform 1 0 4040 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_96
timestamp 1569543463
transform 1 0 4040 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_97
timestamp 1569543463
transform 1 0 3912 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_98
timestamp 1569543463
transform 1 0 3848 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_99
timestamp 1569543463
transform 1 0 3976 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_100
timestamp 1569543463
transform 1 0 3784 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_101
timestamp 1569543463
transform 1 0 3912 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_102
timestamp 1569543463
transform 1 0 4040 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_103
timestamp 1569543463
transform 1 0 3976 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_104
timestamp 1569543463
transform 1 0 4040 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_105
timestamp 1569543463
transform 1 0 3848 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_106
timestamp 1569543463
transform 1 0 3848 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_107
timestamp 1569543463
transform 1 0 3912 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_108
timestamp 1569543463
transform 1 0 4040 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_109
timestamp 1569543463
transform 1 0 3976 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_110
timestamp 1569543463
transform 1 0 3912 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_111
timestamp 1569543463
transform 1 0 3784 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_112
timestamp 1569543463
transform 1 0 3848 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_113
timestamp 1569543463
transform 1 0 3784 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_114
timestamp 1569543463
transform 1 0 3784 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_115
timestamp 1569543463
transform 1 0 3976 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_116
timestamp 1569543463
transform 1 0 3976 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_117
timestamp 1569543463
transform 1 0 3784 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_118
timestamp 1569543463
transform 1 0 3912 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_119
timestamp 1569543463
transform 1 0 3976 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_120
timestamp 1569543463
transform 1 0 3848 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_121
timestamp 1569543463
transform 1 0 4040 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_122
timestamp 1569543463
transform 1 0 3912 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_123
timestamp 1569543463
transform 1 0 4040 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_124
timestamp 1569543463
transform 1 0 3976 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_125
timestamp 1569543463
transform 1 0 3976 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_126
timestamp 1569543463
transform 1 0 3912 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_127
timestamp 1569543463
transform 1 0 3976 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_128
timestamp 1569543463
transform 1 0 3848 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_129
timestamp 1569543463
transform 1 0 3784 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_130
timestamp 1569543463
transform 1 0 4040 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_131
timestamp 1569543463
transform 1 0 3912 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_132
timestamp 1569543463
transform 1 0 3784 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_133
timestamp 1569543463
transform 1 0 3848 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_134
timestamp 1569543463
transform 1 0 4040 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_135
timestamp 1569543463
transform 1 0 3848 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_136
timestamp 1569543463
transform 1 0 3784 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_137
timestamp 1569543463
transform 1 0 4104 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_138
timestamp 1569543463
transform 1 0 4296 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_139
timestamp 1569543463
transform 1 0 4168 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_140
timestamp 1569543463
transform 1 0 4168 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_141
timestamp 1569543463
transform 1 0 4104 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_142
timestamp 1569543463
transform 1 0 4104 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_143
timestamp 1569543463
transform 1 0 4232 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_144
timestamp 1569543463
transform 1 0 4232 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_145
timestamp 1569543463
transform 1 0 4232 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_146
timestamp 1569543463
transform 1 0 4168 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_147
timestamp 1569543463
transform 1 0 4168 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_148
timestamp 1569543463
transform 1 0 4232 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_149
timestamp 1569543463
transform 1 0 4104 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_150
timestamp 1569543463
transform 1 0 4296 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_151
timestamp 1569543463
transform 1 0 4296 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_152
timestamp 1569543463
transform 1 0 4296 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_153
timestamp 1569543463
transform 1 0 4232 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_154
timestamp 1569543463
transform 1 0 4104 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_155
timestamp 1569543463
transform 1 0 4232 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_156
timestamp 1569543463
transform 1 0 4168 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_157
timestamp 1569543463
transform 1 0 4168 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_158
timestamp 1569543463
transform 1 0 4168 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_159
timestamp 1569543463
transform 1 0 4168 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_160
timestamp 1569543463
transform 1 0 4232 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_161
timestamp 1569543463
transform 1 0 4104 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_162
timestamp 1569543463
transform 1 0 4296 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_163
timestamp 1569543463
transform 1 0 4296 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_164
timestamp 1569543463
transform 1 0 4232 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_165
timestamp 1569543463
transform 1 0 4296 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_166
timestamp 1569543463
transform 1 0 4104 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_167
timestamp 1569543463
transform 1 0 4296 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_168
timestamp 1569543463
transform 1 0 4104 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_169
timestamp 1569543463
transform 1 0 3976 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_170
timestamp 1569543463
transform 1 0 3976 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_171
timestamp 1569543463
transform 1 0 3912 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_172
timestamp 1569543463
transform 1 0 4040 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_173
timestamp 1569543463
transform 1 0 3848 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_174
timestamp 1569543463
transform 1 0 3848 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_175
timestamp 1569543463
transform 1 0 3784 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_176
timestamp 1569543463
transform 1 0 3784 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_177
timestamp 1569543463
transform 1 0 3912 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_178
timestamp 1569543463
transform 1 0 3848 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_179
timestamp 1569543463
transform 1 0 4040 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_180
timestamp 1569543463
transform 1 0 3784 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_181
timestamp 1569543463
transform 1 0 3912 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_182
timestamp 1569543463
transform 1 0 3976 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_183
timestamp 1569543463
transform 1 0 3912 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_184
timestamp 1569543463
transform 1 0 3976 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_185
timestamp 1569543463
transform 1 0 4040 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_186
timestamp 1569543463
transform 1 0 3784 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_187
timestamp 1569543463
transform 1 0 4040 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_188
timestamp 1569543463
transform 1 0 3848 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_189
timestamp 1569543463
transform 1 0 3848 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_190
timestamp 1569543463
transform 1 0 4040 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_191
timestamp 1569543463
transform 1 0 3848 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_192
timestamp 1569543463
transform 1 0 3784 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_193
timestamp 1569543463
transform 1 0 4040 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_194
timestamp 1569543463
transform 1 0 4040 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_195
timestamp 1569543463
transform 1 0 3848 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_196
timestamp 1569543463
transform 1 0 3976 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_197
timestamp 1569543463
transform 1 0 3848 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_198
timestamp 1569543463
transform 1 0 3976 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_199
timestamp 1569543463
transform 1 0 3784 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_200
timestamp 1569543463
transform 1 0 3976 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_201
timestamp 1569543463
transform 1 0 3912 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_202
timestamp 1569543463
transform 1 0 3784 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_203
timestamp 1569543463
transform 1 0 3912 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_204
timestamp 1569543463
transform 1 0 3784 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_205
timestamp 1569543463
transform 1 0 3912 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_206
timestamp 1569543463
transform 1 0 4040 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_207
timestamp 1569543463
transform 1 0 3976 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_208
timestamp 1569543463
transform 1 0 3912 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_209
timestamp 1569543463
transform 1 0 3784 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_210
timestamp 1569543463
transform 1 0 3848 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_211
timestamp 1569543463
transform 1 0 4040 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_212
timestamp 1569543463
transform 1 0 3976 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_213
timestamp 1569543463
transform 1 0 3912 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_214
timestamp 1569543463
transform 1 0 4104 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_215
timestamp 1569543463
transform 1 0 4104 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_216
timestamp 1569543463
transform 1 0 4296 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_217
timestamp 1569543463
transform 1 0 4104 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_218
timestamp 1569543463
transform 1 0 4104 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_219
timestamp 1569543463
transform 1 0 4104 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_220
timestamp 1569543463
transform 1 0 4296 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_221
timestamp 1569543463
transform 1 0 4296 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_222
timestamp 1569543463
transform 1 0 4168 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_223
timestamp 1569543463
transform 1 0 4296 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_224
timestamp 1569543463
transform 1 0 4168 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_225
timestamp 1569543463
transform 1 0 4168 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_226
timestamp 1569543463
transform 1 0 4168 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_227
timestamp 1569543463
transform 1 0 4168 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_228
timestamp 1569543463
transform 1 0 4296 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_229
timestamp 1569543463
transform 1 0 4232 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_230
timestamp 1569543463
transform 1 0 4232 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_231
timestamp 1569543463
transform 1 0 4232 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_232
timestamp 1569543463
transform 1 0 4232 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_233
timestamp 1569543463
transform 1 0 4232 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_234
timestamp 1569543463
transform 1 0 4680 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_235
timestamp 1569543463
transform 1 0 4744 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_236
timestamp 1569543463
transform 1 0 4808 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_237
timestamp 1569543463
transform 1 0 4808 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_238
timestamp 1569543463
transform 1 0 4808 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_239
timestamp 1569543463
transform 1 0 4744 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_240
timestamp 1569543463
transform 1 0 4872 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_241
timestamp 1569543463
transform 1 0 4680 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_242
timestamp 1569543463
transform 1 0 4744 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_243
timestamp 1569543463
transform 1 0 4744 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_244
timestamp 1569543463
transform 1 0 4872 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_245
timestamp 1569543463
transform 1 0 4808 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_246
timestamp 1569543463
transform 1 0 4680 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_247
timestamp 1569543463
transform 1 0 4872 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_248
timestamp 1569543463
transform 1 0 4872 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_249
timestamp 1569543463
transform 1 0 4680 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_250
timestamp 1569543463
transform 1 0 4616 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_251
timestamp 1569543463
transform 1 0 4488 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_252
timestamp 1569543463
transform 1 0 4552 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_253
timestamp 1569543463
transform 1 0 4424 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_254
timestamp 1569543463
transform 1 0 4424 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_255
timestamp 1569543463
transform 1 0 4424 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_256
timestamp 1569543463
transform 1 0 4488 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_257
timestamp 1569543463
transform 1 0 4616 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_258
timestamp 1569543463
transform 1 0 4616 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_259
timestamp 1569543463
transform 1 0 4552 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_260
timestamp 1569543463
transform 1 0 4616 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_261
timestamp 1569543463
transform 1 0 4488 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_262
timestamp 1569543463
transform 1 0 4552 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_263
timestamp 1569543463
transform 1 0 4424 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_264
timestamp 1569543463
transform 1 0 4552 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_265
timestamp 1569543463
transform 1 0 4488 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_266
timestamp 1569543463
transform 1 0 4488 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_267
timestamp 1569543463
transform 1 0 4488 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_268
timestamp 1569543463
transform 1 0 4488 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_269
timestamp 1569543463
transform 1 0 4552 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_270
timestamp 1569543463
transform 1 0 4424 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_271
timestamp 1569543463
transform 1 0 4424 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_272
timestamp 1569543463
transform 1 0 4616 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_273
timestamp 1569543463
transform 1 0 4424 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_274
timestamp 1569543463
transform 1 0 4488 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_275
timestamp 1569543463
transform 1 0 4616 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_276
timestamp 1569543463
transform 1 0 4488 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_277
timestamp 1569543463
transform 1 0 4424 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_278
timestamp 1569543463
transform 1 0 4616 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_279
timestamp 1569543463
transform 1 0 4552 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_280
timestamp 1569543463
transform 1 0 4552 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_281
timestamp 1569543463
transform 1 0 4552 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_282
timestamp 1569543463
transform 1 0 4424 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_283
timestamp 1569543463
transform 1 0 4552 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_284
timestamp 1569543463
transform 1 0 4616 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_285
timestamp 1569543463
transform 1 0 4616 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_286
timestamp 1569543463
transform 1 0 4680 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_287
timestamp 1569543463
transform 1 0 4680 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_288
timestamp 1569543463
transform 1 0 4680 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_289
timestamp 1569543463
transform 1 0 4680 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_290
timestamp 1569543463
transform 1 0 4744 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_291
timestamp 1569543463
transform 1 0 4744 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_292
timestamp 1569543463
transform 1 0 4744 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_293
timestamp 1569543463
transform 1 0 4744 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_294
timestamp 1569543463
transform 1 0 4744 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_295
timestamp 1569543463
transform 1 0 4808 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_296
timestamp 1569543463
transform 1 0 4808 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_297
timestamp 1569543463
transform 1 0 4808 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_298
timestamp 1569543463
transform 1 0 4808 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_299
timestamp 1569543463
transform 1 0 4808 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_300
timestamp 1569543463
transform 1 0 4872 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_301
timestamp 1569543463
transform 1 0 4872 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_302
timestamp 1569543463
transform 1 0 4872 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_303
timestamp 1569543463
transform 1 0 4872 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_304
timestamp 1569543463
transform 1 0 4872 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_305
timestamp 1569543463
transform 1 0 4680 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_306
timestamp 1569543463
transform 1 0 3976 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_307
timestamp 1569543463
transform 1 0 3784 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_308
timestamp 1569543463
transform 1 0 4424 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_309
timestamp 1569543463
transform 1 0 4616 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_310
timestamp 1569543463
transform 1 0 4360 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_311
timestamp 1569543463
transform 1 0 3848 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_312
timestamp 1569543463
transform 1 0 4488 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_313
timestamp 1569543463
transform 1 0 4104 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_314
timestamp 1569543463
transform 1 0 4744 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_315
timestamp 1569543463
transform 1 0 4360 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_316
timestamp 1569543463
transform 1 0 3912 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_317
timestamp 1569543463
transform 1 0 4552 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_318
timestamp 1569543463
transform 1 0 4232 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_319
timestamp 1569543463
transform 1 0 4872 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_320
timestamp 1569543463
transform 1 0 4360 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_321
timestamp 1569543463
transform 1 0 4040 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_322
timestamp 1569543463
transform 1 0 4680 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_323
timestamp 1569543463
transform 1 0 4360 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_324
timestamp 1569543463
transform 1 0 4296 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_325
timestamp 1569543463
transform 1 0 4360 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_326
timestamp 1569543463
transform 1 0 4360 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_327
timestamp 1569543463
transform 1 0 4360 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_328
timestamp 1569543463
transform 1 0 4360 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_329
timestamp 1569543463
transform 1 0 4360 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_330
timestamp 1569543463
transform 1 0 4360 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_331
timestamp 1569543463
transform 1 0 4360 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_332
timestamp 1569543463
transform 1 0 4360 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_333
timestamp 1569543463
transform 1 0 4360 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_334
timestamp 1569543463
transform 1 0 4360 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_335
timestamp 1569543463
transform 1 0 4360 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_336
timestamp 1569543463
transform 1 0 4168 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_337
timestamp 1569543463
transform 1 0 4360 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_338
timestamp 1569543463
transform 1 0 4360 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_339
timestamp 1569543463
transform 1 0 4808 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_340
timestamp 1569543463
transform 1 0 4360 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_341
timestamp 1569543463
transform 1 0 4360 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_342
timestamp 1569543463
transform 1 0 3592 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_343
timestamp 1569543463
transform 1 0 3656 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_344
timestamp 1569543463
transform 1 0 3592 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_345
timestamp 1569543463
transform 1 0 3592 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_346
timestamp 1569543463
transform 1 0 3464 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_347
timestamp 1569543463
transform 1 0 3592 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_348
timestamp 1569543463
transform 1 0 3656 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_349
timestamp 1569543463
transform 1 0 3720 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_350
timestamp 1569543463
transform 1 0 3656 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_351
timestamp 1569543463
transform 1 0 3720 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_352
timestamp 1569543463
transform 1 0 3720 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_353
timestamp 1569543463
transform 1 0 3656 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_354
timestamp 1569543463
transform 1 0 3592 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_355
timestamp 1569543463
transform 1 0 3528 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_356
timestamp 1569543463
transform 1 0 3528 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_357
timestamp 1569543463
transform 1 0 3464 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_358
timestamp 1569543463
transform 1 0 3720 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_359
timestamp 1569543463
transform 1 0 3528 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_360
timestamp 1569543463
transform 1 0 3464 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_361
timestamp 1569543463
transform 1 0 3464 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_362
timestamp 1569543463
transform 1 0 3528 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_363
timestamp 1569543463
transform 1 0 3656 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_364
timestamp 1569543463
transform 1 0 3720 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_365
timestamp 1569543463
transform 1 0 3464 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_366
timestamp 1569543463
transform 1 0 3528 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_367
timestamp 1569543463
transform 1 0 3400 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_368
timestamp 1569543463
transform 1 0 3336 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_369
timestamp 1569543463
transform 1 0 3336 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_370
timestamp 1569543463
transform 1 0 3272 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_371
timestamp 1569543463
transform 1 0 3400 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_372
timestamp 1569543463
transform 1 0 3400 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_373
timestamp 1569543463
transform 1 0 3144 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_374
timestamp 1569543463
transform 1 0 3144 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_375
timestamp 1569543463
transform 1 0 3272 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_376
timestamp 1569543463
transform 1 0 3336 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_377
timestamp 1569543463
transform 1 0 3144 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_378
timestamp 1569543463
transform 1 0 3144 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_379
timestamp 1569543463
transform 1 0 3144 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_380
timestamp 1569543463
transform 1 0 3272 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_381
timestamp 1569543463
transform 1 0 3272 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_382
timestamp 1569543463
transform 1 0 3400 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_383
timestamp 1569543463
transform 1 0 3208 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_384
timestamp 1569543463
transform 1 0 3336 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_385
timestamp 1569543463
transform 1 0 3208 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_386
timestamp 1569543463
transform 1 0 3208 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_387
timestamp 1569543463
transform 1 0 3336 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_388
timestamp 1569543463
transform 1 0 3400 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_389
timestamp 1569543463
transform 1 0 3208 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_390
timestamp 1569543463
transform 1 0 3208 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_391
timestamp 1569543463
transform 1 0 3272 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_392
timestamp 1569543463
transform 1 0 3336 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_393
timestamp 1569543463
transform 1 0 3272 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_394
timestamp 1569543463
transform 1 0 3272 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_395
timestamp 1569543463
transform 1 0 3208 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_396
timestamp 1569543463
transform 1 0 3272 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_397
timestamp 1569543463
transform 1 0 3336 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_398
timestamp 1569543463
transform 1 0 3144 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_399
timestamp 1569543463
transform 1 0 3208 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_400
timestamp 1569543463
transform 1 0 3208 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_401
timestamp 1569543463
transform 1 0 3400 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_402
timestamp 1569543463
transform 1 0 3208 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_403
timestamp 1569543463
transform 1 0 3272 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_404
timestamp 1569543463
transform 1 0 3400 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_405
timestamp 1569543463
transform 1 0 3144 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_406
timestamp 1569543463
transform 1 0 3144 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_407
timestamp 1569543463
transform 1 0 3336 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_408
timestamp 1569543463
transform 1 0 3400 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_409
timestamp 1569543463
transform 1 0 3336 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_410
timestamp 1569543463
transform 1 0 3400 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_411
timestamp 1569543463
transform 1 0 3144 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_412
timestamp 1569543463
transform 1 0 3656 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_413
timestamp 1569543463
transform 1 0 3720 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_414
timestamp 1569543463
transform 1 0 3656 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_415
timestamp 1569543463
transform 1 0 3656 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_416
timestamp 1569543463
transform 1 0 3656 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_417
timestamp 1569543463
transform 1 0 3464 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_418
timestamp 1569543463
transform 1 0 3464 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_419
timestamp 1569543463
transform 1 0 3528 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_420
timestamp 1569543463
transform 1 0 3592 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_421
timestamp 1569543463
transform 1 0 3528 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_422
timestamp 1569543463
transform 1 0 3464 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_423
timestamp 1569543463
transform 1 0 3592 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_424
timestamp 1569543463
transform 1 0 3528 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_425
timestamp 1569543463
transform 1 0 3528 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_426
timestamp 1569543463
transform 1 0 3592 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_427
timestamp 1569543463
transform 1 0 3720 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_428
timestamp 1569543463
transform 1 0 3720 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_429
timestamp 1569543463
transform 1 0 3592 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_430
timestamp 1569543463
transform 1 0 3464 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_431
timestamp 1569543463
transform 1 0 3720 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_432
timestamp 1569543463
transform 1 0 2824 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_433
timestamp 1569543463
transform 1 0 3016 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_434
timestamp 1569543463
transform 1 0 2888 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_435
timestamp 1569543463
transform 1 0 3080 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_436
timestamp 1569543463
transform 1 0 3016 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_437
timestamp 1569543463
transform 1 0 3016 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_438
timestamp 1569543463
transform 1 0 3080 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_439
timestamp 1569543463
transform 1 0 2888 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_440
timestamp 1569543463
transform 1 0 2952 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_441
timestamp 1569543463
transform 1 0 2888 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_442
timestamp 1569543463
transform 1 0 2824 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_443
timestamp 1569543463
transform 1 0 2888 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_444
timestamp 1569543463
transform 1 0 2952 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_445
timestamp 1569543463
transform 1 0 2952 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_446
timestamp 1569543463
transform 1 0 2888 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_447
timestamp 1569543463
transform 1 0 2824 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_448
timestamp 1569543463
transform 1 0 2824 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_449
timestamp 1569543463
transform 1 0 3080 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_450
timestamp 1569543463
transform 1 0 2824 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_451
timestamp 1569543463
transform 1 0 3016 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_452
timestamp 1569543463
transform 1 0 2952 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_453
timestamp 1569543463
transform 1 0 3080 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_454
timestamp 1569543463
transform 1 0 3080 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_455
timestamp 1569543463
transform 1 0 3016 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_456
timestamp 1569543463
transform 1 0 2952 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_457
timestamp 1569543463
transform 1 0 2760 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_458
timestamp 1569543463
transform 1 0 2632 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_459
timestamp 1569543463
transform 1 0 2568 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_460
timestamp 1569543463
transform 1 0 2568 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_461
timestamp 1569543463
transform 1 0 2632 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_462
timestamp 1569543463
transform 1 0 2760 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_463
timestamp 1569543463
transform 1 0 2696 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_464
timestamp 1569543463
transform 1 0 2696 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_465
timestamp 1569543463
transform 1 0 2696 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_466
timestamp 1569543463
transform 1 0 2760 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_467
timestamp 1569543463
transform 1 0 2696 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_468
timestamp 1569543463
transform 1 0 2760 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_469
timestamp 1569543463
transform 1 0 2632 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_470
timestamp 1569543463
transform 1 0 2568 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_471
timestamp 1569543463
transform 1 0 2696 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_472
timestamp 1569543463
transform 1 0 2632 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_473
timestamp 1569543463
transform 1 0 2632 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_474
timestamp 1569543463
transform 1 0 2760 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_475
timestamp 1569543463
transform 1 0 2568 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_476
timestamp 1569543463
transform 1 0 2568 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_477
timestamp 1569543463
transform 1 0 2696 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_478
timestamp 1569543463
transform 1 0 2760 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_479
timestamp 1569543463
transform 1 0 2568 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_480
timestamp 1569543463
transform 1 0 2568 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_481
timestamp 1569543463
transform 1 0 2632 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_482
timestamp 1569543463
transform 1 0 2568 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_483
timestamp 1569543463
transform 1 0 2568 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_484
timestamp 1569543463
transform 1 0 2696 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_485
timestamp 1569543463
transform 1 0 2632 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_486
timestamp 1569543463
transform 1 0 2696 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_487
timestamp 1569543463
transform 1 0 2760 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_488
timestamp 1569543463
transform 1 0 2632 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_489
timestamp 1569543463
transform 1 0 2760 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_490
timestamp 1569543463
transform 1 0 2696 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_491
timestamp 1569543463
transform 1 0 2760 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_492
timestamp 1569543463
transform 1 0 2632 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_493
timestamp 1569543463
transform 1 0 2888 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_494
timestamp 1569543463
transform 1 0 2824 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_495
timestamp 1569543463
transform 1 0 3016 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_496
timestamp 1569543463
transform 1 0 3016 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_497
timestamp 1569543463
transform 1 0 2824 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_498
timestamp 1569543463
transform 1 0 2952 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_499
timestamp 1569543463
transform 1 0 2952 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_500
timestamp 1569543463
transform 1 0 2824 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_501
timestamp 1569543463
transform 1 0 3016 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_502
timestamp 1569543463
transform 1 0 2952 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_503
timestamp 1569543463
transform 1 0 3080 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_504
timestamp 1569543463
transform 1 0 2952 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_505
timestamp 1569543463
transform 1 0 3016 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_506
timestamp 1569543463
transform 1 0 3080 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_507
timestamp 1569543463
transform 1 0 3080 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_508
timestamp 1569543463
transform 1 0 3080 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_509
timestamp 1569543463
transform 1 0 2888 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_510
timestamp 1569543463
transform 1 0 2824 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_511
timestamp 1569543463
transform 1 0 2888 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_512
timestamp 1569543463
transform 1 0 2888 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_513
timestamp 1569543463
transform 1 0 2888 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_514
timestamp 1569543463
transform 1 0 2888 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_515
timestamp 1569543463
transform 1 0 3016 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_516
timestamp 1569543463
transform 1 0 2952 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_517
timestamp 1569543463
transform 1 0 3080 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_518
timestamp 1569543463
transform 1 0 3080 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_519
timestamp 1569543463
transform 1 0 3080 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_520
timestamp 1569543463
transform 1 0 3080 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_521
timestamp 1569543463
transform 1 0 2952 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_522
timestamp 1569543463
transform 1 0 2824 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_523
timestamp 1569543463
transform 1 0 2824 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_524
timestamp 1569543463
transform 1 0 2824 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_525
timestamp 1569543463
transform 1 0 2952 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_526
timestamp 1569543463
transform 1 0 3016 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_527
timestamp 1569543463
transform 1 0 3016 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_528
timestamp 1569543463
transform 1 0 3016 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_529
timestamp 1569543463
transform 1 0 2888 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_530
timestamp 1569543463
transform 1 0 2824 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_531
timestamp 1569543463
transform 1 0 2888 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_532
timestamp 1569543463
transform 1 0 2952 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_533
timestamp 1569543463
transform 1 0 2568 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_534
timestamp 1569543463
transform 1 0 2696 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_535
timestamp 1569543463
transform 1 0 2632 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_536
timestamp 1569543463
transform 1 0 2760 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_537
timestamp 1569543463
transform 1 0 2760 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_538
timestamp 1569543463
transform 1 0 2696 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_539
timestamp 1569543463
transform 1 0 2632 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_540
timestamp 1569543463
transform 1 0 2568 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_541
timestamp 1569543463
transform 1 0 2696 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_542
timestamp 1569543463
transform 1 0 2568 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_543
timestamp 1569543463
transform 1 0 2632 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_544
timestamp 1569543463
transform 1 0 2760 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_545
timestamp 1569543463
transform 1 0 2632 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_546
timestamp 1569543463
transform 1 0 2696 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_547
timestamp 1569543463
transform 1 0 2568 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_548
timestamp 1569543463
transform 1 0 2760 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_549
timestamp 1569543463
transform 1 0 2760 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_550
timestamp 1569543463
transform 1 0 2632 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_551
timestamp 1569543463
transform 1 0 2760 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_552
timestamp 1569543463
transform 1 0 2760 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_553
timestamp 1569543463
transform 1 0 2696 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_554
timestamp 1569543463
transform 1 0 2696 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_555
timestamp 1569543463
transform 1 0 2568 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_556
timestamp 1569543463
transform 1 0 2632 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_557
timestamp 1569543463
transform 1 0 2632 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_558
timestamp 1569543463
transform 1 0 2760 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_559
timestamp 1569543463
transform 1 0 2568 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_560
timestamp 1569543463
transform 1 0 2696 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_561
timestamp 1569543463
transform 1 0 2568 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_562
timestamp 1569543463
transform 1 0 2696 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_563
timestamp 1569543463
transform 1 0 2568 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_564
timestamp 1569543463
transform 1 0 2632 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_565
timestamp 1569543463
transform 1 0 2696 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_566
timestamp 1569543463
transform 1 0 2568 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_567
timestamp 1569543463
transform 1 0 2760 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_568
timestamp 1569543463
transform 1 0 2632 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_569
timestamp 1569543463
transform 1 0 3080 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_570
timestamp 1569543463
transform 1 0 2824 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_571
timestamp 1569543463
transform 1 0 3080 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_572
timestamp 1569543463
transform 1 0 2824 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_573
timestamp 1569543463
transform 1 0 2824 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_574
timestamp 1569543463
transform 1 0 3080 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_575
timestamp 1569543463
transform 1 0 2824 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_576
timestamp 1569543463
transform 1 0 2824 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_577
timestamp 1569543463
transform 1 0 3080 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_578
timestamp 1569543463
transform 1 0 3080 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_579
timestamp 1569543463
transform 1 0 2888 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_580
timestamp 1569543463
transform 1 0 2888 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_581
timestamp 1569543463
transform 1 0 2888 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_582
timestamp 1569543463
transform 1 0 2888 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_583
timestamp 1569543463
transform 1 0 2888 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_584
timestamp 1569543463
transform 1 0 2952 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_585
timestamp 1569543463
transform 1 0 2952 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_586
timestamp 1569543463
transform 1 0 2952 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_587
timestamp 1569543463
transform 1 0 2952 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_588
timestamp 1569543463
transform 1 0 2952 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_589
timestamp 1569543463
transform 1 0 3016 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_590
timestamp 1569543463
transform 1 0 3016 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_591
timestamp 1569543463
transform 1 0 3016 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_592
timestamp 1569543463
transform 1 0 3016 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_593
timestamp 1569543463
transform 1 0 3016 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_594
timestamp 1569543463
transform 1 0 3656 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_595
timestamp 1569543463
transform 1 0 3592 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_596
timestamp 1569543463
transform 1 0 3592 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_597
timestamp 1569543463
transform 1 0 3720 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_598
timestamp 1569543463
transform 1 0 3528 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_599
timestamp 1569543463
transform 1 0 3720 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_600
timestamp 1569543463
transform 1 0 3464 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_601
timestamp 1569543463
transform 1 0 3464 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_602
timestamp 1569543463
transform 1 0 3720 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_603
timestamp 1569543463
transform 1 0 3656 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_604
timestamp 1569543463
transform 1 0 3720 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_605
timestamp 1569543463
transform 1 0 3656 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_606
timestamp 1569543463
transform 1 0 3592 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_607
timestamp 1569543463
transform 1 0 3464 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_608
timestamp 1569543463
transform 1 0 3528 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_609
timestamp 1569543463
transform 1 0 3528 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_610
timestamp 1569543463
transform 1 0 3656 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_611
timestamp 1569543463
transform 1 0 3464 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_612
timestamp 1569543463
transform 1 0 3528 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_613
timestamp 1569543463
transform 1 0 3592 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_614
timestamp 1569543463
transform 1 0 3272 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_615
timestamp 1569543463
transform 1 0 3336 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_616
timestamp 1569543463
transform 1 0 3400 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_617
timestamp 1569543463
transform 1 0 3400 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_618
timestamp 1569543463
transform 1 0 3336 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_619
timestamp 1569543463
transform 1 0 3208 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_620
timestamp 1569543463
transform 1 0 3144 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_621
timestamp 1569543463
transform 1 0 3144 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_622
timestamp 1569543463
transform 1 0 3272 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_623
timestamp 1569543463
transform 1 0 3400 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_624
timestamp 1569543463
transform 1 0 3144 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_625
timestamp 1569543463
transform 1 0 3208 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_626
timestamp 1569543463
transform 1 0 3144 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_627
timestamp 1569543463
transform 1 0 3208 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_628
timestamp 1569543463
transform 1 0 3272 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_629
timestamp 1569543463
transform 1 0 3208 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_630
timestamp 1569543463
transform 1 0 3400 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_631
timestamp 1569543463
transform 1 0 3336 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_632
timestamp 1569543463
transform 1 0 3272 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_633
timestamp 1569543463
transform 1 0 3336 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_634
timestamp 1569543463
transform 1 0 3400 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_635
timestamp 1569543463
transform 1 0 3400 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_636
timestamp 1569543463
transform 1 0 3400 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_637
timestamp 1569543463
transform 1 0 3208 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_638
timestamp 1569543463
transform 1 0 3208 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_639
timestamp 1569543463
transform 1 0 3208 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_640
timestamp 1569543463
transform 1 0 3272 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_641
timestamp 1569543463
transform 1 0 3336 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_642
timestamp 1569543463
transform 1 0 3272 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_643
timestamp 1569543463
transform 1 0 3144 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_644
timestamp 1569543463
transform 1 0 3144 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_645
timestamp 1569543463
transform 1 0 3144 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_646
timestamp 1569543463
transform 1 0 3144 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_647
timestamp 1569543463
transform 1 0 3272 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_648
timestamp 1569543463
transform 1 0 3208 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_649
timestamp 1569543463
transform 1 0 3144 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_650
timestamp 1569543463
transform 1 0 3272 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_651
timestamp 1569543463
transform 1 0 3336 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_652
timestamp 1569543463
transform 1 0 3336 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_653
timestamp 1569543463
transform 1 0 3336 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_654
timestamp 1569543463
transform 1 0 3272 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_655
timestamp 1569543463
transform 1 0 3400 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_656
timestamp 1569543463
transform 1 0 3336 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_657
timestamp 1569543463
transform 1 0 3208 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_658
timestamp 1569543463
transform 1 0 3400 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_659
timestamp 1569543463
transform 1 0 3464 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_660
timestamp 1569543463
transform 1 0 3464 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_661
timestamp 1569543463
transform 1 0 3464 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_662
timestamp 1569543463
transform 1 0 3464 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_663
timestamp 1569543463
transform 1 0 3464 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_664
timestamp 1569543463
transform 1 0 3528 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_665
timestamp 1569543463
transform 1 0 3528 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_666
timestamp 1569543463
transform 1 0 3528 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_667
timestamp 1569543463
transform 1 0 3528 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_668
timestamp 1569543463
transform 1 0 3528 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_669
timestamp 1569543463
transform 1 0 3592 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_670
timestamp 1569543463
transform 1 0 3592 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_671
timestamp 1569543463
transform 1 0 3592 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_672
timestamp 1569543463
transform 1 0 3592 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_673
timestamp 1569543463
transform 1 0 3592 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_674
timestamp 1569543463
transform 1 0 3656 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_675
timestamp 1569543463
transform 1 0 3656 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_676
timestamp 1569543463
transform 1 0 3656 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_677
timestamp 1569543463
transform 1 0 3656 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_678
timestamp 1569543463
transform 1 0 3656 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_679
timestamp 1569543463
transform 1 0 3720 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_680
timestamp 1569543463
transform 1 0 3720 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_681
timestamp 1569543463
transform 1 0 3720 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_682
timestamp 1569543463
transform 1 0 3720 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_683
timestamp 1569543463
transform 1 0 3720 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_684
timestamp 1569543463
transform 1 0 3080 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_685
timestamp 1569543463
transform 1 0 3720 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_686
timestamp 1569543463
transform 1 0 3144 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_687
timestamp 1569543463
transform 1 0 2568 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_688
timestamp 1569543463
transform 1 0 3208 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_689
timestamp 1569543463
transform 1 0 2632 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_690
timestamp 1569543463
transform 1 0 3272 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_691
timestamp 1569543463
transform 1 0 2888 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_692
timestamp 1569543463
transform 1 0 3528 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_693
timestamp 1569543463
transform 1 0 2696 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_694
timestamp 1569543463
transform 1 0 3336 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_695
timestamp 1569543463
transform 1 0 2760 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_696
timestamp 1569543463
transform 1 0 3400 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_697
timestamp 1569543463
transform 1 0 2952 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_698
timestamp 1569543463
transform 1 0 3592 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_699
timestamp 1569543463
transform 1 0 3016 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_700
timestamp 1569543463
transform 1 0 3656 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_701
timestamp 1569543463
transform 1 0 2824 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_702
timestamp 1569543463
transform 1 0 3464 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_703
timestamp 1569543463
transform 1 0 3144 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_704
timestamp 1569543463
transform 1 0 3208 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_705
timestamp 1569543463
transform 1 0 3400 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_706
timestamp 1569543463
transform 1 0 3592 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_707
timestamp 1569543463
transform 1 0 3144 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_708
timestamp 1569543463
transform 1 0 3400 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_709
timestamp 1569543463
transform 1 0 3656 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_710
timestamp 1569543463
transform 1 0 3592 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_711
timestamp 1569543463
transform 1 0 3720 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_712
timestamp 1569543463
transform 1 0 3400 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_713
timestamp 1569543463
transform 1 0 3208 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_714
timestamp 1569543463
transform 1 0 3272 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_715
timestamp 1569543463
transform 1 0 3400 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_716
timestamp 1569543463
transform 1 0 3656 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_717
timestamp 1569543463
transform 1 0 3144 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_718
timestamp 1569543463
transform 1 0 3144 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_719
timestamp 1569543463
transform 1 0 3336 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_720
timestamp 1569543463
transform 1 0 3336 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_721
timestamp 1569543463
transform 1 0 3464 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_722
timestamp 1569543463
transform 1 0 3656 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_723
timestamp 1569543463
transform 1 0 3592 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_724
timestamp 1569543463
transform 1 0 3464 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_725
timestamp 1569543463
transform 1 0 3720 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_726
timestamp 1569543463
transform 1 0 3272 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_727
timestamp 1569543463
transform 1 0 3464 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_728
timestamp 1569543463
transform 1 0 3464 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_729
timestamp 1569543463
transform 1 0 3208 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_730
timestamp 1569543463
transform 1 0 3528 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_731
timestamp 1569543463
transform 1 0 3592 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_732
timestamp 1569543463
transform 1 0 3528 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_733
timestamp 1569543463
transform 1 0 3272 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_734
timestamp 1569543463
transform 1 0 3528 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_735
timestamp 1569543463
transform 1 0 3528 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_736
timestamp 1569543463
transform 1 0 3720 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_737
timestamp 1569543463
transform 1 0 3272 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_738
timestamp 1569543463
transform 1 0 3336 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_739
timestamp 1569543463
transform 1 0 3656 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_740
timestamp 1569543463
transform 1 0 3720 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_741
timestamp 1569543463
transform 1 0 3336 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_742
timestamp 1569543463
transform 1 0 3208 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_743
timestamp 1569543463
transform 1 0 2824 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_744
timestamp 1569543463
transform 1 0 3016 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_745
timestamp 1569543463
transform 1 0 2888 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_746
timestamp 1569543463
transform 1 0 2952 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_747
timestamp 1569543463
transform 1 0 2952 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_748
timestamp 1569543463
transform 1 0 2952 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_749
timestamp 1569543463
transform 1 0 3016 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_750
timestamp 1569543463
transform 1 0 2888 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_751
timestamp 1569543463
transform 1 0 3080 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_752
timestamp 1569543463
transform 1 0 3080 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_753
timestamp 1569543463
transform 1 0 3016 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_754
timestamp 1569543463
transform 1 0 2824 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_755
timestamp 1569543463
transform 1 0 2824 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_756
timestamp 1569543463
transform 1 0 2824 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_757
timestamp 1569543463
transform 1 0 2888 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_758
timestamp 1569543463
transform 1 0 3016 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_759
timestamp 1569543463
transform 1 0 2888 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_760
timestamp 1569543463
transform 1 0 2888 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_761
timestamp 1569543463
transform 1 0 3080 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_762
timestamp 1569543463
transform 1 0 3080 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_763
timestamp 1569543463
transform 1 0 2952 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_764
timestamp 1569543463
transform 1 0 2824 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_765
timestamp 1569543463
transform 1 0 2696 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_766
timestamp 1569543463
transform 1 0 2760 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_767
timestamp 1569543463
transform 1 0 2760 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_768
timestamp 1569543463
transform 1 0 2632 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_769
timestamp 1569543463
transform 1 0 2760 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_770
timestamp 1569543463
transform 1 0 2568 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_771
timestamp 1569543463
transform 1 0 2568 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_772
timestamp 1569543463
transform 1 0 2632 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_773
timestamp 1569543463
transform 1 0 2632 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_774
timestamp 1569543463
transform 1 0 2568 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_775
timestamp 1569543463
transform 1 0 2696 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_776
timestamp 1569543463
transform 1 0 2696 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_777
timestamp 1569543463
transform 1 0 2696 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_778
timestamp 1569543463
transform 1 0 2632 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_779
timestamp 1569543463
transform 1 0 2568 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_780
timestamp 1569543463
transform 1 0 2696 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_781
timestamp 1569543463
transform 1 0 2760 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_782
timestamp 1569543463
transform 1 0 2760 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_783
timestamp 1569543463
transform 1 0 2568 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_784
timestamp 1569543463
transform 1 0 2632 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_785
timestamp 1569543463
transform 1 0 2568 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_786
timestamp 1569543463
transform 1 0 2632 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_787
timestamp 1569543463
transform 1 0 2632 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_788
timestamp 1569543463
transform 1 0 2632 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_789
timestamp 1569543463
transform 1 0 2632 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_790
timestamp 1569543463
transform 1 0 2568 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_791
timestamp 1569543463
transform 1 0 2568 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_792
timestamp 1569543463
transform 1 0 2696 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_793
timestamp 1569543463
transform 1 0 2696 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_794
timestamp 1569543463
transform 1 0 2696 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_795
timestamp 1569543463
transform 1 0 2760 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_796
timestamp 1569543463
transform 1 0 2760 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_797
timestamp 1569543463
transform 1 0 2568 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_798
timestamp 1569543463
transform 1 0 2568 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_799
timestamp 1569543463
transform 1 0 2824 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_800
timestamp 1569543463
transform 1 0 3400 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_801
timestamp 1569543463
transform 1 0 3720 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_802
timestamp 1569543463
transform 1 0 3464 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_803
timestamp 1569543463
transform 1 0 3528 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_804
timestamp 1569543463
transform 1 0 3272 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_805
timestamp 1569543463
transform 1 0 3592 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_806
timestamp 1569543463
transform 1 0 3656 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_807
timestamp 1569543463
transform 1 0 3336 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_808
timestamp 1569543463
transform 1 0 3592 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_809
timestamp 1569543463
transform 1 0 3336 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_810
timestamp 1569543463
transform 1 0 3656 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_811
timestamp 1569543463
transform 1 0 3400 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_812
timestamp 1569543463
transform 1 0 3720 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_813
timestamp 1569543463
transform 1 0 3464 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_814
timestamp 1569543463
transform 1 0 3464 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_815
timestamp 1569543463
transform 1 0 3528 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_816
timestamp 1569543463
transform 1 0 3592 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_817
timestamp 1569543463
transform 1 0 3528 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_818
timestamp 1569543463
transform 1 0 3400 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_819
timestamp 1569543463
transform 1 0 3656 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_820
timestamp 1569543463
transform 1 0 3720 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_821
timestamp 1569543463
transform 1 0 4744 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_822
timestamp 1569543463
transform 1 0 4680 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_823
timestamp 1569543463
transform 1 0 4680 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_824
timestamp 1569543463
transform 1 0 4872 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_825
timestamp 1569543463
transform 1 0 4552 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_826
timestamp 1569543463
transform 1 0 4424 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_827
timestamp 1569543463
transform 1 0 4616 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_828
timestamp 1569543463
transform 1 0 4488 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_829
timestamp 1569543463
transform 1 0 4424 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_830
timestamp 1569543463
transform 1 0 4744 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_831
timestamp 1569543463
transform 1 0 4744 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_832
timestamp 1569543463
transform 1 0 4680 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_833
timestamp 1569543463
transform 1 0 4808 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_834
timestamp 1569543463
transform 1 0 4488 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_835
timestamp 1569543463
transform 1 0 4808 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_836
timestamp 1569543463
transform 1 0 4424 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_837
timestamp 1569543463
transform 1 0 4808 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_838
timestamp 1569543463
transform 1 0 4552 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_839
timestamp 1569543463
transform 1 0 4616 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_840
timestamp 1569543463
transform 1 0 4616 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_841
timestamp 1569543463
transform 1 0 4552 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_842
timestamp 1569543463
transform 1 0 4680 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_843
timestamp 1569543463
transform 1 0 4744 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_844
timestamp 1569543463
transform 1 0 4616 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_845
timestamp 1569543463
transform 1 0 4488 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_846
timestamp 1569543463
transform 1 0 4808 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_847
timestamp 1569543463
transform 1 0 4552 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_848
timestamp 1569543463
transform 1 0 4872 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_849
timestamp 1569543463
transform 1 0 4488 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_850
timestamp 1569543463
transform 1 0 4872 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_851
timestamp 1569543463
transform 1 0 4424 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_852
timestamp 1569543463
transform 1 0 4872 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_853
timestamp 1569543463
transform 1 0 3848 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_854
timestamp 1569543463
transform 1 0 4040 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_855
timestamp 1569543463
transform 1 0 4040 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_856
timestamp 1569543463
transform 1 0 4232 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_857
timestamp 1569543463
transform 1 0 4040 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_858
timestamp 1569543463
transform 1 0 4232 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_859
timestamp 1569543463
transform 1 0 4232 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_860
timestamp 1569543463
transform 1 0 3848 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_861
timestamp 1569543463
transform 1 0 3848 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_862
timestamp 1569543463
transform 1 0 4232 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_863
timestamp 1569543463
transform 1 0 4104 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_864
timestamp 1569543463
transform 1 0 4104 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_865
timestamp 1569543463
transform 1 0 4104 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_866
timestamp 1569543463
transform 1 0 4168 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_867
timestamp 1569543463
transform 1 0 4168 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_868
timestamp 1569543463
transform 1 0 4168 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_869
timestamp 1569543463
transform 1 0 3912 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_870
timestamp 1569543463
transform 1 0 3976 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_871
timestamp 1569543463
transform 1 0 4040 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_872
timestamp 1569543463
transform 1 0 4104 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_873
timestamp 1569543463
transform 1 0 4168 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_874
timestamp 1569543463
transform 1 0 4296 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_875
timestamp 1569543463
transform 1 0 4296 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_876
timestamp 1569543463
transform 1 0 4296 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_877
timestamp 1569543463
transform 1 0 4296 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_878
timestamp 1569543463
transform 1 0 3976 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_879
timestamp 1569543463
transform 1 0 3976 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_880
timestamp 1569543463
transform 1 0 3912 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_881
timestamp 1569543463
transform 1 0 3784 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_882
timestamp 1569543463
transform 1 0 3848 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_883
timestamp 1569543463
transform 1 0 3912 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_884
timestamp 1569543463
transform 1 0 3784 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_885
timestamp 1569543463
transform 1 0 3784 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_886
timestamp 1569543463
transform 1 0 3784 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_887
timestamp 1569543463
transform 1 0 3912 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_888
timestamp 1569543463
transform 1 0 3976 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_889
timestamp 1569543463
transform 1 0 4168 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_890
timestamp 1569543463
transform 1 0 3912 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_891
timestamp 1569543463
transform 1 0 4296 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_892
timestamp 1569543463
transform 1 0 4232 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_893
timestamp 1569543463
transform 1 0 3976 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_894
timestamp 1569543463
transform 1 0 3784 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_895
timestamp 1569543463
transform 1 0 4296 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_896
timestamp 1569543463
transform 1 0 4040 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_897
timestamp 1569543463
transform 1 0 3848 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_898
timestamp 1569543463
transform 1 0 4040 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_899
timestamp 1569543463
transform 1 0 4104 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_900
timestamp 1569543463
transform 1 0 3912 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_901
timestamp 1569543463
transform 1 0 3848 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_902
timestamp 1569543463
transform 1 0 4168 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_903
timestamp 1569543463
transform 1 0 3976 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_904
timestamp 1569543463
transform 1 0 4232 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_905
timestamp 1569543463
transform 1 0 4040 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_906
timestamp 1569543463
transform 1 0 3784 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_907
timestamp 1569543463
transform 1 0 4296 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_908
timestamp 1569543463
transform 1 0 4104 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_909
timestamp 1569543463
transform 1 0 3848 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_910
timestamp 1569543463
transform 1 0 4232 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_911
timestamp 1569543463
transform 1 0 3784 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_912
timestamp 1569543463
transform 1 0 4168 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_913
timestamp 1569543463
transform 1 0 3912 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_914
timestamp 1569543463
transform 1 0 3976 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_915
timestamp 1569543463
transform 1 0 4104 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_916
timestamp 1569543463
transform 1 0 4680 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_917
timestamp 1569543463
transform 1 0 4488 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_918
timestamp 1569543463
transform 1 0 4744 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_919
timestamp 1569543463
transform 1 0 4552 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_920
timestamp 1569543463
transform 1 0 4808 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_921
timestamp 1569543463
transform 1 0 4616 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_922
timestamp 1569543463
transform 1 0 4552 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_923
timestamp 1569543463
transform 1 0 4872 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_924
timestamp 1569543463
transform 1 0 4680 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_925
timestamp 1569543463
transform 1 0 4424 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_926
timestamp 1569543463
transform 1 0 4744 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_927
timestamp 1569543463
transform 1 0 4488 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_928
timestamp 1569543463
transform 1 0 4808 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_929
timestamp 1569543463
transform 1 0 4552 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_930
timestamp 1569543463
transform 1 0 4872 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_931
timestamp 1569543463
transform 1 0 4616 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_932
timestamp 1569543463
transform 1 0 4680 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_933
timestamp 1569543463
transform 1 0 4424 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_934
timestamp 1569543463
transform 1 0 4424 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_935
timestamp 1569543463
transform 1 0 4872 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_936
timestamp 1569543463
transform 1 0 4616 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_937
timestamp 1569543463
transform 1 0 4744 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_938
timestamp 1569543463
transform 1 0 4488 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_939
timestamp 1569543463
transform 1 0 4808 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_940
timestamp 1569543463
transform 1 0 4360 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_941
timestamp 1569543463
transform 1 0 4360 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_942
timestamp 1569543463
transform 1 0 4360 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_943
timestamp 1569543463
transform 1 0 4360 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_944
timestamp 1569543463
transform 1 0 4360 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_945
timestamp 1569543463
transform 1 0 4360 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_946
timestamp 1569543463
transform 1 0 4360 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_947
timestamp 1569543463
transform 1 0 2376 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_948
timestamp 1569543463
transform 1 0 2312 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_949
timestamp 1569543463
transform 1 0 2440 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_950
timestamp 1569543463
transform 1 0 2248 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_951
timestamp 1569543463
transform 1 0 2312 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_952
timestamp 1569543463
transform 1 0 2248 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_953
timestamp 1569543463
transform 1 0 2312 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_954
timestamp 1569543463
transform 1 0 2376 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_955
timestamp 1569543463
transform 1 0 2312 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_956
timestamp 1569543463
transform 1 0 2440 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_957
timestamp 1569543463
transform 1 0 2376 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_958
timestamp 1569543463
transform 1 0 2440 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_959
timestamp 1569543463
transform 1 0 2248 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_960
timestamp 1569543463
transform 1 0 2312 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_961
timestamp 1569543463
transform 1 0 2248 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_962
timestamp 1569543463
transform 1 0 2376 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_963
timestamp 1569543463
transform 1 0 2440 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_964
timestamp 1569543463
transform 1 0 2376 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_965
timestamp 1569543463
transform 1 0 2440 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_966
timestamp 1569543463
transform 1 0 2248 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_967
timestamp 1569543463
transform 1 0 2184 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_968
timestamp 1569543463
transform 1 0 2056 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_969
timestamp 1569543463
transform 1 0 1928 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_970
timestamp 1569543463
transform 1 0 2120 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_971
timestamp 1569543463
transform 1 0 2120 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_972
timestamp 1569543463
transform 1 0 2120 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_973
timestamp 1569543463
transform 1 0 1928 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_974
timestamp 1569543463
transform 1 0 2120 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_975
timestamp 1569543463
transform 1 0 1928 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_976
timestamp 1569543463
transform 1 0 1992 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_977
timestamp 1569543463
transform 1 0 2120 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_978
timestamp 1569543463
transform 1 0 1928 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_979
timestamp 1569543463
transform 1 0 1992 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_980
timestamp 1569543463
transform 1 0 1992 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_981
timestamp 1569543463
transform 1 0 2184 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_982
timestamp 1569543463
transform 1 0 1992 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_983
timestamp 1569543463
transform 1 0 2184 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_984
timestamp 1569543463
transform 1 0 1992 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_985
timestamp 1569543463
transform 1 0 1928 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_986
timestamp 1569543463
transform 1 0 2056 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_987
timestamp 1569543463
transform 1 0 2056 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_988
timestamp 1569543463
transform 1 0 2184 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_989
timestamp 1569543463
transform 1 0 2056 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_990
timestamp 1569543463
transform 1 0 2056 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_991
timestamp 1569543463
transform 1 0 2184 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_992
timestamp 1569543463
transform 1 0 1928 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_993
timestamp 1569543463
transform 1 0 2120 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_994
timestamp 1569543463
transform 1 0 2184 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_995
timestamp 1569543463
transform 1 0 2120 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_996
timestamp 1569543463
transform 1 0 2120 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_997
timestamp 1569543463
transform 1 0 1928 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_998
timestamp 1569543463
transform 1 0 2120 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_999
timestamp 1569543463
transform 1 0 2056 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1000
timestamp 1569543463
transform 1 0 1928 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1001
timestamp 1569543463
transform 1 0 2056 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1002
timestamp 1569543463
transform 1 0 1992 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1003
timestamp 1569543463
transform 1 0 1992 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1004
timestamp 1569543463
transform 1 0 1992 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1005
timestamp 1569543463
transform 1 0 1928 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1006
timestamp 1569543463
transform 1 0 2184 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1007
timestamp 1569543463
transform 1 0 1992 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1008
timestamp 1569543463
transform 1 0 2184 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1009
timestamp 1569543463
transform 1 0 2056 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1010
timestamp 1569543463
transform 1 0 2056 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1011
timestamp 1569543463
transform 1 0 2184 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1012
timestamp 1569543463
transform 1 0 2376 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1013
timestamp 1569543463
transform 1 0 2440 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1014
timestamp 1569543463
transform 1 0 2376 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1015
timestamp 1569543463
transform 1 0 2376 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1016
timestamp 1569543463
transform 1 0 2376 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1017
timestamp 1569543463
transform 1 0 2312 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1018
timestamp 1569543463
transform 1 0 2312 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1019
timestamp 1569543463
transform 1 0 2312 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1020
timestamp 1569543463
transform 1 0 2312 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1021
timestamp 1569543463
transform 1 0 2440 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1022
timestamp 1569543463
transform 1 0 2440 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1023
timestamp 1569543463
transform 1 0 2248 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1024
timestamp 1569543463
transform 1 0 2248 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1025
timestamp 1569543463
transform 1 0 2248 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1026
timestamp 1569543463
transform 1 0 2248 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1027
timestamp 1569543463
transform 1 0 2440 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1028
timestamp 1569543463
transform 1 0 1864 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1029
timestamp 1569543463
transform 1 0 1864 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_1030
timestamp 1569543463
transform 1 0 1736 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1031
timestamp 1569543463
transform 1 0 1736 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_1032
timestamp 1569543463
transform 1 0 1864 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_1033
timestamp 1569543463
transform 1 0 1800 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_1034
timestamp 1569543463
transform 1 0 1672 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_1035
timestamp 1569543463
transform 1 0 1672 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_1036
timestamp 1569543463
transform 1 0 1672 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1037
timestamp 1569543463
transform 1 0 1672 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1038
timestamp 1569543463
transform 1 0 1736 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1039
timestamp 1569543463
transform 1 0 1800 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_1040
timestamp 1569543463
transform 1 0 1800 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_1041
timestamp 1569543463
transform 1 0 1864 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1042
timestamp 1569543463
transform 1 0 1608 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_1043
timestamp 1569543463
transform 1 0 1608 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1044
timestamp 1569543463
transform 1 0 1608 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1045
timestamp 1569543463
transform 1 0 1736 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_1046
timestamp 1569543463
transform 1 0 1864 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_1047
timestamp 1569543463
transform 1 0 1800 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1048
timestamp 1569543463
transform 1 0 1800 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1049
timestamp 1569543463
transform 1 0 1736 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_1050
timestamp 1569543463
transform 1 0 1544 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_1051
timestamp 1569543463
transform 1 0 1544 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1052
timestamp 1569543463
transform 1 0 1480 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_1053
timestamp 1569543463
transform 1 0 1544 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1054
timestamp 1569543463
transform 1 0 1544 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1055
timestamp 1569543463
transform 1 0 1544 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1056
timestamp 1569543463
transform 1 0 1544 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1057
timestamp 1569543463
transform 1 0 1288 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1058
timestamp 1569543463
transform 1 0 1416 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1059
timestamp 1569543463
transform 1 0 1416 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1060
timestamp 1569543463
transform 1 0 1416 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1061
timestamp 1569543463
transform 1 0 1416 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1062
timestamp 1569543463
transform 1 0 1480 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1063
timestamp 1569543463
transform 1 0 1480 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1064
timestamp 1569543463
transform 1 0 1480 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1065
timestamp 1569543463
transform 1 0 1352 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1066
timestamp 1569543463
transform 1 0 1352 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1067
timestamp 1569543463
transform 1 0 1352 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1068
timestamp 1569543463
transform 1 0 1480 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1069
timestamp 1569543463
transform 1 0 1288 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1070
timestamp 1569543463
transform 1 0 1736 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1071
timestamp 1569543463
transform 1 0 1608 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1072
timestamp 1569543463
transform 1 0 1608 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1073
timestamp 1569543463
transform 1 0 1608 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1074
timestamp 1569543463
transform 1 0 1608 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1075
timestamp 1569543463
transform 1 0 1800 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1076
timestamp 1569543463
transform 1 0 1736 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1077
timestamp 1569543463
transform 1 0 1800 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1078
timestamp 1569543463
transform 1 0 1736 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1079
timestamp 1569543463
transform 1 0 1736 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1080
timestamp 1569543463
transform 1 0 1672 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1081
timestamp 1569543463
transform 1 0 1672 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1082
timestamp 1569543463
transform 1 0 1672 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1083
timestamp 1569543463
transform 1 0 1672 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1084
timestamp 1569543463
transform 1 0 1864 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_1085
timestamp 1569543463
transform 1 0 1864 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_1086
timestamp 1569543463
transform 1 0 1864 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1087
timestamp 1569543463
transform 1 0 1800 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_1088
timestamp 1569543463
transform 1 0 1864 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1089
timestamp 1569543463
transform 1 0 1800 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1090
timestamp 1569543463
transform 1 0 1736 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1091
timestamp 1569543463
transform 1 0 1800 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1092
timestamp 1569543463
transform 1 0 1736 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1093
timestamp 1569543463
transform 1 0 1864 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1094
timestamp 1569543463
transform 1 0 1672 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1095
timestamp 1569543463
transform 1 0 1864 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1096
timestamp 1569543463
transform 1 0 1672 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1097
timestamp 1569543463
transform 1 0 1736 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1098
timestamp 1569543463
transform 1 0 1864 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1099
timestamp 1569543463
transform 1 0 1864 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1100
timestamp 1569543463
transform 1 0 1608 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1101
timestamp 1569543463
transform 1 0 1800 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1102
timestamp 1569543463
transform 1 0 1672 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1103
timestamp 1569543463
transform 1 0 1736 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1104
timestamp 1569543463
transform 1 0 1608 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1105
timestamp 1569543463
transform 1 0 1608 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1106
timestamp 1569543463
transform 1 0 1800 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1107
timestamp 1569543463
transform 1 0 1800 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1108
timestamp 1569543463
transform 1 0 1672 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1109
timestamp 1569543463
transform 1 0 1608 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1110
timestamp 1569543463
transform 1 0 1544 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1111
timestamp 1569543463
transform 1 0 1416 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1112
timestamp 1569543463
transform 1 0 1480 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1113
timestamp 1569543463
transform 1 0 1544 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1114
timestamp 1569543463
transform 1 0 1288 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1115
timestamp 1569543463
transform 1 0 1416 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1116
timestamp 1569543463
transform 1 0 1544 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1117
timestamp 1569543463
transform 1 0 1416 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1118
timestamp 1569543463
transform 1 0 1480 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1119
timestamp 1569543463
transform 1 0 1352 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1120
timestamp 1569543463
transform 1 0 1352 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1121
timestamp 1569543463
transform 1 0 1288 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1122
timestamp 1569543463
transform 1 0 1480 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1123
timestamp 1569543463
transform 1 0 1352 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1124
timestamp 1569543463
transform 1 0 1544 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1125
timestamp 1569543463
transform 1 0 1352 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1126
timestamp 1569543463
transform 1 0 1480 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1127
timestamp 1569543463
transform 1 0 1288 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1128
timestamp 1569543463
transform 1 0 1288 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1129
timestamp 1569543463
transform 1 0 1416 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1130
timestamp 1569543463
transform 1 0 1352 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1131
timestamp 1569543463
transform 1 0 1544 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1132
timestamp 1569543463
transform 1 0 1544 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1133
timestamp 1569543463
transform 1 0 1416 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1134
timestamp 1569543463
transform 1 0 1288 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1135
timestamp 1569543463
transform 1 0 1480 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1136
timestamp 1569543463
transform 1 0 1288 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1137
timestamp 1569543463
transform 1 0 1288 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1138
timestamp 1569543463
transform 1 0 1416 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1139
timestamp 1569543463
transform 1 0 1480 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1140
timestamp 1569543463
transform 1 0 1416 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1141
timestamp 1569543463
transform 1 0 1544 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1142
timestamp 1569543463
transform 1 0 1288 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1143
timestamp 1569543463
transform 1 0 1416 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1144
timestamp 1569543463
transform 1 0 1480 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1145
timestamp 1569543463
transform 1 0 1544 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1146
timestamp 1569543463
transform 1 0 1288 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1147
timestamp 1569543463
transform 1 0 1352 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1148
timestamp 1569543463
transform 1 0 1416 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1149
timestamp 1569543463
transform 1 0 1352 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1150
timestamp 1569543463
transform 1 0 1352 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1151
timestamp 1569543463
transform 1 0 1480 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1152
timestamp 1569543463
transform 1 0 1480 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1153
timestamp 1569543463
transform 1 0 1544 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1154
timestamp 1569543463
transform 1 0 1352 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1155
timestamp 1569543463
transform 1 0 1672 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1156
timestamp 1569543463
transform 1 0 1672 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1157
timestamp 1569543463
transform 1 0 1736 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1158
timestamp 1569543463
transform 1 0 1736 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1159
timestamp 1569543463
transform 1 0 1736 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1160
timestamp 1569543463
transform 1 0 1736 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1161
timestamp 1569543463
transform 1 0 1736 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1162
timestamp 1569543463
transform 1 0 1800 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1163
timestamp 1569543463
transform 1 0 1800 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1164
timestamp 1569543463
transform 1 0 1800 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1165
timestamp 1569543463
transform 1 0 1800 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1166
timestamp 1569543463
transform 1 0 1800 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1167
timestamp 1569543463
transform 1 0 1672 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1168
timestamp 1569543463
transform 1 0 1608 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1169
timestamp 1569543463
transform 1 0 1864 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1170
timestamp 1569543463
transform 1 0 1864 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1171
timestamp 1569543463
transform 1 0 1608 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1172
timestamp 1569543463
transform 1 0 1864 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1173
timestamp 1569543463
transform 1 0 1672 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1174
timestamp 1569543463
transform 1 0 1608 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1175
timestamp 1569543463
transform 1 0 1864 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1176
timestamp 1569543463
transform 1 0 1864 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1177
timestamp 1569543463
transform 1 0 1608 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1178
timestamp 1569543463
transform 1 0 1672 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1179
timestamp 1569543463
transform 1 0 1608 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1180
timestamp 1569543463
transform 1 0 2248 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1181
timestamp 1569543463
transform 1 0 2376 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1182
timestamp 1569543463
transform 1 0 2440 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1183
timestamp 1569543463
transform 1 0 2376 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1184
timestamp 1569543463
transform 1 0 2440 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1185
timestamp 1569543463
transform 1 0 2376 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1186
timestamp 1569543463
transform 1 0 2312 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1187
timestamp 1569543463
transform 1 0 2312 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1188
timestamp 1569543463
transform 1 0 2376 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1189
timestamp 1569543463
transform 1 0 2248 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1190
timestamp 1569543463
transform 1 0 2312 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1191
timestamp 1569543463
transform 1 0 2312 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1192
timestamp 1569543463
transform 1 0 2248 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1193
timestamp 1569543463
transform 1 0 2248 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1194
timestamp 1569543463
transform 1 0 2440 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1195
timestamp 1569543463
transform 1 0 2440 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1196
timestamp 1569543463
transform 1 0 1992 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1197
timestamp 1569543463
transform 1 0 1992 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1198
timestamp 1569543463
transform 1 0 2056 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1199
timestamp 1569543463
transform 1 0 2120 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1200
timestamp 1569543463
transform 1 0 2184 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1201
timestamp 1569543463
transform 1 0 2184 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1202
timestamp 1569543463
transform 1 0 1992 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1203
timestamp 1569543463
transform 1 0 1992 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1204
timestamp 1569543463
transform 1 0 1928 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1205
timestamp 1569543463
transform 1 0 1928 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1206
timestamp 1569543463
transform 1 0 2120 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1207
timestamp 1569543463
transform 1 0 2056 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1208
timestamp 1569543463
transform 1 0 2056 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1209
timestamp 1569543463
transform 1 0 2056 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1210
timestamp 1569543463
transform 1 0 1928 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1211
timestamp 1569543463
transform 1 0 1928 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1212
timestamp 1569543463
transform 1 0 2120 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1213
timestamp 1569543463
transform 1 0 2120 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1214
timestamp 1569543463
transform 1 0 2184 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1215
timestamp 1569543463
transform 1 0 2184 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1216
timestamp 1569543463
transform 1 0 1928 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1217
timestamp 1569543463
transform 1 0 2120 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1218
timestamp 1569543463
transform 1 0 1928 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1219
timestamp 1569543463
transform 1 0 2120 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1220
timestamp 1569543463
transform 1 0 2120 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1221
timestamp 1569543463
transform 1 0 2120 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1222
timestamp 1569543463
transform 1 0 2120 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1223
timestamp 1569543463
transform 1 0 2184 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1224
timestamp 1569543463
transform 1 0 2184 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1225
timestamp 1569543463
transform 1 0 2184 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1226
timestamp 1569543463
transform 1 0 1992 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1227
timestamp 1569543463
transform 1 0 1992 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1228
timestamp 1569543463
transform 1 0 1992 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1229
timestamp 1569543463
transform 1 0 1992 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1230
timestamp 1569543463
transform 1 0 1992 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1231
timestamp 1569543463
transform 1 0 2056 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1232
timestamp 1569543463
transform 1 0 2056 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1233
timestamp 1569543463
transform 1 0 2056 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1234
timestamp 1569543463
transform 1 0 2056 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1235
timestamp 1569543463
transform 1 0 2056 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1236
timestamp 1569543463
transform 1 0 2184 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1237
timestamp 1569543463
transform 1 0 2184 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1238
timestamp 1569543463
transform 1 0 1928 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1239
timestamp 1569543463
transform 1 0 1928 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1240
timestamp 1569543463
transform 1 0 1928 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1241
timestamp 1569543463
transform 1 0 2376 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1242
timestamp 1569543463
transform 1 0 2376 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1243
timestamp 1569543463
transform 1 0 2376 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1244
timestamp 1569543463
transform 1 0 2376 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1245
timestamp 1569543463
transform 1 0 2376 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1246
timestamp 1569543463
transform 1 0 2440 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1247
timestamp 1569543463
transform 1 0 2440 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1248
timestamp 1569543463
transform 1 0 2440 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1249
timestamp 1569543463
transform 1 0 2440 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1250
timestamp 1569543463
transform 1 0 2440 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1251
timestamp 1569543463
transform 1 0 2248 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1252
timestamp 1569543463
transform 1 0 2312 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1253
timestamp 1569543463
transform 1 0 2312 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1254
timestamp 1569543463
transform 1 0 2312 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1255
timestamp 1569543463
transform 1 0 2312 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1256
timestamp 1569543463
transform 1 0 2312 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1257
timestamp 1569543463
transform 1 0 2248 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1258
timestamp 1569543463
transform 1 0 2248 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1259
timestamp 1569543463
transform 1 0 2248 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1260
timestamp 1569543463
transform 1 0 2248 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1261
timestamp 1569543463
transform 1 0 1672 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1262
timestamp 1569543463
transform 1 0 2312 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1263
timestamp 1569543463
transform 1 0 1352 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1264
timestamp 1569543463
transform 1 0 1992 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1265
timestamp 1569543463
transform 1 0 1416 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1266
timestamp 1569543463
transform 1 0 2056 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1267
timestamp 1569543463
transform 1 0 1480 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1268
timestamp 1569543463
transform 1 0 2120 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1269
timestamp 1569543463
transform 1 0 1544 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1270
timestamp 1569543463
transform 1 0 2184 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1271
timestamp 1569543463
transform 1 0 1608 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1272
timestamp 1569543463
transform 1 0 2248 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1273
timestamp 1569543463
transform 1 0 1736 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1274
timestamp 1569543463
transform 1 0 2376 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1275
timestamp 1569543463
transform 1 0 1800 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1276
timestamp 1569543463
transform 1 0 2440 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1277
timestamp 1569543463
transform 1 0 1864 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1278
timestamp 1569543463
transform 1 0 1288 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1279
timestamp 1569543463
transform 1 0 1928 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1280
timestamp 1569543463
transform 1 0 1224 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_1281
timestamp 1569543463
transform 1 0 584 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1282
timestamp 1569543463
transform 1 0 968 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1283
timestamp 1569543463
transform 1 0 968 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1284
timestamp 1569543463
transform 1 0 1160 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1285
timestamp 1569543463
transform 1 0 1224 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1286
timestamp 1569543463
transform 1 0 1224 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1287
timestamp 1569543463
transform 1 0 1032 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1288
timestamp 1569543463
transform 1 0 1096 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1289
timestamp 1569543463
transform 1 0 1096 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_1290
timestamp 1569543463
transform 1 0 1032 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1291
timestamp 1569543463
transform 1 0 1032 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1292
timestamp 1569543463
transform 1 0 1096 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1293
timestamp 1569543463
transform 1 0 1096 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1294
timestamp 1569543463
transform 1 0 1224 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1295
timestamp 1569543463
transform 1 0 1160 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_1296
timestamp 1569543463
transform 1 0 1224 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1297
timestamp 1569543463
transform 1 0 1160 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_1298
timestamp 1569543463
transform 1 0 1160 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1299
timestamp 1569543463
transform 1 0 904 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_1300
timestamp 1569543463
transform 1 0 904 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1301
timestamp 1569543463
transform 1 0 904 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1302
timestamp 1569543463
transform 1 0 904 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1303
timestamp 1569543463
transform 1 0 904 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1304
timestamp 1569543463
transform 1 0 904 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1305
timestamp 1569543463
transform 1 0 840 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1306
timestamp 1569543463
transform 1 0 840 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1307
timestamp 1569543463
transform 1 0 840 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1308
timestamp 1569543463
transform 1 0 840 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1309
timestamp 1569543463
transform 1 0 840 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1310
timestamp 1569543463
transform 1 0 712 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1311
timestamp 1569543463
transform 1 0 712 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1312
timestamp 1569543463
transform 1 0 712 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1313
timestamp 1569543463
transform 1 0 776 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1314
timestamp 1569543463
transform 1 0 776 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1315
timestamp 1569543463
transform 1 0 776 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1316
timestamp 1569543463
transform 1 0 776 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1317
timestamp 1569543463
transform 1 0 1032 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1318
timestamp 1569543463
transform 1 0 1032 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1319
timestamp 1569543463
transform 1 0 1032 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1320
timestamp 1569543463
transform 1 0 1096 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1321
timestamp 1569543463
transform 1 0 1096 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1322
timestamp 1569543463
transform 1 0 1096 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1323
timestamp 1569543463
transform 1 0 1096 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1324
timestamp 1569543463
transform 1 0 1096 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1325
timestamp 1569543463
transform 1 0 1160 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1326
timestamp 1569543463
transform 1 0 1160 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1327
timestamp 1569543463
transform 1 0 1160 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1328
timestamp 1569543463
transform 1 0 1160 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1329
timestamp 1569543463
transform 1 0 1160 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1330
timestamp 1569543463
transform 1 0 968 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1331
timestamp 1569543463
transform 1 0 968 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1332
timestamp 1569543463
transform 1 0 968 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1333
timestamp 1569543463
transform 1 0 968 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1334
timestamp 1569543463
transform 1 0 968 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1335
timestamp 1569543463
transform 1 0 1224 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1336
timestamp 1569543463
transform 1 0 1224 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1337
timestamp 1569543463
transform 1 0 1224 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_1338
timestamp 1569543463
transform 1 0 1224 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1339
timestamp 1569543463
transform 1 0 1224 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1340
timestamp 1569543463
transform 1 0 1032 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_1341
timestamp 1569543463
transform 1 0 1032 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_1342
timestamp 1569543463
transform 1 0 648 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_1343
timestamp 1569543463
transform 1 0 648 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_1344
timestamp 1569543463
transform 1 0 1160 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1345
timestamp 1569543463
transform 1 0 1224 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_1346
timestamp 1569543463
transform 1 0 1160 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1347
timestamp 1569543463
transform 1 0 1096 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1348
timestamp 1569543463
transform 1 0 1160 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1349
timestamp 1569543463
transform 1 0 1096 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1350
timestamp 1569543463
transform 1 0 1032 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1351
timestamp 1569543463
transform 1 0 968 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1352
timestamp 1569543463
transform 1 0 1160 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1353
timestamp 1569543463
transform 1 0 1160 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1354
timestamp 1569543463
transform 1 0 1096 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1355
timestamp 1569543463
transform 1 0 968 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1356
timestamp 1569543463
transform 1 0 1096 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1357
timestamp 1569543463
transform 1 0 1096 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1358
timestamp 1569543463
transform 1 0 1032 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1359
timestamp 1569543463
transform 1 0 968 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1360
timestamp 1569543463
transform 1 0 1224 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1361
timestamp 1569543463
transform 1 0 1032 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1362
timestamp 1569543463
transform 1 0 968 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1363
timestamp 1569543463
transform 1 0 1224 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1364
timestamp 1569543463
transform 1 0 968 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1365
timestamp 1569543463
transform 1 0 1224 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1366
timestamp 1569543463
transform 1 0 1032 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1367
timestamp 1569543463
transform 1 0 1224 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1368
timestamp 1569543463
transform 1 0 1224 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1369
timestamp 1569543463
transform 1 0 1160 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1370
timestamp 1569543463
transform 1 0 1032 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1371
timestamp 1569543463
transform 1 0 776 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1372
timestamp 1569543463
transform 1 0 840 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1373
timestamp 1569543463
transform 1 0 904 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1374
timestamp 1569543463
transform 1 0 840 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1375
timestamp 1569543463
transform 1 0 712 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1376
timestamp 1569543463
transform 1 0 904 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1377
timestamp 1569543463
transform 1 0 776 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1378
timestamp 1569543463
transform 1 0 712 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1379
timestamp 1569543463
transform 1 0 904 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1380
timestamp 1569543463
transform 1 0 712 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1381
timestamp 1569543463
transform 1 0 840 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1382
timestamp 1569543463
transform 1 0 904 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1383
timestamp 1569543463
transform 1 0 712 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1384
timestamp 1569543463
transform 1 0 840 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1385
timestamp 1569543463
transform 1 0 904 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1386
timestamp 1569543463
transform 1 0 712 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1387
timestamp 1569543463
transform 1 0 840 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1388
timestamp 1569543463
transform 1 0 776 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1389
timestamp 1569543463
transform 1 0 776 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1390
timestamp 1569543463
transform 1 0 776 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1391
timestamp 1569543463
transform 1 0 776 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1392
timestamp 1569543463
transform 1 0 904 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1393
timestamp 1569543463
transform 1 0 776 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1394
timestamp 1569543463
transform 1 0 840 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1395
timestamp 1569543463
transform 1 0 904 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1396
timestamp 1569543463
transform 1 0 776 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1397
timestamp 1569543463
transform 1 0 840 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1398
timestamp 1569543463
transform 1 0 712 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1399
timestamp 1569543463
transform 1 0 840 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1400
timestamp 1569543463
transform 1 0 776 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1401
timestamp 1569543463
transform 1 0 712 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1402
timestamp 1569543463
transform 1 0 904 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1403
timestamp 1569543463
transform 1 0 840 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1404
timestamp 1569543463
transform 1 0 712 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1405
timestamp 1569543463
transform 1 0 904 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1406
timestamp 1569543463
transform 1 0 712 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1407
timestamp 1569543463
transform 1 0 840 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1408
timestamp 1569543463
transform 1 0 712 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1409
timestamp 1569543463
transform 1 0 776 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1410
timestamp 1569543463
transform 1 0 904 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1411
timestamp 1569543463
transform 1 0 1224 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1412
timestamp 1569543463
transform 1 0 1096 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1413
timestamp 1569543463
transform 1 0 1096 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1414
timestamp 1569543463
transform 1 0 1224 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1415
timestamp 1569543463
transform 1 0 1096 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1416
timestamp 1569543463
transform 1 0 1096 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1417
timestamp 1569543463
transform 1 0 1224 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1418
timestamp 1569543463
transform 1 0 1224 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1419
timestamp 1569543463
transform 1 0 1096 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1420
timestamp 1569543463
transform 1 0 1032 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1421
timestamp 1569543463
transform 1 0 1160 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1422
timestamp 1569543463
transform 1 0 968 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1423
timestamp 1569543463
transform 1 0 1032 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1424
timestamp 1569543463
transform 1 0 1160 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1425
timestamp 1569543463
transform 1 0 968 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1426
timestamp 1569543463
transform 1 0 1160 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1427
timestamp 1569543463
transform 1 0 1032 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1428
timestamp 1569543463
transform 1 0 1160 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1429
timestamp 1569543463
transform 1 0 968 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1430
timestamp 1569543463
transform 1 0 1160 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1431
timestamp 1569543463
transform 1 0 968 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1432
timestamp 1569543463
transform 1 0 1224 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1433
timestamp 1569543463
transform 1 0 968 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1434
timestamp 1569543463
transform 1 0 1032 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1435
timestamp 1569543463
transform 1 0 1032 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1436
timestamp 1569543463
transform 1 0 392 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1437
timestamp 1569543463
transform 1 0 584 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1438
timestamp 1569543463
transform 1 0 520 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1439
timestamp 1569543463
transform 1 0 520 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1440
timestamp 1569543463
transform 1 0 392 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1441
timestamp 1569543463
transform 1 0 456 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1442
timestamp 1569543463
transform 1 0 584 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1443
timestamp 1569543463
transform 1 0 520 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1444
timestamp 1569543463
transform 1 0 456 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1445
timestamp 1569543463
transform 1 0 520 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1446
timestamp 1569543463
transform 1 0 456 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1447
timestamp 1569543463
transform 1 0 584 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1448
timestamp 1569543463
transform 1 0 584 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1449
timestamp 1569543463
transform 1 0 584 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1450
timestamp 1569543463
transform 1 0 392 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1451
timestamp 1569543463
transform 1 0 456 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1452
timestamp 1569543463
transform 1 0 520 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1453
timestamp 1569543463
transform 1 0 328 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1454
timestamp 1569543463
transform 1 0 264 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1455
timestamp 1569543463
transform 1 0 328 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1456
timestamp 1569543463
transform 1 0 328 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1457
timestamp 1569543463
transform 1 0 200 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1458
timestamp 1569543463
transform 1 0 136 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1459
timestamp 1569543463
transform 1 0 264 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1460
timestamp 1569543463
transform 1 0 200 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1461
timestamp 1569543463
transform 1 0 72 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1462
timestamp 1569543463
transform 1 0 72 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1463
timestamp 1569543463
transform 1 0 200 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1464
timestamp 1569543463
transform 1 0 136 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1465
timestamp 1569543463
transform 1 0 328 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1466
timestamp 1569543463
transform 1 0 72 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1467
timestamp 1569543463
transform 1 0 200 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1468
timestamp 1569543463
transform 1 0 328 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1469
timestamp 1569543463
transform 1 0 264 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1470
timestamp 1569543463
transform 1 0 136 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1471
timestamp 1569543463
transform 1 0 264 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1472
timestamp 1569543463
transform 1 0 328 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1473
timestamp 1569543463
transform 1 0 328 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1474
timestamp 1569543463
transform 1 0 264 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1475
timestamp 1569543463
transform 1 0 136 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1476
timestamp 1569543463
transform 1 0 264 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1477
timestamp 1569543463
transform 1 0 200 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1478
timestamp 1569543463
transform 1 0 456 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1479
timestamp 1569543463
transform 1 0 584 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1480
timestamp 1569543463
transform 1 0 456 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1481
timestamp 1569543463
transform 1 0 456 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1482
timestamp 1569543463
transform 1 0 456 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1483
timestamp 1569543463
transform 1 0 584 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1484
timestamp 1569543463
transform 1 0 456 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1485
timestamp 1569543463
transform 1 0 392 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1486
timestamp 1569543463
transform 1 0 392 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1487
timestamp 1569543463
transform 1 0 520 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1488
timestamp 1569543463
transform 1 0 584 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1489
timestamp 1569543463
transform 1 0 520 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1490
timestamp 1569543463
transform 1 0 520 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1491
timestamp 1569543463
transform 1 0 392 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1492
timestamp 1569543463
transform 1 0 520 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1493
timestamp 1569543463
transform 1 0 520 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1494
timestamp 1569543463
transform 1 0 392 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1495
timestamp 1569543463
transform 1 0 584 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1496
timestamp 1569543463
transform 1 0 584 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1497
timestamp 1569543463
transform 1 0 392 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1498
timestamp 1569543463
transform 1 0 392 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1499
timestamp 1569543463
transform 1 0 392 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1500
timestamp 1569543463
transform 1 0 456 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1501
timestamp 1569543463
transform 1 0 520 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1502
timestamp 1569543463
transform 1 0 456 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1503
timestamp 1569543463
transform 1 0 520 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1504
timestamp 1569543463
transform 1 0 456 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1505
timestamp 1569543463
transform 1 0 456 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1506
timestamp 1569543463
transform 1 0 392 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1507
timestamp 1569543463
transform 1 0 584 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1508
timestamp 1569543463
transform 1 0 520 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1509
timestamp 1569543463
transform 1 0 584 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1510
timestamp 1569543463
transform 1 0 520 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1511
timestamp 1569543463
transform 1 0 584 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1512
timestamp 1569543463
transform 1 0 456 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1513
timestamp 1569543463
transform 1 0 392 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1514
timestamp 1569543463
transform 1 0 520 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1515
timestamp 1569543463
transform 1 0 584 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1516
timestamp 1569543463
transform 1 0 392 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1517
timestamp 1569543463
transform 1 0 584 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1518
timestamp 1569543463
transform 1 0 200 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1519
timestamp 1569543463
transform 1 0 200 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1520
timestamp 1569543463
transform 1 0 328 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1521
timestamp 1569543463
transform 1 0 72 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1522
timestamp 1569543463
transform 1 0 136 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1523
timestamp 1569543463
transform 1 0 72 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1524
timestamp 1569543463
transform 1 0 264 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1525
timestamp 1569543463
transform 1 0 200 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1526
timestamp 1569543463
transform 1 0 136 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1527
timestamp 1569543463
transform 1 0 328 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1528
timestamp 1569543463
transform 1 0 328 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1529
timestamp 1569543463
transform 1 0 136 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1530
timestamp 1569543463
transform 1 0 72 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1531
timestamp 1569543463
transform 1 0 136 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1532
timestamp 1569543463
transform 1 0 72 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1533
timestamp 1569543463
transform 1 0 328 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1534
timestamp 1569543463
transform 1 0 264 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1535
timestamp 1569543463
transform 1 0 264 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1536
timestamp 1569543463
transform 1 0 200 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1537
timestamp 1569543463
transform 1 0 72 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1538
timestamp 1569543463
transform 1 0 328 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1539
timestamp 1569543463
transform 1 0 200 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1540
timestamp 1569543463
transform 1 0 264 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1541
timestamp 1569543463
transform 1 0 264 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1542
timestamp 1569543463
transform 1 0 136 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1543
timestamp 1569543463
transform 1 0 136 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1544
timestamp 1569543463
transform 1 0 200 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1545
timestamp 1569543463
transform 1 0 264 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1546
timestamp 1569543463
transform 1 0 72 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1547
timestamp 1569543463
transform 1 0 136 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1548
timestamp 1569543463
transform 1 0 328 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1549
timestamp 1569543463
transform 1 0 264 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1550
timestamp 1569543463
transform 1 0 200 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1551
timestamp 1569543463
transform 1 0 328 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1552
timestamp 1569543463
transform 1 0 72 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1553
timestamp 1569543463
transform 1 0 328 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1554
timestamp 1569543463
transform 1 0 200 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1555
timestamp 1569543463
transform 1 0 136 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1556
timestamp 1569543463
transform 1 0 264 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1557
timestamp 1569543463
transform 1 0 328 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1558
timestamp 1569543463
transform 1 0 264 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1559
timestamp 1569543463
transform 1 0 72 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1560
timestamp 1569543463
transform 1 0 72 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1561
timestamp 1569543463
transform 1 0 136 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1562
timestamp 1569543463
transform 1 0 200 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1563
timestamp 1569543463
transform 1 0 392 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1564
timestamp 1569543463
transform 1 0 456 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1565
timestamp 1569543463
transform 1 0 456 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1566
timestamp 1569543463
transform 1 0 584 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1567
timestamp 1569543463
transform 1 0 456 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1568
timestamp 1569543463
transform 1 0 584 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1569
timestamp 1569543463
transform 1 0 520 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1570
timestamp 1569543463
transform 1 0 456 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1571
timestamp 1569543463
transform 1 0 584 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1572
timestamp 1569543463
transform 1 0 392 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1573
timestamp 1569543463
transform 1 0 584 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1574
timestamp 1569543463
transform 1 0 392 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1575
timestamp 1569543463
transform 1 0 520 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1576
timestamp 1569543463
transform 1 0 392 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1577
timestamp 1569543463
transform 1 0 520 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1578
timestamp 1569543463
transform 1 0 520 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1579
timestamp 1569543463
transform 1 0 968 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1580
timestamp 1569543463
transform 1 0 1096 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1581
timestamp 1569543463
transform 1 0 1096 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1582
timestamp 1569543463
transform 1 0 1096 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1583
timestamp 1569543463
transform 1 0 968 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1584
timestamp 1569543463
transform 1 0 1160 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1585
timestamp 1569543463
transform 1 0 1160 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1586
timestamp 1569543463
transform 1 0 1224 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1587
timestamp 1569543463
transform 1 0 1160 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1588
timestamp 1569543463
transform 1 0 1032 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1589
timestamp 1569543463
transform 1 0 968 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1590
timestamp 1569543463
transform 1 0 1096 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1591
timestamp 1569543463
transform 1 0 1032 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1592
timestamp 1569543463
transform 1 0 1160 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1593
timestamp 1569543463
transform 1 0 1032 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1594
timestamp 1569543463
transform 1 0 968 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1595
timestamp 1569543463
transform 1 0 1224 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1596
timestamp 1569543463
transform 1 0 1096 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1597
timestamp 1569543463
transform 1 0 1032 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1598
timestamp 1569543463
transform 1 0 1224 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1599
timestamp 1569543463
transform 1 0 1160 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1600
timestamp 1569543463
transform 1 0 1224 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1601
timestamp 1569543463
transform 1 0 1224 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1602
timestamp 1569543463
transform 1 0 968 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1603
timestamp 1569543463
transform 1 0 1032 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1604
timestamp 1569543463
transform 1 0 840 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1605
timestamp 1569543463
transform 1 0 776 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1606
timestamp 1569543463
transform 1 0 840 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1607
timestamp 1569543463
transform 1 0 776 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1608
timestamp 1569543463
transform 1 0 712 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1609
timestamp 1569543463
transform 1 0 712 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1610
timestamp 1569543463
transform 1 0 840 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1611
timestamp 1569543463
transform 1 0 712 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1612
timestamp 1569543463
transform 1 0 712 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1613
timestamp 1569543463
transform 1 0 904 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1614
timestamp 1569543463
transform 1 0 776 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1615
timestamp 1569543463
transform 1 0 712 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1616
timestamp 1569543463
transform 1 0 776 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1617
timestamp 1569543463
transform 1 0 904 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1618
timestamp 1569543463
transform 1 0 776 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1619
timestamp 1569543463
transform 1 0 840 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1620
timestamp 1569543463
transform 1 0 904 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1621
timestamp 1569543463
transform 1 0 904 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1622
timestamp 1569543463
transform 1 0 840 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1623
timestamp 1569543463
transform 1 0 904 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1624
timestamp 1569543463
transform 1 0 904 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1625
timestamp 1569543463
transform 1 0 776 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1626
timestamp 1569543463
transform 1 0 840 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1627
timestamp 1569543463
transform 1 0 840 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1628
timestamp 1569543463
transform 1 0 840 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1629
timestamp 1569543463
transform 1 0 776 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1630
timestamp 1569543463
transform 1 0 712 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1631
timestamp 1569543463
transform 1 0 904 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1632
timestamp 1569543463
transform 1 0 840 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1633
timestamp 1569543463
transform 1 0 776 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1634
timestamp 1569543463
transform 1 0 904 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1635
timestamp 1569543463
transform 1 0 712 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1636
timestamp 1569543463
transform 1 0 904 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1637
timestamp 1569543463
transform 1 0 712 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1638
timestamp 1569543463
transform 1 0 712 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1639
timestamp 1569543463
transform 1 0 776 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1640
timestamp 1569543463
transform 1 0 1224 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1641
timestamp 1569543463
transform 1 0 968 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1642
timestamp 1569543463
transform 1 0 1160 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1643
timestamp 1569543463
transform 1 0 1032 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1644
timestamp 1569543463
transform 1 0 1224 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1645
timestamp 1569543463
transform 1 0 968 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1646
timestamp 1569543463
transform 1 0 1096 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1647
timestamp 1569543463
transform 1 0 1032 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1648
timestamp 1569543463
transform 1 0 1096 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1649
timestamp 1569543463
transform 1 0 1032 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1650
timestamp 1569543463
transform 1 0 1032 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1651
timestamp 1569543463
transform 1 0 1096 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1652
timestamp 1569543463
transform 1 0 1096 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1653
timestamp 1569543463
transform 1 0 1160 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1654
timestamp 1569543463
transform 1 0 1160 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1655
timestamp 1569543463
transform 1 0 1160 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1656
timestamp 1569543463
transform 1 0 1224 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1657
timestamp 1569543463
transform 1 0 968 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1658
timestamp 1569543463
transform 1 0 1224 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1659
timestamp 1569543463
transform 1 0 968 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1660
timestamp 1569543463
transform 1 0 648 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1661
timestamp 1569543463
transform 1 0 648 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1662
timestamp 1569543463
transform 1 0 648 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1663
timestamp 1569543463
transform 1 0 648 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1664
timestamp 1569543463
transform 1 0 648 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1665
timestamp 1569543463
transform 1 0 648 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1666
timestamp 1569543463
transform 1 0 648 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1667
timestamp 1569543463
transform 1 0 648 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1668
timestamp 1569543463
transform 1 0 648 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1669
timestamp 1569543463
transform 1 0 648 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1670
timestamp 1569543463
transform 1 0 648 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1671
timestamp 1569543463
transform 1 0 648 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1672
timestamp 1569543463
transform 1 0 648 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1673
timestamp 1569543463
transform 1 0 648 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1674
timestamp 1569543463
transform 1 0 648 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1675
timestamp 1569543463
transform 1 0 648 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1676
timestamp 1569543463
transform 1 0 648 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1677
timestamp 1569543463
transform 1 0 648 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1678
timestamp 1569543463
transform 1 0 648 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1679
timestamp 1569543463
transform 1 0 2248 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1680
timestamp 1569543463
transform 1 0 2376 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1681
timestamp 1569543463
transform 1 0 2376 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1682
timestamp 1569543463
transform 1 0 2312 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1683
timestamp 1569543463
transform 1 0 2248 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1684
timestamp 1569543463
transform 1 0 2440 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1685
timestamp 1569543463
transform 1 0 2248 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1686
timestamp 1569543463
transform 1 0 2312 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1687
timestamp 1569543463
transform 1 0 2248 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1688
timestamp 1569543463
transform 1 0 2440 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1689
timestamp 1569543463
transform 1 0 2312 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1690
timestamp 1569543463
transform 1 0 2376 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1691
timestamp 1569543463
transform 1 0 2440 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1692
timestamp 1569543463
transform 1 0 2312 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1693
timestamp 1569543463
transform 1 0 2376 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1694
timestamp 1569543463
transform 1 0 2440 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1695
timestamp 1569543463
transform 1 0 2376 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1696
timestamp 1569543463
transform 1 0 2248 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1697
timestamp 1569543463
transform 1 0 2312 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1698
timestamp 1569543463
transform 1 0 2440 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1699
timestamp 1569543463
transform 1 0 2056 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1700
timestamp 1569543463
transform 1 0 1928 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1701
timestamp 1569543463
transform 1 0 2056 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1702
timestamp 1569543463
transform 1 0 2056 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1703
timestamp 1569543463
transform 1 0 2056 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1704
timestamp 1569543463
transform 1 0 1928 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1705
timestamp 1569543463
transform 1 0 2120 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1706
timestamp 1569543463
transform 1 0 2120 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1707
timestamp 1569543463
transform 1 0 2184 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1708
timestamp 1569543463
transform 1 0 2120 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1709
timestamp 1569543463
transform 1 0 1992 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1710
timestamp 1569543463
transform 1 0 2120 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1711
timestamp 1569543463
transform 1 0 2120 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1712
timestamp 1569543463
transform 1 0 2184 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1713
timestamp 1569543463
transform 1 0 2184 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1714
timestamp 1569543463
transform 1 0 2056 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1715
timestamp 1569543463
transform 1 0 2184 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1716
timestamp 1569543463
transform 1 0 2184 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1717
timestamp 1569543463
transform 1 0 1928 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1718
timestamp 1569543463
transform 1 0 1992 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1719
timestamp 1569543463
transform 1 0 1992 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1720
timestamp 1569543463
transform 1 0 1928 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1721
timestamp 1569543463
transform 1 0 1928 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1722
timestamp 1569543463
transform 1 0 1992 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1723
timestamp 1569543463
transform 1 0 1992 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1724
timestamp 1569543463
transform 1 0 2056 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1725
timestamp 1569543463
transform 1 0 2184 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1726
timestamp 1569543463
transform 1 0 2056 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1727
timestamp 1569543463
transform 1 0 2056 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1728
timestamp 1569543463
transform 1 0 1928 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1729
timestamp 1569543463
transform 1 0 2056 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1730
timestamp 1569543463
transform 1 0 2056 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1731
timestamp 1569543463
transform 1 0 2184 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1732
timestamp 1569543463
transform 1 0 2184 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1733
timestamp 1569543463
transform 1 0 2184 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1734
timestamp 1569543463
transform 1 0 2184 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1735
timestamp 1569543463
transform 1 0 2120 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1736
timestamp 1569543463
transform 1 0 1992 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1737
timestamp 1569543463
transform 1 0 2120 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1738
timestamp 1569543463
transform 1 0 2120 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1739
timestamp 1569543463
transform 1 0 1928 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1740
timestamp 1569543463
transform 1 0 2120 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1741
timestamp 1569543463
transform 1 0 2120 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1742
timestamp 1569543463
transform 1 0 1928 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1743
timestamp 1569543463
transform 1 0 1928 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1744
timestamp 1569543463
transform 1 0 1928 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1745
timestamp 1569543463
transform 1 0 1992 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1746
timestamp 1569543463
transform 1 0 1992 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1747
timestamp 1569543463
transform 1 0 1992 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1748
timestamp 1569543463
transform 1 0 1992 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1749
timestamp 1569543463
transform 1 0 2376 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1750
timestamp 1569543463
transform 1 0 2440 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1751
timestamp 1569543463
transform 1 0 2440 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1752
timestamp 1569543463
transform 1 0 2376 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1753
timestamp 1569543463
transform 1 0 2440 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1754
timestamp 1569543463
transform 1 0 2440 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1755
timestamp 1569543463
transform 1 0 2440 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1756
timestamp 1569543463
transform 1 0 2312 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1757
timestamp 1569543463
transform 1 0 2248 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1758
timestamp 1569543463
transform 1 0 2248 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1759
timestamp 1569543463
transform 1 0 2312 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1760
timestamp 1569543463
transform 1 0 2248 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1761
timestamp 1569543463
transform 1 0 2248 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1762
timestamp 1569543463
transform 1 0 2312 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1763
timestamp 1569543463
transform 1 0 2248 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1764
timestamp 1569543463
transform 1 0 2312 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1765
timestamp 1569543463
transform 1 0 2312 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1766
timestamp 1569543463
transform 1 0 2376 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1767
timestamp 1569543463
transform 1 0 2376 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1768
timestamp 1569543463
transform 1 0 2376 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1769
timestamp 1569543463
transform 1 0 1672 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1770
timestamp 1569543463
transform 1 0 1672 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1771
timestamp 1569543463
transform 1 0 1608 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1772
timestamp 1569543463
transform 1 0 1608 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1773
timestamp 1569543463
transform 1 0 1800 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1774
timestamp 1569543463
transform 1 0 1800 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1775
timestamp 1569543463
transform 1 0 1672 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1776
timestamp 1569543463
transform 1 0 1672 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1777
timestamp 1569543463
transform 1 0 1672 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1778
timestamp 1569543463
transform 1 0 1736 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1779
timestamp 1569543463
transform 1 0 1864 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1780
timestamp 1569543463
transform 1 0 1736 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1781
timestamp 1569543463
transform 1 0 1736 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1782
timestamp 1569543463
transform 1 0 1800 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1783
timestamp 1569543463
transform 1 0 1800 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1784
timestamp 1569543463
transform 1 0 1800 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1785
timestamp 1569543463
transform 1 0 1736 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1786
timestamp 1569543463
transform 1 0 1736 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1787
timestamp 1569543463
transform 1 0 1864 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1788
timestamp 1569543463
transform 1 0 1864 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1789
timestamp 1569543463
transform 1 0 1864 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1790
timestamp 1569543463
transform 1 0 1864 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1791
timestamp 1569543463
transform 1 0 1608 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1792
timestamp 1569543463
transform 1 0 1608 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1793
timestamp 1569543463
transform 1 0 1608 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1794
timestamp 1569543463
transform 1 0 1544 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1795
timestamp 1569543463
transform 1 0 1544 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1796
timestamp 1569543463
transform 1 0 1288 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1797
timestamp 1569543463
transform 1 0 1288 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1798
timestamp 1569543463
transform 1 0 1288 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1799
timestamp 1569543463
transform 1 0 1288 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1800
timestamp 1569543463
transform 1 0 1288 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1801
timestamp 1569543463
transform 1 0 1480 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1802
timestamp 1569543463
transform 1 0 1416 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1803
timestamp 1569543463
transform 1 0 1416 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1804
timestamp 1569543463
transform 1 0 1480 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1805
timestamp 1569543463
transform 1 0 1352 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1806
timestamp 1569543463
transform 1 0 1352 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1807
timestamp 1569543463
transform 1 0 1352 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1808
timestamp 1569543463
transform 1 0 1416 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1809
timestamp 1569543463
transform 1 0 1416 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1810
timestamp 1569543463
transform 1 0 1416 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1811
timestamp 1569543463
transform 1 0 1480 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1812
timestamp 1569543463
transform 1 0 1480 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1813
timestamp 1569543463
transform 1 0 1480 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1814
timestamp 1569543463
transform 1 0 1544 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_1815
timestamp 1569543463
transform 1 0 1544 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_1816
timestamp 1569543463
transform 1 0 1544 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_1817
timestamp 1569543463
transform 1 0 1352 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_1818
timestamp 1569543463
transform 1 0 1352 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_1819
timestamp 1569543463
transform 1 0 1544 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1820
timestamp 1569543463
transform 1 0 1352 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1821
timestamp 1569543463
transform 1 0 1352 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1822
timestamp 1569543463
transform 1 0 1352 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1823
timestamp 1569543463
transform 1 0 1352 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1824
timestamp 1569543463
transform 1 0 1352 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1825
timestamp 1569543463
transform 1 0 1544 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1826
timestamp 1569543463
transform 1 0 1544 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1827
timestamp 1569543463
transform 1 0 1544 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1828
timestamp 1569543463
transform 1 0 1416 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1829
timestamp 1569543463
transform 1 0 1416 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1830
timestamp 1569543463
transform 1 0 1288 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1831
timestamp 1569543463
transform 1 0 1416 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1832
timestamp 1569543463
transform 1 0 1416 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1833
timestamp 1569543463
transform 1 0 1416 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1834
timestamp 1569543463
transform 1 0 1288 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1835
timestamp 1569543463
transform 1 0 1288 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1836
timestamp 1569543463
transform 1 0 1480 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1837
timestamp 1569543463
transform 1 0 1480 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1838
timestamp 1569543463
transform 1 0 1480 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1839
timestamp 1569543463
transform 1 0 1480 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1840
timestamp 1569543463
transform 1 0 1480 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1841
timestamp 1569543463
transform 1 0 1288 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1842
timestamp 1569543463
transform 1 0 1288 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1843
timestamp 1569543463
transform 1 0 1544 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1844
timestamp 1569543463
transform 1 0 1800 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1845
timestamp 1569543463
transform 1 0 1800 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1846
timestamp 1569543463
transform 1 0 1608 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1847
timestamp 1569543463
transform 1 0 1608 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1848
timestamp 1569543463
transform 1 0 1608 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1849
timestamp 1569543463
transform 1 0 1608 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1850
timestamp 1569543463
transform 1 0 1608 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1851
timestamp 1569543463
transform 1 0 1800 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1852
timestamp 1569543463
transform 1 0 1800 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1853
timestamp 1569543463
transform 1 0 1864 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1854
timestamp 1569543463
transform 1 0 1864 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1855
timestamp 1569543463
transform 1 0 1864 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1856
timestamp 1569543463
transform 1 0 1672 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1857
timestamp 1569543463
transform 1 0 1672 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1858
timestamp 1569543463
transform 1 0 1672 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1859
timestamp 1569543463
transform 1 0 1672 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1860
timestamp 1569543463
transform 1 0 1672 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1861
timestamp 1569543463
transform 1 0 1864 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1862
timestamp 1569543463
transform 1 0 1736 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1863
timestamp 1569543463
transform 1 0 1736 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_1864
timestamp 1569543463
transform 1 0 1736 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_1865
timestamp 1569543463
transform 1 0 1736 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1866
timestamp 1569543463
transform 1 0 1736 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_1867
timestamp 1569543463
transform 1 0 1864 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_1868
timestamp 1569543463
transform 1 0 1800 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_1869
timestamp 1569543463
transform 1 0 1800 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1870
timestamp 1569543463
transform 1 0 1608 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1871
timestamp 1569543463
transform 1 0 1864 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1872
timestamp 1569543463
transform 1 0 1608 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1873
timestamp 1569543463
transform 1 0 1800 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1874
timestamp 1569543463
transform 1 0 1672 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1875
timestamp 1569543463
transform 1 0 1864 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1876
timestamp 1569543463
transform 1 0 1672 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1877
timestamp 1569543463
transform 1 0 1864 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1878
timestamp 1569543463
transform 1 0 1672 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1879
timestamp 1569543463
transform 1 0 1864 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1880
timestamp 1569543463
transform 1 0 1672 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1881
timestamp 1569543463
transform 1 0 1672 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1882
timestamp 1569543463
transform 1 0 1736 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1883
timestamp 1569543463
transform 1 0 1800 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1884
timestamp 1569543463
transform 1 0 1736 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1885
timestamp 1569543463
transform 1 0 1736 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1886
timestamp 1569543463
transform 1 0 1608 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1887
timestamp 1569543463
transform 1 0 1736 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1888
timestamp 1569543463
transform 1 0 1608 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1889
timestamp 1569543463
transform 1 0 1736 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1890
timestamp 1569543463
transform 1 0 1608 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1891
timestamp 1569543463
transform 1 0 1864 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1892
timestamp 1569543463
transform 1 0 1800 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1893
timestamp 1569543463
transform 1 0 1800 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1894
timestamp 1569543463
transform 1 0 1352 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1895
timestamp 1569543463
transform 1 0 1480 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1896
timestamp 1569543463
transform 1 0 1480 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1897
timestamp 1569543463
transform 1 0 1544 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1898
timestamp 1569543463
transform 1 0 1544 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1899
timestamp 1569543463
transform 1 0 1416 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1900
timestamp 1569543463
transform 1 0 1288 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1901
timestamp 1569543463
transform 1 0 1544 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1902
timestamp 1569543463
transform 1 0 1416 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1903
timestamp 1569543463
transform 1 0 1544 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1904
timestamp 1569543463
transform 1 0 1288 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1905
timestamp 1569543463
transform 1 0 1544 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1906
timestamp 1569543463
transform 1 0 1480 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1907
timestamp 1569543463
transform 1 0 1288 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1908
timestamp 1569543463
transform 1 0 1480 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1909
timestamp 1569543463
transform 1 0 1288 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1910
timestamp 1569543463
transform 1 0 1352 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1911
timestamp 1569543463
transform 1 0 1352 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1912
timestamp 1569543463
transform 1 0 1352 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1913
timestamp 1569543463
transform 1 0 1288 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1914
timestamp 1569543463
transform 1 0 1352 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1915
timestamp 1569543463
transform 1 0 1416 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1916
timestamp 1569543463
transform 1 0 1416 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1917
timestamp 1569543463
transform 1 0 1416 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1918
timestamp 1569543463
transform 1 0 1480 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1919
timestamp 1569543463
transform 1 0 1352 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1920
timestamp 1569543463
transform 1 0 1288 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1921
timestamp 1569543463
transform 1 0 1544 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1922
timestamp 1569543463
transform 1 0 1352 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1923
timestamp 1569543463
transform 1 0 1288 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1924
timestamp 1569543463
transform 1 0 1416 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1925
timestamp 1569543463
transform 1 0 1416 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1926
timestamp 1569543463
transform 1 0 1480 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1927
timestamp 1569543463
transform 1 0 1480 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1928
timestamp 1569543463
transform 1 0 1480 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1929
timestamp 1569543463
transform 1 0 1352 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1930
timestamp 1569543463
transform 1 0 1480 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1931
timestamp 1569543463
transform 1 0 1544 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1932
timestamp 1569543463
transform 1 0 1416 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1933
timestamp 1569543463
transform 1 0 1544 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1934
timestamp 1569543463
transform 1 0 1288 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1935
timestamp 1569543463
transform 1 0 1544 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1936
timestamp 1569543463
transform 1 0 1416 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1937
timestamp 1569543463
transform 1 0 1288 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1938
timestamp 1569543463
transform 1 0 1352 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1939
timestamp 1569543463
transform 1 0 1608 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1940
timestamp 1569543463
transform 1 0 1864 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1941
timestamp 1569543463
transform 1 0 1608 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1942
timestamp 1569543463
transform 1 0 1672 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1943
timestamp 1569543463
transform 1 0 1672 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1944
timestamp 1569543463
transform 1 0 1672 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1945
timestamp 1569543463
transform 1 0 1736 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1946
timestamp 1569543463
transform 1 0 1736 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1947
timestamp 1569543463
transform 1 0 1800 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1948
timestamp 1569543463
transform 1 0 1736 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1949
timestamp 1569543463
transform 1 0 1800 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1950
timestamp 1569543463
transform 1 0 1864 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1951
timestamp 1569543463
transform 1 0 1800 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1952
timestamp 1569543463
transform 1 0 1608 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1953
timestamp 1569543463
transform 1 0 1800 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1954
timestamp 1569543463
transform 1 0 1864 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_1955
timestamp 1569543463
transform 1 0 1608 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1956
timestamp 1569543463
transform 1 0 1864 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_1957
timestamp 1569543463
transform 1 0 1672 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1958
timestamp 1569543463
transform 1 0 1736 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_1959
timestamp 1569543463
transform 1 0 2376 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1960
timestamp 1569543463
transform 1 0 2376 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1961
timestamp 1569543463
transform 1 0 2248 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1962
timestamp 1569543463
transform 1 0 2440 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1963
timestamp 1569543463
transform 1 0 2440 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1964
timestamp 1569543463
transform 1 0 2312 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1965
timestamp 1569543463
transform 1 0 2376 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1966
timestamp 1569543463
transform 1 0 2248 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1967
timestamp 1569543463
transform 1 0 2248 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1968
timestamp 1569543463
transform 1 0 2312 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1969
timestamp 1569543463
transform 1 0 2312 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1970
timestamp 1569543463
transform 1 0 2248 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1971
timestamp 1569543463
transform 1 0 2248 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1972
timestamp 1569543463
transform 1 0 2312 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1973
timestamp 1569543463
transform 1 0 1992 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1974
timestamp 1569543463
transform 1 0 1992 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1975
timestamp 1569543463
transform 1 0 1928 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1976
timestamp 1569543463
transform 1 0 2056 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1977
timestamp 1569543463
transform 1 0 2056 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1978
timestamp 1569543463
transform 1 0 1992 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1979
timestamp 1569543463
transform 1 0 2120 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1980
timestamp 1569543463
transform 1 0 2120 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1981
timestamp 1569543463
transform 1 0 2056 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1982
timestamp 1569543463
transform 1 0 2184 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1983
timestamp 1569543463
transform 1 0 2184 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1984
timestamp 1569543463
transform 1 0 2120 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1985
timestamp 1569543463
transform 1 0 2056 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1986
timestamp 1569543463
transform 1 0 2056 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1987
timestamp 1569543463
transform 1 0 2120 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1988
timestamp 1569543463
transform 1 0 2120 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1989
timestamp 1569543463
transform 1 0 2184 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1990
timestamp 1569543463
transform 1 0 1928 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1991
timestamp 1569543463
transform 1 0 2184 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1992
timestamp 1569543463
transform 1 0 1992 0 1 2184
box -8 -8 8 8
use VIA1$5  VIA1$5_1993
timestamp 1569543463
transform 1 0 2184 0 1 2056
box -8 -8 8 8
use VIA1$5  VIA1$5_1994
timestamp 1569543463
transform 1 0 1928 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_1995
timestamp 1569543463
transform 1 0 1928 0 1 1992
box -8 -8 8 8
use VIA1$5  VIA1$5_1996
timestamp 1569543463
transform 1 0 1928 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1997
timestamp 1569543463
transform 1 0 1992 0 1 2120
box -8 -8 8 8
use VIA1$5  VIA1$5_1998
timestamp 1569543463
transform 1 0 2056 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_1999
timestamp 1569543463
transform 1 0 1928 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_2000
timestamp 1569543463
transform 1 0 1928 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_2001
timestamp 1569543463
transform 1 0 1992 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_2002
timestamp 1569543463
transform 1 0 1992 0 1 2440
box -8 -8 8 8
use VIA1$5  VIA1$5_2003
timestamp 1569543463
transform 1 0 2184 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_2004
timestamp 1569543463
transform 1 0 1928 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_2005
timestamp 1569543463
transform 1 0 2056 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_2006
timestamp 1569543463
transform 1 0 1992 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_2007
timestamp 1569543463
transform 1 0 2120 0 1 2248
box -8 -8 8 8
use VIA1$5  VIA1$5_2008
timestamp 1569543463
transform 1 0 2056 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_2009
timestamp 1569543463
transform 1 0 2120 0 1 2312
box -8 -8 8 8
use VIA1$5  VIA1$5_2010
timestamp 1569543463
transform 1 0 1928 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_2011
timestamp 1569543463
transform 1 0 1992 0 1 2376
box -8 -8 8 8
use VIA1$5  VIA1$5_2012
timestamp 1569543463
transform 1 0 1864 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2013
timestamp 1569543463
transform 1 0 1672 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2014
timestamp 1569543463
transform 1 0 1672 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2015
timestamp 1569543463
transform 1 0 1608 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2016
timestamp 1569543463
transform 1 0 1736 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2017
timestamp 1569543463
transform 1 0 1608 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2018
timestamp 1569543463
transform 1 0 1800 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2019
timestamp 1569543463
transform 1 0 1672 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2020
timestamp 1569543463
transform 1 0 1800 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2021
timestamp 1569543463
transform 1 0 1672 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2022
timestamp 1569543463
transform 1 0 1736 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2023
timestamp 1569543463
transform 1 0 1608 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2024
timestamp 1569543463
transform 1 0 1608 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2025
timestamp 1569543463
transform 1 0 1480 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2026
timestamp 1569543463
transform 1 0 1416 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2027
timestamp 1569543463
transform 1 0 1352 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2028
timestamp 1569543463
transform 1 0 1416 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2029
timestamp 1569543463
transform 1 0 1416 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2030
timestamp 1569543463
transform 1 0 1416 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2031
timestamp 1569543463
transform 1 0 1352 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2032
timestamp 1569543463
transform 1 0 1352 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2033
timestamp 1569543463
transform 1 0 1288 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2034
timestamp 1569543463
transform 1 0 1544 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2035
timestamp 1569543463
transform 1 0 1288 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2036
timestamp 1569543463
transform 1 0 1544 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2037
timestamp 1569543463
transform 1 0 1288 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2038
timestamp 1569543463
transform 1 0 1352 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2039
timestamp 1569543463
transform 1 0 1480 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2040
timestamp 1569543463
transform 1 0 1544 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2041
timestamp 1569543463
transform 1 0 1480 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2042
timestamp 1569543463
transform 1 0 1544 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2043
timestamp 1569543463
transform 1 0 1480 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2044
timestamp 1569543463
transform 1 0 1288 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2045
timestamp 1569543463
transform 1 0 1288 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2046
timestamp 1569543463
transform 1 0 1288 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2047
timestamp 1569543463
transform 1 0 1288 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2048
timestamp 1569543463
transform 1 0 1544 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2049
timestamp 1569543463
transform 1 0 1544 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2050
timestamp 1569543463
transform 1 0 1416 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2051
timestamp 1569543463
transform 1 0 1288 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2052
timestamp 1569543463
transform 1 0 1416 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2053
timestamp 1569543463
transform 1 0 1352 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2054
timestamp 1569543463
transform 1 0 1352 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2055
timestamp 1569543463
transform 1 0 1416 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2056
timestamp 1569543463
transform 1 0 1480 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2057
timestamp 1569543463
transform 1 0 1288 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2058
timestamp 1569543463
transform 1 0 1416 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2059
timestamp 1569543463
transform 1 0 1480 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2060
timestamp 1569543463
transform 1 0 1352 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2061
timestamp 1569543463
transform 1 0 1480 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2062
timestamp 1569543463
transform 1 0 1352 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2063
timestamp 1569543463
transform 1 0 1416 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2064
timestamp 1569543463
transform 1 0 1352 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2065
timestamp 1569543463
transform 1 0 1480 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2066
timestamp 1569543463
transform 1 0 1480 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2067
timestamp 1569543463
transform 1 0 1608 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2068
timestamp 1569543463
transform 1 0 1480 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2069
timestamp 1569543463
transform 1 0 1480 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2070
timestamp 1569543463
transform 1 0 1480 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2071
timestamp 1569543463
transform 1 0 1352 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2072
timestamp 1569543463
transform 1 0 1288 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2073
timestamp 1569543463
transform 1 0 1480 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2074
timestamp 1569543463
transform 1 0 1480 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2075
timestamp 1569543463
transform 1 0 1352 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2076
timestamp 1569543463
transform 1 0 1416 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2077
timestamp 1569543463
transform 1 0 1480 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2078
timestamp 1569543463
transform 1 0 1288 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2079
timestamp 1569543463
transform 1 0 1288 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2080
timestamp 1569543463
transform 1 0 1416 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2081
timestamp 1569543463
transform 1 0 1480 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2082
timestamp 1569543463
transform 1 0 1480 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2083
timestamp 1569543463
transform 1 0 1352 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2084
timestamp 1569543463
transform 1 0 1352 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2085
timestamp 1569543463
transform 1 0 1352 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2086
timestamp 1569543463
transform 1 0 1288 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2087
timestamp 1569543463
transform 1 0 1288 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2088
timestamp 1569543463
transform 1 0 1352 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2089
timestamp 1569543463
transform 1 0 1352 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2090
timestamp 1569543463
transform 1 0 1288 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2091
timestamp 1569543463
transform 1 0 1416 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2092
timestamp 1569543463
transform 1 0 1352 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2093
timestamp 1569543463
transform 1 0 1416 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2094
timestamp 1569543463
transform 1 0 1480 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2095
timestamp 1569543463
transform 1 0 1288 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2096
timestamp 1569543463
transform 1 0 1416 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2097
timestamp 1569543463
transform 1 0 1416 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2098
timestamp 1569543463
transform 1 0 1352 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2099
timestamp 1569543463
transform 1 0 1288 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2100
timestamp 1569543463
transform 1 0 1352 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2101
timestamp 1569543463
transform 1 0 1416 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2102
timestamp 1569543463
transform 1 0 1480 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2103
timestamp 1569543463
transform 1 0 1288 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2104
timestamp 1569543463
transform 1 0 1416 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2105
timestamp 1569543463
transform 1 0 1416 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2106
timestamp 1569543463
transform 1 0 1288 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2107
timestamp 1569543463
transform 1 0 1416 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2108
timestamp 1569543463
transform 1 0 2440 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2109
timestamp 1569543463
transform 1 0 2440 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2110
timestamp 1569543463
transform 1 0 2440 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2111
timestamp 1569543463
transform 1 0 2376 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2112
timestamp 1569543463
transform 1 0 2376 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2113
timestamp 1569543463
transform 1 0 2440 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2114
timestamp 1569543463
transform 1 0 2376 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2115
timestamp 1569543463
transform 1 0 2312 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2116
timestamp 1569543463
transform 1 0 2376 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2117
timestamp 1569543463
transform 1 0 2440 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2118
timestamp 1569543463
transform 1 0 2376 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2119
timestamp 1569543463
transform 1 0 2376 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2120
timestamp 1569543463
transform 1 0 2376 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2121
timestamp 1569543463
transform 1 0 2312 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2122
timestamp 1569543463
transform 1 0 2312 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2123
timestamp 1569543463
transform 1 0 2312 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2124
timestamp 1569543463
transform 1 0 2312 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2125
timestamp 1569543463
transform 1 0 2312 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2126
timestamp 1569543463
transform 1 0 2440 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2127
timestamp 1569543463
transform 1 0 2440 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2128
timestamp 1569543463
transform 1 0 2440 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2129
timestamp 1569543463
transform 1 0 1096 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2130
timestamp 1569543463
transform 1 0 1160 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2131
timestamp 1569543463
transform 1 0 968 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2132
timestamp 1569543463
transform 1 0 1096 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2133
timestamp 1569543463
transform 1 0 1032 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2134
timestamp 1569543463
transform 1 0 968 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2135
timestamp 1569543463
transform 1 0 1160 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2136
timestamp 1569543463
transform 1 0 1224 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2137
timestamp 1569543463
transform 1 0 1032 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2138
timestamp 1569543463
transform 1 0 1160 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2139
timestamp 1569543463
transform 1 0 1224 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2140
timestamp 1569543463
transform 1 0 1160 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2141
timestamp 1569543463
transform 1 0 968 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2142
timestamp 1569543463
transform 1 0 1096 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2143
timestamp 1569543463
transform 1 0 1032 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2144
timestamp 1569543463
transform 1 0 1096 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2145
timestamp 1569543463
transform 1 0 1032 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2146
timestamp 1569543463
transform 1 0 1224 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2147
timestamp 1569543463
transform 1 0 1224 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2148
timestamp 1569543463
transform 1 0 968 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2149
timestamp 1569543463
transform 1 0 904 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2150
timestamp 1569543463
transform 1 0 904 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2151
timestamp 1569543463
transform 1 0 840 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2152
timestamp 1569543463
transform 1 0 776 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2153
timestamp 1569543463
transform 1 0 840 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2154
timestamp 1569543463
transform 1 0 712 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2155
timestamp 1569543463
transform 1 0 904 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2156
timestamp 1569543463
transform 1 0 712 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2157
timestamp 1569543463
transform 1 0 776 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2158
timestamp 1569543463
transform 1 0 712 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2159
timestamp 1569543463
transform 1 0 776 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2160
timestamp 1569543463
transform 1 0 776 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2161
timestamp 1569543463
transform 1 0 840 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2162
timestamp 1569543463
transform 1 0 904 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2163
timestamp 1569543463
transform 1 0 712 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2164
timestamp 1569543463
transform 1 0 840 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2165
timestamp 1569543463
transform 1 0 840 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2166
timestamp 1569543463
transform 1 0 712 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2167
timestamp 1569543463
transform 1 0 904 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2168
timestamp 1569543463
transform 1 0 776 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2169
timestamp 1569543463
transform 1 0 712 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2170
timestamp 1569543463
transform 1 0 904 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2171
timestamp 1569543463
transform 1 0 904 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2172
timestamp 1569543463
transform 1 0 840 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2173
timestamp 1569543463
transform 1 0 904 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2174
timestamp 1569543463
transform 1 0 840 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2175
timestamp 1569543463
transform 1 0 712 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2176
timestamp 1569543463
transform 1 0 712 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2177
timestamp 1569543463
transform 1 0 776 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2178
timestamp 1569543463
transform 1 0 840 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2179
timestamp 1569543463
transform 1 0 776 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2180
timestamp 1569543463
transform 1 0 840 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2181
timestamp 1569543463
transform 1 0 712 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2182
timestamp 1569543463
transform 1 0 776 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2183
timestamp 1569543463
transform 1 0 776 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2184
timestamp 1569543463
transform 1 0 904 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2185
timestamp 1569543463
transform 1 0 1160 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2186
timestamp 1569543463
transform 1 0 1032 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2187
timestamp 1569543463
transform 1 0 1160 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2188
timestamp 1569543463
transform 1 0 1160 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2189
timestamp 1569543463
transform 1 0 1096 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2190
timestamp 1569543463
transform 1 0 968 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2191
timestamp 1569543463
transform 1 0 1032 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2192
timestamp 1569543463
transform 1 0 1096 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2193
timestamp 1569543463
transform 1 0 1160 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2194
timestamp 1569543463
transform 1 0 968 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2195
timestamp 1569543463
transform 1 0 1224 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2196
timestamp 1569543463
transform 1 0 1224 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2197
timestamp 1569543463
transform 1 0 968 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2198
timestamp 1569543463
transform 1 0 1032 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2199
timestamp 1569543463
transform 1 0 1224 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2200
timestamp 1569543463
transform 1 0 968 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2201
timestamp 1569543463
transform 1 0 1032 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2202
timestamp 1569543463
transform 1 0 1096 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2203
timestamp 1569543463
transform 1 0 1160 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2204
timestamp 1569543463
transform 1 0 1032 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2205
timestamp 1569543463
transform 1 0 968 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2206
timestamp 1569543463
transform 1 0 1096 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2207
timestamp 1569543463
transform 1 0 1224 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2208
timestamp 1569543463
transform 1 0 1096 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2209
timestamp 1569543463
transform 1 0 1224 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2210
timestamp 1569543463
transform 1 0 584 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2211
timestamp 1569543463
transform 1 0 520 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2212
timestamp 1569543463
transform 1 0 392 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2213
timestamp 1569543463
transform 1 0 584 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2214
timestamp 1569543463
transform 1 0 520 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2215
timestamp 1569543463
transform 1 0 392 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2216
timestamp 1569543463
transform 1 0 584 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2217
timestamp 1569543463
transform 1 0 456 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2218
timestamp 1569543463
transform 1 0 392 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2219
timestamp 1569543463
transform 1 0 456 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2220
timestamp 1569543463
transform 1 0 520 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2221
timestamp 1569543463
transform 1 0 520 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2222
timestamp 1569543463
transform 1 0 392 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2223
timestamp 1569543463
transform 1 0 456 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2224
timestamp 1569543463
transform 1 0 456 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2225
timestamp 1569543463
transform 1 0 584 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2226
timestamp 1569543463
transform 1 0 72 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2227
timestamp 1569543463
transform 1 0 328 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2228
timestamp 1569543463
transform 1 0 72 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2229
timestamp 1569543463
transform 1 0 264 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2230
timestamp 1569543463
transform 1 0 264 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2231
timestamp 1569543463
transform 1 0 136 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2232
timestamp 1569543463
transform 1 0 328 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2233
timestamp 1569543463
transform 1 0 200 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2234
timestamp 1569543463
transform 1 0 136 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2235
timestamp 1569543463
transform 1 0 264 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2236
timestamp 1569543463
transform 1 0 328 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2237
timestamp 1569543463
transform 1 0 72 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2238
timestamp 1569543463
transform 1 0 200 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2239
timestamp 1569543463
transform 1 0 72 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2240
timestamp 1569543463
transform 1 0 200 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2241
timestamp 1569543463
transform 1 0 136 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2242
timestamp 1569543463
transform 1 0 264 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2243
timestamp 1569543463
transform 1 0 136 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2244
timestamp 1569543463
transform 1 0 328 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2245
timestamp 1569543463
transform 1 0 200 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2246
timestamp 1569543463
transform 1 0 264 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2247
timestamp 1569543463
transform 1 0 264 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2248
timestamp 1569543463
transform 1 0 136 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2249
timestamp 1569543463
transform 1 0 264 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2250
timestamp 1569543463
transform 1 0 264 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2251
timestamp 1569543463
transform 1 0 200 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2252
timestamp 1569543463
transform 1 0 136 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2253
timestamp 1569543463
transform 1 0 328 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2254
timestamp 1569543463
transform 1 0 136 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2255
timestamp 1569543463
transform 1 0 72 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2256
timestamp 1569543463
transform 1 0 200 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2257
timestamp 1569543463
transform 1 0 136 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2258
timestamp 1569543463
transform 1 0 72 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2259
timestamp 1569543463
transform 1 0 328 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2260
timestamp 1569543463
transform 1 0 328 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2261
timestamp 1569543463
transform 1 0 328 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2262
timestamp 1569543463
transform 1 0 72 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2263
timestamp 1569543463
transform 1 0 328 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2264
timestamp 1569543463
transform 1 0 72 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2265
timestamp 1569543463
transform 1 0 200 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2266
timestamp 1569543463
transform 1 0 200 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2267
timestamp 1569543463
transform 1 0 136 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2268
timestamp 1569543463
transform 1 0 264 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2269
timestamp 1569543463
transform 1 0 200 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2270
timestamp 1569543463
transform 1 0 72 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2271
timestamp 1569543463
transform 1 0 520 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2272
timestamp 1569543463
transform 1 0 392 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2273
timestamp 1569543463
transform 1 0 392 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2274
timestamp 1569543463
transform 1 0 392 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2275
timestamp 1569543463
transform 1 0 520 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2276
timestamp 1569543463
transform 1 0 584 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2277
timestamp 1569543463
transform 1 0 584 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2278
timestamp 1569543463
transform 1 0 456 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2279
timestamp 1569543463
transform 1 0 456 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2280
timestamp 1569543463
transform 1 0 520 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2281
timestamp 1569543463
transform 1 0 520 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2282
timestamp 1569543463
transform 1 0 520 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2283
timestamp 1569543463
transform 1 0 456 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2284
timestamp 1569543463
transform 1 0 392 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2285
timestamp 1569543463
transform 1 0 584 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2286
timestamp 1569543463
transform 1 0 584 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2287
timestamp 1569543463
transform 1 0 584 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2288
timestamp 1569543463
transform 1 0 456 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2289
timestamp 1569543463
transform 1 0 456 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2290
timestamp 1569543463
transform 1 0 392 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2291
timestamp 1569543463
transform 1 0 392 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2292
timestamp 1569543463
transform 1 0 584 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2293
timestamp 1569543463
transform 1 0 520 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2294
timestamp 1569543463
transform 1 0 392 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2295
timestamp 1569543463
transform 1 0 584 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2296
timestamp 1569543463
transform 1 0 392 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2297
timestamp 1569543463
transform 1 0 456 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2298
timestamp 1569543463
transform 1 0 456 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2299
timestamp 1569543463
transform 1 0 456 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2300
timestamp 1569543463
transform 1 0 392 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2301
timestamp 1569543463
transform 1 0 584 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2302
timestamp 1569543463
transform 1 0 520 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2303
timestamp 1569543463
transform 1 0 520 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2304
timestamp 1569543463
transform 1 0 456 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2305
timestamp 1569543463
transform 1 0 584 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2306
timestamp 1569543463
transform 1 0 520 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2307
timestamp 1569543463
transform 1 0 584 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2308
timestamp 1569543463
transform 1 0 520 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2309
timestamp 1569543463
transform 1 0 456 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2310
timestamp 1569543463
transform 1 0 392 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2311
timestamp 1569543463
transform 1 0 264 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2312
timestamp 1569543463
transform 1 0 200 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2313
timestamp 1569543463
transform 1 0 72 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2314
timestamp 1569543463
transform 1 0 72 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2315
timestamp 1569543463
transform 1 0 264 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2316
timestamp 1569543463
transform 1 0 264 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2317
timestamp 1569543463
transform 1 0 200 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2318
timestamp 1569543463
transform 1 0 200 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2319
timestamp 1569543463
transform 1 0 72 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2320
timestamp 1569543463
transform 1 0 328 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2321
timestamp 1569543463
transform 1 0 200 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2322
timestamp 1569543463
transform 1 0 136 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2323
timestamp 1569543463
transform 1 0 136 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2324
timestamp 1569543463
transform 1 0 328 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2325
timestamp 1569543463
transform 1 0 72 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2326
timestamp 1569543463
transform 1 0 136 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2327
timestamp 1569543463
transform 1 0 328 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2328
timestamp 1569543463
transform 1 0 72 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2329
timestamp 1569543463
transform 1 0 136 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2330
timestamp 1569543463
transform 1 0 136 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2331
timestamp 1569543463
transform 1 0 328 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2332
timestamp 1569543463
transform 1 0 200 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2333
timestamp 1569543463
transform 1 0 264 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2334
timestamp 1569543463
transform 1 0 264 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2335
timestamp 1569543463
transform 1 0 328 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2336
timestamp 1569543463
transform 1 0 328 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2337
timestamp 1569543463
transform 1 0 328 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2338
timestamp 1569543463
transform 1 0 72 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2339
timestamp 1569543463
transform 1 0 200 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2340
timestamp 1569543463
transform 1 0 72 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2341
timestamp 1569543463
transform 1 0 136 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2342
timestamp 1569543463
transform 1 0 136 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2343
timestamp 1569543463
transform 1 0 72 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2344
timestamp 1569543463
transform 1 0 136 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2345
timestamp 1569543463
transform 1 0 72 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2346
timestamp 1569543463
transform 1 0 136 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2347
timestamp 1569543463
transform 1 0 328 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2348
timestamp 1569543463
transform 1 0 200 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2349
timestamp 1569543463
transform 1 0 136 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2350
timestamp 1569543463
transform 1 0 72 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2351
timestamp 1569543463
transform 1 0 200 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2352
timestamp 1569543463
transform 1 0 328 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2353
timestamp 1569543463
transform 1 0 264 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2354
timestamp 1569543463
transform 1 0 264 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2355
timestamp 1569543463
transform 1 0 264 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2356
timestamp 1569543463
transform 1 0 264 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2357
timestamp 1569543463
transform 1 0 264 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2358
timestamp 1569543463
transform 1 0 200 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2359
timestamp 1569543463
transform 1 0 200 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2360
timestamp 1569543463
transform 1 0 328 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2361
timestamp 1569543463
transform 1 0 392 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2362
timestamp 1569543463
transform 1 0 456 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2363
timestamp 1569543463
transform 1 0 392 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2364
timestamp 1569543463
transform 1 0 456 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2365
timestamp 1569543463
transform 1 0 584 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2366
timestamp 1569543463
transform 1 0 456 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2367
timestamp 1569543463
transform 1 0 456 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2368
timestamp 1569543463
transform 1 0 456 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2369
timestamp 1569543463
transform 1 0 584 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2370
timestamp 1569543463
transform 1 0 584 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2371
timestamp 1569543463
transform 1 0 520 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2372
timestamp 1569543463
transform 1 0 520 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2373
timestamp 1569543463
transform 1 0 520 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2374
timestamp 1569543463
transform 1 0 520 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2375
timestamp 1569543463
transform 1 0 584 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2376
timestamp 1569543463
transform 1 0 392 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2377
timestamp 1569543463
transform 1 0 584 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2378
timestamp 1569543463
transform 1 0 520 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2379
timestamp 1569543463
transform 1 0 392 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2380
timestamp 1569543463
transform 1 0 392 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2381
timestamp 1569543463
transform 1 0 1224 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2382
timestamp 1569543463
transform 1 0 968 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2383
timestamp 1569543463
transform 1 0 1096 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2384
timestamp 1569543463
transform 1 0 968 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2385
timestamp 1569543463
transform 1 0 968 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2386
timestamp 1569543463
transform 1 0 968 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2387
timestamp 1569543463
transform 1 0 1224 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2388
timestamp 1569543463
transform 1 0 1160 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2389
timestamp 1569543463
transform 1 0 1032 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2390
timestamp 1569543463
transform 1 0 1160 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2391
timestamp 1569543463
transform 1 0 1160 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2392
timestamp 1569543463
transform 1 0 1096 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2393
timestamp 1569543463
transform 1 0 1160 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2394
timestamp 1569543463
transform 1 0 1032 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2395
timestamp 1569543463
transform 1 0 1032 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2396
timestamp 1569543463
transform 1 0 1160 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2397
timestamp 1569543463
transform 1 0 1032 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2398
timestamp 1569543463
transform 1 0 1224 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2399
timestamp 1569543463
transform 1 0 968 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2400
timestamp 1569543463
transform 1 0 1096 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2401
timestamp 1569543463
transform 1 0 1096 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2402
timestamp 1569543463
transform 1 0 1224 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2403
timestamp 1569543463
transform 1 0 1032 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2404
timestamp 1569543463
transform 1 0 1224 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2405
timestamp 1569543463
transform 1 0 1096 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2406
timestamp 1569543463
transform 1 0 840 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2407
timestamp 1569543463
transform 1 0 840 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2408
timestamp 1569543463
transform 1 0 840 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2409
timestamp 1569543463
transform 1 0 712 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2410
timestamp 1569543463
transform 1 0 904 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2411
timestamp 1569543463
transform 1 0 904 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2412
timestamp 1569543463
transform 1 0 904 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2413
timestamp 1569543463
transform 1 0 904 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2414
timestamp 1569543463
transform 1 0 712 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2415
timestamp 1569543463
transform 1 0 776 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2416
timestamp 1569543463
transform 1 0 840 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2417
timestamp 1569543463
transform 1 0 776 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2418
timestamp 1569543463
transform 1 0 776 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2419
timestamp 1569543463
transform 1 0 776 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2420
timestamp 1569543463
transform 1 0 776 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2421
timestamp 1569543463
transform 1 0 712 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2422
timestamp 1569543463
transform 1 0 904 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2423
timestamp 1569543463
transform 1 0 712 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2424
timestamp 1569543463
transform 1 0 840 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2425
timestamp 1569543463
transform 1 0 712 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2426
timestamp 1569543463
transform 1 0 712 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2427
timestamp 1569543463
transform 1 0 712 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2428
timestamp 1569543463
transform 1 0 712 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2429
timestamp 1569543463
transform 1 0 712 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2430
timestamp 1569543463
transform 1 0 776 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2431
timestamp 1569543463
transform 1 0 776 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2432
timestamp 1569543463
transform 1 0 712 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2433
timestamp 1569543463
transform 1 0 840 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2434
timestamp 1569543463
transform 1 0 840 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2435
timestamp 1569543463
transform 1 0 776 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2436
timestamp 1569543463
transform 1 0 776 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2437
timestamp 1569543463
transform 1 0 776 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2438
timestamp 1569543463
transform 1 0 904 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2439
timestamp 1569543463
transform 1 0 840 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2440
timestamp 1569543463
transform 1 0 840 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2441
timestamp 1569543463
transform 1 0 904 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2442
timestamp 1569543463
transform 1 0 840 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2443
timestamp 1569543463
transform 1 0 904 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2444
timestamp 1569543463
transform 1 0 904 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2445
timestamp 1569543463
transform 1 0 904 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2446
timestamp 1569543463
transform 1 0 1096 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2447
timestamp 1569543463
transform 1 0 1096 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2448
timestamp 1569543463
transform 1 0 1096 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2449
timestamp 1569543463
transform 1 0 1224 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2450
timestamp 1569543463
transform 1 0 1096 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2451
timestamp 1569543463
transform 1 0 1096 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2452
timestamp 1569543463
transform 1 0 1224 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2453
timestamp 1569543463
transform 1 0 1160 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2454
timestamp 1569543463
transform 1 0 1160 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2455
timestamp 1569543463
transform 1 0 1160 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2456
timestamp 1569543463
transform 1 0 968 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2457
timestamp 1569543463
transform 1 0 968 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2458
timestamp 1569543463
transform 1 0 968 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2459
timestamp 1569543463
transform 1 0 1032 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2460
timestamp 1569543463
transform 1 0 1032 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2461
timestamp 1569543463
transform 1 0 1032 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2462
timestamp 1569543463
transform 1 0 1224 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2463
timestamp 1569543463
transform 1 0 1224 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2464
timestamp 1569543463
transform 1 0 1224 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2465
timestamp 1569543463
transform 1 0 1160 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2466
timestamp 1569543463
transform 1 0 968 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2467
timestamp 1569543463
transform 1 0 968 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2468
timestamp 1569543463
transform 1 0 1160 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2469
timestamp 1569543463
transform 1 0 1032 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2470
timestamp 1569543463
transform 1 0 1032 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2471
timestamp 1569543463
transform 1 0 648 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2472
timestamp 1569543463
transform 1 0 648 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_2473
timestamp 1569543463
transform 1 0 648 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2474
timestamp 1569543463
transform 1 0 648 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2475
timestamp 1569543463
transform 1 0 648 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2476
timestamp 1569543463
transform 1 0 648 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2477
timestamp 1569543463
transform 1 0 648 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_2478
timestamp 1569543463
transform 1 0 648 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_2479
timestamp 1569543463
transform 1 0 648 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2480
timestamp 1569543463
transform 1 0 648 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_2481
timestamp 1569543463
transform 1 0 648 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2482
timestamp 1569543463
transform 1 0 648 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2483
timestamp 1569543463
transform 1 0 648 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_2484
timestamp 1569543463
transform 1 0 648 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_2485
timestamp 1569543463
transform 1 0 648 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_2486
timestamp 1569543463
transform 1 0 648 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_2487
timestamp 1569543463
transform 1 0 648 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2488
timestamp 1569543463
transform 1 0 648 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_2489
timestamp 1569543463
transform 1 0 648 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_2490
timestamp 1569543463
transform 1 0 1096 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2491
timestamp 1569543463
transform 1 0 1032 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2492
timestamp 1569543463
transform 1 0 1096 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2493
timestamp 1569543463
transform 1 0 1032 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2494
timestamp 1569543463
transform 1 0 968 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2495
timestamp 1569543463
transform 1 0 1160 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2496
timestamp 1569543463
transform 1 0 1160 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2497
timestamp 1569543463
transform 1 0 1096 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2498
timestamp 1569543463
transform 1 0 1096 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2499
timestamp 1569543463
transform 1 0 1224 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2500
timestamp 1569543463
transform 1 0 1224 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2501
timestamp 1569543463
transform 1 0 1224 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2502
timestamp 1569543463
transform 1 0 1160 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2503
timestamp 1569543463
transform 1 0 1224 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2504
timestamp 1569543463
transform 1 0 1224 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2505
timestamp 1569543463
transform 1 0 968 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2506
timestamp 1569543463
transform 1 0 968 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2507
timestamp 1569543463
transform 1 0 968 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2508
timestamp 1569543463
transform 1 0 1032 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2509
timestamp 1569543463
transform 1 0 968 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2510
timestamp 1569543463
transform 1 0 1160 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2511
timestamp 1569543463
transform 1 0 1160 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2512
timestamp 1569543463
transform 1 0 1032 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2513
timestamp 1569543463
transform 1 0 1096 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2514
timestamp 1569543463
transform 1 0 1032 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2515
timestamp 1569543463
transform 1 0 712 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2516
timestamp 1569543463
transform 1 0 840 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2517
timestamp 1569543463
transform 1 0 840 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2518
timestamp 1569543463
transform 1 0 776 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2519
timestamp 1569543463
transform 1 0 776 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2520
timestamp 1569543463
transform 1 0 840 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2521
timestamp 1569543463
transform 1 0 712 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2522
timestamp 1569543463
transform 1 0 904 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2523
timestamp 1569543463
transform 1 0 904 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2524
timestamp 1569543463
transform 1 0 712 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2525
timestamp 1569543463
transform 1 0 904 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2526
timestamp 1569543463
transform 1 0 904 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2527
timestamp 1569543463
transform 1 0 776 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2528
timestamp 1569543463
transform 1 0 712 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2529
timestamp 1569543463
transform 1 0 840 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2530
timestamp 1569543463
transform 1 0 904 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2531
timestamp 1569543463
transform 1 0 776 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2532
timestamp 1569543463
transform 1 0 712 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2533
timestamp 1569543463
transform 1 0 776 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2534
timestamp 1569543463
transform 1 0 840 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2535
timestamp 1569543463
transform 1 0 840 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2536
timestamp 1569543463
transform 1 0 840 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2537
timestamp 1569543463
transform 1 0 712 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2538
timestamp 1569543463
transform 1 0 840 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2539
timestamp 1569543463
transform 1 0 840 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2540
timestamp 1569543463
transform 1 0 712 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2541
timestamp 1569543463
transform 1 0 712 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2542
timestamp 1569543463
transform 1 0 776 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2543
timestamp 1569543463
transform 1 0 776 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2544
timestamp 1569543463
transform 1 0 776 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2545
timestamp 1569543463
transform 1 0 904 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2546
timestamp 1569543463
transform 1 0 776 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2547
timestamp 1569543463
transform 1 0 904 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2548
timestamp 1569543463
transform 1 0 904 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2549
timestamp 1569543463
transform 1 0 712 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2550
timestamp 1569543463
transform 1 0 904 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2551
timestamp 1569543463
transform 1 0 1032 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2552
timestamp 1569543463
transform 1 0 1032 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2553
timestamp 1569543463
transform 1 0 1160 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2554
timestamp 1569543463
transform 1 0 1160 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2555
timestamp 1569543463
transform 1 0 1224 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2556
timestamp 1569543463
transform 1 0 1160 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2557
timestamp 1569543463
transform 1 0 1096 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2558
timestamp 1569543463
transform 1 0 1160 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2559
timestamp 1569543463
transform 1 0 1224 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2560
timestamp 1569543463
transform 1 0 1096 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2561
timestamp 1569543463
transform 1 0 1224 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2562
timestamp 1569543463
transform 1 0 1096 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2563
timestamp 1569543463
transform 1 0 1224 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2564
timestamp 1569543463
transform 1 0 1096 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2565
timestamp 1569543463
transform 1 0 968 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2566
timestamp 1569543463
transform 1 0 968 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2567
timestamp 1569543463
transform 1 0 968 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2568
timestamp 1569543463
transform 1 0 968 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2569
timestamp 1569543463
transform 1 0 1032 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2570
timestamp 1569543463
transform 1 0 1032 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2571
timestamp 1569543463
transform 1 0 392 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2572
timestamp 1569543463
transform 1 0 584 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2573
timestamp 1569543463
transform 1 0 584 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2574
timestamp 1569543463
transform 1 0 392 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2575
timestamp 1569543463
transform 1 0 456 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2576
timestamp 1569543463
transform 1 0 584 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2577
timestamp 1569543463
transform 1 0 392 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2578
timestamp 1569543463
transform 1 0 520 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2579
timestamp 1569543463
transform 1 0 520 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2580
timestamp 1569543463
transform 1 0 392 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2581
timestamp 1569543463
transform 1 0 584 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2582
timestamp 1569543463
transform 1 0 520 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2583
timestamp 1569543463
transform 1 0 456 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2584
timestamp 1569543463
transform 1 0 392 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2585
timestamp 1569543463
transform 1 0 584 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2586
timestamp 1569543463
transform 1 0 520 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2587
timestamp 1569543463
transform 1 0 456 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2588
timestamp 1569543463
transform 1 0 520 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2589
timestamp 1569543463
transform 1 0 456 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2590
timestamp 1569543463
transform 1 0 456 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2591
timestamp 1569543463
transform 1 0 200 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2592
timestamp 1569543463
transform 1 0 72 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2593
timestamp 1569543463
transform 1 0 200 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2594
timestamp 1569543463
transform 1 0 72 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2595
timestamp 1569543463
transform 1 0 72 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2596
timestamp 1569543463
transform 1 0 136 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2597
timestamp 1569543463
transform 1 0 264 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2598
timestamp 1569543463
transform 1 0 136 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2599
timestamp 1569543463
transform 1 0 72 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2600
timestamp 1569543463
transform 1 0 328 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2601
timestamp 1569543463
transform 1 0 264 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2602
timestamp 1569543463
transform 1 0 136 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2603
timestamp 1569543463
transform 1 0 72 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2604
timestamp 1569543463
transform 1 0 136 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2605
timestamp 1569543463
transform 1 0 264 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2606
timestamp 1569543463
transform 1 0 264 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2607
timestamp 1569543463
transform 1 0 136 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2608
timestamp 1569543463
transform 1 0 264 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2609
timestamp 1569543463
transform 1 0 200 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2610
timestamp 1569543463
transform 1 0 328 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2611
timestamp 1569543463
transform 1 0 328 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2612
timestamp 1569543463
transform 1 0 200 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2613
timestamp 1569543463
transform 1 0 200 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2614
timestamp 1569543463
transform 1 0 328 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2615
timestamp 1569543463
transform 1 0 328 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2616
timestamp 1569543463
transform 1 0 136 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2617
timestamp 1569543463
transform 1 0 136 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2618
timestamp 1569543463
transform 1 0 136 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2619
timestamp 1569543463
transform 1 0 136 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2620
timestamp 1569543463
transform 1 0 72 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2621
timestamp 1569543463
transform 1 0 72 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2622
timestamp 1569543463
transform 1 0 200 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2623
timestamp 1569543463
transform 1 0 200 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2624
timestamp 1569543463
transform 1 0 200 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2625
timestamp 1569543463
transform 1 0 200 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2626
timestamp 1569543463
transform 1 0 72 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2627
timestamp 1569543463
transform 1 0 264 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2628
timestamp 1569543463
transform 1 0 264 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2629
timestamp 1569543463
transform 1 0 264 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2630
timestamp 1569543463
transform 1 0 264 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2631
timestamp 1569543463
transform 1 0 328 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2632
timestamp 1569543463
transform 1 0 328 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2633
timestamp 1569543463
transform 1 0 328 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2634
timestamp 1569543463
transform 1 0 328 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2635
timestamp 1569543463
transform 1 0 72 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2636
timestamp 1569543463
transform 1 0 520 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2637
timestamp 1569543463
transform 1 0 520 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2638
timestamp 1569543463
transform 1 0 456 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2639
timestamp 1569543463
transform 1 0 456 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2640
timestamp 1569543463
transform 1 0 392 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2641
timestamp 1569543463
transform 1 0 392 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2642
timestamp 1569543463
transform 1 0 392 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2643
timestamp 1569543463
transform 1 0 392 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2644
timestamp 1569543463
transform 1 0 456 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2645
timestamp 1569543463
transform 1 0 456 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2646
timestamp 1569543463
transform 1 0 584 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2647
timestamp 1569543463
transform 1 0 584 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2648
timestamp 1569543463
transform 1 0 584 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2649
timestamp 1569543463
transform 1 0 520 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2650
timestamp 1569543463
transform 1 0 520 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2651
timestamp 1569543463
transform 1 0 584 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2652
timestamp 1569543463
transform 1 0 584 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2653
timestamp 1569543463
transform 1 0 392 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2654
timestamp 1569543463
transform 1 0 520 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2655
timestamp 1569543463
transform 1 0 520 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2656
timestamp 1569543463
transform 1 0 584 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2657
timestamp 1569543463
transform 1 0 520 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2658
timestamp 1569543463
transform 1 0 456 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2659
timestamp 1569543463
transform 1 0 456 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2660
timestamp 1569543463
transform 1 0 584 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2661
timestamp 1569543463
transform 1 0 520 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2662
timestamp 1569543463
transform 1 0 392 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2663
timestamp 1569543463
transform 1 0 584 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2664
timestamp 1569543463
transform 1 0 392 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2665
timestamp 1569543463
transform 1 0 456 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2666
timestamp 1569543463
transform 1 0 456 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2667
timestamp 1569543463
transform 1 0 392 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2668
timestamp 1569543463
transform 1 0 136 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2669
timestamp 1569543463
transform 1 0 328 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2670
timestamp 1569543463
transform 1 0 264 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2671
timestamp 1569543463
transform 1 0 264 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2672
timestamp 1569543463
transform 1 0 72 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2673
timestamp 1569543463
transform 1 0 200 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2674
timestamp 1569543463
transform 1 0 328 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2675
timestamp 1569543463
transform 1 0 136 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2676
timestamp 1569543463
transform 1 0 328 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2677
timestamp 1569543463
transform 1 0 72 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2678
timestamp 1569543463
transform 1 0 264 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2679
timestamp 1569543463
transform 1 0 328 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2680
timestamp 1569543463
transform 1 0 136 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2681
timestamp 1569543463
transform 1 0 264 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2682
timestamp 1569543463
transform 1 0 136 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2683
timestamp 1569543463
transform 1 0 72 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2684
timestamp 1569543463
transform 1 0 200 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2685
timestamp 1569543463
transform 1 0 200 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2686
timestamp 1569543463
transform 1 0 200 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2687
timestamp 1569543463
transform 1 0 72 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2688
timestamp 1569543463
transform 1 0 264 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2689
timestamp 1569543463
transform 1 0 264 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2690
timestamp 1569543463
transform 1 0 200 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2691
timestamp 1569543463
transform 1 0 136 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2692
timestamp 1569543463
transform 1 0 136 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2693
timestamp 1569543463
transform 1 0 136 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2694
timestamp 1569543463
transform 1 0 136 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2695
timestamp 1569543463
transform 1 0 72 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2696
timestamp 1569543463
transform 1 0 328 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2697
timestamp 1569543463
transform 1 0 328 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2698
timestamp 1569543463
transform 1 0 328 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2699
timestamp 1569543463
transform 1 0 328 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2700
timestamp 1569543463
transform 1 0 72 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2701
timestamp 1569543463
transform 1 0 72 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2702
timestamp 1569543463
transform 1 0 264 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2703
timestamp 1569543463
transform 1 0 200 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2704
timestamp 1569543463
transform 1 0 200 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2705
timestamp 1569543463
transform 1 0 200 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2706
timestamp 1569543463
transform 1 0 264 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2707
timestamp 1569543463
transform 1 0 72 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2708
timestamp 1569543463
transform 1 0 392 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2709
timestamp 1569543463
transform 1 0 392 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2710
timestamp 1569543463
transform 1 0 392 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2711
timestamp 1569543463
transform 1 0 392 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2712
timestamp 1569543463
transform 1 0 456 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2713
timestamp 1569543463
transform 1 0 456 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2714
timestamp 1569543463
transform 1 0 456 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2715
timestamp 1569543463
transform 1 0 456 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2716
timestamp 1569543463
transform 1 0 520 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2717
timestamp 1569543463
transform 1 0 520 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2718
timestamp 1569543463
transform 1 0 520 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2719
timestamp 1569543463
transform 1 0 520 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2720
timestamp 1569543463
transform 1 0 584 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2721
timestamp 1569543463
transform 1 0 584 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2722
timestamp 1569543463
transform 1 0 584 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2723
timestamp 1569543463
transform 1 0 584 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2724
timestamp 1569543463
transform 1 0 1096 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2725
timestamp 1569543463
transform 1 0 1160 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2726
timestamp 1569543463
transform 1 0 968 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2727
timestamp 1569543463
transform 1 0 1096 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2728
timestamp 1569543463
transform 1 0 1224 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2729
timestamp 1569543463
transform 1 0 968 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2730
timestamp 1569543463
transform 1 0 1096 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2731
timestamp 1569543463
transform 1 0 1224 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2732
timestamp 1569543463
transform 1 0 1096 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2733
timestamp 1569543463
transform 1 0 1224 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2734
timestamp 1569543463
transform 1 0 968 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2735
timestamp 1569543463
transform 1 0 968 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2736
timestamp 1569543463
transform 1 0 1160 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2737
timestamp 1569543463
transform 1 0 1160 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2738
timestamp 1569543463
transform 1 0 1032 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2739
timestamp 1569543463
transform 1 0 1032 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2740
timestamp 1569543463
transform 1 0 1032 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2741
timestamp 1569543463
transform 1 0 1032 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2742
timestamp 1569543463
transform 1 0 1224 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2743
timestamp 1569543463
transform 1 0 1160 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2744
timestamp 1569543463
transform 1 0 712 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2745
timestamp 1569543463
transform 1 0 840 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2746
timestamp 1569543463
transform 1 0 776 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2747
timestamp 1569543463
transform 1 0 776 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2748
timestamp 1569543463
transform 1 0 904 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2749
timestamp 1569543463
transform 1 0 776 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2750
timestamp 1569543463
transform 1 0 904 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2751
timestamp 1569543463
transform 1 0 840 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2752
timestamp 1569543463
transform 1 0 840 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2753
timestamp 1569543463
transform 1 0 840 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2754
timestamp 1569543463
transform 1 0 904 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2755
timestamp 1569543463
transform 1 0 776 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2756
timestamp 1569543463
transform 1 0 904 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2757
timestamp 1569543463
transform 1 0 712 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2758
timestamp 1569543463
transform 1 0 712 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2759
timestamp 1569543463
transform 1 0 712 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2760
timestamp 1569543463
transform 1 0 904 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2761
timestamp 1569543463
transform 1 0 904 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2762
timestamp 1569543463
transform 1 0 904 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2763
timestamp 1569543463
transform 1 0 776 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2764
timestamp 1569543463
transform 1 0 840 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2765
timestamp 1569543463
transform 1 0 776 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2766
timestamp 1569543463
transform 1 0 776 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2767
timestamp 1569543463
transform 1 0 776 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2768
timestamp 1569543463
transform 1 0 840 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2769
timestamp 1569543463
transform 1 0 712 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2770
timestamp 1569543463
transform 1 0 712 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2771
timestamp 1569543463
transform 1 0 840 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2772
timestamp 1569543463
transform 1 0 712 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2773
timestamp 1569543463
transform 1 0 712 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2774
timestamp 1569543463
transform 1 0 904 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2775
timestamp 1569543463
transform 1 0 840 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2776
timestamp 1569543463
transform 1 0 968 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2777
timestamp 1569543463
transform 1 0 968 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2778
timestamp 1569543463
transform 1 0 968 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2779
timestamp 1569543463
transform 1 0 968 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2780
timestamp 1569543463
transform 1 0 1032 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2781
timestamp 1569543463
transform 1 0 1032 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2782
timestamp 1569543463
transform 1 0 1032 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2783
timestamp 1569543463
transform 1 0 1032 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2784
timestamp 1569543463
transform 1 0 1096 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2785
timestamp 1569543463
transform 1 0 1096 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2786
timestamp 1569543463
transform 1 0 1096 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2787
timestamp 1569543463
transform 1 0 1096 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2788
timestamp 1569543463
transform 1 0 1160 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2789
timestamp 1569543463
transform 1 0 1160 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2790
timestamp 1569543463
transform 1 0 1160 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2791
timestamp 1569543463
transform 1 0 1160 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2792
timestamp 1569543463
transform 1 0 1224 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2793
timestamp 1569543463
transform 1 0 1224 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2794
timestamp 1569543463
transform 1 0 1224 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2795
timestamp 1569543463
transform 1 0 1224 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2796
timestamp 1569543463
transform 1 0 456 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2797
timestamp 1569543463
transform 1 0 1096 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2798
timestamp 1569543463
transform 1 0 136 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2799
timestamp 1569543463
transform 1 0 776 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2800
timestamp 1569543463
transform 1 0 520 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2801
timestamp 1569543463
transform 1 0 1160 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2802
timestamp 1569543463
transform 1 0 200 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2803
timestamp 1569543463
transform 1 0 840 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2804
timestamp 1569543463
transform 1 0 264 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2805
timestamp 1569543463
transform 1 0 904 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2806
timestamp 1569543463
transform 1 0 328 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2807
timestamp 1569543463
transform 1 0 968 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2808
timestamp 1569543463
transform 1 0 392 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2809
timestamp 1569543463
transform 1 0 1032 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2810
timestamp 1569543463
transform 1 0 648 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2811
timestamp 1569543463
transform 1 0 584 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2812
timestamp 1569543463
transform 1 0 1224 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2813
timestamp 1569543463
transform 1 0 648 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2814
timestamp 1569543463
transform 1 0 648 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2815
timestamp 1569543463
transform 1 0 648 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2816
timestamp 1569543463
transform 1 0 648 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2817
timestamp 1569543463
transform 1 0 648 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2818
timestamp 1569543463
transform 1 0 648 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2819
timestamp 1569543463
transform 1 0 648 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2820
timestamp 1569543463
transform 1 0 648 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2821
timestamp 1569543463
transform 1 0 648 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2822
timestamp 1569543463
transform 1 0 648 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2823
timestamp 1569543463
transform 1 0 648 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2824
timestamp 1569543463
transform 1 0 648 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2825
timestamp 1569543463
transform 1 0 72 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2826
timestamp 1569543463
transform 1 0 712 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2827
timestamp 1569543463
transform 1 0 648 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2828
timestamp 1569543463
transform 1 0 648 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2829
timestamp 1569543463
transform 1 0 648 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2830
timestamp 1569543463
transform 1 0 648 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2831
timestamp 1569543463
transform 1 0 648 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2832
timestamp 1569543463
transform 1 0 2376 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2833
timestamp 1569543463
transform 1 0 2440 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2834
timestamp 1569543463
transform 1 0 2376 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2835
timestamp 1569543463
transform 1 0 2376 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2836
timestamp 1569543463
transform 1 0 2376 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2837
timestamp 1569543463
transform 1 0 2376 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2838
timestamp 1569543463
transform 1 0 2376 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2839
timestamp 1569543463
transform 1 0 2376 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2840
timestamp 1569543463
transform 1 0 2440 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2841
timestamp 1569543463
transform 1 0 2440 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2842
timestamp 1569543463
transform 1 0 2312 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2843
timestamp 1569543463
transform 1 0 2312 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2844
timestamp 1569543463
transform 1 0 2312 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2845
timestamp 1569543463
transform 1 0 2312 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2846
timestamp 1569543463
transform 1 0 2312 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2847
timestamp 1569543463
transform 1 0 2440 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2848
timestamp 1569543463
transform 1 0 2440 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2849
timestamp 1569543463
transform 1 0 2440 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2850
timestamp 1569543463
transform 1 0 2440 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2851
timestamp 1569543463
transform 1 0 2440 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2852
timestamp 1569543463
transform 1 0 2312 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2853
timestamp 1569543463
transform 1 0 2312 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2854
timestamp 1569543463
transform 1 0 2312 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2855
timestamp 1569543463
transform 1 0 2312 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2856
timestamp 1569543463
transform 1 0 2440 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2857
timestamp 1569543463
transform 1 0 2376 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2858
timestamp 1569543463
transform 1 0 2376 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2859
timestamp 1569543463
transform 1 0 1352 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2860
timestamp 1569543463
transform 1 0 1352 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2861
timestamp 1569543463
transform 1 0 1352 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2862
timestamp 1569543463
transform 1 0 1352 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2863
timestamp 1569543463
transform 1 0 1288 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2864
timestamp 1569543463
transform 1 0 1352 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2865
timestamp 1569543463
transform 1 0 1352 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2866
timestamp 1569543463
transform 1 0 1416 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2867
timestamp 1569543463
transform 1 0 1352 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2868
timestamp 1569543463
transform 1 0 1416 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2869
timestamp 1569543463
transform 1 0 1416 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2870
timestamp 1569543463
transform 1 0 1416 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2871
timestamp 1569543463
transform 1 0 1416 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2872
timestamp 1569543463
transform 1 0 1480 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2873
timestamp 1569543463
transform 1 0 1480 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2874
timestamp 1569543463
transform 1 0 1288 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2875
timestamp 1569543463
transform 1 0 1480 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2876
timestamp 1569543463
transform 1 0 1480 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2877
timestamp 1569543463
transform 1 0 1352 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2878
timestamp 1569543463
transform 1 0 1288 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2879
timestamp 1569543463
transform 1 0 1416 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2880
timestamp 1569543463
transform 1 0 1416 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2881
timestamp 1569543463
transform 1 0 1416 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2882
timestamp 1569543463
transform 1 0 1416 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2883
timestamp 1569543463
transform 1 0 1288 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2884
timestamp 1569543463
transform 1 0 1480 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_2885
timestamp 1569543463
transform 1 0 1480 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_2886
timestamp 1569543463
transform 1 0 1480 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_2887
timestamp 1569543463
transform 1 0 1480 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_2888
timestamp 1569543463
transform 1 0 1352 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2889
timestamp 1569543463
transform 1 0 1288 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2890
timestamp 1569543463
transform 1 0 1480 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_2891
timestamp 1569543463
transform 1 0 1288 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_2892
timestamp 1569543463
transform 1 0 1288 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_2893
timestamp 1569543463
transform 1 0 1288 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_2894
timestamp 1569543463
transform 1 0 1288 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_2895
timestamp 1569543463
transform 1 0 1352 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2896
timestamp 1569543463
transform 1 0 1480 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2897
timestamp 1569543463
transform 1 0 1480 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2898
timestamp 1569543463
transform 1 0 1416 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2899
timestamp 1569543463
transform 1 0 1416 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2900
timestamp 1569543463
transform 1 0 1480 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2901
timestamp 1569543463
transform 1 0 1480 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2902
timestamp 1569543463
transform 1 0 1352 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2903
timestamp 1569543463
transform 1 0 1352 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2904
timestamp 1569543463
transform 1 0 1352 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2905
timestamp 1569543463
transform 1 0 1352 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2906
timestamp 1569543463
transform 1 0 1352 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2907
timestamp 1569543463
transform 1 0 1480 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2908
timestamp 1569543463
transform 1 0 1352 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2909
timestamp 1569543463
transform 1 0 1480 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2910
timestamp 1569543463
transform 1 0 1352 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2911
timestamp 1569543463
transform 1 0 1416 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2912
timestamp 1569543463
transform 1 0 1416 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2913
timestamp 1569543463
transform 1 0 1480 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2914
timestamp 1569543463
transform 1 0 1416 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2915
timestamp 1569543463
transform 1 0 1416 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2916
timestamp 1569543463
transform 1 0 1416 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2917
timestamp 1569543463
transform 1 0 1288 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2918
timestamp 1569543463
transform 1 0 1288 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2919
timestamp 1569543463
transform 1 0 1416 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2920
timestamp 1569543463
transform 1 0 1288 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2921
timestamp 1569543463
transform 1 0 1288 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2922
timestamp 1569543463
transform 1 0 1288 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2923
timestamp 1569543463
transform 1 0 1288 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2924
timestamp 1569543463
transform 1 0 1288 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2925
timestamp 1569543463
transform 1 0 1288 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2926
timestamp 1569543463
transform 1 0 1480 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2927
timestamp 1569543463
transform 1 0 2376 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2928
timestamp 1569543463
transform 1 0 2312 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2929
timestamp 1569543463
transform 1 0 2312 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2930
timestamp 1569543463
transform 1 0 2312 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2931
timestamp 1569543463
transform 1 0 2312 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2932
timestamp 1569543463
transform 1 0 2312 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2933
timestamp 1569543463
transform 1 0 2312 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2934
timestamp 1569543463
transform 1 0 2376 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2935
timestamp 1569543463
transform 1 0 2376 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2936
timestamp 1569543463
transform 1 0 2376 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2937
timestamp 1569543463
transform 1 0 2376 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2938
timestamp 1569543463
transform 1 0 2376 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2939
timestamp 1569543463
transform 1 0 2440 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_2940
timestamp 1569543463
transform 1 0 2440 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_2941
timestamp 1569543463
transform 1 0 2440 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_2942
timestamp 1569543463
transform 1 0 2440 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_2943
timestamp 1569543463
transform 1 0 2440 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_2944
timestamp 1569543463
transform 1 0 2312 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2945
timestamp 1569543463
transform 1 0 2440 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_2946
timestamp 1569543463
transform 1 0 2376 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2947
timestamp 1569543463
transform 1 0 2312 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2948
timestamp 1569543463
transform 1 0 2440 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_2949
timestamp 1569543463
transform 1 0 2376 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2950
timestamp 1569543463
transform 1 0 2440 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_2951
timestamp 1569543463
transform 1 0 1416 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2952
timestamp 1569543463
transform 1 0 1480 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2953
timestamp 1569543463
transform 1 0 2312 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2954
timestamp 1569543463
transform 1 0 2376 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2955
timestamp 1569543463
transform 1 0 2440 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2956
timestamp 1569543463
transform 1 0 1288 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2957
timestamp 1569543463
transform 1 0 1352 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_2958
timestamp 1569543463
transform 1 0 4680 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2959
timestamp 1569543463
transform 1 0 4744 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2960
timestamp 1569543463
transform 1 0 4872 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2961
timestamp 1569543463
transform 1 0 4872 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2962
timestamp 1569543463
transform 1 0 4744 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2963
timestamp 1569543463
transform 1 0 4680 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2964
timestamp 1569543463
transform 1 0 4680 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2965
timestamp 1569543463
transform 1 0 4744 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2966
timestamp 1569543463
transform 1 0 4680 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2967
timestamp 1569543463
transform 1 0 4808 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2968
timestamp 1569543463
transform 1 0 4744 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2969
timestamp 1569543463
transform 1 0 4872 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2970
timestamp 1569543463
transform 1 0 4808 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2971
timestamp 1569543463
transform 1 0 4808 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2972
timestamp 1569543463
transform 1 0 4808 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2973
timestamp 1569543463
transform 1 0 4872 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2974
timestamp 1569543463
transform 1 0 4616 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2975
timestamp 1569543463
transform 1 0 4488 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2976
timestamp 1569543463
transform 1 0 4424 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2977
timestamp 1569543463
transform 1 0 4424 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2978
timestamp 1569543463
transform 1 0 4488 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2979
timestamp 1569543463
transform 1 0 4616 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2980
timestamp 1569543463
transform 1 0 4488 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2981
timestamp 1569543463
transform 1 0 4616 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2982
timestamp 1569543463
transform 1 0 4616 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2983
timestamp 1569543463
transform 1 0 4552 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2984
timestamp 1569543463
transform 1 0 4552 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_2985
timestamp 1569543463
transform 1 0 4552 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2986
timestamp 1569543463
transform 1 0 4424 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2987
timestamp 1569543463
transform 1 0 4552 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_2988
timestamp 1569543463
transform 1 0 4424 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_2989
timestamp 1569543463
transform 1 0 4488 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_2990
timestamp 1569543463
transform 1 0 4616 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_2991
timestamp 1569543463
transform 1 0 4552 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2992
timestamp 1569543463
transform 1 0 4424 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2993
timestamp 1569543463
transform 1 0 4616 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_2994
timestamp 1569543463
transform 1 0 4488 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_2995
timestamp 1569543463
transform 1 0 4616 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2996
timestamp 1569543463
transform 1 0 4616 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2997
timestamp 1569543463
transform 1 0 4488 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_2998
timestamp 1569543463
transform 1 0 4488 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_2999
timestamp 1569543463
transform 1 0 4488 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3000
timestamp 1569543463
transform 1 0 4552 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3001
timestamp 1569543463
transform 1 0 4424 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3002
timestamp 1569543463
transform 1 0 4424 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3003
timestamp 1569543463
transform 1 0 4488 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3004
timestamp 1569543463
transform 1 0 4424 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3005
timestamp 1569543463
transform 1 0 4552 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3006
timestamp 1569543463
transform 1 0 4424 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3007
timestamp 1569543463
transform 1 0 4552 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3008
timestamp 1569543463
transform 1 0 4552 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3009
timestamp 1569543463
transform 1 0 4616 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3010
timestamp 1569543463
transform 1 0 4872 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3011
timestamp 1569543463
transform 1 0 4744 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3012
timestamp 1569543463
transform 1 0 4872 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3013
timestamp 1569543463
transform 1 0 4744 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3014
timestamp 1569543463
transform 1 0 4872 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3015
timestamp 1569543463
transform 1 0 4808 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3016
timestamp 1569543463
transform 1 0 4744 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3017
timestamp 1569543463
transform 1 0 4680 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3018
timestamp 1569543463
transform 1 0 4808 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3019
timestamp 1569543463
transform 1 0 4680 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3020
timestamp 1569543463
transform 1 0 4808 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3021
timestamp 1569543463
transform 1 0 4808 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3022
timestamp 1569543463
transform 1 0 4680 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3023
timestamp 1569543463
transform 1 0 4872 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3024
timestamp 1569543463
transform 1 0 4872 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3025
timestamp 1569543463
transform 1 0 4680 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3026
timestamp 1569543463
transform 1 0 4680 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3027
timestamp 1569543463
transform 1 0 4744 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3028
timestamp 1569543463
transform 1 0 4808 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3029
timestamp 1569543463
transform 1 0 4744 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3030
timestamp 1569543463
transform 1 0 4104 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3031
timestamp 1569543463
transform 1 0 4232 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3032
timestamp 1569543463
transform 1 0 4104 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3033
timestamp 1569543463
transform 1 0 4232 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3034
timestamp 1569543463
transform 1 0 4168 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3035
timestamp 1569543463
transform 1 0 4296 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3036
timestamp 1569543463
transform 1 0 4296 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3037
timestamp 1569543463
transform 1 0 4168 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3038
timestamp 1569543463
transform 1 0 4296 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3039
timestamp 1569543463
transform 1 0 4104 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3040
timestamp 1569543463
transform 1 0 4232 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3041
timestamp 1569543463
transform 1 0 4168 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3042
timestamp 1569543463
transform 1 0 4168 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3043
timestamp 1569543463
transform 1 0 4232 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3044
timestamp 1569543463
transform 1 0 4104 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3045
timestamp 1569543463
transform 1 0 4296 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3046
timestamp 1569543463
transform 1 0 3848 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3047
timestamp 1569543463
transform 1 0 3976 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3048
timestamp 1569543463
transform 1 0 3912 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3049
timestamp 1569543463
transform 1 0 3976 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3050
timestamp 1569543463
transform 1 0 3784 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3051
timestamp 1569543463
transform 1 0 3848 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3052
timestamp 1569543463
transform 1 0 3976 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3053
timestamp 1569543463
transform 1 0 3784 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3054
timestamp 1569543463
transform 1 0 4040 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3055
timestamp 1569543463
transform 1 0 3976 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3056
timestamp 1569543463
transform 1 0 3912 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3057
timestamp 1569543463
transform 1 0 3912 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3058
timestamp 1569543463
transform 1 0 3848 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3059
timestamp 1569543463
transform 1 0 3848 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3060
timestamp 1569543463
transform 1 0 3784 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3061
timestamp 1569543463
transform 1 0 4040 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3062
timestamp 1569543463
transform 1 0 4040 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3063
timestamp 1569543463
transform 1 0 3912 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3064
timestamp 1569543463
transform 1 0 4040 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3065
timestamp 1569543463
transform 1 0 3784 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3066
timestamp 1569543463
transform 1 0 3912 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3067
timestamp 1569543463
transform 1 0 3784 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3068
timestamp 1569543463
transform 1 0 3848 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3069
timestamp 1569543463
transform 1 0 4040 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3070
timestamp 1569543463
transform 1 0 3848 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3071
timestamp 1569543463
transform 1 0 3976 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3072
timestamp 1569543463
transform 1 0 3976 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3073
timestamp 1569543463
transform 1 0 3848 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3074
timestamp 1569543463
transform 1 0 3976 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3075
timestamp 1569543463
transform 1 0 3912 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3076
timestamp 1569543463
transform 1 0 3784 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3077
timestamp 1569543463
transform 1 0 3976 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3078
timestamp 1569543463
transform 1 0 4040 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3079
timestamp 1569543463
transform 1 0 3784 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3080
timestamp 1569543463
transform 1 0 3912 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3081
timestamp 1569543463
transform 1 0 4040 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3082
timestamp 1569543463
transform 1 0 3784 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3083
timestamp 1569543463
transform 1 0 3848 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3084
timestamp 1569543463
transform 1 0 4040 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3085
timestamp 1569543463
transform 1 0 4040 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3086
timestamp 1569543463
transform 1 0 3912 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3087
timestamp 1569543463
transform 1 0 3848 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3088
timestamp 1569543463
transform 1 0 3784 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3089
timestamp 1569543463
transform 1 0 3976 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3090
timestamp 1569543463
transform 1 0 3912 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3091
timestamp 1569543463
transform 1 0 4104 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3092
timestamp 1569543463
transform 1 0 4104 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3093
timestamp 1569543463
transform 1 0 4232 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3094
timestamp 1569543463
transform 1 0 4104 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3095
timestamp 1569543463
transform 1 0 4232 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3096
timestamp 1569543463
transform 1 0 4168 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3097
timestamp 1569543463
transform 1 0 4296 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3098
timestamp 1569543463
transform 1 0 4168 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3099
timestamp 1569543463
transform 1 0 4232 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3100
timestamp 1569543463
transform 1 0 4296 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3101
timestamp 1569543463
transform 1 0 4168 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3102
timestamp 1569543463
transform 1 0 4104 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3103
timestamp 1569543463
transform 1 0 4104 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3104
timestamp 1569543463
transform 1 0 4168 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3105
timestamp 1569543463
transform 1 0 4168 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3106
timestamp 1569543463
transform 1 0 4232 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3107
timestamp 1569543463
transform 1 0 4232 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3108
timestamp 1569543463
transform 1 0 4296 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3109
timestamp 1569543463
transform 1 0 4296 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3110
timestamp 1569543463
transform 1 0 4296 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3111
timestamp 1569543463
transform 1 0 4168 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3112
timestamp 1569543463
transform 1 0 4232 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3113
timestamp 1569543463
transform 1 0 4104 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3114
timestamp 1569543463
transform 1 0 4104 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3115
timestamp 1569543463
transform 1 0 4232 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3116
timestamp 1569543463
transform 1 0 4168 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3117
timestamp 1569543463
transform 1 0 4232 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3118
timestamp 1569543463
transform 1 0 4104 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3119
timestamp 1569543463
transform 1 0 4104 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3120
timestamp 1569543463
transform 1 0 4168 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3121
timestamp 1569543463
transform 1 0 4104 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3122
timestamp 1569543463
transform 1 0 4296 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3123
timestamp 1569543463
transform 1 0 4232 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3124
timestamp 1569543463
transform 1 0 4168 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3125
timestamp 1569543463
transform 1 0 4232 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3126
timestamp 1569543463
transform 1 0 4296 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3127
timestamp 1569543463
transform 1 0 4296 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3128
timestamp 1569543463
transform 1 0 4296 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3129
timestamp 1569543463
transform 1 0 4296 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3130
timestamp 1569543463
transform 1 0 4168 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3131
timestamp 1569543463
transform 1 0 3848 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3132
timestamp 1569543463
transform 1 0 4040 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3133
timestamp 1569543463
transform 1 0 3912 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3134
timestamp 1569543463
transform 1 0 3848 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3135
timestamp 1569543463
transform 1 0 3784 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3136
timestamp 1569543463
transform 1 0 3784 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3137
timestamp 1569543463
transform 1 0 3848 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3138
timestamp 1569543463
transform 1 0 3784 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3139
timestamp 1569543463
transform 1 0 3912 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3140
timestamp 1569543463
transform 1 0 3976 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3141
timestamp 1569543463
transform 1 0 3912 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3142
timestamp 1569543463
transform 1 0 3848 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3143
timestamp 1569543463
transform 1 0 3976 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3144
timestamp 1569543463
transform 1 0 3976 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3145
timestamp 1569543463
transform 1 0 3784 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3146
timestamp 1569543463
transform 1 0 3976 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3147
timestamp 1569543463
transform 1 0 3976 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3148
timestamp 1569543463
transform 1 0 3784 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3149
timestamp 1569543463
transform 1 0 4040 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3150
timestamp 1569543463
transform 1 0 3912 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3151
timestamp 1569543463
transform 1 0 4040 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3152
timestamp 1569543463
transform 1 0 3848 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3153
timestamp 1569543463
transform 1 0 4040 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3154
timestamp 1569543463
transform 1 0 3912 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3155
timestamp 1569543463
transform 1 0 4040 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3156
timestamp 1569543463
transform 1 0 4040 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3157
timestamp 1569543463
transform 1 0 3784 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3158
timestamp 1569543463
transform 1 0 3784 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3159
timestamp 1569543463
transform 1 0 3784 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3160
timestamp 1569543463
transform 1 0 3784 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3161
timestamp 1569543463
transform 1 0 4040 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3162
timestamp 1569543463
transform 1 0 3912 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3163
timestamp 1569543463
transform 1 0 3912 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3164
timestamp 1569543463
transform 1 0 3976 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3165
timestamp 1569543463
transform 1 0 3976 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3166
timestamp 1569543463
transform 1 0 3976 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3167
timestamp 1569543463
transform 1 0 3848 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3168
timestamp 1569543463
transform 1 0 3976 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3169
timestamp 1569543463
transform 1 0 3976 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3170
timestamp 1569543463
transform 1 0 3848 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3171
timestamp 1569543463
transform 1 0 3848 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3172
timestamp 1569543463
transform 1 0 3848 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3173
timestamp 1569543463
transform 1 0 4040 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3174
timestamp 1569543463
transform 1 0 3912 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3175
timestamp 1569543463
transform 1 0 4040 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3176
timestamp 1569543463
transform 1 0 3912 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3177
timestamp 1569543463
transform 1 0 3912 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3178
timestamp 1569543463
transform 1 0 3848 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3179
timestamp 1569543463
transform 1 0 4040 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3180
timestamp 1569543463
transform 1 0 3784 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3181
timestamp 1569543463
transform 1 0 4232 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3182
timestamp 1569543463
transform 1 0 4232 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3183
timestamp 1569543463
transform 1 0 4232 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3184
timestamp 1569543463
transform 1 0 4104 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3185
timestamp 1569543463
transform 1 0 4296 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3186
timestamp 1569543463
transform 1 0 4296 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3187
timestamp 1569543463
transform 1 0 4296 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3188
timestamp 1569543463
transform 1 0 4104 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3189
timestamp 1569543463
transform 1 0 4168 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3190
timestamp 1569543463
transform 1 0 4104 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3191
timestamp 1569543463
transform 1 0 4104 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3192
timestamp 1569543463
transform 1 0 4296 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3193
timestamp 1569543463
transform 1 0 4296 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3194
timestamp 1569543463
transform 1 0 4168 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3195
timestamp 1569543463
transform 1 0 4168 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3196
timestamp 1569543463
transform 1 0 4232 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3197
timestamp 1569543463
transform 1 0 4232 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3198
timestamp 1569543463
transform 1 0 4168 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3199
timestamp 1569543463
transform 1 0 4168 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3200
timestamp 1569543463
transform 1 0 4104 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3201
timestamp 1569543463
transform 1 0 4744 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3202
timestamp 1569543463
transform 1 0 4744 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3203
timestamp 1569543463
transform 1 0 4744 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3204
timestamp 1569543463
transform 1 0 4744 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3205
timestamp 1569543463
transform 1 0 4744 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3206
timestamp 1569543463
transform 1 0 4808 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3207
timestamp 1569543463
transform 1 0 4808 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3208
timestamp 1569543463
transform 1 0 4808 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3209
timestamp 1569543463
transform 1 0 4872 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3210
timestamp 1569543463
transform 1 0 4680 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3211
timestamp 1569543463
transform 1 0 4808 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3212
timestamp 1569543463
transform 1 0 4808 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3213
timestamp 1569543463
transform 1 0 4872 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3214
timestamp 1569543463
transform 1 0 4680 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3215
timestamp 1569543463
transform 1 0 4680 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3216
timestamp 1569543463
transform 1 0 4872 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3217
timestamp 1569543463
transform 1 0 4680 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3218
timestamp 1569543463
transform 1 0 4680 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3219
timestamp 1569543463
transform 1 0 4872 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3220
timestamp 1569543463
transform 1 0 4872 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3221
timestamp 1569543463
transform 1 0 4552 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3222
timestamp 1569543463
transform 1 0 4488 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3223
timestamp 1569543463
transform 1 0 4488 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3224
timestamp 1569543463
transform 1 0 4488 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3225
timestamp 1569543463
transform 1 0 4616 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3226
timestamp 1569543463
transform 1 0 4552 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3227
timestamp 1569543463
transform 1 0 4424 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3228
timestamp 1569543463
transform 1 0 4616 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3229
timestamp 1569543463
transform 1 0 4616 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3230
timestamp 1569543463
transform 1 0 4616 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3231
timestamp 1569543463
transform 1 0 4616 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3232
timestamp 1569543463
transform 1 0 4552 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3233
timestamp 1569543463
transform 1 0 4552 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3234
timestamp 1569543463
transform 1 0 4552 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3235
timestamp 1569543463
transform 1 0 4424 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3236
timestamp 1569543463
transform 1 0 4424 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3237
timestamp 1569543463
transform 1 0 4424 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3238
timestamp 1569543463
transform 1 0 4424 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3239
timestamp 1569543463
transform 1 0 4488 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3240
timestamp 1569543463
transform 1 0 4488 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3241
timestamp 1569543463
transform 1 0 4552 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3242
timestamp 1569543463
transform 1 0 4616 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3243
timestamp 1569543463
transform 1 0 4616 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3244
timestamp 1569543463
transform 1 0 4424 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3245
timestamp 1569543463
transform 1 0 4424 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3246
timestamp 1569543463
transform 1 0 4424 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3247
timestamp 1569543463
transform 1 0 4424 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3248
timestamp 1569543463
transform 1 0 4424 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3249
timestamp 1569543463
transform 1 0 4488 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3250
timestamp 1569543463
transform 1 0 4616 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3251
timestamp 1569543463
transform 1 0 4616 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3252
timestamp 1569543463
transform 1 0 4616 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3253
timestamp 1569543463
transform 1 0 4488 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3254
timestamp 1569543463
transform 1 0 4488 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3255
timestamp 1569543463
transform 1 0 4488 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3256
timestamp 1569543463
transform 1 0 4488 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3257
timestamp 1569543463
transform 1 0 4552 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3258
timestamp 1569543463
transform 1 0 4552 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3259
timestamp 1569543463
transform 1 0 4552 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3260
timestamp 1569543463
transform 1 0 4552 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3261
timestamp 1569543463
transform 1 0 4680 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3262
timestamp 1569543463
transform 1 0 4680 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3263
timestamp 1569543463
transform 1 0 4744 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3264
timestamp 1569543463
transform 1 0 4744 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3265
timestamp 1569543463
transform 1 0 4808 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3266
timestamp 1569543463
transform 1 0 4808 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3267
timestamp 1569543463
transform 1 0 4872 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3268
timestamp 1569543463
transform 1 0 4872 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3269
timestamp 1569543463
transform 1 0 4680 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3270
timestamp 1569543463
transform 1 0 4680 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3271
timestamp 1569543463
transform 1 0 4680 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3272
timestamp 1569543463
transform 1 0 4744 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3273
timestamp 1569543463
transform 1 0 4744 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3274
timestamp 1569543463
transform 1 0 4744 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3275
timestamp 1569543463
transform 1 0 4808 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3276
timestamp 1569543463
transform 1 0 4808 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3277
timestamp 1569543463
transform 1 0 4808 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3278
timestamp 1569543463
transform 1 0 4872 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3279
timestamp 1569543463
transform 1 0 4872 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3280
timestamp 1569543463
transform 1 0 4872 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3281
timestamp 1569543463
transform 1 0 4360 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3282
timestamp 1569543463
transform 1 0 4360 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3283
timestamp 1569543463
transform 1 0 4360 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3284
timestamp 1569543463
transform 1 0 4360 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3285
timestamp 1569543463
transform 1 0 4360 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3286
timestamp 1569543463
transform 1 0 4360 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3287
timestamp 1569543463
transform 1 0 4360 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3288
timestamp 1569543463
transform 1 0 4360 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3289
timestamp 1569543463
transform 1 0 4360 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3290
timestamp 1569543463
transform 1 0 4360 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3291
timestamp 1569543463
transform 1 0 4360 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3292
timestamp 1569543463
transform 1 0 4360 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3293
timestamp 1569543463
transform 1 0 4360 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3294
timestamp 1569543463
transform 1 0 4360 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3295
timestamp 1569543463
transform 1 0 4360 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3296
timestamp 1569543463
transform 1 0 4360 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3297
timestamp 1569543463
transform 1 0 4360 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3298
timestamp 1569543463
transform 1 0 4360 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3299
timestamp 1569543463
transform 1 0 4360 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3300
timestamp 1569543463
transform 1 0 3464 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3301
timestamp 1569543463
transform 1 0 3720 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3302
timestamp 1569543463
transform 1 0 3592 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3303
timestamp 1569543463
transform 1 0 3720 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3304
timestamp 1569543463
transform 1 0 3464 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3305
timestamp 1569543463
transform 1 0 3592 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3306
timestamp 1569543463
transform 1 0 3464 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3307
timestamp 1569543463
transform 1 0 3656 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3308
timestamp 1569543463
transform 1 0 3528 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3309
timestamp 1569543463
transform 1 0 3656 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3310
timestamp 1569543463
transform 1 0 3720 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3311
timestamp 1569543463
transform 1 0 3528 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3312
timestamp 1569543463
transform 1 0 3592 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3313
timestamp 1569543463
transform 1 0 3528 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3314
timestamp 1569543463
transform 1 0 3528 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3315
timestamp 1569543463
transform 1 0 3656 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3316
timestamp 1569543463
transform 1 0 3656 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3317
timestamp 1569543463
transform 1 0 3592 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3318
timestamp 1569543463
transform 1 0 3464 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3319
timestamp 1569543463
transform 1 0 3720 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3320
timestamp 1569543463
transform 1 0 3336 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3321
timestamp 1569543463
transform 1 0 3336 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3322
timestamp 1569543463
transform 1 0 3208 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3323
timestamp 1569543463
transform 1 0 3336 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3324
timestamp 1569543463
transform 1 0 3400 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3325
timestamp 1569543463
transform 1 0 3144 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3326
timestamp 1569543463
transform 1 0 3400 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3327
timestamp 1569543463
transform 1 0 3208 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3328
timestamp 1569543463
transform 1 0 3272 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3329
timestamp 1569543463
transform 1 0 3400 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3330
timestamp 1569543463
transform 1 0 3144 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3331
timestamp 1569543463
transform 1 0 3144 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3332
timestamp 1569543463
transform 1 0 3208 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3333
timestamp 1569543463
transform 1 0 3144 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3334
timestamp 1569543463
transform 1 0 3400 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3335
timestamp 1569543463
transform 1 0 3272 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3336
timestamp 1569543463
transform 1 0 3208 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3337
timestamp 1569543463
transform 1 0 3272 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3338
timestamp 1569543463
transform 1 0 3336 0 1 2568
box -8 -8 8 8
use VIA1$5  VIA1$5_3339
timestamp 1569543463
transform 1 0 3272 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3340
timestamp 1569543463
transform 1 0 3336 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3341
timestamp 1569543463
transform 1 0 3208 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3342
timestamp 1569543463
transform 1 0 3272 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3343
timestamp 1569543463
transform 1 0 3208 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3344
timestamp 1569543463
transform 1 0 3144 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3345
timestamp 1569543463
transform 1 0 3400 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3346
timestamp 1569543463
transform 1 0 3400 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3347
timestamp 1569543463
transform 1 0 3272 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3348
timestamp 1569543463
transform 1 0 3336 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3349
timestamp 1569543463
transform 1 0 3272 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3350
timestamp 1569543463
transform 1 0 3208 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3351
timestamp 1569543463
transform 1 0 3336 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3352
timestamp 1569543463
transform 1 0 3272 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3353
timestamp 1569543463
transform 1 0 3336 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3354
timestamp 1569543463
transform 1 0 3208 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3355
timestamp 1569543463
transform 1 0 3400 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3356
timestamp 1569543463
transform 1 0 3400 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3357
timestamp 1569543463
transform 1 0 3144 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3358
timestamp 1569543463
transform 1 0 3144 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3359
timestamp 1569543463
transform 1 0 3400 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3360
timestamp 1569543463
transform 1 0 3144 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3361
timestamp 1569543463
transform 1 0 3336 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3362
timestamp 1569543463
transform 1 0 3144 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3363
timestamp 1569543463
transform 1 0 3272 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3364
timestamp 1569543463
transform 1 0 3208 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3365
timestamp 1569543463
transform 1 0 3592 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3366
timestamp 1569543463
transform 1 0 3720 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3367
timestamp 1569543463
transform 1 0 3464 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3368
timestamp 1569543463
transform 1 0 3720 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3369
timestamp 1569543463
transform 1 0 3464 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3370
timestamp 1569543463
transform 1 0 3656 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3371
timestamp 1569543463
transform 1 0 3528 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3372
timestamp 1569543463
transform 1 0 3528 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3373
timestamp 1569543463
transform 1 0 3592 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3374
timestamp 1569543463
transform 1 0 3592 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3375
timestamp 1569543463
transform 1 0 3528 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3376
timestamp 1569543463
transform 1 0 3656 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3377
timestamp 1569543463
transform 1 0 3656 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3378
timestamp 1569543463
transform 1 0 3656 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3379
timestamp 1569543463
transform 1 0 3528 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3380
timestamp 1569543463
transform 1 0 3528 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3381
timestamp 1569543463
transform 1 0 3464 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3382
timestamp 1569543463
transform 1 0 3720 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3383
timestamp 1569543463
transform 1 0 3592 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3384
timestamp 1569543463
transform 1 0 3464 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3385
timestamp 1569543463
transform 1 0 3720 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3386
timestamp 1569543463
transform 1 0 3464 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3387
timestamp 1569543463
transform 1 0 3720 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3388
timestamp 1569543463
transform 1 0 3656 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3389
timestamp 1569543463
transform 1 0 3592 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3390
timestamp 1569543463
transform 1 0 3080 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3391
timestamp 1569543463
transform 1 0 3080 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3392
timestamp 1569543463
transform 1 0 2952 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3393
timestamp 1569543463
transform 1 0 2696 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3394
timestamp 1569543463
transform 1 0 2952 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3395
timestamp 1569543463
transform 1 0 3016 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3396
timestamp 1569543463
transform 1 0 2888 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3397
timestamp 1569543463
transform 1 0 3016 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3398
timestamp 1569543463
transform 1 0 2760 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3399
timestamp 1569543463
transform 1 0 3016 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3400
timestamp 1569543463
transform 1 0 2952 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3401
timestamp 1569543463
transform 1 0 3080 0 1 2696
box -8 -8 8 8
use VIA1$5  VIA1$5_3402
timestamp 1569543463
transform 1 0 2824 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3403
timestamp 1569543463
transform 1 0 3080 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3404
timestamp 1569543463
transform 1 0 2824 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3405
timestamp 1569543463
transform 1 0 3080 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3406
timestamp 1569543463
transform 1 0 2952 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3407
timestamp 1569543463
transform 1 0 2952 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3408
timestamp 1569543463
transform 1 0 2888 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3409
timestamp 1569543463
transform 1 0 2888 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3410
timestamp 1569543463
transform 1 0 2632 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3411
timestamp 1569543463
transform 1 0 2952 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3412
timestamp 1569543463
transform 1 0 2696 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3413
timestamp 1569543463
transform 1 0 2888 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3414
timestamp 1569543463
transform 1 0 3016 0 1 2760
box -8 -8 8 8
use VIA1$5  VIA1$5_3415
timestamp 1569543463
transform 1 0 3016 0 1 2824
box -8 -8 8 8
use VIA1$5  VIA1$5_3416
timestamp 1569543463
transform 1 0 3016 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3417
timestamp 1569543463
transform 1 0 2760 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3418
timestamp 1569543463
transform 1 0 3016 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3419
timestamp 1569543463
transform 1 0 2760 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3420
timestamp 1569543463
transform 1 0 2888 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3421
timestamp 1569543463
transform 1 0 3080 0 1 2888
box -8 -8 8 8
use VIA1$5  VIA1$5_3422
timestamp 1569543463
transform 1 0 2824 0 1 2952
box -8 -8 8 8
use VIA1$5  VIA1$5_3423
timestamp 1569543463
transform 1 0 3080 0 1 3016
box -8 -8 8 8
use VIA1$5  VIA1$5_3424
timestamp 1569543463
transform 1 0 2824 0 1 3080
box -8 -8 8 8
use VIA1$5  VIA1$5_3425
timestamp 1569543463
transform 1 0 3080 0 1 2632
box -8 -8 8 8
use VIA1$5  VIA1$5_3426
timestamp 1569543463
transform 1 0 2888 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3427
timestamp 1569543463
transform 1 0 3016 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3428
timestamp 1569543463
transform 1 0 3080 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3429
timestamp 1569543463
transform 1 0 2888 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3430
timestamp 1569543463
transform 1 0 2824 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3431
timestamp 1569543463
transform 1 0 2888 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3432
timestamp 1569543463
transform 1 0 2888 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3433
timestamp 1569543463
transform 1 0 2888 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3434
timestamp 1569543463
transform 1 0 3016 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3435
timestamp 1569543463
transform 1 0 3080 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3436
timestamp 1569543463
transform 1 0 3080 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3437
timestamp 1569543463
transform 1 0 2952 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3438
timestamp 1569543463
transform 1 0 2952 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3439
timestamp 1569543463
transform 1 0 2952 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3440
timestamp 1569543463
transform 1 0 2952 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3441
timestamp 1569543463
transform 1 0 3016 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3442
timestamp 1569543463
transform 1 0 3016 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3443
timestamp 1569543463
transform 1 0 3080 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3444
timestamp 1569543463
transform 1 0 2824 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3445
timestamp 1569543463
transform 1 0 2824 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3446
timestamp 1569543463
transform 1 0 3016 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3447
timestamp 1569543463
transform 1 0 2824 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3448
timestamp 1569543463
transform 1 0 2824 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3449
timestamp 1569543463
transform 1 0 2952 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3450
timestamp 1569543463
transform 1 0 3080 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3451
timestamp 1569543463
transform 1 0 2696 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3452
timestamp 1569543463
transform 1 0 2568 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3453
timestamp 1569543463
transform 1 0 2760 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3454
timestamp 1569543463
transform 1 0 2632 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3455
timestamp 1569543463
transform 1 0 2696 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3456
timestamp 1569543463
transform 1 0 2696 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3457
timestamp 1569543463
transform 1 0 2696 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3458
timestamp 1569543463
transform 1 0 2696 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3459
timestamp 1569543463
transform 1 0 2632 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3460
timestamp 1569543463
transform 1 0 2632 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3461
timestamp 1569543463
transform 1 0 2568 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3462
timestamp 1569543463
transform 1 0 2760 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3463
timestamp 1569543463
transform 1 0 2760 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3464
timestamp 1569543463
transform 1 0 2760 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3465
timestamp 1569543463
transform 1 0 2632 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3466
timestamp 1569543463
transform 1 0 2760 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3467
timestamp 1569543463
transform 1 0 2568 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3468
timestamp 1569543463
transform 1 0 2568 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3469
timestamp 1569543463
transform 1 0 2568 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3470
timestamp 1569543463
transform 1 0 2632 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3471
timestamp 1569543463
transform 1 0 2568 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3472
timestamp 1569543463
transform 1 0 2632 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3473
timestamp 1569543463
transform 1 0 2632 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3474
timestamp 1569543463
transform 1 0 2632 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3475
timestamp 1569543463
transform 1 0 2760 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3476
timestamp 1569543463
transform 1 0 2760 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3477
timestamp 1569543463
transform 1 0 2696 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3478
timestamp 1569543463
transform 1 0 2696 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3479
timestamp 1569543463
transform 1 0 2760 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3480
timestamp 1569543463
transform 1 0 2760 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3481
timestamp 1569543463
transform 1 0 2760 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3482
timestamp 1569543463
transform 1 0 2632 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3483
timestamp 1569543463
transform 1 0 2568 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3484
timestamp 1569543463
transform 1 0 2632 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3485
timestamp 1569543463
transform 1 0 2568 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3486
timestamp 1569543463
transform 1 0 2568 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3487
timestamp 1569543463
transform 1 0 2568 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3488
timestamp 1569543463
transform 1 0 2696 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3489
timestamp 1569543463
transform 1 0 2696 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3490
timestamp 1569543463
transform 1 0 2696 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3491
timestamp 1569543463
transform 1 0 3080 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3492
timestamp 1569543463
transform 1 0 3016 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3493
timestamp 1569543463
transform 1 0 3080 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3494
timestamp 1569543463
transform 1 0 3016 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3495
timestamp 1569543463
transform 1 0 2824 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3496
timestamp 1569543463
transform 1 0 2824 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3497
timestamp 1569543463
transform 1 0 2888 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3498
timestamp 1569543463
transform 1 0 2888 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3499
timestamp 1569543463
transform 1 0 3080 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3500
timestamp 1569543463
transform 1 0 2952 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3501
timestamp 1569543463
transform 1 0 2952 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3502
timestamp 1569543463
transform 1 0 3080 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3503
timestamp 1569543463
transform 1 0 3016 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3504
timestamp 1569543463
transform 1 0 3080 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3505
timestamp 1569543463
transform 1 0 2824 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3506
timestamp 1569543463
transform 1 0 2824 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3507
timestamp 1569543463
transform 1 0 2824 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3508
timestamp 1569543463
transform 1 0 2888 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3509
timestamp 1569543463
transform 1 0 2888 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3510
timestamp 1569543463
transform 1 0 2888 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3511
timestamp 1569543463
transform 1 0 3016 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3512
timestamp 1569543463
transform 1 0 2952 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3513
timestamp 1569543463
transform 1 0 2952 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3514
timestamp 1569543463
transform 1 0 2952 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3515
timestamp 1569543463
transform 1 0 3016 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3516
timestamp 1569543463
transform 1 0 3656 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3517
timestamp 1569543463
transform 1 0 3720 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3518
timestamp 1569543463
transform 1 0 3720 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3519
timestamp 1569543463
transform 1 0 3720 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3520
timestamp 1569543463
transform 1 0 3720 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3521
timestamp 1569543463
transform 1 0 3720 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3522
timestamp 1569543463
transform 1 0 3464 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3523
timestamp 1569543463
transform 1 0 3464 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3524
timestamp 1569543463
transform 1 0 3464 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3525
timestamp 1569543463
transform 1 0 3464 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3526
timestamp 1569543463
transform 1 0 3464 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3527
timestamp 1569543463
transform 1 0 3528 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3528
timestamp 1569543463
transform 1 0 3528 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3529
timestamp 1569543463
transform 1 0 3528 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3530
timestamp 1569543463
transform 1 0 3528 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3531
timestamp 1569543463
transform 1 0 3528 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3532
timestamp 1569543463
transform 1 0 3592 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3533
timestamp 1569543463
transform 1 0 3592 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3534
timestamp 1569543463
transform 1 0 3592 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3535
timestamp 1569543463
transform 1 0 3592 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3536
timestamp 1569543463
transform 1 0 3592 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3537
timestamp 1569543463
transform 1 0 3656 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3538
timestamp 1569543463
transform 1 0 3656 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3539
timestamp 1569543463
transform 1 0 3656 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3540
timestamp 1569543463
transform 1 0 3656 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3541
timestamp 1569543463
transform 1 0 3208 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3542
timestamp 1569543463
transform 1 0 3272 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3543
timestamp 1569543463
transform 1 0 3336 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3544
timestamp 1569543463
transform 1 0 3400 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3545
timestamp 1569543463
transform 1 0 3336 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3546
timestamp 1569543463
transform 1 0 3336 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3547
timestamp 1569543463
transform 1 0 3336 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3548
timestamp 1569543463
transform 1 0 3336 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3549
timestamp 1569543463
transform 1 0 3144 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3550
timestamp 1569543463
transform 1 0 3400 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3551
timestamp 1569543463
transform 1 0 3400 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3552
timestamp 1569543463
transform 1 0 3400 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3553
timestamp 1569543463
transform 1 0 3400 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3554
timestamp 1569543463
transform 1 0 3208 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3555
timestamp 1569543463
transform 1 0 3208 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3556
timestamp 1569543463
transform 1 0 3208 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3557
timestamp 1569543463
transform 1 0 3208 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3558
timestamp 1569543463
transform 1 0 3144 0 1 3144
box -8 -8 8 8
use VIA1$5  VIA1$5_3559
timestamp 1569543463
transform 1 0 3272 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3560
timestamp 1569543463
transform 1 0 3272 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3561
timestamp 1569543463
transform 1 0 3272 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3562
timestamp 1569543463
transform 1 0 3272 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_3563
timestamp 1569543463
transform 1 0 3144 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_3564
timestamp 1569543463
transform 1 0 3144 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_3565
timestamp 1569543463
transform 1 0 3144 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_3566
timestamp 1569543463
transform 1 0 3336 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3567
timestamp 1569543463
transform 1 0 3336 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3568
timestamp 1569543463
transform 1 0 3400 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3569
timestamp 1569543463
transform 1 0 3400 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3570
timestamp 1569543463
transform 1 0 3272 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3571
timestamp 1569543463
transform 1 0 3272 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3572
timestamp 1569543463
transform 1 0 3336 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3573
timestamp 1569543463
transform 1 0 3336 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3574
timestamp 1569543463
transform 1 0 3336 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3575
timestamp 1569543463
transform 1 0 3272 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3576
timestamp 1569543463
transform 1 0 3272 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3577
timestamp 1569543463
transform 1 0 3400 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3578
timestamp 1569543463
transform 1 0 3400 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3579
timestamp 1569543463
transform 1 0 3400 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3580
timestamp 1569543463
transform 1 0 3272 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3581
timestamp 1569543463
transform 1 0 3144 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3582
timestamp 1569543463
transform 1 0 3144 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3583
timestamp 1569543463
transform 1 0 3144 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3584
timestamp 1569543463
transform 1 0 3208 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3585
timestamp 1569543463
transform 1 0 3208 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3586
timestamp 1569543463
transform 1 0 3208 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3587
timestamp 1569543463
transform 1 0 3144 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3588
timestamp 1569543463
transform 1 0 3144 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3589
timestamp 1569543463
transform 1 0 3208 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3590
timestamp 1569543463
transform 1 0 3208 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3591
timestamp 1569543463
transform 1 0 3464 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3592
timestamp 1569543463
transform 1 0 3464 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3593
timestamp 1569543463
transform 1 0 3528 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3594
timestamp 1569543463
transform 1 0 3528 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3595
timestamp 1569543463
transform 1 0 3592 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3596
timestamp 1569543463
transform 1 0 3592 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3597
timestamp 1569543463
transform 1 0 3720 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3598
timestamp 1569543463
transform 1 0 3464 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3599
timestamp 1569543463
transform 1 0 3464 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3600
timestamp 1569543463
transform 1 0 3464 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3601
timestamp 1569543463
transform 1 0 3528 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3602
timestamp 1569543463
transform 1 0 3528 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3603
timestamp 1569543463
transform 1 0 3528 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3604
timestamp 1569543463
transform 1 0 3592 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3605
timestamp 1569543463
transform 1 0 3592 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3606
timestamp 1569543463
transform 1 0 3592 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3607
timestamp 1569543463
transform 1 0 3720 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3608
timestamp 1569543463
transform 1 0 3720 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3609
timestamp 1569543463
transform 1 0 3656 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3610
timestamp 1569543463
transform 1 0 3656 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3611
timestamp 1569543463
transform 1 0 3720 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_3612
timestamp 1569543463
transform 1 0 3720 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_3613
timestamp 1569543463
transform 1 0 3656 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_3614
timestamp 1569543463
transform 1 0 3656 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_3615
timestamp 1569543463
transform 1 0 3656 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_3616
timestamp 1569543463
transform 1 0 3592 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3617
timestamp 1569543463
transform 1 0 3720 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3618
timestamp 1569543463
transform 1 0 3720 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3619
timestamp 1569543463
transform 1 0 3720 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3620
timestamp 1569543463
transform 1 0 3592 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3621
timestamp 1569543463
transform 1 0 3592 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3622
timestamp 1569543463
transform 1 0 3656 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3623
timestamp 1569543463
transform 1 0 3720 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3624
timestamp 1569543463
transform 1 0 3656 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3625
timestamp 1569543463
transform 1 0 3592 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3626
timestamp 1569543463
transform 1 0 3528 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3627
timestamp 1569543463
transform 1 0 3464 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3628
timestamp 1569543463
transform 1 0 3464 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3629
timestamp 1569543463
transform 1 0 3464 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3630
timestamp 1569543463
transform 1 0 3656 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3631
timestamp 1569543463
transform 1 0 3464 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3632
timestamp 1569543463
transform 1 0 3656 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3633
timestamp 1569543463
transform 1 0 3464 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3634
timestamp 1569543463
transform 1 0 3528 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3635
timestamp 1569543463
transform 1 0 3720 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3636
timestamp 1569543463
transform 1 0 3528 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3637
timestamp 1569543463
transform 1 0 3528 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3638
timestamp 1569543463
transform 1 0 3528 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3639
timestamp 1569543463
transform 1 0 3656 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3640
timestamp 1569543463
transform 1 0 3592 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3641
timestamp 1569543463
transform 1 0 3336 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3642
timestamp 1569543463
transform 1 0 3336 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3643
timestamp 1569543463
transform 1 0 3336 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3644
timestamp 1569543463
transform 1 0 3272 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3645
timestamp 1569543463
transform 1 0 3336 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3646
timestamp 1569543463
transform 1 0 3272 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3647
timestamp 1569543463
transform 1 0 3400 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3648
timestamp 1569543463
transform 1 0 3144 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3649
timestamp 1569543463
transform 1 0 3400 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3650
timestamp 1569543463
transform 1 0 3400 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3651
timestamp 1569543463
transform 1 0 3272 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3652
timestamp 1569543463
transform 1 0 3144 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3653
timestamp 1569543463
transform 1 0 3400 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3654
timestamp 1569543463
transform 1 0 3400 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3655
timestamp 1569543463
transform 1 0 3144 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3656
timestamp 1569543463
transform 1 0 3144 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3657
timestamp 1569543463
transform 1 0 3272 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3658
timestamp 1569543463
transform 1 0 3208 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3659
timestamp 1569543463
transform 1 0 3208 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3660
timestamp 1569543463
transform 1 0 3336 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3661
timestamp 1569543463
transform 1 0 3208 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3662
timestamp 1569543463
transform 1 0 3208 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3663
timestamp 1569543463
transform 1 0 3208 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3664
timestamp 1569543463
transform 1 0 3272 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3665
timestamp 1569543463
transform 1 0 3144 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3666
timestamp 1569543463
transform 1 0 3272 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3667
timestamp 1569543463
transform 1 0 3272 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3668
timestamp 1569543463
transform 1 0 3272 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3669
timestamp 1569543463
transform 1 0 3272 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3670
timestamp 1569543463
transform 1 0 3144 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3671
timestamp 1569543463
transform 1 0 3336 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3672
timestamp 1569543463
transform 1 0 3336 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3673
timestamp 1569543463
transform 1 0 3336 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3674
timestamp 1569543463
transform 1 0 3336 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3675
timestamp 1569543463
transform 1 0 3208 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3676
timestamp 1569543463
transform 1 0 3144 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3677
timestamp 1569543463
transform 1 0 3400 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3678
timestamp 1569543463
transform 1 0 3400 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3679
timestamp 1569543463
transform 1 0 3400 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3680
timestamp 1569543463
transform 1 0 3400 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3681
timestamp 1569543463
transform 1 0 3208 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3682
timestamp 1569543463
transform 1 0 3208 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3683
timestamp 1569543463
transform 1 0 3144 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3684
timestamp 1569543463
transform 1 0 3144 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3685
timestamp 1569543463
transform 1 0 3208 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3686
timestamp 1569543463
transform 1 0 3592 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3687
timestamp 1569543463
transform 1 0 3656 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3688
timestamp 1569543463
transform 1 0 3656 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3689
timestamp 1569543463
transform 1 0 3656 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3690
timestamp 1569543463
transform 1 0 3464 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3691
timestamp 1569543463
transform 1 0 3656 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3692
timestamp 1569543463
transform 1 0 3464 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3693
timestamp 1569543463
transform 1 0 3464 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3694
timestamp 1569543463
transform 1 0 3464 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3695
timestamp 1569543463
transform 1 0 3720 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3696
timestamp 1569543463
transform 1 0 3528 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3697
timestamp 1569543463
transform 1 0 3720 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3698
timestamp 1569543463
transform 1 0 3528 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3699
timestamp 1569543463
transform 1 0 3528 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3700
timestamp 1569543463
transform 1 0 3720 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3701
timestamp 1569543463
transform 1 0 3528 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3702
timestamp 1569543463
transform 1 0 3720 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3703
timestamp 1569543463
transform 1 0 3592 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3704
timestamp 1569543463
transform 1 0 3592 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3705
timestamp 1569543463
transform 1 0 3592 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3706
timestamp 1569543463
transform 1 0 2824 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3707
timestamp 1569543463
transform 1 0 3080 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3708
timestamp 1569543463
transform 1 0 2824 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3709
timestamp 1569543463
transform 1 0 2824 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3710
timestamp 1569543463
transform 1 0 2824 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3711
timestamp 1569543463
transform 1 0 2824 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3712
timestamp 1569543463
transform 1 0 2888 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3713
timestamp 1569543463
transform 1 0 2888 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3714
timestamp 1569543463
transform 1 0 2888 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3715
timestamp 1569543463
transform 1 0 2888 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3716
timestamp 1569543463
transform 1 0 2952 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3717
timestamp 1569543463
transform 1 0 2952 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3718
timestamp 1569543463
transform 1 0 2952 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3719
timestamp 1569543463
transform 1 0 2952 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3720
timestamp 1569543463
transform 1 0 2888 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3721
timestamp 1569543463
transform 1 0 3016 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3722
timestamp 1569543463
transform 1 0 3016 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3723
timestamp 1569543463
transform 1 0 3016 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3724
timestamp 1569543463
transform 1 0 3016 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3725
timestamp 1569543463
transform 1 0 3016 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3726
timestamp 1569543463
transform 1 0 3080 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3727
timestamp 1569543463
transform 1 0 3080 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3728
timestamp 1569543463
transform 1 0 2952 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3729
timestamp 1569543463
transform 1 0 3080 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3730
timestamp 1569543463
transform 1 0 3080 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3731
timestamp 1569543463
transform 1 0 2696 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3732
timestamp 1569543463
transform 1 0 2696 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3733
timestamp 1569543463
transform 1 0 2696 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3734
timestamp 1569543463
transform 1 0 2696 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3735
timestamp 1569543463
transform 1 0 2760 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3736
timestamp 1569543463
transform 1 0 2760 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3737
timestamp 1569543463
transform 1 0 2760 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3738
timestamp 1569543463
transform 1 0 2760 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3739
timestamp 1569543463
transform 1 0 2696 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3740
timestamp 1569543463
transform 1 0 2568 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3741
timestamp 1569543463
transform 1 0 2568 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3742
timestamp 1569543463
transform 1 0 2760 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3743
timestamp 1569543463
transform 1 0 2568 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3744
timestamp 1569543463
transform 1 0 2568 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3745
timestamp 1569543463
transform 1 0 2632 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3746
timestamp 1569543463
transform 1 0 2568 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3747
timestamp 1569543463
transform 1 0 2632 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3748
timestamp 1569543463
transform 1 0 2632 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3749
timestamp 1569543463
transform 1 0 2632 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3750
timestamp 1569543463
transform 1 0 2632 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3751
timestamp 1569543463
transform 1 0 2696 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3752
timestamp 1569543463
transform 1 0 2696 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3753
timestamp 1569543463
transform 1 0 2696 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3754
timestamp 1569543463
transform 1 0 2696 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3755
timestamp 1569543463
transform 1 0 2760 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3756
timestamp 1569543463
transform 1 0 2760 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3757
timestamp 1569543463
transform 1 0 2760 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3758
timestamp 1569543463
transform 1 0 2760 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3759
timestamp 1569543463
transform 1 0 2632 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3760
timestamp 1569543463
transform 1 0 2632 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3761
timestamp 1569543463
transform 1 0 2632 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3762
timestamp 1569543463
transform 1 0 2632 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3763
timestamp 1569543463
transform 1 0 2568 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3764
timestamp 1569543463
transform 1 0 2568 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3765
timestamp 1569543463
transform 1 0 2568 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3766
timestamp 1569543463
transform 1 0 2568 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3767
timestamp 1569543463
transform 1 0 2824 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3768
timestamp 1569543463
transform 1 0 2824 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3769
timestamp 1569543463
transform 1 0 2824 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3770
timestamp 1569543463
transform 1 0 2824 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3771
timestamp 1569543463
transform 1 0 2888 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3772
timestamp 1569543463
transform 1 0 2888 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3773
timestamp 1569543463
transform 1 0 2888 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3774
timestamp 1569543463
transform 1 0 2888 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3775
timestamp 1569543463
transform 1 0 2952 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3776
timestamp 1569543463
transform 1 0 2952 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3777
timestamp 1569543463
transform 1 0 2952 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3778
timestamp 1569543463
transform 1 0 2952 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3779
timestamp 1569543463
transform 1 0 3016 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3780
timestamp 1569543463
transform 1 0 3016 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3781
timestamp 1569543463
transform 1 0 3016 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3782
timestamp 1569543463
transform 1 0 3016 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3783
timestamp 1569543463
transform 1 0 3080 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3784
timestamp 1569543463
transform 1 0 3080 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3785
timestamp 1569543463
transform 1 0 3080 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_3786
timestamp 1569543463
transform 1 0 3080 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3787
timestamp 1569543463
transform 1 0 3016 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3788
timestamp 1569543463
transform 1 0 2888 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3789
timestamp 1569543463
transform 1 0 3080 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3790
timestamp 1569543463
transform 1 0 2952 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3791
timestamp 1569543463
transform 1 0 2824 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3792
timestamp 1569543463
transform 1 0 2824 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3793
timestamp 1569543463
transform 1 0 3080 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3794
timestamp 1569543463
transform 1 0 3080 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3795
timestamp 1569543463
transform 1 0 3016 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3796
timestamp 1569543463
transform 1 0 2888 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3797
timestamp 1569543463
transform 1 0 2824 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3798
timestamp 1569543463
transform 1 0 2888 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3799
timestamp 1569543463
transform 1 0 3016 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3800
timestamp 1569543463
transform 1 0 2952 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3801
timestamp 1569543463
transform 1 0 2952 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3802
timestamp 1569543463
transform 1 0 2888 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3803
timestamp 1569543463
transform 1 0 2824 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3804
timestamp 1569543463
transform 1 0 2952 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3805
timestamp 1569543463
transform 1 0 3016 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3806
timestamp 1569543463
transform 1 0 3080 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3807
timestamp 1569543463
transform 1 0 2760 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3808
timestamp 1569543463
transform 1 0 2696 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3809
timestamp 1569543463
transform 1 0 2632 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3810
timestamp 1569543463
transform 1 0 2568 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3811
timestamp 1569543463
transform 1 0 2632 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3812
timestamp 1569543463
transform 1 0 2760 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3813
timestamp 1569543463
transform 1 0 2632 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3814
timestamp 1569543463
transform 1 0 2696 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3815
timestamp 1569543463
transform 1 0 2760 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3816
timestamp 1569543463
transform 1 0 2568 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3817
timestamp 1569543463
transform 1 0 2568 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3818
timestamp 1569543463
transform 1 0 2696 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3819
timestamp 1569543463
transform 1 0 2696 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3820
timestamp 1569543463
transform 1 0 2760 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3821
timestamp 1569543463
transform 1 0 2568 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3822
timestamp 1569543463
transform 1 0 2632 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3823
timestamp 1569543463
transform 1 0 2696 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3824
timestamp 1569543463
transform 1 0 2632 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3825
timestamp 1569543463
transform 1 0 2760 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3826
timestamp 1569543463
transform 1 0 2760 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3827
timestamp 1569543463
transform 1 0 2760 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3828
timestamp 1569543463
transform 1 0 2696 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3829
timestamp 1569543463
transform 1 0 2696 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3830
timestamp 1569543463
transform 1 0 2760 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3831
timestamp 1569543463
transform 1 0 2696 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3832
timestamp 1569543463
transform 1 0 2568 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3833
timestamp 1569543463
transform 1 0 2568 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3834
timestamp 1569543463
transform 1 0 2568 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3835
timestamp 1569543463
transform 1 0 2632 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3836
timestamp 1569543463
transform 1 0 2568 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3837
timestamp 1569543463
transform 1 0 2632 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3838
timestamp 1569543463
transform 1 0 2632 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3839
timestamp 1569543463
transform 1 0 2824 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3840
timestamp 1569543463
transform 1 0 2952 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3841
timestamp 1569543463
transform 1 0 2952 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3842
timestamp 1569543463
transform 1 0 2824 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3843
timestamp 1569543463
transform 1 0 2952 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3844
timestamp 1569543463
transform 1 0 2952 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3845
timestamp 1569543463
transform 1 0 2824 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3846
timestamp 1569543463
transform 1 0 3016 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3847
timestamp 1569543463
transform 1 0 3016 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3848
timestamp 1569543463
transform 1 0 2824 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3849
timestamp 1569543463
transform 1 0 3016 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3850
timestamp 1569543463
transform 1 0 3016 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3851
timestamp 1569543463
transform 1 0 3080 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3852
timestamp 1569543463
transform 1 0 3080 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3853
timestamp 1569543463
transform 1 0 3080 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3854
timestamp 1569543463
transform 1 0 3080 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3855
timestamp 1569543463
transform 1 0 2888 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3856
timestamp 1569543463
transform 1 0 2888 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3857
timestamp 1569543463
transform 1 0 2888 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3858
timestamp 1569543463
transform 1 0 2888 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3859
timestamp 1569543463
transform 1 0 3464 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3860
timestamp 1569543463
transform 1 0 3656 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3861
timestamp 1569543463
transform 1 0 3464 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3862
timestamp 1569543463
transform 1 0 3464 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3863
timestamp 1569543463
transform 1 0 3528 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3864
timestamp 1569543463
transform 1 0 3592 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3865
timestamp 1569543463
transform 1 0 3720 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3866
timestamp 1569543463
transform 1 0 3592 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3867
timestamp 1569543463
transform 1 0 3592 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3868
timestamp 1569543463
transform 1 0 3720 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3869
timestamp 1569543463
transform 1 0 3528 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3870
timestamp 1569543463
transform 1 0 3464 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3871
timestamp 1569543463
transform 1 0 3592 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3872
timestamp 1569543463
transform 1 0 3528 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3873
timestamp 1569543463
transform 1 0 3656 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3874
timestamp 1569543463
transform 1 0 3656 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3875
timestamp 1569543463
transform 1 0 3720 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3876
timestamp 1569543463
transform 1 0 3656 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3877
timestamp 1569543463
transform 1 0 3528 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3878
timestamp 1569543463
transform 1 0 3720 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3879
timestamp 1569543463
transform 1 0 3336 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3880
timestamp 1569543463
transform 1 0 3208 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3881
timestamp 1569543463
transform 1 0 3400 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3882
timestamp 1569543463
transform 1 0 3336 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3883
timestamp 1569543463
transform 1 0 3208 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3884
timestamp 1569543463
transform 1 0 3336 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3885
timestamp 1569543463
transform 1 0 3208 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3886
timestamp 1569543463
transform 1 0 3272 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3887
timestamp 1569543463
transform 1 0 3400 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3888
timestamp 1569543463
transform 1 0 3144 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3889
timestamp 1569543463
transform 1 0 3272 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3890
timestamp 1569543463
transform 1 0 3272 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3891
timestamp 1569543463
transform 1 0 3272 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3892
timestamp 1569543463
transform 1 0 3144 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3893
timestamp 1569543463
transform 1 0 3400 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3894
timestamp 1569543463
transform 1 0 3400 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3895
timestamp 1569543463
transform 1 0 3144 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_3896
timestamp 1569543463
transform 1 0 3336 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3897
timestamp 1569543463
transform 1 0 3208 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_3898
timestamp 1569543463
transform 1 0 3144 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3899
timestamp 1569543463
transform 1 0 3272 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3900
timestamp 1569543463
transform 1 0 3272 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3901
timestamp 1569543463
transform 1 0 3272 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3902
timestamp 1569543463
transform 1 0 3336 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3903
timestamp 1569543463
transform 1 0 3336 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3904
timestamp 1569543463
transform 1 0 3336 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3905
timestamp 1569543463
transform 1 0 3336 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3906
timestamp 1569543463
transform 1 0 3400 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3907
timestamp 1569543463
transform 1 0 3400 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3908
timestamp 1569543463
transform 1 0 3400 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3909
timestamp 1569543463
transform 1 0 3144 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3910
timestamp 1569543463
transform 1 0 3144 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3911
timestamp 1569543463
transform 1 0 3400 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3912
timestamp 1569543463
transform 1 0 3144 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3913
timestamp 1569543463
transform 1 0 3144 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3914
timestamp 1569543463
transform 1 0 3208 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3915
timestamp 1569543463
transform 1 0 3208 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3916
timestamp 1569543463
transform 1 0 3208 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3917
timestamp 1569543463
transform 1 0 3208 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3918
timestamp 1569543463
transform 1 0 3272 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3919
timestamp 1569543463
transform 1 0 3464 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3920
timestamp 1569543463
transform 1 0 3592 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3921
timestamp 1569543463
transform 1 0 3592 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3922
timestamp 1569543463
transform 1 0 3592 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3923
timestamp 1569543463
transform 1 0 3592 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3924
timestamp 1569543463
transform 1 0 3656 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3925
timestamp 1569543463
transform 1 0 3656 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3926
timestamp 1569543463
transform 1 0 3656 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3927
timestamp 1569543463
transform 1 0 3656 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3928
timestamp 1569543463
transform 1 0 3720 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3929
timestamp 1569543463
transform 1 0 3720 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3930
timestamp 1569543463
transform 1 0 3720 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3931
timestamp 1569543463
transform 1 0 3464 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3932
timestamp 1569543463
transform 1 0 3720 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3933
timestamp 1569543463
transform 1 0 3464 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3934
timestamp 1569543463
transform 1 0 3528 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3935
timestamp 1569543463
transform 1 0 3528 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3936
timestamp 1569543463
transform 1 0 3528 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3937
timestamp 1569543463
transform 1 0 3528 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3938
timestamp 1569543463
transform 1 0 3464 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3939
timestamp 1569543463
transform 1 0 2696 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3940
timestamp 1569543463
transform 1 0 3336 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3941
timestamp 1569543463
transform 1 0 2760 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3942
timestamp 1569543463
transform 1 0 3400 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3943
timestamp 1569543463
transform 1 0 2824 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3944
timestamp 1569543463
transform 1 0 3464 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3945
timestamp 1569543463
transform 1 0 2888 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3946
timestamp 1569543463
transform 1 0 3528 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3947
timestamp 1569543463
transform 1 0 2952 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3948
timestamp 1569543463
transform 1 0 3592 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3949
timestamp 1569543463
transform 1 0 3016 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3950
timestamp 1569543463
transform 1 0 3656 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3951
timestamp 1569543463
transform 1 0 3080 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3952
timestamp 1569543463
transform 1 0 3720 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3953
timestamp 1569543463
transform 1 0 3144 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3954
timestamp 1569543463
transform 1 0 2568 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3955
timestamp 1569543463
transform 1 0 3208 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3956
timestamp 1569543463
transform 1 0 2632 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3957
timestamp 1569543463
transform 1 0 3272 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_3958
timestamp 1569543463
transform 1 0 4616 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3959
timestamp 1569543463
transform 1 0 4680 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3960
timestamp 1569543463
transform 1 0 4744 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3961
timestamp 1569543463
transform 1 0 4808 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3962
timestamp 1569543463
transform 1 0 4872 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3963
timestamp 1569543463
transform 1 0 4488 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3964
timestamp 1569543463
transform 1 0 4552 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_3965
timestamp 1569543463
transform 1 0 3976 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3966
timestamp 1569543463
transform 1 0 3976 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3967
timestamp 1569543463
transform 1 0 3976 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3968
timestamp 1569543463
transform 1 0 3976 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3969
timestamp 1569543463
transform 1 0 4040 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3970
timestamp 1569543463
transform 1 0 4040 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3971
timestamp 1569543463
transform 1 0 4040 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3972
timestamp 1569543463
transform 1 0 4104 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3973
timestamp 1569543463
transform 1 0 4104 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3974
timestamp 1569543463
transform 1 0 4168 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3975
timestamp 1569543463
transform 1 0 3848 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3976
timestamp 1569543463
transform 1 0 3848 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3977
timestamp 1569543463
transform 1 0 3912 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3978
timestamp 1569543463
transform 1 0 3912 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3979
timestamp 1569543463
transform 1 0 3912 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3980
timestamp 1569543463
transform 1 0 3912 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3981
timestamp 1569543463
transform 1 0 3784 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3982
timestamp 1569543463
transform 1 0 3784 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3983
timestamp 1569543463
transform 1 0 3784 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_3984
timestamp 1569543463
transform 1 0 3848 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3985
timestamp 1569543463
transform 1 0 3848 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_3986
timestamp 1569543463
transform 1 0 3912 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_3987
timestamp 1569543463
transform 1 0 3784 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3988
timestamp 1569543463
transform 1 0 3784 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3989
timestamp 1569543463
transform 1 0 3784 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_3990
timestamp 1569543463
transform 1 0 3784 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_3991
timestamp 1569543463
transform 1 0 3848 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_3992
timestamp 1569543463
transform 1 0 3848 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_3993
timestamp 1569543463
transform 1 0 4296 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_3994
timestamp 1569543463
transform 1 0 4296 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_3995
timestamp 1569543463
transform 1 0 4296 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_3996
timestamp 1569543463
transform 1 0 4296 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_3997
timestamp 1569543463
transform 1 0 4296 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_3998
timestamp 1569543463
transform 1 0 4296 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_3999
timestamp 1569543463
transform 1 0 4296 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4000
timestamp 1569543463
transform 1 0 4616 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4001
timestamp 1569543463
transform 1 0 4680 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4002
timestamp 1569543463
transform 1 0 4744 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4003
timestamp 1569543463
transform 1 0 4808 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4004
timestamp 1569543463
transform 1 0 4872 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4005
timestamp 1569543463
transform 1 0 4936 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4006
timestamp 1569543463
transform 1 0 4936 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4007
timestamp 1569543463
transform 1 0 4936 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4008
timestamp 1569543463
transform 1 0 4936 0 1 4936
box -8 -8 8 8
use VIA1$5  VIA1$5_4009
timestamp 1569543463
transform 1 0 4424 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4010
timestamp 1569543463
transform 1 0 4488 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4011
timestamp 1569543463
transform 1 0 4424 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_4012
timestamp 1569543463
transform 1 0 4424 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_4013
timestamp 1569543463
transform 1 0 4424 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4014
timestamp 1569543463
transform 1 0 4424 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4015
timestamp 1569543463
transform 1 0 4424 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4016
timestamp 1569543463
transform 1 0 4488 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4017
timestamp 1569543463
transform 1 0 4616 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4018
timestamp 1569543463
transform 1 0 4552 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4019
timestamp 1569543463
transform 1 0 4488 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_4020
timestamp 1569543463
transform 1 0 4424 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4021
timestamp 1569543463
transform 1 0 4488 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4022
timestamp 1569543463
transform 1 0 4552 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4023
timestamp 1569543463
transform 1 0 4744 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4024
timestamp 1569543463
transform 1 0 4744 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4025
timestamp 1569543463
transform 1 0 4744 0 1 4936
box -8 -8 8 8
use VIA1$5  VIA1$5_4026
timestamp 1569543463
transform 1 0 4808 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4027
timestamp 1569543463
transform 1 0 4808 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4028
timestamp 1569543463
transform 1 0 4808 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4029
timestamp 1569543463
transform 1 0 4808 0 1 4936
box -8 -8 8 8
use VIA1$5  VIA1$5_4030
timestamp 1569543463
transform 1 0 4424 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4031
timestamp 1569543463
transform 1 0 4552 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4032
timestamp 1569543463
transform 1 0 4872 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4033
timestamp 1569543463
transform 1 0 4872 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4034
timestamp 1569543463
transform 1 0 4872 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4035
timestamp 1569543463
transform 1 0 4872 0 1 4936
box -8 -8 8 8
use VIA1$5  VIA1$5_4036
timestamp 1569543463
transform 1 0 4616 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4037
timestamp 1569543463
transform 1 0 4680 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4038
timestamp 1569543463
transform 1 0 4744 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4039
timestamp 1569543463
transform 1 0 4808 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4040
timestamp 1569543463
transform 1 0 4872 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4041
timestamp 1569543463
transform 1 0 4360 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4042
timestamp 1569543463
transform 1 0 4360 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_4043
timestamp 1569543463
transform 1 0 4360 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_4044
timestamp 1569543463
transform 1 0 4360 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4045
timestamp 1569543463
transform 1 0 4360 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4046
timestamp 1569543463
transform 1 0 4360 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4047
timestamp 1569543463
transform 1 0 4360 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4048
timestamp 1569543463
transform 1 0 4360 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4049
timestamp 1569543463
transform 1 0 4424 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4050
timestamp 1569543463
transform 1 0 4488 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4051
timestamp 1569543463
transform 1 0 4552 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4052
timestamp 1569543463
transform 1 0 2504 0 1 4616
box -8 -8 8 8
use VIA1$5  VIA1$5_4053
timestamp 1569543463
transform 1 0 2504 0 1 4680
box -8 -8 8 8
use VIA1$5  VIA1$5_4054
timestamp 1569543463
transform 1 0 2504 0 1 4744
box -8 -8 8 8
use VIA1$5  VIA1$5_4055
timestamp 1569543463
transform 1 0 2504 0 1 4808
box -8 -8 8 8
use VIA1$5  VIA1$5_4056
timestamp 1569543463
transform 1 0 2504 0 1 4872
box -8 -8 8 8
use VIA1$5  VIA1$5_4057
timestamp 1569543463
transform 1 0 2504 0 1 136
box -8 -8 8 8
use VIA1$5  VIA1$5_4058
timestamp 1569543463
transform 1 0 2504 0 1 200
box -8 -8 8 8
use VIA1$5  VIA1$5_4059
timestamp 1569543463
transform 1 0 2504 0 1 264
box -8 -8 8 8
use VIA1$5  VIA1$5_4060
timestamp 1569543463
transform 1 0 2504 0 1 328
box -8 -8 8 8
use VIA1$5  VIA1$5_4061
timestamp 1569543463
transform 1 0 2504 0 1 392
box -8 -8 8 8
use VIA1$5  VIA1$5_4062
timestamp 1569543463
transform 1 0 2504 0 1 456
box -8 -8 8 8
use VIA1$5  VIA1$5_4063
timestamp 1569543463
transform 1 0 2504 0 1 520
box -8 -8 8 8
use VIA1$5  VIA1$5_4064
timestamp 1569543463
transform 1 0 2504 0 1 584
box -8 -8 8 8
use VIA1$5  VIA1$5_4065
timestamp 1569543463
transform 1 0 2504 0 1 648
box -8 -8 8 8
use VIA1$5  VIA1$5_4066
timestamp 1569543463
transform 1 0 2504 0 1 712
box -8 -8 8 8
use VIA1$5  VIA1$5_4067
timestamp 1569543463
transform 1 0 2504 0 1 776
box -8 -8 8 8
use VIA1$5  VIA1$5_4068
timestamp 1569543463
transform 1 0 2504 0 1 840
box -8 -8 8 8
use VIA1$5  VIA1$5_4069
timestamp 1569543463
transform 1 0 2504 0 1 904
box -8 -8 8 8
use VIA1$5  VIA1$5_4070
timestamp 1569543463
transform 1 0 2504 0 1 968
box -8 -8 8 8
use VIA1$5  VIA1$5_4071
timestamp 1569543463
transform 1 0 2504 0 1 1032
box -8 -8 8 8
use VIA1$5  VIA1$5_4072
timestamp 1569543463
transform 1 0 2504 0 1 1096
box -8 -8 8 8
use VIA1$5  VIA1$5_4073
timestamp 1569543463
transform 1 0 2504 0 1 1160
box -8 -8 8 8
use VIA1$5  VIA1$5_4074
timestamp 1569543463
transform 1 0 2504 0 1 1224
box -8 -8 8 8
use VIA1$5  VIA1$5_4075
timestamp 1569543463
transform 1 0 2504 0 1 1288
box -8 -8 8 8
use VIA1$5  VIA1$5_4076
timestamp 1569543463
transform 1 0 2504 0 1 1352
box -8 -8 8 8
use VIA1$5  VIA1$5_4077
timestamp 1569543463
transform 1 0 2504 0 1 1416
box -8 -8 8 8
use VIA1$5  VIA1$5_4078
timestamp 1569543463
transform 1 0 2504 0 1 1480
box -8 -8 8 8
use VIA1$5  VIA1$5_4079
timestamp 1569543463
transform 1 0 2504 0 1 1544
box -8 -8 8 8
use VIA1$5  VIA1$5_4080
timestamp 1569543463
transform 1 0 2504 0 1 1608
box -8 -8 8 8
use VIA1$5  VIA1$5_4081
timestamp 1569543463
transform 1 0 2504 0 1 1672
box -8 -8 8 8
use VIA1$5  VIA1$5_4082
timestamp 1569543463
transform 1 0 2504 0 1 1736
box -8 -8 8 8
use VIA1$5  VIA1$5_4083
timestamp 1569543463
transform 1 0 2504 0 1 1800
box -8 -8 8 8
use VIA1$5  VIA1$5_4084
timestamp 1569543463
transform 1 0 2504 0 1 1864
box -8 -8 8 8
use VIA1$5  VIA1$5_4085
timestamp 1569543463
transform 1 0 2504 0 1 1928
box -8 -8 8 8
use VIA1$5  VIA1$5_4086
timestamp 1569543463
transform 1 0 392 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4087
timestamp 1569543463
transform 1 0 1160 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4088
timestamp 1569543463
transform 1 0 1928 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4089
timestamp 1569543463
transform 1 0 3464 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4090
timestamp 1569543463
transform 1 0 4232 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4091
timestamp 1569543463
transform 1 0 456 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4092
timestamp 1569543463
transform 1 0 1224 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4093
timestamp 1569543463
transform 1 0 3528 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4094
timestamp 1569543463
transform 1 0 4296 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4095
timestamp 1569543463
transform 1 0 520 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4096
timestamp 1569543463
transform 1 0 1288 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4097
timestamp 1569543463
transform 1 0 3592 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4098
timestamp 1569543463
transform 1 0 4360 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4099
timestamp 1569543463
transform 1 0 584 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4100
timestamp 1569543463
transform 1 0 1352 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4101
timestamp 1569543463
transform 1 0 3656 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4102
timestamp 1569543463
transform 1 0 4424 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4103
timestamp 1569543463
transform 1 0 648 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4104
timestamp 1569543463
transform 1 0 1416 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4105
timestamp 1569543463
transform 1 0 3720 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4106
timestamp 1569543463
transform 1 0 4488 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4107
timestamp 1569543463
transform 1 0 712 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4108
timestamp 1569543463
transform 1 0 1480 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4109
timestamp 1569543463
transform 1 0 3784 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4110
timestamp 1569543463
transform 1 0 4552 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4111
timestamp 1569543463
transform 1 0 2504 0 1 3208
box -8 -8 8 8
use VIA1$5  VIA1$5_4112
timestamp 1569543463
transform 1 0 2504 0 1 3272
box -8 -8 8 8
use VIA1$5  VIA1$5_4113
timestamp 1569543463
transform 1 0 2504 0 1 3336
box -8 -8 8 8
use VIA1$5  VIA1$5_4114
timestamp 1569543463
transform 1 0 2504 0 1 3400
box -8 -8 8 8
use VIA1$5  VIA1$5_4115
timestamp 1569543463
transform 1 0 2504 0 1 3464
box -8 -8 8 8
use VIA1$5  VIA1$5_4116
timestamp 1569543463
transform 1 0 2504 0 1 3528
box -8 -8 8 8
use VIA1$5  VIA1$5_4117
timestamp 1569543463
transform 1 0 2504 0 1 3592
box -8 -8 8 8
use VIA1$5  VIA1$5_4118
timestamp 1569543463
transform 1 0 2504 0 1 3656
box -8 -8 8 8
use VIA1$5  VIA1$5_4119
timestamp 1569543463
transform 1 0 2504 0 1 3720
box -8 -8 8 8
use VIA1$5  VIA1$5_4120
timestamp 1569543463
transform 1 0 2504 0 1 3784
box -8 -8 8 8
use VIA1$5  VIA1$5_4121
timestamp 1569543463
transform 1 0 2504 0 1 3848
box -8 -8 8 8
use VIA1$5  VIA1$5_4122
timestamp 1569543463
transform 1 0 2504 0 1 3912
box -8 -8 8 8
use VIA1$5  VIA1$5_4123
timestamp 1569543463
transform 1 0 2504 0 1 3976
box -8 -8 8 8
use VIA1$5  VIA1$5_4124
timestamp 1569543463
transform 1 0 2504 0 1 4040
box -8 -8 8 8
use VIA1$5  VIA1$5_4125
timestamp 1569543463
transform 1 0 2504 0 1 4104
box -8 -8 8 8
use VIA1$5  VIA1$5_4126
timestamp 1569543463
transform 1 0 2504 0 1 4168
box -8 -8 8 8
use VIA1$5  VIA1$5_4127
timestamp 1569543463
transform 1 0 2504 0 1 4232
box -8 -8 8 8
use VIA1$5  VIA1$5_4128
timestamp 1569543463
transform 1 0 2504 0 1 4296
box -8 -8 8 8
use VIA1$5  VIA1$5_4129
timestamp 1569543463
transform 1 0 2504 0 1 4360
box -8 -8 8 8
use VIA1$5  VIA1$5_4130
timestamp 1569543463
transform 1 0 2504 0 1 4424
box -8 -8 8 8
use VIA1$5  VIA1$5_4131
timestamp 1569543463
transform 1 0 2504 0 1 4488
box -8 -8 8 8
use VIA1$5  VIA1$5_4132
timestamp 1569543463
transform 1 0 2504 0 1 4552
box -8 -8 8 8
use VIA1$5  VIA1$5_4133
timestamp 1569543463
transform 1 0 2504 0 1 72
box -8 -8 8 8
use VIA1$5  VIA1$5_4134
timestamp 1569543463
transform 1 0 776 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4135
timestamp 1569543463
transform 1 0 1544 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4136
timestamp 1569543463
transform 1 0 3848 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4137
timestamp 1569543463
transform 1 0 4616 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4138
timestamp 1569543463
transform 1 0 72 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4139
timestamp 1569543463
transform 1 0 840 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4140
timestamp 1569543463
transform 1 0 1608 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4141
timestamp 1569543463
transform 1 0 3912 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4142
timestamp 1569543463
transform 1 0 4680 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4143
timestamp 1569543463
transform 1 0 136 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4144
timestamp 1569543463
transform 1 0 904 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4145
timestamp 1569543463
transform 1 0 1672 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4146
timestamp 1569543463
transform 1 0 3208 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4147
timestamp 1569543463
transform 1 0 3976 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4148
timestamp 1569543463
transform 1 0 4744 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4149
timestamp 1569543463
transform 1 0 200 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4150
timestamp 1569543463
transform 1 0 968 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4151
timestamp 1569543463
transform 1 0 1736 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4152
timestamp 1569543463
transform 1 0 3272 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4153
timestamp 1569543463
transform 1 0 4040 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4154
timestamp 1569543463
transform 1 0 4808 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4155
timestamp 1569543463
transform 1 0 264 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4156
timestamp 1569543463
transform 1 0 1032 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4157
timestamp 1569543463
transform 1 0 1800 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4158
timestamp 1569543463
transform 1 0 3336 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4159
timestamp 1569543463
transform 1 0 4104 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4160
timestamp 1569543463
transform 1 0 4872 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4161
timestamp 1569543463
transform 1 0 328 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4162
timestamp 1569543463
transform 1 0 1096 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4163
timestamp 1569543463
transform 1 0 1864 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4164
timestamp 1569543463
transform 1 0 3400 0 1 2504
box -8 -8 8 8
use VIA1$5  VIA1$5_4165
timestamp 1569543463
transform 1 0 4168 0 1 2504
box -8 -8 8 8
use VIA2$5  VIA2$5_0
timestamp 1569543463
transform 1 0 4840 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1
timestamp 1569543463
transform 1 0 4776 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_2
timestamp 1569543463
transform 1 0 4712 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_3
timestamp 1569543463
transform 1 0 4712 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_4
timestamp 1569543463
transform 1 0 4712 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_5
timestamp 1569543463
transform 1 0 4776 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_6
timestamp 1569543463
transform 1 0 4904 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_7
timestamp 1569543463
transform 1 0 4776 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_8
timestamp 1569543463
transform 1 0 4904 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_9
timestamp 1569543463
transform 1 0 4712 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_10
timestamp 1569543463
transform 1 0 4904 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_11
timestamp 1569543463
transform 1 0 4840 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_12
timestamp 1569543463
transform 1 0 4712 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_13
timestamp 1569543463
transform 1 0 4776 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_14
timestamp 1569543463
transform 1 0 4904 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_15
timestamp 1569543463
transform 1 0 4840 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_16
timestamp 1569543463
transform 1 0 4904 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_17
timestamp 1569543463
transform 1 0 4776 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_18
timestamp 1569543463
transform 1 0 4840 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_19
timestamp 1569543463
transform 1 0 4840 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_20
timestamp 1569543463
transform 1 0 4584 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_21
timestamp 1569543463
transform 1 0 4520 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_22
timestamp 1569543463
transform 1 0 4584 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_23
timestamp 1569543463
transform 1 0 4456 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_24
timestamp 1569543463
transform 1 0 4648 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_25
timestamp 1569543463
transform 1 0 4648 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_26
timestamp 1569543463
transform 1 0 4456 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_27
timestamp 1569543463
transform 1 0 4456 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_28
timestamp 1569543463
transform 1 0 4584 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_29
timestamp 1569543463
transform 1 0 4392 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_30
timestamp 1569543463
transform 1 0 4520 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_31
timestamp 1569543463
transform 1 0 4648 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_32
timestamp 1569543463
transform 1 0 4584 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_33
timestamp 1569543463
transform 1 0 4520 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_34
timestamp 1569543463
transform 1 0 4520 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_35
timestamp 1569543463
transform 1 0 4584 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_36
timestamp 1569543463
transform 1 0 4392 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_37
timestamp 1569543463
transform 1 0 4456 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_38
timestamp 1569543463
transform 1 0 4392 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_39
timestamp 1569543463
transform 1 0 4392 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_40
timestamp 1569543463
transform 1 0 4648 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_41
timestamp 1569543463
transform 1 0 4520 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_42
timestamp 1569543463
transform 1 0 4648 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_43
timestamp 1569543463
transform 1 0 4456 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_44
timestamp 1569543463
transform 1 0 4392 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_45
timestamp 1569543463
transform 1 0 4584 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_46
timestamp 1569543463
transform 1 0 4456 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_47
timestamp 1569543463
transform 1 0 4520 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_48
timestamp 1569543463
transform 1 0 4456 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_49
timestamp 1569543463
transform 1 0 4584 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_50
timestamp 1569543463
transform 1 0 4392 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_51
timestamp 1569543463
transform 1 0 4584 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_52
timestamp 1569543463
transform 1 0 4648 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_53
timestamp 1569543463
transform 1 0 4520 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_54
timestamp 1569543463
transform 1 0 4456 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_55
timestamp 1569543463
transform 1 0 4520 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_56
timestamp 1569543463
transform 1 0 4456 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_57
timestamp 1569543463
transform 1 0 4648 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_58
timestamp 1569543463
transform 1 0 4648 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_59
timestamp 1569543463
transform 1 0 4520 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_60
timestamp 1569543463
transform 1 0 4584 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_61
timestamp 1569543463
transform 1 0 4648 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_62
timestamp 1569543463
transform 1 0 4392 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_63
timestamp 1569543463
transform 1 0 4520 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_64
timestamp 1569543463
transform 1 0 4392 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_65
timestamp 1569543463
transform 1 0 4648 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_66
timestamp 1569543463
transform 1 0 4392 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_67
timestamp 1569543463
transform 1 0 4456 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_68
timestamp 1569543463
transform 1 0 4392 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_69
timestamp 1569543463
transform 1 0 4584 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_70
timestamp 1569543463
transform 1 0 4776 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_71
timestamp 1569543463
transform 1 0 4712 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_72
timestamp 1569543463
transform 1 0 4840 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_73
timestamp 1569543463
transform 1 0 4904 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_74
timestamp 1569543463
transform 1 0 4904 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_75
timestamp 1569543463
transform 1 0 4904 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_76
timestamp 1569543463
transform 1 0 4840 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_77
timestamp 1569543463
transform 1 0 4776 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_78
timestamp 1569543463
transform 1 0 4904 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_79
timestamp 1569543463
transform 1 0 4776 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_80
timestamp 1569543463
transform 1 0 4840 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_81
timestamp 1569543463
transform 1 0 4712 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_82
timestamp 1569543463
transform 1 0 4712 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_83
timestamp 1569543463
transform 1 0 4840 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_84
timestamp 1569543463
transform 1 0 4904 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_85
timestamp 1569543463
transform 1 0 4776 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_86
timestamp 1569543463
transform 1 0 4712 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_87
timestamp 1569543463
transform 1 0 4840 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_88
timestamp 1569543463
transform 1 0 4712 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_89
timestamp 1569543463
transform 1 0 4776 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_90
timestamp 1569543463
transform 1 0 4136 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_91
timestamp 1569543463
transform 1 0 4264 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_92
timestamp 1569543463
transform 1 0 4200 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_93
timestamp 1569543463
transform 1 0 4200 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_94
timestamp 1569543463
transform 1 0 4200 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_95
timestamp 1569543463
transform 1 0 4072 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_96
timestamp 1569543463
transform 1 0 4072 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_97
timestamp 1569543463
transform 1 0 4136 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_98
timestamp 1569543463
transform 1 0 4200 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_99
timestamp 1569543463
transform 1 0 4072 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_100
timestamp 1569543463
transform 1 0 4072 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_101
timestamp 1569543463
transform 1 0 4328 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_102
timestamp 1569543463
transform 1 0 4136 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_103
timestamp 1569543463
transform 1 0 4328 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_104
timestamp 1569543463
transform 1 0 4264 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_105
timestamp 1569543463
transform 1 0 4200 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_106
timestamp 1569543463
transform 1 0 4136 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_107
timestamp 1569543463
transform 1 0 4328 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_108
timestamp 1569543463
transform 1 0 4328 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_109
timestamp 1569543463
transform 1 0 4264 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_110
timestamp 1569543463
transform 1 0 4264 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_111
timestamp 1569543463
transform 1 0 4264 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_112
timestamp 1569543463
transform 1 0 4072 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_113
timestamp 1569543463
transform 1 0 4136 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_114
timestamp 1569543463
transform 1 0 4328 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_115
timestamp 1569543463
transform 1 0 3816 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_116
timestamp 1569543463
transform 1 0 3880 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_117
timestamp 1569543463
transform 1 0 4008 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_118
timestamp 1569543463
transform 1 0 3816 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_119
timestamp 1569543463
transform 1 0 3944 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_120
timestamp 1569543463
transform 1 0 3752 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_121
timestamp 1569543463
transform 1 0 3944 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_122
timestamp 1569543463
transform 1 0 3880 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_123
timestamp 1569543463
transform 1 0 4008 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_124
timestamp 1569543463
transform 1 0 3944 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_125
timestamp 1569543463
transform 1 0 3944 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_126
timestamp 1569543463
transform 1 0 3880 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_127
timestamp 1569543463
transform 1 0 3752 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_128
timestamp 1569543463
transform 1 0 4008 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_129
timestamp 1569543463
transform 1 0 3752 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_130
timestamp 1569543463
transform 1 0 4008 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_131
timestamp 1569543463
transform 1 0 3944 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_132
timestamp 1569543463
transform 1 0 3880 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_133
timestamp 1569543463
transform 1 0 3816 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_134
timestamp 1569543463
transform 1 0 4008 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_135
timestamp 1569543463
transform 1 0 3752 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_136
timestamp 1569543463
transform 1 0 3752 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_137
timestamp 1569543463
transform 1 0 3816 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_138
timestamp 1569543463
transform 1 0 3880 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_139
timestamp 1569543463
transform 1 0 3816 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_140
timestamp 1569543463
transform 1 0 3752 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_141
timestamp 1569543463
transform 1 0 3880 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_142
timestamp 1569543463
transform 1 0 3944 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_143
timestamp 1569543463
transform 1 0 3752 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_144
timestamp 1569543463
transform 1 0 3816 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_145
timestamp 1569543463
transform 1 0 3752 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_146
timestamp 1569543463
transform 1 0 3944 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_147
timestamp 1569543463
transform 1 0 4008 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_148
timestamp 1569543463
transform 1 0 4008 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_149
timestamp 1569543463
transform 1 0 3880 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_150
timestamp 1569543463
transform 1 0 4008 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_151
timestamp 1569543463
transform 1 0 3944 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_152
timestamp 1569543463
transform 1 0 3880 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_153
timestamp 1569543463
transform 1 0 4008 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_154
timestamp 1569543463
transform 1 0 3880 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_155
timestamp 1569543463
transform 1 0 3752 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_156
timestamp 1569543463
transform 1 0 3816 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_157
timestamp 1569543463
transform 1 0 4008 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_158
timestamp 1569543463
transform 1 0 3944 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_159
timestamp 1569543463
transform 1 0 3816 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_160
timestamp 1569543463
transform 1 0 3816 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_161
timestamp 1569543463
transform 1 0 3944 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_162
timestamp 1569543463
transform 1 0 3752 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_163
timestamp 1569543463
transform 1 0 3816 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_164
timestamp 1569543463
transform 1 0 3880 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_165
timestamp 1569543463
transform 1 0 4200 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_166
timestamp 1569543463
transform 1 0 4072 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_167
timestamp 1569543463
transform 1 0 4200 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_168
timestamp 1569543463
transform 1 0 4264 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_169
timestamp 1569543463
transform 1 0 4072 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_170
timestamp 1569543463
transform 1 0 4136 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_171
timestamp 1569543463
transform 1 0 4200 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_172
timestamp 1569543463
transform 1 0 4264 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_173
timestamp 1569543463
transform 1 0 4328 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_174
timestamp 1569543463
transform 1 0 4136 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_175
timestamp 1569543463
transform 1 0 4136 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_176
timestamp 1569543463
transform 1 0 4328 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_177
timestamp 1569543463
transform 1 0 4072 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_178
timestamp 1569543463
transform 1 0 4328 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_179
timestamp 1569543463
transform 1 0 4200 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_180
timestamp 1569543463
transform 1 0 4328 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_181
timestamp 1569543463
transform 1 0 4264 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_182
timestamp 1569543463
transform 1 0 4328 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_183
timestamp 1569543463
transform 1 0 4200 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_184
timestamp 1569543463
transform 1 0 4264 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_185
timestamp 1569543463
transform 1 0 4072 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_186
timestamp 1569543463
transform 1 0 4136 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_187
timestamp 1569543463
transform 1 0 4264 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_188
timestamp 1569543463
transform 1 0 4072 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_189
timestamp 1569543463
transform 1 0 4136 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_190
timestamp 1569543463
transform 1 0 4136 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_191
timestamp 1569543463
transform 1 0 4264 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_192
timestamp 1569543463
transform 1 0 4200 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_193
timestamp 1569543463
transform 1 0 4072 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_194
timestamp 1569543463
transform 1 0 4264 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_195
timestamp 1569543463
transform 1 0 4328 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_196
timestamp 1569543463
transform 1 0 4072 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_197
timestamp 1569543463
transform 1 0 4328 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_198
timestamp 1569543463
transform 1 0 4136 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_199
timestamp 1569543463
transform 1 0 4200 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_200
timestamp 1569543463
transform 1 0 4136 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_201
timestamp 1569543463
transform 1 0 4264 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_202
timestamp 1569543463
transform 1 0 4328 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_203
timestamp 1569543463
transform 1 0 4200 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_204
timestamp 1569543463
transform 1 0 4072 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_205
timestamp 1569543463
transform 1 0 4136 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_206
timestamp 1569543463
transform 1 0 4200 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_207
timestamp 1569543463
transform 1 0 4264 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_208
timestamp 1569543463
transform 1 0 4072 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_209
timestamp 1569543463
transform 1 0 4136 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_210
timestamp 1569543463
transform 1 0 4328 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_211
timestamp 1569543463
transform 1 0 4264 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_212
timestamp 1569543463
transform 1 0 4328 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_213
timestamp 1569543463
transform 1 0 4072 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_214
timestamp 1569543463
transform 1 0 4200 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_215
timestamp 1569543463
transform 1 0 3816 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_216
timestamp 1569543463
transform 1 0 4008 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_217
timestamp 1569543463
transform 1 0 4008 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_218
timestamp 1569543463
transform 1 0 3752 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_219
timestamp 1569543463
transform 1 0 3880 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_220
timestamp 1569543463
transform 1 0 3816 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_221
timestamp 1569543463
transform 1 0 3944 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_222
timestamp 1569543463
transform 1 0 3752 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_223
timestamp 1569543463
transform 1 0 3944 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_224
timestamp 1569543463
transform 1 0 3816 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_225
timestamp 1569543463
transform 1 0 3816 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_226
timestamp 1569543463
transform 1 0 3752 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_227
timestamp 1569543463
transform 1 0 3752 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_228
timestamp 1569543463
transform 1 0 3944 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_229
timestamp 1569543463
transform 1 0 4008 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_230
timestamp 1569543463
transform 1 0 3880 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_231
timestamp 1569543463
transform 1 0 4008 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_232
timestamp 1569543463
transform 1 0 4008 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_233
timestamp 1569543463
transform 1 0 3816 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_234
timestamp 1569543463
transform 1 0 3880 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_235
timestamp 1569543463
transform 1 0 3944 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_236
timestamp 1569543463
transform 1 0 3944 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_237
timestamp 1569543463
transform 1 0 3880 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_238
timestamp 1569543463
transform 1 0 3752 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_239
timestamp 1569543463
transform 1 0 3880 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_240
timestamp 1569543463
transform 1 0 3816 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_241
timestamp 1569543463
transform 1 0 4008 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_242
timestamp 1569543463
transform 1 0 3880 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_243
timestamp 1569543463
transform 1 0 3944 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_244
timestamp 1569543463
transform 1 0 3944 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_245
timestamp 1569543463
transform 1 0 3816 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_246
timestamp 1569543463
transform 1 0 3880 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_247
timestamp 1569543463
transform 1 0 4008 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_248
timestamp 1569543463
transform 1 0 3880 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_249
timestamp 1569543463
transform 1 0 3816 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_250
timestamp 1569543463
transform 1 0 3816 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_251
timestamp 1569543463
transform 1 0 4008 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_252
timestamp 1569543463
transform 1 0 3944 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_253
timestamp 1569543463
transform 1 0 3944 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_254
timestamp 1569543463
transform 1 0 3944 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_255
timestamp 1569543463
transform 1 0 3752 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_256
timestamp 1569543463
transform 1 0 3816 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_257
timestamp 1569543463
transform 1 0 3752 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_258
timestamp 1569543463
transform 1 0 4008 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_259
timestamp 1569543463
transform 1 0 3752 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_260
timestamp 1569543463
transform 1 0 3752 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_261
timestamp 1569543463
transform 1 0 3752 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_262
timestamp 1569543463
transform 1 0 4008 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_263
timestamp 1569543463
transform 1 0 3880 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_264
timestamp 1569543463
transform 1 0 3880 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_265
timestamp 1569543463
transform 1 0 4328 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_266
timestamp 1569543463
transform 1 0 4200 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_267
timestamp 1569543463
transform 1 0 4264 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_268
timestamp 1569543463
transform 1 0 4200 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_269
timestamp 1569543463
transform 1 0 4328 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_270
timestamp 1569543463
transform 1 0 4072 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_271
timestamp 1569543463
transform 1 0 4136 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_272
timestamp 1569543463
transform 1 0 4328 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_273
timestamp 1569543463
transform 1 0 4072 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_274
timestamp 1569543463
transform 1 0 4264 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_275
timestamp 1569543463
transform 1 0 4136 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_276
timestamp 1569543463
transform 1 0 4072 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_277
timestamp 1569543463
transform 1 0 4264 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_278
timestamp 1569543463
transform 1 0 4200 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_279
timestamp 1569543463
transform 1 0 4136 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_280
timestamp 1569543463
transform 1 0 4136 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_281
timestamp 1569543463
transform 1 0 4328 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_282
timestamp 1569543463
transform 1 0 4136 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_283
timestamp 1569543463
transform 1 0 4200 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_284
timestamp 1569543463
transform 1 0 4072 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_285
timestamp 1569543463
transform 1 0 4328 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_286
timestamp 1569543463
transform 1 0 4264 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_287
timestamp 1569543463
transform 1 0 4200 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_288
timestamp 1569543463
transform 1 0 4264 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_289
timestamp 1569543463
transform 1 0 4072 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_290
timestamp 1569543463
transform 1 0 4712 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_291
timestamp 1569543463
transform 1 0 4712 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_292
timestamp 1569543463
transform 1 0 4904 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_293
timestamp 1569543463
transform 1 0 4776 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_294
timestamp 1569543463
transform 1 0 4776 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_295
timestamp 1569543463
transform 1 0 4904 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_296
timestamp 1569543463
transform 1 0 4840 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_297
timestamp 1569543463
transform 1 0 4904 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_298
timestamp 1569543463
transform 1 0 4840 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_299
timestamp 1569543463
transform 1 0 4904 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_300
timestamp 1569543463
transform 1 0 4840 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_301
timestamp 1569543463
transform 1 0 4776 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_302
timestamp 1569543463
transform 1 0 4840 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_303
timestamp 1569543463
transform 1 0 4776 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_304
timestamp 1569543463
transform 1 0 4904 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_305
timestamp 1569543463
transform 1 0 4712 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_306
timestamp 1569543463
transform 1 0 4712 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_307
timestamp 1569543463
transform 1 0 4776 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_308
timestamp 1569543463
transform 1 0 4712 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_309
timestamp 1569543463
transform 1 0 4840 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_310
timestamp 1569543463
transform 1 0 4520 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_311
timestamp 1569543463
transform 1 0 4520 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_312
timestamp 1569543463
transform 1 0 4520 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_313
timestamp 1569543463
transform 1 0 4520 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_314
timestamp 1569543463
transform 1 0 4392 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_315
timestamp 1569543463
transform 1 0 4392 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_316
timestamp 1569543463
transform 1 0 4392 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_317
timestamp 1569543463
transform 1 0 4392 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_318
timestamp 1569543463
transform 1 0 4392 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_319
timestamp 1569543463
transform 1 0 4584 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_320
timestamp 1569543463
transform 1 0 4584 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_321
timestamp 1569543463
transform 1 0 4648 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_322
timestamp 1569543463
transform 1 0 4648 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_323
timestamp 1569543463
transform 1 0 4648 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_324
timestamp 1569543463
transform 1 0 4584 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_325
timestamp 1569543463
transform 1 0 4456 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_326
timestamp 1569543463
transform 1 0 4456 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_327
timestamp 1569543463
transform 1 0 4456 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_328
timestamp 1569543463
transform 1 0 4648 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_329
timestamp 1569543463
transform 1 0 4584 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_330
timestamp 1569543463
transform 1 0 4456 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_331
timestamp 1569543463
transform 1 0 4456 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_332
timestamp 1569543463
transform 1 0 4648 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_333
timestamp 1569543463
transform 1 0 4584 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_334
timestamp 1569543463
transform 1 0 4520 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_335
timestamp 1569543463
transform 1 0 4648 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_336
timestamp 1569543463
transform 1 0 4456 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_337
timestamp 1569543463
transform 1 0 4520 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_338
timestamp 1569543463
transform 1 0 4584 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_339
timestamp 1569543463
transform 1 0 4456 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_340
timestamp 1569543463
transform 1 0 4520 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_341
timestamp 1569543463
transform 1 0 4392 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_342
timestamp 1569543463
transform 1 0 4520 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_343
timestamp 1569543463
transform 1 0 4648 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_344
timestamp 1569543463
transform 1 0 4456 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_345
timestamp 1569543463
transform 1 0 4520 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_346
timestamp 1569543463
transform 1 0 4584 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_347
timestamp 1569543463
transform 1 0 4392 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_348
timestamp 1569543463
transform 1 0 4648 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_349
timestamp 1569543463
transform 1 0 4520 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_350
timestamp 1569543463
transform 1 0 4392 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_351
timestamp 1569543463
transform 1 0 4392 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_352
timestamp 1569543463
transform 1 0 4584 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_353
timestamp 1569543463
transform 1 0 4456 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_354
timestamp 1569543463
transform 1 0 4648 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_355
timestamp 1569543463
transform 1 0 4584 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_356
timestamp 1569543463
transform 1 0 4392 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_357
timestamp 1569543463
transform 1 0 4456 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_358
timestamp 1569543463
transform 1 0 4584 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_359
timestamp 1569543463
transform 1 0 4648 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_360
timestamp 1569543463
transform 1 0 4712 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_361
timestamp 1569543463
transform 1 0 4840 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_362
timestamp 1569543463
transform 1 0 4904 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_363
timestamp 1569543463
transform 1 0 4776 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_364
timestamp 1569543463
transform 1 0 4776 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_365
timestamp 1569543463
transform 1 0 4712 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_366
timestamp 1569543463
transform 1 0 4904 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_367
timestamp 1569543463
transform 1 0 4840 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_368
timestamp 1569543463
transform 1 0 4776 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_369
timestamp 1569543463
transform 1 0 4712 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_370
timestamp 1569543463
transform 1 0 4904 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_371
timestamp 1569543463
transform 1 0 4840 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_372
timestamp 1569543463
transform 1 0 4840 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_373
timestamp 1569543463
transform 1 0 4712 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_374
timestamp 1569543463
transform 1 0 4840 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_375
timestamp 1569543463
transform 1 0 4712 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_376
timestamp 1569543463
transform 1 0 4904 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_377
timestamp 1569543463
transform 1 0 4776 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_378
timestamp 1569543463
transform 1 0 4776 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_379
timestamp 1569543463
transform 1 0 4904 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_380
timestamp 1569543463
transform 1 0 3688 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_381
timestamp 1569543463
transform 1 0 3560 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_382
timestamp 1569543463
transform 1 0 3624 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_383
timestamp 1569543463
transform 1 0 3496 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_384
timestamp 1569543463
transform 1 0 3560 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_385
timestamp 1569543463
transform 1 0 3560 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_386
timestamp 1569543463
transform 1 0 3496 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_387
timestamp 1569543463
transform 1 0 3624 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_388
timestamp 1569543463
transform 1 0 3688 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_389
timestamp 1569543463
transform 1 0 3688 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_390
timestamp 1569543463
transform 1 0 3688 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_391
timestamp 1569543463
transform 1 0 3496 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_392
timestamp 1569543463
transform 1 0 3496 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_393
timestamp 1569543463
transform 1 0 3688 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_394
timestamp 1569543463
transform 1 0 3560 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_395
timestamp 1569543463
transform 1 0 3624 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_396
timestamp 1569543463
transform 1 0 3624 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_397
timestamp 1569543463
transform 1 0 3496 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_398
timestamp 1569543463
transform 1 0 3624 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_399
timestamp 1569543463
transform 1 0 3560 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_400
timestamp 1569543463
transform 1 0 3368 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_401
timestamp 1569543463
transform 1 0 3240 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_402
timestamp 1569543463
transform 1 0 3176 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_403
timestamp 1569543463
transform 1 0 3368 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_404
timestamp 1569543463
transform 1 0 3304 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_405
timestamp 1569543463
transform 1 0 3240 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_406
timestamp 1569543463
transform 1 0 3304 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_407
timestamp 1569543463
transform 1 0 3368 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_408
timestamp 1569543463
transform 1 0 3176 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_409
timestamp 1569543463
transform 1 0 3240 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_410
timestamp 1569543463
transform 1 0 3176 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_411
timestamp 1569543463
transform 1 0 3304 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_412
timestamp 1569543463
transform 1 0 3176 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_413
timestamp 1569543463
transform 1 0 3368 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_414
timestamp 1569543463
transform 1 0 3304 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_415
timestamp 1569543463
transform 1 0 3304 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_416
timestamp 1569543463
transform 1 0 3176 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_417
timestamp 1569543463
transform 1 0 3240 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_418
timestamp 1569543463
transform 1 0 3368 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_419
timestamp 1569543463
transform 1 0 3240 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_420
timestamp 1569543463
transform 1 0 3240 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_421
timestamp 1569543463
transform 1 0 3240 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_422
timestamp 1569543463
transform 1 0 3176 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_423
timestamp 1569543463
transform 1 0 3176 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_424
timestamp 1569543463
transform 1 0 3368 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_425
timestamp 1569543463
transform 1 0 3176 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_426
timestamp 1569543463
transform 1 0 3240 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_427
timestamp 1569543463
transform 1 0 3176 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_428
timestamp 1569543463
transform 1 0 3176 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_429
timestamp 1569543463
transform 1 0 3368 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_430
timestamp 1569543463
transform 1 0 3240 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_431
timestamp 1569543463
transform 1 0 3368 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_432
timestamp 1569543463
transform 1 0 3368 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_433
timestamp 1569543463
transform 1 0 3368 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_434
timestamp 1569543463
transform 1 0 3304 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_435
timestamp 1569543463
transform 1 0 3304 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_436
timestamp 1569543463
transform 1 0 3304 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_437
timestamp 1569543463
transform 1 0 3240 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_438
timestamp 1569543463
transform 1 0 3304 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_439
timestamp 1569543463
transform 1 0 3304 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_440
timestamp 1569543463
transform 1 0 3560 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_441
timestamp 1569543463
transform 1 0 3624 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_442
timestamp 1569543463
transform 1 0 3496 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_443
timestamp 1569543463
transform 1 0 3560 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_444
timestamp 1569543463
transform 1 0 3688 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_445
timestamp 1569543463
transform 1 0 3688 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_446
timestamp 1569543463
transform 1 0 3624 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_447
timestamp 1569543463
transform 1 0 3560 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_448
timestamp 1569543463
transform 1 0 3688 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_449
timestamp 1569543463
transform 1 0 3560 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_450
timestamp 1569543463
transform 1 0 3624 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_451
timestamp 1569543463
transform 1 0 3688 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_452
timestamp 1569543463
transform 1 0 3688 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_453
timestamp 1569543463
transform 1 0 3496 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_454
timestamp 1569543463
transform 1 0 3560 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_455
timestamp 1569543463
transform 1 0 3624 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_456
timestamp 1569543463
transform 1 0 3496 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_457
timestamp 1569543463
transform 1 0 3496 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_458
timestamp 1569543463
transform 1 0 3624 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_459
timestamp 1569543463
transform 1 0 3496 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_460
timestamp 1569543463
transform 1 0 3432 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_461
timestamp 1569543463
transform 1 0 3432 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_462
timestamp 1569543463
transform 1 0 3432 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_463
timestamp 1569543463
transform 1 0 3432 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_464
timestamp 1569543463
transform 1 0 3432 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_465
timestamp 1569543463
transform 1 0 3432 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_466
timestamp 1569543463
transform 1 0 3432 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_467
timestamp 1569543463
transform 1 0 3432 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_468
timestamp 1569543463
transform 1 0 3432 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_469
timestamp 1569543463
transform 1 0 3432 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_470
timestamp 1569543463
transform 1 0 3048 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_471
timestamp 1569543463
transform 1 0 2920 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_472
timestamp 1569543463
transform 1 0 3048 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_473
timestamp 1569543463
transform 1 0 3048 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_474
timestamp 1569543463
transform 1 0 2920 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_475
timestamp 1569543463
transform 1 0 2984 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_476
timestamp 1569543463
transform 1 0 2984 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_477
timestamp 1569543463
transform 1 0 2920 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_478
timestamp 1569543463
transform 1 0 2984 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_479
timestamp 1569543463
transform 1 0 2920 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_480
timestamp 1569543463
transform 1 0 2856 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_481
timestamp 1569543463
transform 1 0 3048 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_482
timestamp 1569543463
transform 1 0 3112 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_483
timestamp 1569543463
transform 1 0 2856 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_484
timestamp 1569543463
transform 1 0 3048 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_485
timestamp 1569543463
transform 1 0 3112 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_486
timestamp 1569543463
transform 1 0 2920 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_487
timestamp 1569543463
transform 1 0 3112 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_488
timestamp 1569543463
transform 1 0 3112 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_489
timestamp 1569543463
transform 1 0 2856 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_490
timestamp 1569543463
transform 1 0 2984 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_491
timestamp 1569543463
transform 1 0 2856 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_492
timestamp 1569543463
transform 1 0 3112 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_493
timestamp 1569543463
transform 1 0 2984 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_494
timestamp 1569543463
transform 1 0 2856 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_495
timestamp 1569543463
transform 1 0 2792 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_496
timestamp 1569543463
transform 1 0 2664 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_497
timestamp 1569543463
transform 1 0 2728 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_498
timestamp 1569543463
transform 1 0 2792 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_499
timestamp 1569543463
transform 1 0 2728 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_500
timestamp 1569543463
transform 1 0 2664 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_501
timestamp 1569543463
transform 1 0 2536 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_502
timestamp 1569543463
transform 1 0 2536 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_503
timestamp 1569543463
transform 1 0 2664 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_504
timestamp 1569543463
transform 1 0 2664 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_505
timestamp 1569543463
transform 1 0 2536 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_506
timestamp 1569543463
transform 1 0 2792 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_507
timestamp 1569543463
transform 1 0 2728 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_508
timestamp 1569543463
transform 1 0 2600 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_509
timestamp 1569543463
transform 1 0 2664 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_510
timestamp 1569543463
transform 1 0 2792 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_511
timestamp 1569543463
transform 1 0 2728 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_512
timestamp 1569543463
transform 1 0 2600 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_513
timestamp 1569543463
transform 1 0 2600 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_514
timestamp 1569543463
transform 1 0 2536 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_515
timestamp 1569543463
transform 1 0 2600 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_516
timestamp 1569543463
transform 1 0 2600 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_517
timestamp 1569543463
transform 1 0 2728 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_518
timestamp 1569543463
transform 1 0 2536 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_519
timestamp 1569543463
transform 1 0 2792 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_520
timestamp 1569543463
transform 1 0 2728 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_521
timestamp 1569543463
transform 1 0 2792 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_522
timestamp 1569543463
transform 1 0 2728 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_523
timestamp 1569543463
transform 1 0 2792 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_524
timestamp 1569543463
transform 1 0 2728 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_525
timestamp 1569543463
transform 1 0 2792 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_526
timestamp 1569543463
transform 1 0 2664 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_527
timestamp 1569543463
transform 1 0 2664 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_528
timestamp 1569543463
transform 1 0 2792 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_529
timestamp 1569543463
transform 1 0 2792 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_530
timestamp 1569543463
transform 1 0 2664 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_531
timestamp 1569543463
transform 1 0 2536 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_532
timestamp 1569543463
transform 1 0 2664 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_533
timestamp 1569543463
transform 1 0 2664 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_534
timestamp 1569543463
transform 1 0 2536 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_535
timestamp 1569543463
transform 1 0 2536 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_536
timestamp 1569543463
transform 1 0 2536 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_537
timestamp 1569543463
transform 1 0 2600 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_538
timestamp 1569543463
transform 1 0 2728 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_539
timestamp 1569543463
transform 1 0 2600 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_540
timestamp 1569543463
transform 1 0 2728 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_541
timestamp 1569543463
transform 1 0 2600 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_542
timestamp 1569543463
transform 1 0 2600 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_543
timestamp 1569543463
transform 1 0 2600 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_544
timestamp 1569543463
transform 1 0 2536 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_545
timestamp 1569543463
transform 1 0 2856 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_546
timestamp 1569543463
transform 1 0 3048 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_547
timestamp 1569543463
transform 1 0 3048 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_548
timestamp 1569543463
transform 1 0 3048 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_549
timestamp 1569543463
transform 1 0 3048 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_550
timestamp 1569543463
transform 1 0 3048 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_551
timestamp 1569543463
transform 1 0 2856 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_552
timestamp 1569543463
transform 1 0 2984 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_553
timestamp 1569543463
transform 1 0 2856 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_554
timestamp 1569543463
transform 1 0 2856 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_555
timestamp 1569543463
transform 1 0 3112 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_556
timestamp 1569543463
transform 1 0 3112 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_557
timestamp 1569543463
transform 1 0 2920 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_558
timestamp 1569543463
transform 1 0 3112 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_559
timestamp 1569543463
transform 1 0 3112 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_560
timestamp 1569543463
transform 1 0 2984 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_561
timestamp 1569543463
transform 1 0 3112 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_562
timestamp 1569543463
transform 1 0 2920 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_563
timestamp 1569543463
transform 1 0 2984 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_564
timestamp 1569543463
transform 1 0 2856 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_565
timestamp 1569543463
transform 1 0 2920 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_566
timestamp 1569543463
transform 1 0 2984 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_567
timestamp 1569543463
transform 1 0 2920 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_568
timestamp 1569543463
transform 1 0 2920 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_569
timestamp 1569543463
transform 1 0 2984 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_570
timestamp 1569543463
transform 1 0 3048 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_571
timestamp 1569543463
transform 1 0 2920 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_572
timestamp 1569543463
transform 1 0 3112 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_573
timestamp 1569543463
transform 1 0 2984 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_574
timestamp 1569543463
transform 1 0 3048 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_575
timestamp 1569543463
transform 1 0 3112 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_576
timestamp 1569543463
transform 1 0 2856 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_577
timestamp 1569543463
transform 1 0 2920 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_578
timestamp 1569543463
transform 1 0 2856 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_579
timestamp 1569543463
transform 1 0 3112 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_580
timestamp 1569543463
transform 1 0 2984 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_581
timestamp 1569543463
transform 1 0 3048 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_582
timestamp 1569543463
transform 1 0 2984 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_583
timestamp 1569543463
transform 1 0 2920 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_584
timestamp 1569543463
transform 1 0 2856 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_585
timestamp 1569543463
transform 1 0 3112 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_586
timestamp 1569543463
transform 1 0 2856 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_587
timestamp 1569543463
transform 1 0 2920 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_588
timestamp 1569543463
transform 1 0 3048 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_589
timestamp 1569543463
transform 1 0 2920 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_590
timestamp 1569543463
transform 1 0 3112 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_591
timestamp 1569543463
transform 1 0 2984 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_592
timestamp 1569543463
transform 1 0 3048 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_593
timestamp 1569543463
transform 1 0 2856 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_594
timestamp 1569543463
transform 1 0 2984 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_595
timestamp 1569543463
transform 1 0 2728 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_596
timestamp 1569543463
transform 1 0 2664 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_597
timestamp 1569543463
transform 1 0 2536 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_598
timestamp 1569543463
transform 1 0 2728 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_599
timestamp 1569543463
transform 1 0 2728 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_600
timestamp 1569543463
transform 1 0 2600 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_601
timestamp 1569543463
transform 1 0 2792 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_602
timestamp 1569543463
transform 1 0 2600 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_603
timestamp 1569543463
transform 1 0 2792 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_604
timestamp 1569543463
transform 1 0 2600 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_605
timestamp 1569543463
transform 1 0 2664 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_606
timestamp 1569543463
transform 1 0 2600 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_607
timestamp 1569543463
transform 1 0 2728 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_608
timestamp 1569543463
transform 1 0 2792 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_609
timestamp 1569543463
transform 1 0 2728 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_610
timestamp 1569543463
transform 1 0 2600 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_611
timestamp 1569543463
transform 1 0 2664 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_612
timestamp 1569543463
transform 1 0 2792 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_613
timestamp 1569543463
transform 1 0 2536 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_614
timestamp 1569543463
transform 1 0 2664 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_615
timestamp 1569543463
transform 1 0 2536 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_616
timestamp 1569543463
transform 1 0 2664 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_617
timestamp 1569543463
transform 1 0 2536 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_618
timestamp 1569543463
transform 1 0 2792 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_619
timestamp 1569543463
transform 1 0 2536 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_620
timestamp 1569543463
transform 1 0 2792 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_621
timestamp 1569543463
transform 1 0 2664 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_622
timestamp 1569543463
transform 1 0 2536 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_623
timestamp 1569543463
transform 1 0 2664 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_624
timestamp 1569543463
transform 1 0 2792 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_625
timestamp 1569543463
transform 1 0 2536 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_626
timestamp 1569543463
transform 1 0 2600 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_627
timestamp 1569543463
transform 1 0 2792 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_628
timestamp 1569543463
transform 1 0 2792 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_629
timestamp 1569543463
transform 1 0 2536 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_630
timestamp 1569543463
transform 1 0 2728 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_631
timestamp 1569543463
transform 1 0 2600 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_632
timestamp 1569543463
transform 1 0 2600 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_633
timestamp 1569543463
transform 1 0 2664 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_634
timestamp 1569543463
transform 1 0 2536 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_635
timestamp 1569543463
transform 1 0 2728 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_636
timestamp 1569543463
transform 1 0 2664 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_637
timestamp 1569543463
transform 1 0 2728 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_638
timestamp 1569543463
transform 1 0 2792 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_639
timestamp 1569543463
transform 1 0 2664 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_640
timestamp 1569543463
transform 1 0 2728 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_641
timestamp 1569543463
transform 1 0 2600 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_642
timestamp 1569543463
transform 1 0 2600 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_643
timestamp 1569543463
transform 1 0 2536 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_644
timestamp 1569543463
transform 1 0 2728 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_645
timestamp 1569543463
transform 1 0 2920 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_646
timestamp 1569543463
transform 1 0 2856 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_647
timestamp 1569543463
transform 1 0 2920 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_648
timestamp 1569543463
transform 1 0 2920 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_649
timestamp 1569543463
transform 1 0 2856 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_650
timestamp 1569543463
transform 1 0 3112 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_651
timestamp 1569543463
transform 1 0 3112 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_652
timestamp 1569543463
transform 1 0 3048 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_653
timestamp 1569543463
transform 1 0 2856 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_654
timestamp 1569543463
transform 1 0 3112 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_655
timestamp 1569543463
transform 1 0 2856 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_656
timestamp 1569543463
transform 1 0 3112 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_657
timestamp 1569543463
transform 1 0 2984 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_658
timestamp 1569543463
transform 1 0 3048 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_659
timestamp 1569543463
transform 1 0 2856 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_660
timestamp 1569543463
transform 1 0 2984 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_661
timestamp 1569543463
transform 1 0 2984 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_662
timestamp 1569543463
transform 1 0 2984 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_663
timestamp 1569543463
transform 1 0 2920 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_664
timestamp 1569543463
transform 1 0 2984 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_665
timestamp 1569543463
transform 1 0 2920 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_666
timestamp 1569543463
transform 1 0 3048 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_667
timestamp 1569543463
transform 1 0 3112 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_668
timestamp 1569543463
transform 1 0 3048 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_669
timestamp 1569543463
transform 1 0 3048 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_670
timestamp 1569543463
transform 1 0 3496 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_671
timestamp 1569543463
transform 1 0 3624 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_672
timestamp 1569543463
transform 1 0 3560 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_673
timestamp 1569543463
transform 1 0 3496 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_674
timestamp 1569543463
transform 1 0 3624 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_675
timestamp 1569543463
transform 1 0 3560 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_676
timestamp 1569543463
transform 1 0 3496 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_677
timestamp 1569543463
transform 1 0 3560 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_678
timestamp 1569543463
transform 1 0 3688 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_679
timestamp 1569543463
transform 1 0 3496 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_680
timestamp 1569543463
transform 1 0 3688 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_681
timestamp 1569543463
transform 1 0 3624 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_682
timestamp 1569543463
transform 1 0 3688 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_683
timestamp 1569543463
transform 1 0 3496 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_684
timestamp 1569543463
transform 1 0 3560 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_685
timestamp 1569543463
transform 1 0 3688 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_686
timestamp 1569543463
transform 1 0 3560 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_687
timestamp 1569543463
transform 1 0 3688 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_688
timestamp 1569543463
transform 1 0 3624 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_689
timestamp 1569543463
transform 1 0 3624 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_690
timestamp 1569543463
transform 1 0 3240 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_691
timestamp 1569543463
transform 1 0 3240 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_692
timestamp 1569543463
transform 1 0 3368 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_693
timestamp 1569543463
transform 1 0 3304 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_694
timestamp 1569543463
transform 1 0 3304 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_695
timestamp 1569543463
transform 1 0 3304 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_696
timestamp 1569543463
transform 1 0 3304 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_697
timestamp 1569543463
transform 1 0 3304 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_698
timestamp 1569543463
transform 1 0 3368 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_699
timestamp 1569543463
transform 1 0 3368 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_700
timestamp 1569543463
transform 1 0 3368 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_701
timestamp 1569543463
transform 1 0 3176 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_702
timestamp 1569543463
transform 1 0 3176 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_703
timestamp 1569543463
transform 1 0 3176 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_704
timestamp 1569543463
transform 1 0 3176 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_705
timestamp 1569543463
transform 1 0 3176 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_706
timestamp 1569543463
transform 1 0 3368 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_707
timestamp 1569543463
transform 1 0 3240 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_708
timestamp 1569543463
transform 1 0 3240 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_709
timestamp 1569543463
transform 1 0 3240 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_710
timestamp 1569543463
transform 1 0 3368 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_711
timestamp 1569543463
transform 1 0 3176 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_712
timestamp 1569543463
transform 1 0 3368 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_713
timestamp 1569543463
transform 1 0 3176 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_714
timestamp 1569543463
transform 1 0 3368 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_715
timestamp 1569543463
transform 1 0 3368 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_716
timestamp 1569543463
transform 1 0 3240 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_717
timestamp 1569543463
transform 1 0 3304 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_718
timestamp 1569543463
transform 1 0 3176 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_719
timestamp 1569543463
transform 1 0 3240 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_720
timestamp 1569543463
transform 1 0 3368 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_721
timestamp 1569543463
transform 1 0 3240 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_722
timestamp 1569543463
transform 1 0 3304 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_723
timestamp 1569543463
transform 1 0 3176 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_724
timestamp 1569543463
transform 1 0 3304 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_725
timestamp 1569543463
transform 1 0 3240 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_726
timestamp 1569543463
transform 1 0 3304 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_727
timestamp 1569543463
transform 1 0 3240 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_728
timestamp 1569543463
transform 1 0 3304 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_729
timestamp 1569543463
transform 1 0 3176 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_730
timestamp 1569543463
transform 1 0 3624 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_731
timestamp 1569543463
transform 1 0 3624 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_732
timestamp 1569543463
transform 1 0 3496 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_733
timestamp 1569543463
transform 1 0 3624 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_734
timestamp 1569543463
transform 1 0 3560 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_735
timestamp 1569543463
transform 1 0 3688 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_736
timestamp 1569543463
transform 1 0 3560 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_737
timestamp 1569543463
transform 1 0 3560 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_738
timestamp 1569543463
transform 1 0 3688 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_739
timestamp 1569543463
transform 1 0 3624 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_740
timestamp 1569543463
transform 1 0 3688 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_741
timestamp 1569543463
transform 1 0 3624 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_742
timestamp 1569543463
transform 1 0 3496 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_743
timestamp 1569543463
transform 1 0 3560 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_744
timestamp 1569543463
transform 1 0 3496 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_745
timestamp 1569543463
transform 1 0 3496 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_746
timestamp 1569543463
transform 1 0 3688 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_747
timestamp 1569543463
transform 1 0 3496 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_748
timestamp 1569543463
transform 1 0 3560 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_749
timestamp 1569543463
transform 1 0 3688 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_750
timestamp 1569543463
transform 1 0 3432 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_751
timestamp 1569543463
transform 1 0 3432 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_752
timestamp 1569543463
transform 1 0 3432 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_753
timestamp 1569543463
transform 1 0 3432 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_754
timestamp 1569543463
transform 1 0 3432 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_755
timestamp 1569543463
transform 1 0 3432 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_756
timestamp 1569543463
transform 1 0 3432 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_757
timestamp 1569543463
transform 1 0 3432 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_758
timestamp 1569543463
transform 1 0 3432 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_759
timestamp 1569543463
transform 1 0 3432 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_760
timestamp 1569543463
transform 1 0 3688 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_761
timestamp 1569543463
transform 1 0 3368 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_762
timestamp 1569543463
transform 1 0 3624 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_763
timestamp 1569543463
transform 1 0 3496 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_764
timestamp 1569543463
transform 1 0 3432 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_765
timestamp 1569543463
transform 1 0 3304 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_766
timestamp 1569543463
transform 1 0 3176 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_767
timestamp 1569543463
transform 1 0 3688 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_768
timestamp 1569543463
transform 1 0 3432 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_769
timestamp 1569543463
transform 1 0 3432 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_770
timestamp 1569543463
transform 1 0 3624 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_771
timestamp 1569543463
transform 1 0 3176 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_772
timestamp 1569543463
transform 1 0 3240 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_773
timestamp 1569543463
transform 1 0 3240 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_774
timestamp 1569543463
transform 1 0 3176 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_775
timestamp 1569543463
transform 1 0 3560 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_776
timestamp 1569543463
transform 1 0 3496 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_777
timestamp 1569543463
transform 1 0 3432 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_778
timestamp 1569543463
transform 1 0 3560 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_779
timestamp 1569543463
transform 1 0 3624 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_780
timestamp 1569543463
transform 1 0 3624 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_781
timestamp 1569543463
transform 1 0 3240 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_782
timestamp 1569543463
transform 1 0 3176 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_783
timestamp 1569543463
transform 1 0 3688 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_784
timestamp 1569543463
transform 1 0 3304 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_785
timestamp 1569543463
transform 1 0 3240 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_786
timestamp 1569543463
transform 1 0 3304 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_787
timestamp 1569543463
transform 1 0 3688 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_788
timestamp 1569543463
transform 1 0 3496 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_789
timestamp 1569543463
transform 1 0 3304 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_790
timestamp 1569543463
transform 1 0 3368 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_791
timestamp 1569543463
transform 1 0 3496 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_792
timestamp 1569543463
transform 1 0 3368 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_793
timestamp 1569543463
transform 1 0 3560 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_794
timestamp 1569543463
transform 1 0 3560 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_795
timestamp 1569543463
transform 1 0 3368 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_796
timestamp 1569543463
transform 1 0 3112 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_797
timestamp 1569543463
transform 1 0 3048 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_798
timestamp 1569543463
transform 1 0 2920 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_799
timestamp 1569543463
transform 1 0 3112 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_800
timestamp 1569543463
transform 1 0 2984 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_801
timestamp 1569543463
transform 1 0 2984 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_802
timestamp 1569543463
transform 1 0 2920 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_803
timestamp 1569543463
transform 1 0 2856 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_804
timestamp 1569543463
transform 1 0 3048 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_805
timestamp 1569543463
transform 1 0 2920 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_806
timestamp 1569543463
transform 1 0 2984 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_807
timestamp 1569543463
transform 1 0 2920 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_808
timestamp 1569543463
transform 1 0 3112 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_809
timestamp 1569543463
transform 1 0 2856 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_810
timestamp 1569543463
transform 1 0 3112 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_811
timestamp 1569543463
transform 1 0 3048 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_812
timestamp 1569543463
transform 1 0 2984 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_813
timestamp 1569543463
transform 1 0 2856 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_814
timestamp 1569543463
transform 1 0 3048 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_815
timestamp 1569543463
transform 1 0 2856 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_816
timestamp 1569543463
transform 1 0 2664 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_817
timestamp 1569543463
transform 1 0 2600 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_818
timestamp 1569543463
transform 1 0 2792 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_819
timestamp 1569543463
transform 1 0 2664 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_820
timestamp 1569543463
transform 1 0 2728 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_821
timestamp 1569543463
transform 1 0 2536 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_822
timestamp 1569543463
transform 1 0 2728 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_823
timestamp 1569543463
transform 1 0 2728 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_824
timestamp 1569543463
transform 1 0 2664 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_825
timestamp 1569543463
transform 1 0 2600 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_826
timestamp 1569543463
transform 1 0 2792 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_827
timestamp 1569543463
transform 1 0 2536 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_828
timestamp 1569543463
transform 1 0 2728 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_829
timestamp 1569543463
transform 1 0 2792 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_830
timestamp 1569543463
transform 1 0 2792 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_831
timestamp 1569543463
transform 1 0 2600 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_832
timestamp 1569543463
transform 1 0 2536 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_833
timestamp 1569543463
transform 1 0 2664 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_834
timestamp 1569543463
transform 1 0 2600 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_835
timestamp 1569543463
transform 1 0 2536 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_836
timestamp 1569543463
transform 1 0 2664 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_837
timestamp 1569543463
transform 1 0 2600 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_838
timestamp 1569543463
transform 1 0 2536 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_839
timestamp 1569543463
transform 1 0 2728 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_840
timestamp 1569543463
transform 1 0 2536 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_841
timestamp 1569543463
transform 1 0 2600 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_842
timestamp 1569543463
transform 1 0 2600 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_843
timestamp 1569543463
transform 1 0 2600 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_844
timestamp 1569543463
transform 1 0 2792 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_845
timestamp 1569543463
transform 1 0 2664 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_846
timestamp 1569543463
transform 1 0 2664 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_847
timestamp 1569543463
transform 1 0 2536 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_848
timestamp 1569543463
transform 1 0 2536 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_849
timestamp 1569543463
transform 1 0 2728 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_850
timestamp 1569543463
transform 1 0 2664 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_851
timestamp 1569543463
transform 1 0 2536 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_852
timestamp 1569543463
transform 1 0 2600 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_853
timestamp 1569543463
transform 1 0 2728 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_854
timestamp 1569543463
transform 1 0 2792 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_855
timestamp 1569543463
transform 1 0 2856 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_856
timestamp 1569543463
transform 1 0 2536 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_857
timestamp 1569543463
transform 1 0 3688 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_858
timestamp 1569543463
transform 1 0 3624 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_859
timestamp 1569543463
transform 1 0 3688 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_860
timestamp 1569543463
transform 1 0 3688 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_861
timestamp 1569543463
transform 1 0 3240 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_862
timestamp 1569543463
transform 1 0 3432 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_863
timestamp 1569543463
transform 1 0 3432 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_864
timestamp 1569543463
transform 1 0 3432 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_865
timestamp 1569543463
transform 1 0 3496 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_866
timestamp 1569543463
transform 1 0 3496 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_867
timestamp 1569543463
transform 1 0 3496 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_868
timestamp 1569543463
transform 1 0 3304 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_869
timestamp 1569543463
transform 1 0 3304 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_870
timestamp 1569543463
transform 1 0 3560 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_871
timestamp 1569543463
transform 1 0 3560 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_872
timestamp 1569543463
transform 1 0 3560 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_873
timestamp 1569543463
transform 1 0 3368 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_874
timestamp 1569543463
transform 1 0 3368 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_875
timestamp 1569543463
transform 1 0 3624 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_876
timestamp 1569543463
transform 1 0 3368 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_877
timestamp 1569543463
transform 1 0 3624 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_878
timestamp 1569543463
transform 1 0 4648 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_879
timestamp 1569543463
transform 1 0 4712 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_880
timestamp 1569543463
transform 1 0 4392 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_881
timestamp 1569543463
transform 1 0 4904 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_882
timestamp 1569543463
transform 1 0 4712 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_883
timestamp 1569543463
transform 1 0 4584 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_884
timestamp 1569543463
transform 1 0 4456 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_885
timestamp 1569543463
transform 1 0 4584 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_886
timestamp 1569543463
transform 1 0 4712 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_887
timestamp 1569543463
transform 1 0 4456 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_888
timestamp 1569543463
transform 1 0 4840 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_889
timestamp 1569543463
transform 1 0 4776 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_890
timestamp 1569543463
transform 1 0 4648 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_891
timestamp 1569543463
transform 1 0 4840 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_892
timestamp 1569543463
transform 1 0 4776 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_893
timestamp 1569543463
transform 1 0 4456 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_894
timestamp 1569543463
transform 1 0 4584 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_895
timestamp 1569543463
transform 1 0 4520 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_896
timestamp 1569543463
transform 1 0 4840 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_897
timestamp 1569543463
transform 1 0 4776 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_898
timestamp 1569543463
transform 1 0 4776 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_899
timestamp 1569543463
transform 1 0 4520 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_900
timestamp 1569543463
transform 1 0 4392 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_901
timestamp 1569543463
transform 1 0 4904 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_902
timestamp 1569543463
transform 1 0 4520 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_903
timestamp 1569543463
transform 1 0 4520 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_904
timestamp 1569543463
transform 1 0 4648 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_905
timestamp 1569543463
transform 1 0 4648 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_906
timestamp 1569543463
transform 1 0 4712 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_907
timestamp 1569543463
transform 1 0 4584 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_908
timestamp 1569543463
transform 1 0 4456 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_909
timestamp 1569543463
transform 1 0 4392 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_910
timestamp 1569543463
transform 1 0 4904 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_911
timestamp 1569543463
transform 1 0 4392 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_912
timestamp 1569543463
transform 1 0 4904 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_913
timestamp 1569543463
transform 1 0 4840 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_914
timestamp 1569543463
transform 1 0 4072 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_915
timestamp 1569543463
transform 1 0 3944 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_916
timestamp 1569543463
transform 1 0 3880 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_917
timestamp 1569543463
transform 1 0 4136 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_918
timestamp 1569543463
transform 1 0 3880 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_919
timestamp 1569543463
transform 1 0 3944 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_920
timestamp 1569543463
transform 1 0 4200 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_921
timestamp 1569543463
transform 1 0 4200 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_922
timestamp 1569543463
transform 1 0 3880 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_923
timestamp 1569543463
transform 1 0 3944 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_924
timestamp 1569543463
transform 1 0 4200 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_925
timestamp 1569543463
transform 1 0 3944 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_926
timestamp 1569543463
transform 1 0 3752 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_927
timestamp 1569543463
transform 1 0 4136 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_928
timestamp 1569543463
transform 1 0 4200 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_929
timestamp 1569543463
transform 1 0 4264 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_930
timestamp 1569543463
transform 1 0 4008 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_931
timestamp 1569543463
transform 1 0 4008 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_932
timestamp 1569543463
transform 1 0 3752 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_933
timestamp 1569543463
transform 1 0 4264 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_934
timestamp 1569543463
transform 1 0 3880 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_935
timestamp 1569543463
transform 1 0 4008 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_936
timestamp 1569543463
transform 1 0 3816 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_937
timestamp 1569543463
transform 1 0 3752 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_938
timestamp 1569543463
transform 1 0 4264 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_939
timestamp 1569543463
transform 1 0 4328 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_940
timestamp 1569543463
transform 1 0 4264 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_941
timestamp 1569543463
transform 1 0 3752 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_942
timestamp 1569543463
transform 1 0 4072 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_943
timestamp 1569543463
transform 1 0 4136 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_944
timestamp 1569543463
transform 1 0 3816 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_945
timestamp 1569543463
transform 1 0 4328 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_946
timestamp 1569543463
transform 1 0 4072 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_947
timestamp 1569543463
transform 1 0 3816 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_948
timestamp 1569543463
transform 1 0 4328 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_949
timestamp 1569543463
transform 1 0 4072 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_950
timestamp 1569543463
transform 1 0 3816 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_951
timestamp 1569543463
transform 1 0 4328 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_952
timestamp 1569543463
transform 1 0 4008 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_953
timestamp 1569543463
transform 1 0 4136 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_954
timestamp 1569543463
transform 1 0 4072 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_955
timestamp 1569543463
transform 1 0 4072 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_956
timestamp 1569543463
transform 1 0 3752 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_957
timestamp 1569543463
transform 1 0 4072 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_958
timestamp 1569543463
transform 1 0 3880 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_959
timestamp 1569543463
transform 1 0 3816 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_960
timestamp 1569543463
transform 1 0 3880 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_961
timestamp 1569543463
transform 1 0 4136 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_962
timestamp 1569543463
transform 1 0 3880 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_963
timestamp 1569543463
transform 1 0 3752 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_964
timestamp 1569543463
transform 1 0 4136 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_965
timestamp 1569543463
transform 1 0 4136 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_966
timestamp 1569543463
transform 1 0 3944 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_967
timestamp 1569543463
transform 1 0 4328 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_968
timestamp 1569543463
transform 1 0 4200 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_969
timestamp 1569543463
transform 1 0 3944 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_970
timestamp 1569543463
transform 1 0 4200 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_971
timestamp 1569543463
transform 1 0 3944 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_972
timestamp 1569543463
transform 1 0 4328 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_973
timestamp 1569543463
transform 1 0 4200 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_974
timestamp 1569543463
transform 1 0 4328 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_975
timestamp 1569543463
transform 1 0 4264 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_976
timestamp 1569543463
transform 1 0 3816 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_977
timestamp 1569543463
transform 1 0 4264 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_978
timestamp 1569543463
transform 1 0 4264 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_979
timestamp 1569543463
transform 1 0 4008 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_980
timestamp 1569543463
transform 1 0 4008 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_981
timestamp 1569543463
transform 1 0 3816 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_982
timestamp 1569543463
transform 1 0 4008 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_983
timestamp 1569543463
transform 1 0 3752 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_984
timestamp 1569543463
transform 1 0 4520 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_985
timestamp 1569543463
transform 1 0 4520 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_986
timestamp 1569543463
transform 1 0 4520 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_987
timestamp 1569543463
transform 1 0 4584 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_988
timestamp 1569543463
transform 1 0 4584 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_989
timestamp 1569543463
transform 1 0 4584 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_990
timestamp 1569543463
transform 1 0 4456 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_991
timestamp 1569543463
transform 1 0 4648 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_992
timestamp 1569543463
transform 1 0 4648 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_993
timestamp 1569543463
transform 1 0 4648 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_994
timestamp 1569543463
transform 1 0 4712 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_995
timestamp 1569543463
transform 1 0 4712 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_996
timestamp 1569543463
transform 1 0 4712 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_997
timestamp 1569543463
transform 1 0 4776 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_998
timestamp 1569543463
transform 1 0 4776 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_999
timestamp 1569543463
transform 1 0 4776 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1000
timestamp 1569543463
transform 1 0 4840 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1001
timestamp 1569543463
transform 1 0 4840 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1002
timestamp 1569543463
transform 1 0 4840 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1003
timestamp 1569543463
transform 1 0 4904 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1004
timestamp 1569543463
transform 1 0 4904 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1005
timestamp 1569543463
transform 1 0 4904 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1006
timestamp 1569543463
transform 1 0 4392 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1007
timestamp 1569543463
transform 1 0 4392 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1008
timestamp 1569543463
transform 1 0 4392 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1009
timestamp 1569543463
transform 1 0 4456 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1010
timestamp 1569543463
transform 1 0 4456 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1011
timestamp 1569543463
transform 1 0 2472 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1012
timestamp 1569543463
transform 1 0 2472 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1013
timestamp 1569543463
transform 1 0 2344 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1014
timestamp 1569543463
transform 1 0 2216 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1015
timestamp 1569543463
transform 1 0 2408 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1016
timestamp 1569543463
transform 1 0 2344 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1017
timestamp 1569543463
transform 1 0 2216 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1018
timestamp 1569543463
transform 1 0 2344 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1019
timestamp 1569543463
transform 1 0 2472 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1020
timestamp 1569543463
transform 1 0 2280 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1021
timestamp 1569543463
transform 1 0 2408 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1022
timestamp 1569543463
transform 1 0 2216 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1023
timestamp 1569543463
transform 1 0 2344 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1024
timestamp 1569543463
transform 1 0 2344 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1025
timestamp 1569543463
transform 1 0 2408 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1026
timestamp 1569543463
transform 1 0 2280 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1027
timestamp 1569543463
transform 1 0 2280 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1028
timestamp 1569543463
transform 1 0 2408 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1029
timestamp 1569543463
transform 1 0 2408 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1030
timestamp 1569543463
transform 1 0 2280 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1031
timestamp 1569543463
transform 1 0 2472 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1032
timestamp 1569543463
transform 1 0 2216 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1033
timestamp 1569543463
transform 1 0 2216 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1034
timestamp 1569543463
transform 1 0 2472 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1035
timestamp 1569543463
transform 1 0 2280 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1036
timestamp 1569543463
transform 1 0 2088 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1037
timestamp 1569543463
transform 1 0 2088 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1038
timestamp 1569543463
transform 1 0 1960 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1039
timestamp 1569543463
transform 1 0 2088 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1040
timestamp 1569543463
transform 1 0 2088 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1041
timestamp 1569543463
transform 1 0 2152 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1042
timestamp 1569543463
transform 1 0 2152 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1043
timestamp 1569543463
transform 1 0 1960 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1044
timestamp 1569543463
transform 1 0 2152 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1045
timestamp 1569543463
transform 1 0 1960 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1046
timestamp 1569543463
transform 1 0 1960 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1047
timestamp 1569543463
transform 1 0 1960 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1048
timestamp 1569543463
transform 1 0 2024 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1049
timestamp 1569543463
transform 1 0 2024 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1050
timestamp 1569543463
transform 1 0 2024 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1051
timestamp 1569543463
transform 1 0 1896 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1052
timestamp 1569543463
transform 1 0 2152 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1053
timestamp 1569543463
transform 1 0 1896 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1054
timestamp 1569543463
transform 1 0 2024 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1055
timestamp 1569543463
transform 1 0 2024 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1056
timestamp 1569543463
transform 1 0 1896 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1057
timestamp 1569543463
transform 1 0 2152 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1058
timestamp 1569543463
transform 1 0 1896 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1059
timestamp 1569543463
transform 1 0 2088 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1060
timestamp 1569543463
transform 1 0 1896 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1061
timestamp 1569543463
transform 1 0 1896 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1062
timestamp 1569543463
transform 1 0 2152 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1063
timestamp 1569543463
transform 1 0 1960 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1064
timestamp 1569543463
transform 1 0 1960 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1065
timestamp 1569543463
transform 1 0 1960 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1066
timestamp 1569543463
transform 1 0 1960 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1067
timestamp 1569543463
transform 1 0 2152 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1068
timestamp 1569543463
transform 1 0 1960 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1069
timestamp 1569543463
transform 1 0 2152 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1070
timestamp 1569543463
transform 1 0 2024 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1071
timestamp 1569543463
transform 1 0 2024 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1072
timestamp 1569543463
transform 1 0 2024 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1073
timestamp 1569543463
transform 1 0 2024 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1074
timestamp 1569543463
transform 1 0 2024 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1075
timestamp 1569543463
transform 1 0 2152 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1076
timestamp 1569543463
transform 1 0 2152 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1077
timestamp 1569543463
transform 1 0 1896 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1078
timestamp 1569543463
transform 1 0 2088 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1079
timestamp 1569543463
transform 1 0 1896 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1080
timestamp 1569543463
transform 1 0 1896 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1081
timestamp 1569543463
transform 1 0 2088 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1082
timestamp 1569543463
transform 1 0 2088 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1083
timestamp 1569543463
transform 1 0 2088 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1084
timestamp 1569543463
transform 1 0 1896 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1085
timestamp 1569543463
transform 1 0 2088 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1086
timestamp 1569543463
transform 1 0 2344 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1087
timestamp 1569543463
transform 1 0 2344 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1088
timestamp 1569543463
transform 1 0 2344 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1089
timestamp 1569543463
transform 1 0 2472 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1090
timestamp 1569543463
transform 1 0 2472 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1091
timestamp 1569543463
transform 1 0 2472 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1092
timestamp 1569543463
transform 1 0 2472 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1093
timestamp 1569543463
transform 1 0 2472 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1094
timestamp 1569543463
transform 1 0 2344 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1095
timestamp 1569543463
transform 1 0 2216 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1096
timestamp 1569543463
transform 1 0 2216 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1097
timestamp 1569543463
transform 1 0 2216 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1098
timestamp 1569543463
transform 1 0 2216 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1099
timestamp 1569543463
transform 1 0 2344 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1100
timestamp 1569543463
transform 1 0 2216 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1101
timestamp 1569543463
transform 1 0 2408 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1102
timestamp 1569543463
transform 1 0 2408 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1103
timestamp 1569543463
transform 1 0 2408 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1104
timestamp 1569543463
transform 1 0 2408 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1105
timestamp 1569543463
transform 1 0 2408 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1106
timestamp 1569543463
transform 1 0 2280 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1107
timestamp 1569543463
transform 1 0 2280 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1108
timestamp 1569543463
transform 1 0 2280 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1109
timestamp 1569543463
transform 1 0 2280 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1110
timestamp 1569543463
transform 1 0 2280 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1111
timestamp 1569543463
transform 1 0 1832 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1112
timestamp 1569543463
transform 1 0 1768 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1113
timestamp 1569543463
transform 1 0 1768 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1114
timestamp 1569543463
transform 1 0 1768 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1115
timestamp 1569543463
transform 1 0 1768 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1116
timestamp 1569543463
transform 1 0 1640 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1117
timestamp 1569543463
transform 1 0 1832 0 1 40
box -8 -8 8 8
use VIA2$5  VIA2$5_1118
timestamp 1569543463
transform 1 0 1832 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1119
timestamp 1569543463
transform 1 0 1832 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1120
timestamp 1569543463
transform 1 0 1768 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1121
timestamp 1569543463
transform 1 0 1832 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1122
timestamp 1569543463
transform 1 0 1704 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1123
timestamp 1569543463
transform 1 0 1704 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1124
timestamp 1569543463
transform 1 0 1640 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1125
timestamp 1569543463
transform 1 0 1640 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1126
timestamp 1569543463
transform 1 0 1704 0 1 104
box -8 -8 8 8
use VIA2$5  VIA2$5_1127
timestamp 1569543463
transform 1 0 1704 0 1 168
box -8 -8 8 8
use VIA2$5  VIA2$5_1128
timestamp 1569543463
transform 1 0 1512 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1129
timestamp 1569543463
transform 1 0 1320 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1130
timestamp 1569543463
transform 1 0 1320 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1131
timestamp 1569543463
transform 1 0 1320 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1132
timestamp 1569543463
transform 1 0 1512 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1133
timestamp 1569543463
transform 1 0 1512 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1134
timestamp 1569543463
transform 1 0 1448 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1135
timestamp 1569543463
transform 1 0 1448 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1136
timestamp 1569543463
transform 1 0 1384 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1137
timestamp 1569543463
transform 1 0 1384 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1138
timestamp 1569543463
transform 1 0 1384 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1139
timestamp 1569543463
transform 1 0 1384 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1140
timestamp 1569543463
transform 1 0 1512 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1141
timestamp 1569543463
transform 1 0 1512 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1142
timestamp 1569543463
transform 1 0 1448 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1143
timestamp 1569543463
transform 1 0 1512 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1144
timestamp 1569543463
transform 1 0 1448 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1145
timestamp 1569543463
transform 1 0 1448 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1146
timestamp 1569543463
transform 1 0 1640 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1147
timestamp 1569543463
transform 1 0 1640 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1148
timestamp 1569543463
transform 1 0 1704 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1149
timestamp 1569543463
transform 1 0 1704 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1150
timestamp 1569543463
transform 1 0 1832 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1151
timestamp 1569543463
transform 1 0 1832 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1152
timestamp 1569543463
transform 1 0 1832 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1153
timestamp 1569543463
transform 1 0 1832 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1154
timestamp 1569543463
transform 1 0 1832 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1155
timestamp 1569543463
transform 1 0 1768 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1156
timestamp 1569543463
transform 1 0 1768 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1157
timestamp 1569543463
transform 1 0 1768 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1158
timestamp 1569543463
transform 1 0 1704 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1159
timestamp 1569543463
transform 1 0 1640 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1160
timestamp 1569543463
transform 1 0 1640 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1161
timestamp 1569543463
transform 1 0 1640 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1162
timestamp 1569543463
transform 1 0 1704 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1163
timestamp 1569543463
transform 1 0 1704 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1164
timestamp 1569543463
transform 1 0 1768 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1165
timestamp 1569543463
transform 1 0 1768 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1166
timestamp 1569543463
transform 1 0 1576 0 1 296
box -8 -8 8 8
use VIA2$5  VIA2$5_1167
timestamp 1569543463
transform 1 0 1576 0 1 360
box -8 -8 8 8
use VIA2$5  VIA2$5_1168
timestamp 1569543463
transform 1 0 1576 0 1 424
box -8 -8 8 8
use VIA2$5  VIA2$5_1169
timestamp 1569543463
transform 1 0 1576 0 1 488
box -8 -8 8 8
use VIA2$5  VIA2$5_1170
timestamp 1569543463
transform 1 0 1576 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1171
timestamp 1569543463
transform 1 0 1576 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1172
timestamp 1569543463
transform 1 0 1576 0 1 232
box -8 -8 8 8
use VIA2$5  VIA2$5_1173
timestamp 1569543463
transform 1 0 1640 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1174
timestamp 1569543463
transform 1 0 1704 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1175
timestamp 1569543463
transform 1 0 1640 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1176
timestamp 1569543463
transform 1 0 1704 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1177
timestamp 1569543463
transform 1 0 1768 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1178
timestamp 1569543463
transform 1 0 1832 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1179
timestamp 1569543463
transform 1 0 1704 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1180
timestamp 1569543463
transform 1 0 1832 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1181
timestamp 1569543463
transform 1 0 1640 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1182
timestamp 1569543463
transform 1 0 1768 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1183
timestamp 1569543463
transform 1 0 1832 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1184
timestamp 1569543463
transform 1 0 1768 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1185
timestamp 1569543463
transform 1 0 1640 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1186
timestamp 1569543463
transform 1 0 1832 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1187
timestamp 1569543463
transform 1 0 1768 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1188
timestamp 1569543463
transform 1 0 1704 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1189
timestamp 1569543463
transform 1 0 1704 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1190
timestamp 1569543463
transform 1 0 1832 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1191
timestamp 1569543463
transform 1 0 1768 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1192
timestamp 1569543463
transform 1 0 1640 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1193
timestamp 1569543463
transform 1 0 1512 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1194
timestamp 1569543463
transform 1 0 1512 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1195
timestamp 1569543463
transform 1 0 1320 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1196
timestamp 1569543463
transform 1 0 1320 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1197
timestamp 1569543463
transform 1 0 1320 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1198
timestamp 1569543463
transform 1 0 1320 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1199
timestamp 1569543463
transform 1 0 1320 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1200
timestamp 1569543463
transform 1 0 1384 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1201
timestamp 1569543463
transform 1 0 1384 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1202
timestamp 1569543463
transform 1 0 1448 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1203
timestamp 1569543463
transform 1 0 1384 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1204
timestamp 1569543463
transform 1 0 1384 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1205
timestamp 1569543463
transform 1 0 1448 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1206
timestamp 1569543463
transform 1 0 1384 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1207
timestamp 1569543463
transform 1 0 1512 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1208
timestamp 1569543463
transform 1 0 1448 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1209
timestamp 1569543463
transform 1 0 1448 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1210
timestamp 1569543463
transform 1 0 1512 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1211
timestamp 1569543463
transform 1 0 1448 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1212
timestamp 1569543463
transform 1 0 1512 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1213
timestamp 1569543463
transform 1 0 1320 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1214
timestamp 1569543463
transform 1 0 1320 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1215
timestamp 1569543463
transform 1 0 1384 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1216
timestamp 1569543463
transform 1 0 1448 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1217
timestamp 1569543463
transform 1 0 1512 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1218
timestamp 1569543463
transform 1 0 1384 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1219
timestamp 1569543463
transform 1 0 1512 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1220
timestamp 1569543463
transform 1 0 1512 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1221
timestamp 1569543463
transform 1 0 1384 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1222
timestamp 1569543463
transform 1 0 1448 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1223
timestamp 1569543463
transform 1 0 1384 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1224
timestamp 1569543463
transform 1 0 1512 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1225
timestamp 1569543463
transform 1 0 1320 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1226
timestamp 1569543463
transform 1 0 1448 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1227
timestamp 1569543463
transform 1 0 1320 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1228
timestamp 1569543463
transform 1 0 1448 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1229
timestamp 1569543463
transform 1 0 1512 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1230
timestamp 1569543463
transform 1 0 1448 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1231
timestamp 1569543463
transform 1 0 1384 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1232
timestamp 1569543463
transform 1 0 1320 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1233
timestamp 1569543463
transform 1 0 1832 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1234
timestamp 1569543463
transform 1 0 1768 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1235
timestamp 1569543463
transform 1 0 1768 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1236
timestamp 1569543463
transform 1 0 1768 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1237
timestamp 1569543463
transform 1 0 1640 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1238
timestamp 1569543463
transform 1 0 1640 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1239
timestamp 1569543463
transform 1 0 1832 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1240
timestamp 1569543463
transform 1 0 1704 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1241
timestamp 1569543463
transform 1 0 1832 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1242
timestamp 1569543463
transform 1 0 1832 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1243
timestamp 1569543463
transform 1 0 1832 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1244
timestamp 1569543463
transform 1 0 1704 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1245
timestamp 1569543463
transform 1 0 1768 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1246
timestamp 1569543463
transform 1 0 1768 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1247
timestamp 1569543463
transform 1 0 1640 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1248
timestamp 1569543463
transform 1 0 1640 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1249
timestamp 1569543463
transform 1 0 1704 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1250
timestamp 1569543463
transform 1 0 1704 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1251
timestamp 1569543463
transform 1 0 1704 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1252
timestamp 1569543463
transform 1 0 1640 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1253
timestamp 1569543463
transform 1 0 1576 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1254
timestamp 1569543463
transform 1 0 1576 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1255
timestamp 1569543463
transform 1 0 1576 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1256
timestamp 1569543463
transform 1 0 1576 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1257
timestamp 1569543463
transform 1 0 1576 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1258
timestamp 1569543463
transform 1 0 1576 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1259
timestamp 1569543463
transform 1 0 1576 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1260
timestamp 1569543463
transform 1 0 1576 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1261
timestamp 1569543463
transform 1 0 1576 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1262
timestamp 1569543463
transform 1 0 1576 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1263
timestamp 1569543463
transform 1 0 2280 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1264
timestamp 1569543463
transform 1 0 2344 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1265
timestamp 1569543463
transform 1 0 2472 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1266
timestamp 1569543463
transform 1 0 2472 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1267
timestamp 1569543463
transform 1 0 2472 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1268
timestamp 1569543463
transform 1 0 2344 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1269
timestamp 1569543463
transform 1 0 2216 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1270
timestamp 1569543463
transform 1 0 2216 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1271
timestamp 1569543463
transform 1 0 2216 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1272
timestamp 1569543463
transform 1 0 2408 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1273
timestamp 1569543463
transform 1 0 2216 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1274
timestamp 1569543463
transform 1 0 2216 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1275
timestamp 1569543463
transform 1 0 2408 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1276
timestamp 1569543463
transform 1 0 2472 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1277
timestamp 1569543463
transform 1 0 2344 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1278
timestamp 1569543463
transform 1 0 2408 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1279
timestamp 1569543463
transform 1 0 2344 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1280
timestamp 1569543463
transform 1 0 2344 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1281
timestamp 1569543463
transform 1 0 2408 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1282
timestamp 1569543463
transform 1 0 2408 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1283
timestamp 1569543463
transform 1 0 2472 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1284
timestamp 1569543463
transform 1 0 2280 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1285
timestamp 1569543463
transform 1 0 2280 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1286
timestamp 1569543463
transform 1 0 2280 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1287
timestamp 1569543463
transform 1 0 2280 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1288
timestamp 1569543463
transform 1 0 1896 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1289
timestamp 1569543463
transform 1 0 1896 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1290
timestamp 1569543463
transform 1 0 1896 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1291
timestamp 1569543463
transform 1 0 1896 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1292
timestamp 1569543463
transform 1 0 2152 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1293
timestamp 1569543463
transform 1 0 1896 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1294
timestamp 1569543463
transform 1 0 1960 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1295
timestamp 1569543463
transform 1 0 1960 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1296
timestamp 1569543463
transform 1 0 1960 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1297
timestamp 1569543463
transform 1 0 1960 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1298
timestamp 1569543463
transform 1 0 1960 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1299
timestamp 1569543463
transform 1 0 2024 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1300
timestamp 1569543463
transform 1 0 2024 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1301
timestamp 1569543463
transform 1 0 2024 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1302
timestamp 1569543463
transform 1 0 2024 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1303
timestamp 1569543463
transform 1 0 2024 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1304
timestamp 1569543463
transform 1 0 2088 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1305
timestamp 1569543463
transform 1 0 2088 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1306
timestamp 1569543463
transform 1 0 2088 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1307
timestamp 1569543463
transform 1 0 2088 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1308
timestamp 1569543463
transform 1 0 2088 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1309
timestamp 1569543463
transform 1 0 2152 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1310
timestamp 1569543463
transform 1 0 2152 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1311
timestamp 1569543463
transform 1 0 2152 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1312
timestamp 1569543463
transform 1 0 2152 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1313
timestamp 1569543463
transform 1 0 2152 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1314
timestamp 1569543463
transform 1 0 1960 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1315
timestamp 1569543463
transform 1 0 2024 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1316
timestamp 1569543463
transform 1 0 2024 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1317
timestamp 1569543463
transform 1 0 1896 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1318
timestamp 1569543463
transform 1 0 2088 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1319
timestamp 1569543463
transform 1 0 2088 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1320
timestamp 1569543463
transform 1 0 2152 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1321
timestamp 1569543463
transform 1 0 1896 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1322
timestamp 1569543463
transform 1 0 2088 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1323
timestamp 1569543463
transform 1 0 2024 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1324
timestamp 1569543463
transform 1 0 2152 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1325
timestamp 1569543463
transform 1 0 2088 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1326
timestamp 1569543463
transform 1 0 2088 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1327
timestamp 1569543463
transform 1 0 2024 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1328
timestamp 1569543463
transform 1 0 2024 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1329
timestamp 1569543463
transform 1 0 1896 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1330
timestamp 1569543463
transform 1 0 2152 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1331
timestamp 1569543463
transform 1 0 1896 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1332
timestamp 1569543463
transform 1 0 2152 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1333
timestamp 1569543463
transform 1 0 1896 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1334
timestamp 1569543463
transform 1 0 1960 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1335
timestamp 1569543463
transform 1 0 1960 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1336
timestamp 1569543463
transform 1 0 1960 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1337
timestamp 1569543463
transform 1 0 1960 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1338
timestamp 1569543463
transform 1 0 2280 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1339
timestamp 1569543463
transform 1 0 2280 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1340
timestamp 1569543463
transform 1 0 2280 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1341
timestamp 1569543463
transform 1 0 2408 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1342
timestamp 1569543463
transform 1 0 2408 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1343
timestamp 1569543463
transform 1 0 2344 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1344
timestamp 1569543463
transform 1 0 2344 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1345
timestamp 1569543463
transform 1 0 2344 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1346
timestamp 1569543463
transform 1 0 2408 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1347
timestamp 1569543463
transform 1 0 2408 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1348
timestamp 1569543463
transform 1 0 2408 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1349
timestamp 1569543463
transform 1 0 2472 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1350
timestamp 1569543463
transform 1 0 2216 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1351
timestamp 1569543463
transform 1 0 2472 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1352
timestamp 1569543463
transform 1 0 2216 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1353
timestamp 1569543463
transform 1 0 2472 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1354
timestamp 1569543463
transform 1 0 2216 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1355
timestamp 1569543463
transform 1 0 2472 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1356
timestamp 1569543463
transform 1 0 2216 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1357
timestamp 1569543463
transform 1 0 2472 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1358
timestamp 1569543463
transform 1 0 2216 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1359
timestamp 1569543463
transform 1 0 2344 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1360
timestamp 1569543463
transform 1 0 2344 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1361
timestamp 1569543463
transform 1 0 2280 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1362
timestamp 1569543463
transform 1 0 2280 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1363
timestamp 1569543463
transform 1 0 1192 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1364
timestamp 1569543463
transform 1 0 1256 0 1 552
box -8 -8 8 8
use VIA2$5  VIA2$5_1365
timestamp 1569543463
transform 1 0 1256 0 1 616
box -8 -8 8 8
use VIA2$5  VIA2$5_1366
timestamp 1569543463
transform 1 0 616 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1367
timestamp 1569543463
transform 1 0 552 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1368
timestamp 1569543463
transform 1 0 616 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1369
timestamp 1569543463
transform 1 0 1256 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1370
timestamp 1569543463
transform 1 0 1256 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1371
timestamp 1569543463
transform 1 0 1256 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1372
timestamp 1569543463
transform 1 0 1256 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1373
timestamp 1569543463
transform 1 0 1256 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1374
timestamp 1569543463
transform 1 0 1064 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1375
timestamp 1569543463
transform 1 0 1064 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1376
timestamp 1569543463
transform 1 0 1192 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1377
timestamp 1569543463
transform 1 0 1192 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1378
timestamp 1569543463
transform 1 0 1192 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1379
timestamp 1569543463
transform 1 0 1192 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1380
timestamp 1569543463
transform 1 0 1064 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1381
timestamp 1569543463
transform 1 0 1128 0 1 744
box -8 -8 8 8
use VIA2$5  VIA2$5_1382
timestamp 1569543463
transform 1 0 1128 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1383
timestamp 1569543463
transform 1 0 1128 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1384
timestamp 1569543463
transform 1 0 1128 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1385
timestamp 1569543463
transform 1 0 1128 0 1 680
box -8 -8 8 8
use VIA2$5  VIA2$5_1386
timestamp 1569543463
transform 1 0 1064 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1387
timestamp 1569543463
transform 1 0 1000 0 1 808
box -8 -8 8 8
use VIA2$5  VIA2$5_1388
timestamp 1569543463
transform 1 0 1192 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1389
timestamp 1569543463
transform 1 0 1000 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1390
timestamp 1569543463
transform 1 0 1000 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1391
timestamp 1569543463
transform 1 0 936 0 1 872
box -8 -8 8 8
use VIA2$5  VIA2$5_1392
timestamp 1569543463
transform 1 0 936 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1393
timestamp 1569543463
transform 1 0 872 0 1 936
box -8 -8 8 8
use VIA2$5  VIA2$5_1394
timestamp 1569543463
transform 1 0 872 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1395
timestamp 1569543463
transform 1 0 744 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1396
timestamp 1569543463
transform 1 0 744 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1397
timestamp 1569543463
transform 1 0 872 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1398
timestamp 1569543463
transform 1 0 808 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1399
timestamp 1569543463
transform 1 0 872 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1400
timestamp 1569543463
transform 1 0 808 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1401
timestamp 1569543463
transform 1 0 936 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1402
timestamp 1569543463
transform 1 0 808 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1403
timestamp 1569543463
transform 1 0 680 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1404
timestamp 1569543463
transform 1 0 744 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1405
timestamp 1569543463
transform 1 0 936 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1406
timestamp 1569543463
transform 1 0 936 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1407
timestamp 1569543463
transform 1 0 808 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1408
timestamp 1569543463
transform 1 0 680 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1409
timestamp 1569543463
transform 1 0 744 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1410
timestamp 1569543463
transform 1 0 808 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1411
timestamp 1569543463
transform 1 0 936 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1412
timestamp 1569543463
transform 1 0 680 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1413
timestamp 1569543463
transform 1 0 872 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1414
timestamp 1569543463
transform 1 0 936 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1415
timestamp 1569543463
transform 1 0 872 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1416
timestamp 1569543463
transform 1 0 1128 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1417
timestamp 1569543463
transform 1 0 1000 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1418
timestamp 1569543463
transform 1 0 1256 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1419
timestamp 1569543463
transform 1 0 1000 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1420
timestamp 1569543463
transform 1 0 1256 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1421
timestamp 1569543463
transform 1 0 1128 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1422
timestamp 1569543463
transform 1 0 1000 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1423
timestamp 1569543463
transform 1 0 1064 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1424
timestamp 1569543463
transform 1 0 1064 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1425
timestamp 1569543463
transform 1 0 1256 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1426
timestamp 1569543463
transform 1 0 1064 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1427
timestamp 1569543463
transform 1 0 1064 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1428
timestamp 1569543463
transform 1 0 1128 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1429
timestamp 1569543463
transform 1 0 1128 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1430
timestamp 1569543463
transform 1 0 1064 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1431
timestamp 1569543463
transform 1 0 1192 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1432
timestamp 1569543463
transform 1 0 1192 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1433
timestamp 1569543463
transform 1 0 1192 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1434
timestamp 1569543463
transform 1 0 1192 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1435
timestamp 1569543463
transform 1 0 1192 0 1 1000
box -8 -8 8 8
use VIA2$5  VIA2$5_1436
timestamp 1569543463
transform 1 0 1128 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1437
timestamp 1569543463
transform 1 0 1256 0 1 1064
box -8 -8 8 8
use VIA2$5  VIA2$5_1438
timestamp 1569543463
transform 1 0 1000 0 1 1128
box -8 -8 8 8
use VIA2$5  VIA2$5_1439
timestamp 1569543463
transform 1 0 1256 0 1 1192
box -8 -8 8 8
use VIA2$5  VIA2$5_1440
timestamp 1569543463
transform 1 0 1000 0 1 1256
box -8 -8 8 8
use VIA2$5  VIA2$5_1441
timestamp 1569543463
transform 1 0 1000 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1442
timestamp 1569543463
transform 1 0 1256 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1443
timestamp 1569543463
transform 1 0 1128 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1444
timestamp 1569543463
transform 1 0 1064 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1445
timestamp 1569543463
transform 1 0 1000 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1446
timestamp 1569543463
transform 1 0 1256 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1447
timestamp 1569543463
transform 1 0 1000 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1448
timestamp 1569543463
transform 1 0 1192 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1449
timestamp 1569543463
transform 1 0 1064 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1450
timestamp 1569543463
transform 1 0 1064 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1451
timestamp 1569543463
transform 1 0 1192 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1452
timestamp 1569543463
transform 1 0 1192 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1453
timestamp 1569543463
transform 1 0 1128 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1454
timestamp 1569543463
transform 1 0 1064 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1455
timestamp 1569543463
transform 1 0 1256 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1456
timestamp 1569543463
transform 1 0 1256 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1457
timestamp 1569543463
transform 1 0 1192 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1458
timestamp 1569543463
transform 1 0 1000 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1459
timestamp 1569543463
transform 1 0 1128 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1460
timestamp 1569543463
transform 1 0 1128 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1461
timestamp 1569543463
transform 1 0 744 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1462
timestamp 1569543463
transform 1 0 680 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1463
timestamp 1569543463
transform 1 0 936 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1464
timestamp 1569543463
transform 1 0 744 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1465
timestamp 1569543463
transform 1 0 680 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1466
timestamp 1569543463
transform 1 0 936 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1467
timestamp 1569543463
transform 1 0 808 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1468
timestamp 1569543463
transform 1 0 936 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1469
timestamp 1569543463
transform 1 0 872 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1470
timestamp 1569543463
transform 1 0 808 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1471
timestamp 1569543463
transform 1 0 744 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1472
timestamp 1569543463
transform 1 0 872 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1473
timestamp 1569543463
transform 1 0 872 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1474
timestamp 1569543463
transform 1 0 808 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1475
timestamp 1569543463
transform 1 0 936 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1476
timestamp 1569543463
transform 1 0 680 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1477
timestamp 1569543463
transform 1 0 872 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1478
timestamp 1569543463
transform 1 0 808 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1479
timestamp 1569543463
transform 1 0 680 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1480
timestamp 1569543463
transform 1 0 744 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1481
timestamp 1569543463
transform 1 0 808 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1482
timestamp 1569543463
transform 1 0 936 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1483
timestamp 1569543463
transform 1 0 872 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1484
timestamp 1569543463
transform 1 0 808 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1485
timestamp 1569543463
transform 1 0 808 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1486
timestamp 1569543463
transform 1 0 936 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1487
timestamp 1569543463
transform 1 0 936 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1488
timestamp 1569543463
transform 1 0 872 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1489
timestamp 1569543463
transform 1 0 680 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1490
timestamp 1569543463
transform 1 0 744 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1491
timestamp 1569543463
transform 1 0 680 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1492
timestamp 1569543463
transform 1 0 680 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1493
timestamp 1569543463
transform 1 0 872 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1494
timestamp 1569543463
transform 1 0 744 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1495
timestamp 1569543463
transform 1 0 744 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1496
timestamp 1569543463
transform 1 0 808 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1497
timestamp 1569543463
transform 1 0 936 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1498
timestamp 1569543463
transform 1 0 744 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1499
timestamp 1569543463
transform 1 0 680 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1500
timestamp 1569543463
transform 1 0 872 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1501
timestamp 1569543463
transform 1 0 1000 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1502
timestamp 1569543463
transform 1 0 1256 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1503
timestamp 1569543463
transform 1 0 1128 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1504
timestamp 1569543463
transform 1 0 1064 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1505
timestamp 1569543463
transform 1 0 1256 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1506
timestamp 1569543463
transform 1 0 1256 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1507
timestamp 1569543463
transform 1 0 1000 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1508
timestamp 1569543463
transform 1 0 1128 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1509
timestamp 1569543463
transform 1 0 1192 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1510
timestamp 1569543463
transform 1 0 1192 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1511
timestamp 1569543463
transform 1 0 1000 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1512
timestamp 1569543463
transform 1 0 1000 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1513
timestamp 1569543463
transform 1 0 1256 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1514
timestamp 1569543463
transform 1 0 1064 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1515
timestamp 1569543463
transform 1 0 1064 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1516
timestamp 1569543463
transform 1 0 1064 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1517
timestamp 1569543463
transform 1 0 1128 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1518
timestamp 1569543463
transform 1 0 1128 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1519
timestamp 1569543463
transform 1 0 1192 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1520
timestamp 1569543463
transform 1 0 1192 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1521
timestamp 1569543463
transform 1 0 872 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1522
timestamp 1569543463
transform 1 0 1128 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1523
timestamp 1569543463
transform 1 0 936 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1524
timestamp 1569543463
transform 1 0 808 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1525
timestamp 1569543463
transform 1 0 1064 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1526
timestamp 1569543463
transform 1 0 680 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1527
timestamp 1569543463
transform 1 0 1000 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1528
timestamp 1569543463
transform 1 0 1192 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1529
timestamp 1569543463
transform 1 0 1256 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1530
timestamp 1569543463
transform 1 0 744 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1531
timestamp 1569543463
transform 1 0 488 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1532
timestamp 1569543463
transform 1 0 488 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1533
timestamp 1569543463
transform 1 0 424 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1534
timestamp 1569543463
transform 1 0 616 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1535
timestamp 1569543463
transform 1 0 552 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1536
timestamp 1569543463
transform 1 0 616 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1537
timestamp 1569543463
transform 1 0 552 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1538
timestamp 1569543463
transform 1 0 424 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1539
timestamp 1569543463
transform 1 0 616 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1540
timestamp 1569543463
transform 1 0 552 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1541
timestamp 1569543463
transform 1 0 616 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1542
timestamp 1569543463
transform 1 0 360 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1543
timestamp 1569543463
transform 1 0 488 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1544
timestamp 1569543463
transform 1 0 360 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1545
timestamp 1569543463
transform 1 0 488 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1546
timestamp 1569543463
transform 1 0 424 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1547
timestamp 1569543463
transform 1 0 552 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1548
timestamp 1569543463
transform 1 0 296 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1549
timestamp 1569543463
transform 1 0 40 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1550
timestamp 1569543463
transform 1 0 296 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1551
timestamp 1569543463
transform 1 0 40 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1552
timestamp 1569543463
transform 1 0 232 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1553
timestamp 1569543463
transform 1 0 168 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1554
timestamp 1569543463
transform 1 0 232 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1555
timestamp 1569543463
transform 1 0 232 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1556
timestamp 1569543463
transform 1 0 104 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1557
timestamp 1569543463
transform 1 0 296 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1558
timestamp 1569543463
transform 1 0 296 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1559
timestamp 1569543463
transform 1 0 168 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1560
timestamp 1569543463
transform 1 0 296 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1561
timestamp 1569543463
transform 1 0 168 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1562
timestamp 1569543463
transform 1 0 104 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1563
timestamp 1569543463
transform 1 0 168 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1564
timestamp 1569543463
transform 1 0 232 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1565
timestamp 1569543463
transform 1 0 104 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1566
timestamp 1569543463
transform 1 0 360 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1567
timestamp 1569543463
transform 1 0 360 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1568
timestamp 1569543463
transform 1 0 616 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1569
timestamp 1569543463
transform 1 0 552 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1570
timestamp 1569543463
transform 1 0 424 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1571
timestamp 1569543463
transform 1 0 360 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1572
timestamp 1569543463
transform 1 0 616 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1573
timestamp 1569543463
transform 1 0 424 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1574
timestamp 1569543463
transform 1 0 488 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1575
timestamp 1569543463
transform 1 0 552 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1576
timestamp 1569543463
transform 1 0 424 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1577
timestamp 1569543463
transform 1 0 424 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1578
timestamp 1569543463
transform 1 0 488 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1579
timestamp 1569543463
transform 1 0 488 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1580
timestamp 1569543463
transform 1 0 360 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1581
timestamp 1569543463
transform 1 0 552 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1582
timestamp 1569543463
transform 1 0 552 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1583
timestamp 1569543463
transform 1 0 488 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1584
timestamp 1569543463
transform 1 0 616 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1585
timestamp 1569543463
transform 1 0 616 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1586
timestamp 1569543463
transform 1 0 488 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1587
timestamp 1569543463
transform 1 0 552 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1588
timestamp 1569543463
transform 1 0 616 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1589
timestamp 1569543463
transform 1 0 232 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1590
timestamp 1569543463
transform 1 0 296 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1591
timestamp 1569543463
transform 1 0 424 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1592
timestamp 1569543463
transform 1 0 360 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1593
timestamp 1569543463
transform 1 0 552 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1594
timestamp 1569543463
transform 1 0 488 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1595
timestamp 1569543463
transform 1 0 424 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1596
timestamp 1569543463
transform 1 0 552 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1597
timestamp 1569543463
transform 1 0 360 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1598
timestamp 1569543463
transform 1 0 616 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1599
timestamp 1569543463
transform 1 0 488 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1600
timestamp 1569543463
transform 1 0 424 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1601
timestamp 1569543463
transform 1 0 360 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1602
timestamp 1569543463
transform 1 0 488 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1603
timestamp 1569543463
transform 1 0 616 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1604
timestamp 1569543463
transform 1 0 360 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1605
timestamp 1569543463
transform 1 0 616 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1606
timestamp 1569543463
transform 1 0 552 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1607
timestamp 1569543463
transform 1 0 424 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1608
timestamp 1569543463
transform 1 0 488 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1609
timestamp 1569543463
transform 1 0 424 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1610
timestamp 1569543463
transform 1 0 488 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1611
timestamp 1569543463
transform 1 0 552 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1612
timestamp 1569543463
transform 1 0 552 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1613
timestamp 1569543463
transform 1 0 360 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1614
timestamp 1569543463
transform 1 0 360 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1615
timestamp 1569543463
transform 1 0 616 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1616
timestamp 1569543463
transform 1 0 424 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1617
timestamp 1569543463
transform 1 0 616 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1618
timestamp 1569543463
transform 1 0 40 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1619
timestamp 1569543463
transform 1 0 168 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1620
timestamp 1569543463
transform 1 0 296 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1621
timestamp 1569543463
transform 1 0 40 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1622
timestamp 1569543463
transform 1 0 232 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1623
timestamp 1569543463
transform 1 0 296 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1624
timestamp 1569543463
transform 1 0 168 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1625
timestamp 1569543463
transform 1 0 296 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1626
timestamp 1569543463
transform 1 0 104 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1627
timestamp 1569543463
transform 1 0 168 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1628
timestamp 1569543463
transform 1 0 168 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1629
timestamp 1569543463
transform 1 0 40 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1630
timestamp 1569543463
transform 1 0 296 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1631
timestamp 1569543463
transform 1 0 168 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1632
timestamp 1569543463
transform 1 0 104 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1633
timestamp 1569543463
transform 1 0 232 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1634
timestamp 1569543463
transform 1 0 104 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1635
timestamp 1569543463
transform 1 0 232 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1636
timestamp 1569543463
transform 1 0 40 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1637
timestamp 1569543463
transform 1 0 296 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1638
timestamp 1569543463
transform 1 0 232 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1639
timestamp 1569543463
transform 1 0 104 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1640
timestamp 1569543463
transform 1 0 232 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1641
timestamp 1569543463
transform 1 0 40 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1642
timestamp 1569543463
transform 1 0 104 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1643
timestamp 1569543463
transform 1 0 296 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1644
timestamp 1569543463
transform 1 0 40 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1645
timestamp 1569543463
transform 1 0 296 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1646
timestamp 1569543463
transform 1 0 296 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1647
timestamp 1569543463
transform 1 0 40 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1648
timestamp 1569543463
transform 1 0 168 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1649
timestamp 1569543463
transform 1 0 232 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1650
timestamp 1569543463
transform 1 0 40 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1651
timestamp 1569543463
transform 1 0 168 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1652
timestamp 1569543463
transform 1 0 104 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1653
timestamp 1569543463
transform 1 0 40 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1654
timestamp 1569543463
transform 1 0 232 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1655
timestamp 1569543463
transform 1 0 104 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1656
timestamp 1569543463
transform 1 0 168 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1657
timestamp 1569543463
transform 1 0 232 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1658
timestamp 1569543463
transform 1 0 40 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1659
timestamp 1569543463
transform 1 0 104 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1660
timestamp 1569543463
transform 1 0 104 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1661
timestamp 1569543463
transform 1 0 296 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1662
timestamp 1569543463
transform 1 0 104 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1663
timestamp 1569543463
transform 1 0 168 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1664
timestamp 1569543463
transform 1 0 232 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1665
timestamp 1569543463
transform 1 0 168 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1666
timestamp 1569543463
transform 1 0 296 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1667
timestamp 1569543463
transform 1 0 232 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1668
timestamp 1569543463
transform 1 0 424 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1669
timestamp 1569543463
transform 1 0 488 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1670
timestamp 1569543463
transform 1 0 424 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1671
timestamp 1569543463
transform 1 0 424 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1672
timestamp 1569543463
transform 1 0 488 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1673
timestamp 1569543463
transform 1 0 616 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1674
timestamp 1569543463
transform 1 0 424 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1675
timestamp 1569543463
transform 1 0 360 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1676
timestamp 1569543463
transform 1 0 616 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1677
timestamp 1569543463
transform 1 0 552 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1678
timestamp 1569543463
transform 1 0 552 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1679
timestamp 1569543463
transform 1 0 616 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1680
timestamp 1569543463
transform 1 0 552 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1681
timestamp 1569543463
transform 1 0 552 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1682
timestamp 1569543463
transform 1 0 488 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1683
timestamp 1569543463
transform 1 0 360 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1684
timestamp 1569543463
transform 1 0 552 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1685
timestamp 1569543463
transform 1 0 616 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1686
timestamp 1569543463
transform 1 0 488 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1687
timestamp 1569543463
transform 1 0 360 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1688
timestamp 1569543463
transform 1 0 616 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1689
timestamp 1569543463
transform 1 0 360 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1690
timestamp 1569543463
transform 1 0 424 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1691
timestamp 1569543463
transform 1 0 360 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1692
timestamp 1569543463
transform 1 0 488 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1693
timestamp 1569543463
transform 1 0 1192 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1694
timestamp 1569543463
transform 1 0 1192 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1695
timestamp 1569543463
transform 1 0 1256 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1696
timestamp 1569543463
transform 1 0 1128 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1697
timestamp 1569543463
transform 1 0 1064 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1698
timestamp 1569543463
transform 1 0 1128 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1699
timestamp 1569543463
transform 1 0 1192 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1700
timestamp 1569543463
transform 1 0 1128 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1701
timestamp 1569543463
transform 1 0 1192 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1702
timestamp 1569543463
transform 1 0 1128 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1703
timestamp 1569543463
transform 1 0 1256 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1704
timestamp 1569543463
transform 1 0 1064 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1705
timestamp 1569543463
transform 1 0 1000 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1706
timestamp 1569543463
transform 1 0 1256 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1707
timestamp 1569543463
transform 1 0 1000 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1708
timestamp 1569543463
transform 1 0 1256 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1709
timestamp 1569543463
transform 1 0 1000 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1710
timestamp 1569543463
transform 1 0 1256 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1711
timestamp 1569543463
transform 1 0 1128 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1712
timestamp 1569543463
transform 1 0 1000 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1713
timestamp 1569543463
transform 1 0 1064 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1714
timestamp 1569543463
transform 1 0 1064 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1715
timestamp 1569543463
transform 1 0 1192 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1716
timestamp 1569543463
transform 1 0 1064 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1717
timestamp 1569543463
transform 1 0 1000 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1718
timestamp 1569543463
transform 1 0 808 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1719
timestamp 1569543463
transform 1 0 680 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1720
timestamp 1569543463
transform 1 0 872 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1721
timestamp 1569543463
transform 1 0 936 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1722
timestamp 1569543463
transform 1 0 872 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1723
timestamp 1569543463
transform 1 0 936 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1724
timestamp 1569543463
transform 1 0 744 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1725
timestamp 1569543463
transform 1 0 744 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1726
timestamp 1569543463
transform 1 0 744 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1727
timestamp 1569543463
transform 1 0 872 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1728
timestamp 1569543463
transform 1 0 744 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1729
timestamp 1569543463
transform 1 0 744 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1730
timestamp 1569543463
transform 1 0 680 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1731
timestamp 1569543463
transform 1 0 808 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1732
timestamp 1569543463
transform 1 0 808 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1733
timestamp 1569543463
transform 1 0 808 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1734
timestamp 1569543463
transform 1 0 808 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1735
timestamp 1569543463
transform 1 0 872 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1736
timestamp 1569543463
transform 1 0 680 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1737
timestamp 1569543463
transform 1 0 680 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1738
timestamp 1569543463
transform 1 0 936 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1739
timestamp 1569543463
transform 1 0 872 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1740
timestamp 1569543463
transform 1 0 936 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1741
timestamp 1569543463
transform 1 0 680 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1742
timestamp 1569543463
transform 1 0 936 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1743
timestamp 1569543463
transform 1 0 936 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1744
timestamp 1569543463
transform 1 0 936 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1745
timestamp 1569543463
transform 1 0 808 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1746
timestamp 1569543463
transform 1 0 680 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1747
timestamp 1569543463
transform 1 0 680 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1748
timestamp 1569543463
transform 1 0 680 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1749
timestamp 1569543463
transform 1 0 872 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1750
timestamp 1569543463
transform 1 0 680 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1751
timestamp 1569543463
transform 1 0 808 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1752
timestamp 1569543463
transform 1 0 744 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1753
timestamp 1569543463
transform 1 0 872 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1754
timestamp 1569543463
transform 1 0 808 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1755
timestamp 1569543463
transform 1 0 872 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1756
timestamp 1569543463
transform 1 0 872 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1757
timestamp 1569543463
transform 1 0 872 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1758
timestamp 1569543463
transform 1 0 936 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1759
timestamp 1569543463
transform 1 0 744 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1760
timestamp 1569543463
transform 1 0 744 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1761
timestamp 1569543463
transform 1 0 936 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1762
timestamp 1569543463
transform 1 0 744 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1763
timestamp 1569543463
transform 1 0 936 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1764
timestamp 1569543463
transform 1 0 808 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1765
timestamp 1569543463
transform 1 0 680 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1766
timestamp 1569543463
transform 1 0 744 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1767
timestamp 1569543463
transform 1 0 808 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1768
timestamp 1569543463
transform 1 0 1064 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1769
timestamp 1569543463
transform 1 0 1064 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1770
timestamp 1569543463
transform 1 0 1128 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1771
timestamp 1569543463
transform 1 0 1000 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1772
timestamp 1569543463
transform 1 0 1192 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1773
timestamp 1569543463
transform 1 0 1192 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1774
timestamp 1569543463
transform 1 0 1192 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1775
timestamp 1569543463
transform 1 0 1192 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1776
timestamp 1569543463
transform 1 0 1192 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1777
timestamp 1569543463
transform 1 0 1064 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1778
timestamp 1569543463
transform 1 0 1000 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1779
timestamp 1569543463
transform 1 0 1064 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1780
timestamp 1569543463
transform 1 0 1000 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1781
timestamp 1569543463
transform 1 0 1064 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1782
timestamp 1569543463
transform 1 0 1128 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1783
timestamp 1569543463
transform 1 0 1000 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1784
timestamp 1569543463
transform 1 0 1128 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1785
timestamp 1569543463
transform 1 0 1000 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1786
timestamp 1569543463
transform 1 0 1256 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1787
timestamp 1569543463
transform 1 0 1256 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1788
timestamp 1569543463
transform 1 0 1256 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_1789
timestamp 1569543463
transform 1 0 1128 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_1790
timestamp 1569543463
transform 1 0 1256 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_1791
timestamp 1569543463
transform 1 0 1256 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_1792
timestamp 1569543463
transform 1 0 1128 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_1793
timestamp 1569543463
transform 1 0 2280 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1794
timestamp 1569543463
transform 1 0 2280 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1795
timestamp 1569543463
transform 1 0 2472 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1796
timestamp 1569543463
transform 1 0 2344 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1797
timestamp 1569543463
transform 1 0 2216 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1798
timestamp 1569543463
transform 1 0 2472 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1799
timestamp 1569543463
transform 1 0 2344 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1800
timestamp 1569543463
transform 1 0 2216 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1801
timestamp 1569543463
transform 1 0 2408 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1802
timestamp 1569543463
transform 1 0 2408 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1803
timestamp 1569543463
transform 1 0 2408 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1804
timestamp 1569543463
transform 1 0 2344 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1805
timestamp 1569543463
transform 1 0 2344 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1806
timestamp 1569543463
transform 1 0 2408 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1807
timestamp 1569543463
transform 1 0 2216 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1808
timestamp 1569543463
transform 1 0 2280 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1809
timestamp 1569543463
transform 1 0 2472 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1810
timestamp 1569543463
transform 1 0 2216 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1811
timestamp 1569543463
transform 1 0 2472 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1812
timestamp 1569543463
transform 1 0 2280 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1813
timestamp 1569543463
transform 1 0 2024 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1814
timestamp 1569543463
transform 1 0 1896 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1815
timestamp 1569543463
transform 1 0 2024 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1816
timestamp 1569543463
transform 1 0 2088 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1817
timestamp 1569543463
transform 1 0 2088 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1818
timestamp 1569543463
transform 1 0 2024 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1819
timestamp 1569543463
transform 1 0 2088 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1820
timestamp 1569543463
transform 1 0 2152 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1821
timestamp 1569543463
transform 1 0 1896 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1822
timestamp 1569543463
transform 1 0 1896 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1823
timestamp 1569543463
transform 1 0 2152 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1824
timestamp 1569543463
transform 1 0 1896 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1825
timestamp 1569543463
transform 1 0 1960 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1826
timestamp 1569543463
transform 1 0 1960 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1827
timestamp 1569543463
transform 1 0 1960 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1828
timestamp 1569543463
transform 1 0 2152 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1829
timestamp 1569543463
transform 1 0 1960 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1830
timestamp 1569543463
transform 1 0 2088 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1831
timestamp 1569543463
transform 1 0 2024 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1832
timestamp 1569543463
transform 1 0 2152 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1833
timestamp 1569543463
transform 1 0 1896 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1834
timestamp 1569543463
transform 1 0 2024 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1835
timestamp 1569543463
transform 1 0 2088 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1836
timestamp 1569543463
transform 1 0 2024 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1837
timestamp 1569543463
transform 1 0 2152 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1838
timestamp 1569543463
transform 1 0 2152 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1839
timestamp 1569543463
transform 1 0 1896 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1840
timestamp 1569543463
transform 1 0 1960 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1841
timestamp 1569543463
transform 1 0 1960 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1842
timestamp 1569543463
transform 1 0 1960 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1843
timestamp 1569543463
transform 1 0 2024 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1844
timestamp 1569543463
transform 1 0 2024 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1845
timestamp 1569543463
transform 1 0 1896 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1846
timestamp 1569543463
transform 1 0 2088 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1847
timestamp 1569543463
transform 1 0 2088 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1848
timestamp 1569543463
transform 1 0 1960 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1849
timestamp 1569543463
transform 1 0 2152 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1850
timestamp 1569543463
transform 1 0 2152 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1851
timestamp 1569543463
transform 1 0 2088 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1852
timestamp 1569543463
transform 1 0 1896 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1853
timestamp 1569543463
transform 1 0 2344 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1854
timestamp 1569543463
transform 1 0 2280 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1855
timestamp 1569543463
transform 1 0 2344 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1856
timestamp 1569543463
transform 1 0 2408 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1857
timestamp 1569543463
transform 1 0 2408 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1858
timestamp 1569543463
transform 1 0 2472 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1859
timestamp 1569543463
transform 1 0 2472 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1860
timestamp 1569543463
transform 1 0 2344 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1861
timestamp 1569543463
transform 1 0 2344 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1862
timestamp 1569543463
transform 1 0 2408 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1863
timestamp 1569543463
transform 1 0 2408 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1864
timestamp 1569543463
transform 1 0 2280 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1865
timestamp 1569543463
transform 1 0 2472 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1866
timestamp 1569543463
transform 1 0 2472 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1867
timestamp 1569543463
transform 1 0 2216 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1868
timestamp 1569543463
transform 1 0 2280 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1869
timestamp 1569543463
transform 1 0 2280 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1870
timestamp 1569543463
transform 1 0 2216 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1871
timestamp 1569543463
transform 1 0 2216 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1872
timestamp 1569543463
transform 1 0 2216 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1873
timestamp 1569543463
transform 1 0 1896 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1874
timestamp 1569543463
transform 1 0 2344 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1875
timestamp 1569543463
transform 1 0 2408 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1876
timestamp 1569543463
transform 1 0 1960 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1877
timestamp 1569543463
transform 1 0 2472 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1878
timestamp 1569543463
transform 1 0 2024 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1879
timestamp 1569543463
transform 1 0 2088 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1880
timestamp 1569543463
transform 1 0 2152 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1881
timestamp 1569543463
transform 1 0 2216 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1882
timestamp 1569543463
transform 1 0 2280 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1883
timestamp 1569543463
transform 1 0 1768 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1884
timestamp 1569543463
transform 1 0 1768 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1885
timestamp 1569543463
transform 1 0 1832 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1886
timestamp 1569543463
transform 1 0 1704 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1887
timestamp 1569543463
transform 1 0 1768 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1888
timestamp 1569543463
transform 1 0 1832 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1889
timestamp 1569543463
transform 1 0 1640 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1890
timestamp 1569543463
transform 1 0 1640 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1891
timestamp 1569543463
transform 1 0 1640 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1892
timestamp 1569543463
transform 1 0 1704 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1893
timestamp 1569543463
transform 1 0 1704 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1894
timestamp 1569543463
transform 1 0 1704 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1895
timestamp 1569543463
transform 1 0 1832 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1896
timestamp 1569543463
transform 1 0 1640 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1897
timestamp 1569543463
transform 1 0 1832 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1898
timestamp 1569543463
transform 1 0 1768 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1899
timestamp 1569543463
transform 1 0 1512 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1900
timestamp 1569543463
transform 1 0 1512 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1901
timestamp 1569543463
transform 1 0 1320 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1902
timestamp 1569543463
transform 1 0 1320 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1903
timestamp 1569543463
transform 1 0 1384 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1904
timestamp 1569543463
transform 1 0 1384 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1905
timestamp 1569543463
transform 1 0 1448 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1906
timestamp 1569543463
transform 1 0 1448 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1907
timestamp 1569543463
transform 1 0 1512 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1908
timestamp 1569543463
transform 1 0 1320 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1909
timestamp 1569543463
transform 1 0 1320 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1910
timestamp 1569543463
transform 1 0 1512 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1911
timestamp 1569543463
transform 1 0 1448 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1912
timestamp 1569543463
transform 1 0 1384 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1913
timestamp 1569543463
transform 1 0 1448 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1914
timestamp 1569543463
transform 1 0 1384 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1915
timestamp 1569543463
transform 1 0 1384 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1916
timestamp 1569543463
transform 1 0 1448 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1917
timestamp 1569543463
transform 1 0 1448 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1918
timestamp 1569543463
transform 1 0 1512 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1919
timestamp 1569543463
transform 1 0 1320 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1920
timestamp 1569543463
transform 1 0 1448 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1921
timestamp 1569543463
transform 1 0 1448 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1922
timestamp 1569543463
transform 1 0 1384 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1923
timestamp 1569543463
transform 1 0 1512 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1924
timestamp 1569543463
transform 1 0 1512 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1925
timestamp 1569543463
transform 1 0 1384 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1926
timestamp 1569543463
transform 1 0 1320 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1927
timestamp 1569543463
transform 1 0 1320 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1928
timestamp 1569543463
transform 1 0 1384 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1929
timestamp 1569543463
transform 1 0 1320 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1930
timestamp 1569543463
transform 1 0 1512 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1931
timestamp 1569543463
transform 1 0 1704 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1932
timestamp 1569543463
transform 1 0 1768 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1933
timestamp 1569543463
transform 1 0 1832 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1934
timestamp 1569543463
transform 1 0 1704 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1935
timestamp 1569543463
transform 1 0 1704 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1936
timestamp 1569543463
transform 1 0 1768 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1937
timestamp 1569543463
transform 1 0 1768 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1938
timestamp 1569543463
transform 1 0 1832 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1939
timestamp 1569543463
transform 1 0 1832 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1940
timestamp 1569543463
transform 1 0 1640 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1941
timestamp 1569543463
transform 1 0 1640 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1942
timestamp 1569543463
transform 1 0 1832 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1943
timestamp 1569543463
transform 1 0 1640 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1944
timestamp 1569543463
transform 1 0 1640 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1945
timestamp 1569543463
transform 1 0 1704 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1946
timestamp 1569543463
transform 1 0 1768 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1947
timestamp 1569543463
transform 1 0 1576 0 1 1320
box -8 -8 8 8
use VIA2$5  VIA2$5_1948
timestamp 1569543463
transform 1 0 1576 0 1 1448
box -8 -8 8 8
use VIA2$5  VIA2$5_1949
timestamp 1569543463
transform 1 0 1320 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1950
timestamp 1569543463
transform 1 0 1640 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1951
timestamp 1569543463
transform 1 0 1448 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1952
timestamp 1569543463
transform 1 0 1704 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1953
timestamp 1569543463
transform 1 0 1576 0 1 1640
box -8 -8 8 8
use VIA2$5  VIA2$5_1954
timestamp 1569543463
transform 1 0 1576 0 1 1768
box -8 -8 8 8
use VIA2$5  VIA2$5_1955
timestamp 1569543463
transform 1 0 1768 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1956
timestamp 1569543463
transform 1 0 1512 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1957
timestamp 1569543463
transform 1 0 1832 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1958
timestamp 1569543463
transform 1 0 1384 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1959
timestamp 1569543463
transform 1 0 1576 0 1 1576
box -8 -8 8 8
use VIA2$5  VIA2$5_1960
timestamp 1569543463
transform 1 0 1576 0 1 1832
box -8 -8 8 8
use VIA2$5  VIA2$5_1961
timestamp 1569543463
transform 1 0 1576 0 1 1384
box -8 -8 8 8
use VIA2$5  VIA2$5_1962
timestamp 1569543463
transform 1 0 1576 0 1 1512
box -8 -8 8 8
use VIA2$5  VIA2$5_1963
timestamp 1569543463
transform 1 0 1576 0 1 1704
box -8 -8 8 8
use VIA2$5  VIA2$5_1964
timestamp 1569543463
transform 1 0 1704 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1965
timestamp 1569543463
transform 1 0 1768 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1966
timestamp 1569543463
transform 1 0 1704 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1967
timestamp 1569543463
transform 1 0 1832 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1968
timestamp 1569543463
transform 1 0 1768 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1969
timestamp 1569543463
transform 1 0 1768 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1970
timestamp 1569543463
transform 1 0 1768 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1971
timestamp 1569543463
transform 1 0 1640 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1972
timestamp 1569543463
transform 1 0 1640 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1973
timestamp 1569543463
transform 1 0 1704 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1974
timestamp 1569543463
transform 1 0 1768 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1975
timestamp 1569543463
transform 1 0 1832 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1976
timestamp 1569543463
transform 1 0 1640 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1977
timestamp 1569543463
transform 1 0 1832 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1978
timestamp 1569543463
transform 1 0 1832 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1979
timestamp 1569543463
transform 1 0 1832 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1980
timestamp 1569543463
transform 1 0 1640 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1981
timestamp 1569543463
transform 1 0 1640 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1982
timestamp 1569543463
transform 1 0 1704 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1983
timestamp 1569543463
transform 1 0 1704 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1984
timestamp 1569543463
transform 1 0 1384 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1985
timestamp 1569543463
transform 1 0 1512 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1986
timestamp 1569543463
transform 1 0 1448 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1987
timestamp 1569543463
transform 1 0 1512 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1988
timestamp 1569543463
transform 1 0 1512 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1989
timestamp 1569543463
transform 1 0 1512 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1990
timestamp 1569543463
transform 1 0 1320 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_1991
timestamp 1569543463
transform 1 0 1320 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1992
timestamp 1569543463
transform 1 0 1384 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1993
timestamp 1569543463
transform 1 0 1320 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1994
timestamp 1569543463
transform 1 0 1384 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_1995
timestamp 1569543463
transform 1 0 1320 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_1996
timestamp 1569543463
transform 1 0 1512 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1997
timestamp 1569543463
transform 1 0 1448 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_1998
timestamp 1569543463
transform 1 0 1448 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_1999
timestamp 1569543463
transform 1 0 1448 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2000
timestamp 1569543463
transform 1 0 1448 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2001
timestamp 1569543463
transform 1 0 1320 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2002
timestamp 1569543463
transform 1 0 1384 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2003
timestamp 1569543463
transform 1 0 1384 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2004
timestamp 1569543463
transform 1 0 1384 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2005
timestamp 1569543463
transform 1 0 1320 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2006
timestamp 1569543463
transform 1 0 1512 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2007
timestamp 1569543463
transform 1 0 1384 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2008
timestamp 1569543463
transform 1 0 1320 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2009
timestamp 1569543463
transform 1 0 1512 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2010
timestamp 1569543463
transform 1 0 1320 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2011
timestamp 1569543463
transform 1 0 1384 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2012
timestamp 1569543463
transform 1 0 1320 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2013
timestamp 1569543463
transform 1 0 1448 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2014
timestamp 1569543463
transform 1 0 1384 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2015
timestamp 1569543463
transform 1 0 1448 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2016
timestamp 1569543463
transform 1 0 1384 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2017
timestamp 1569543463
transform 1 0 1448 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2018
timestamp 1569543463
transform 1 0 1320 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2019
timestamp 1569543463
transform 1 0 1512 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2020
timestamp 1569543463
transform 1 0 1448 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2021
timestamp 1569543463
transform 1 0 1512 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2022
timestamp 1569543463
transform 1 0 1448 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2023
timestamp 1569543463
transform 1 0 1512 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2024
timestamp 1569543463
transform 1 0 1704 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2025
timestamp 1569543463
transform 1 0 1704 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2026
timestamp 1569543463
transform 1 0 1768 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2027
timestamp 1569543463
transform 1 0 1768 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2028
timestamp 1569543463
transform 1 0 1704 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2029
timestamp 1569543463
transform 1 0 1768 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2030
timestamp 1569543463
transform 1 0 1832 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2031
timestamp 1569543463
transform 1 0 1832 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2032
timestamp 1569543463
transform 1 0 1832 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2033
timestamp 1569543463
transform 1 0 1832 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2034
timestamp 1569543463
transform 1 0 1832 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2035
timestamp 1569543463
transform 1 0 1704 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2036
timestamp 1569543463
transform 1 0 1704 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2037
timestamp 1569543463
transform 1 0 1768 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2038
timestamp 1569543463
transform 1 0 1768 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2039
timestamp 1569543463
transform 1 0 1640 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2040
timestamp 1569543463
transform 1 0 1640 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2041
timestamp 1569543463
transform 1 0 1640 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2042
timestamp 1569543463
transform 1 0 1640 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2043
timestamp 1569543463
transform 1 0 1640 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2044
timestamp 1569543463
transform 1 0 1576 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2045
timestamp 1569543463
transform 1 0 1576 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2046
timestamp 1569543463
transform 1 0 1576 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2047
timestamp 1569543463
transform 1 0 1576 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2048
timestamp 1569543463
transform 1 0 1576 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2049
timestamp 1569543463
transform 1 0 1576 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2050
timestamp 1569543463
transform 1 0 1576 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2051
timestamp 1569543463
transform 1 0 1576 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2052
timestamp 1569543463
transform 1 0 1576 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2053
timestamp 1569543463
transform 1 0 1576 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2054
timestamp 1569543463
transform 1 0 2344 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2055
timestamp 1569543463
transform 1 0 2408 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2056
timestamp 1569543463
transform 1 0 2472 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2057
timestamp 1569543463
transform 1 0 2408 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2058
timestamp 1569543463
transform 1 0 2280 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2059
timestamp 1569543463
transform 1 0 2280 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2060
timestamp 1569543463
transform 1 0 2280 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2061
timestamp 1569543463
transform 1 0 2344 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2062
timestamp 1569543463
transform 1 0 2344 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2063
timestamp 1569543463
transform 1 0 2216 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2064
timestamp 1569543463
transform 1 0 2344 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2065
timestamp 1569543463
transform 1 0 2280 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2066
timestamp 1569543463
transform 1 0 2280 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2067
timestamp 1569543463
transform 1 0 2216 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2068
timestamp 1569543463
transform 1 0 2216 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2069
timestamp 1569543463
transform 1 0 2216 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2070
timestamp 1569543463
transform 1 0 2408 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2071
timestamp 1569543463
transform 1 0 2472 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2072
timestamp 1569543463
transform 1 0 2216 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2073
timestamp 1569543463
transform 1 0 1896 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2074
timestamp 1569543463
transform 1 0 2024 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2075
timestamp 1569543463
transform 1 0 2024 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2076
timestamp 1569543463
transform 1 0 2024 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2077
timestamp 1569543463
transform 1 0 1960 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2078
timestamp 1569543463
transform 1 0 2088 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2079
timestamp 1569543463
transform 1 0 2088 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2080
timestamp 1569543463
transform 1 0 2088 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2081
timestamp 1569543463
transform 1 0 1896 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2082
timestamp 1569543463
transform 1 0 1960 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2083
timestamp 1569543463
transform 1 0 2152 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2084
timestamp 1569543463
transform 1 0 2024 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2085
timestamp 1569543463
transform 1 0 2088 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2086
timestamp 1569543463
transform 1 0 2024 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2087
timestamp 1569543463
transform 1 0 1960 0 1 2152
box -8 -8 8 8
use VIA2$5  VIA2$5_2088
timestamp 1569543463
transform 1 0 2088 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2089
timestamp 1569543463
transform 1 0 2152 0 1 1896
box -8 -8 8 8
use VIA2$5  VIA2$5_2090
timestamp 1569543463
transform 1 0 1896 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2091
timestamp 1569543463
transform 1 0 2152 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2092
timestamp 1569543463
transform 1 0 1896 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2093
timestamp 1569543463
transform 1 0 2152 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2094
timestamp 1569543463
transform 1 0 1896 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2095
timestamp 1569543463
transform 1 0 2152 0 1 2088
box -8 -8 8 8
use VIA2$5  VIA2$5_2096
timestamp 1569543463
transform 1 0 1960 0 1 1960
box -8 -8 8 8
use VIA2$5  VIA2$5_2097
timestamp 1569543463
transform 1 0 1960 0 1 2024
box -8 -8 8 8
use VIA2$5  VIA2$5_2098
timestamp 1569543463
transform 1 0 1896 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2099
timestamp 1569543463
transform 1 0 1896 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2100
timestamp 1569543463
transform 1 0 1896 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2101
timestamp 1569543463
transform 1 0 1896 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2102
timestamp 1569543463
transform 1 0 1896 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2103
timestamp 1569543463
transform 1 0 1960 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2104
timestamp 1569543463
transform 1 0 1960 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2105
timestamp 1569543463
transform 1 0 1960 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2106
timestamp 1569543463
transform 1 0 1960 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2107
timestamp 1569543463
transform 1 0 1960 0 1 2472
box -8 -8 8 8
use VIA2$5  VIA2$5_2108
timestamp 1569543463
transform 1 0 2152 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2109
timestamp 1569543463
transform 1 0 2152 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2110
timestamp 1569543463
transform 1 0 2024 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2111
timestamp 1569543463
transform 1 0 2024 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2112
timestamp 1569543463
transform 1 0 2024 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2113
timestamp 1569543463
transform 1 0 2024 0 1 2408
box -8 -8 8 8
use VIA2$5  VIA2$5_2114
timestamp 1569543463
transform 1 0 2088 0 1 2344
box -8 -8 8 8
use VIA2$5  VIA2$5_2115
timestamp 1569543463
transform 1 0 2088 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2116
timestamp 1569543463
transform 1 0 2088 0 1 2280
box -8 -8 8 8
use VIA2$5  VIA2$5_2117
timestamp 1569543463
transform 1 0 2216 0 1 2216
box -8 -8 8 8
use VIA2$5  VIA2$5_2118
timestamp 1569543463
transform 1 0 1896 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2119
timestamp 1569543463
transform 1 0 1640 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2120
timestamp 1569543463
transform 1 0 1768 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2121
timestamp 1569543463
transform 1 0 1704 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2122
timestamp 1569543463
transform 1 0 1768 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2123
timestamp 1569543463
transform 1 0 1832 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2124
timestamp 1569543463
transform 1 0 1704 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2125
timestamp 1569543463
transform 1 0 1640 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2126
timestamp 1569543463
transform 1 0 1704 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2127
timestamp 1569543463
transform 1 0 1768 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2128
timestamp 1569543463
transform 1 0 1640 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2129
timestamp 1569543463
transform 1 0 1640 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2130
timestamp 1569543463
transform 1 0 1704 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2131
timestamp 1569543463
transform 1 0 1832 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2132
timestamp 1569543463
transform 1 0 1640 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2133
timestamp 1569543463
transform 1 0 1384 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2134
timestamp 1569543463
transform 1 0 1448 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2135
timestamp 1569543463
transform 1 0 1512 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2136
timestamp 1569543463
transform 1 0 1512 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2137
timestamp 1569543463
transform 1 0 1448 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2138
timestamp 1569543463
transform 1 0 1384 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2139
timestamp 1569543463
transform 1 0 1320 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2140
timestamp 1569543463
transform 1 0 1448 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2141
timestamp 1569543463
transform 1 0 1320 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2142
timestamp 1569543463
transform 1 0 1448 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2143
timestamp 1569543463
transform 1 0 1320 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2144
timestamp 1569543463
transform 1 0 1384 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2145
timestamp 1569543463
transform 1 0 1512 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2146
timestamp 1569543463
transform 1 0 1512 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2147
timestamp 1569543463
transform 1 0 1448 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2148
timestamp 1569543463
transform 1 0 1384 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2149
timestamp 1569543463
transform 1 0 1384 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2150
timestamp 1569543463
transform 1 0 1320 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2151
timestamp 1569543463
transform 1 0 1320 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2152
timestamp 1569543463
transform 1 0 1512 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2153
timestamp 1569543463
transform 1 0 1512 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2154
timestamp 1569543463
transform 1 0 1448 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2155
timestamp 1569543463
transform 1 0 1384 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2156
timestamp 1569543463
transform 1 0 1512 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2157
timestamp 1569543463
transform 1 0 1512 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2158
timestamp 1569543463
transform 1 0 1384 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2159
timestamp 1569543463
transform 1 0 1384 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2160
timestamp 1569543463
transform 1 0 1448 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2161
timestamp 1569543463
transform 1 0 1512 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2162
timestamp 1569543463
transform 1 0 1512 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2163
timestamp 1569543463
transform 1 0 1384 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2164
timestamp 1569543463
transform 1 0 1320 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2165
timestamp 1569543463
transform 1 0 1320 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2166
timestamp 1569543463
transform 1 0 1384 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2167
timestamp 1569543463
transform 1 0 1448 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2168
timestamp 1569543463
transform 1 0 1448 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2169
timestamp 1569543463
transform 1 0 1448 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2170
timestamp 1569543463
transform 1 0 1320 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2171
timestamp 1569543463
transform 1 0 1320 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2172
timestamp 1569543463
transform 1 0 1320 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2173
timestamp 1569543463
transform 1 0 1576 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2174
timestamp 1569543463
transform 1 0 1576 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2175
timestamp 1569543463
transform 1 0 1576 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2176
timestamp 1569543463
transform 1 0 1576 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2177
timestamp 1569543463
transform 1 0 1576 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2178
timestamp 1569543463
transform 1 0 1576 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2179
timestamp 1569543463
transform 1 0 1320 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2180
timestamp 1569543463
transform 1 0 1384 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2181
timestamp 1569543463
transform 1 0 1320 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2182
timestamp 1569543463
transform 1 0 1512 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2183
timestamp 1569543463
transform 1 0 1384 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2184
timestamp 1569543463
transform 1 0 1320 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2185
timestamp 1569543463
transform 1 0 1512 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2186
timestamp 1569543463
transform 1 0 1384 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2187
timestamp 1569543463
transform 1 0 1320 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2188
timestamp 1569543463
transform 1 0 1512 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2189
timestamp 1569543463
transform 1 0 1448 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2190
timestamp 1569543463
transform 1 0 1512 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2191
timestamp 1569543463
transform 1 0 1384 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2192
timestamp 1569543463
transform 1 0 1320 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2193
timestamp 1569543463
transform 1 0 1448 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2194
timestamp 1569543463
transform 1 0 1384 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2195
timestamp 1569543463
transform 1 0 1320 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2196
timestamp 1569543463
transform 1 0 1384 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2197
timestamp 1569543463
transform 1 0 1384 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2198
timestamp 1569543463
transform 1 0 1384 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2199
timestamp 1569543463
transform 1 0 1320 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2200
timestamp 1569543463
transform 1 0 1512 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2201
timestamp 1569543463
transform 1 0 1448 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2202
timestamp 1569543463
transform 1 0 1512 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2203
timestamp 1569543463
transform 1 0 1320 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2204
timestamp 1569543463
transform 1 0 1384 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2205
timestamp 1569543463
transform 1 0 1448 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2206
timestamp 1569543463
transform 1 0 1448 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2207
timestamp 1569543463
transform 1 0 1512 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2208
timestamp 1569543463
transform 1 0 1512 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2209
timestamp 1569543463
transform 1 0 1448 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2210
timestamp 1569543463
transform 1 0 1320 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2211
timestamp 1569543463
transform 1 0 1512 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2212
timestamp 1569543463
transform 1 0 1448 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2213
timestamp 1569543463
transform 1 0 1448 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2214
timestamp 1569543463
transform 1 0 1448 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2215
timestamp 1569543463
transform 1 0 2472 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2216
timestamp 1569543463
transform 1 0 2344 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2217
timestamp 1569543463
transform 1 0 2344 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2218
timestamp 1569543463
transform 1 0 2472 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2219
timestamp 1569543463
transform 1 0 2472 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2220
timestamp 1569543463
transform 1 0 2472 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2221
timestamp 1569543463
transform 1 0 2472 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2222
timestamp 1569543463
transform 1 0 2344 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2223
timestamp 1569543463
transform 1 0 2408 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2224
timestamp 1569543463
transform 1 0 2472 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2225
timestamp 1569543463
transform 1 0 2408 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2226
timestamp 1569543463
transform 1 0 2472 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2227
timestamp 1569543463
transform 1 0 2408 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2228
timestamp 1569543463
transform 1 0 2344 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2229
timestamp 1569543463
transform 1 0 2408 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2230
timestamp 1569543463
transform 1 0 2408 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2231
timestamp 1569543463
transform 1 0 2408 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2232
timestamp 1569543463
transform 1 0 2344 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2233
timestamp 1569543463
transform 1 0 2408 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2234
timestamp 1569543463
transform 1 0 2344 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2235
timestamp 1569543463
transform 1 0 2472 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2236
timestamp 1569543463
transform 1 0 1256 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2237
timestamp 1569543463
transform 1 0 1064 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2238
timestamp 1569543463
transform 1 0 1000 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2239
timestamp 1569543463
transform 1 0 1256 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2240
timestamp 1569543463
transform 1 0 1000 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2241
timestamp 1569543463
transform 1 0 1128 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2242
timestamp 1569543463
transform 1 0 1064 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2243
timestamp 1569543463
transform 1 0 1192 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2244
timestamp 1569543463
transform 1 0 1064 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2245
timestamp 1569543463
transform 1 0 1192 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2246
timestamp 1569543463
transform 1 0 1256 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2247
timestamp 1569543463
transform 1 0 1064 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2248
timestamp 1569543463
transform 1 0 1000 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2249
timestamp 1569543463
transform 1 0 1128 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2250
timestamp 1569543463
transform 1 0 1000 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2251
timestamp 1569543463
transform 1 0 1192 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2252
timestamp 1569543463
transform 1 0 1128 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2253
timestamp 1569543463
transform 1 0 1256 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2254
timestamp 1569543463
transform 1 0 1192 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2255
timestamp 1569543463
transform 1 0 1256 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2256
timestamp 1569543463
transform 1 0 1064 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2257
timestamp 1569543463
transform 1 0 1128 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2258
timestamp 1569543463
transform 1 0 1128 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2259
timestamp 1569543463
transform 1 0 1192 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2260
timestamp 1569543463
transform 1 0 1000 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2261
timestamp 1569543463
transform 1 0 680 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2262
timestamp 1569543463
transform 1 0 936 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2263
timestamp 1569543463
transform 1 0 808 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2264
timestamp 1569543463
transform 1 0 680 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2265
timestamp 1569543463
transform 1 0 744 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2266
timestamp 1569543463
transform 1 0 744 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2267
timestamp 1569543463
transform 1 0 744 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2268
timestamp 1569543463
transform 1 0 936 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2269
timestamp 1569543463
transform 1 0 680 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2270
timestamp 1569543463
transform 1 0 808 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2271
timestamp 1569543463
transform 1 0 808 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2272
timestamp 1569543463
transform 1 0 808 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2273
timestamp 1569543463
transform 1 0 872 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2274
timestamp 1569543463
transform 1 0 872 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2275
timestamp 1569543463
transform 1 0 936 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2276
timestamp 1569543463
transform 1 0 872 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2277
timestamp 1569543463
transform 1 0 936 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2278
timestamp 1569543463
transform 1 0 680 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2279
timestamp 1569543463
transform 1 0 808 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2280
timestamp 1569543463
transform 1 0 744 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2281
timestamp 1569543463
transform 1 0 680 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2282
timestamp 1569543463
transform 1 0 872 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2283
timestamp 1569543463
transform 1 0 936 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2284
timestamp 1569543463
transform 1 0 744 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2285
timestamp 1569543463
transform 1 0 872 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2286
timestamp 1569543463
transform 1 0 936 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2287
timestamp 1569543463
transform 1 0 808 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2288
timestamp 1569543463
transform 1 0 872 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2289
timestamp 1569543463
transform 1 0 680 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2290
timestamp 1569543463
transform 1 0 872 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2291
timestamp 1569543463
transform 1 0 680 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2292
timestamp 1569543463
transform 1 0 744 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2293
timestamp 1569543463
transform 1 0 744 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2294
timestamp 1569543463
transform 1 0 808 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2295
timestamp 1569543463
transform 1 0 808 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2296
timestamp 1569543463
transform 1 0 936 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2297
timestamp 1569543463
transform 1 0 872 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2298
timestamp 1569543463
transform 1 0 936 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2299
timestamp 1569543463
transform 1 0 808 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2300
timestamp 1569543463
transform 1 0 744 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2301
timestamp 1569543463
transform 1 0 744 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2302
timestamp 1569543463
transform 1 0 808 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2303
timestamp 1569543463
transform 1 0 936 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2304
timestamp 1569543463
transform 1 0 680 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2305
timestamp 1569543463
transform 1 0 680 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2306
timestamp 1569543463
transform 1 0 936 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2307
timestamp 1569543463
transform 1 0 872 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2308
timestamp 1569543463
transform 1 0 744 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2309
timestamp 1569543463
transform 1 0 872 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2310
timestamp 1569543463
transform 1 0 680 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2311
timestamp 1569543463
transform 1 0 1000 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2312
timestamp 1569543463
transform 1 0 1128 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2313
timestamp 1569543463
transform 1 0 1192 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2314
timestamp 1569543463
transform 1 0 1000 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2315
timestamp 1569543463
transform 1 0 1000 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2316
timestamp 1569543463
transform 1 0 1064 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2317
timestamp 1569543463
transform 1 0 1256 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2318
timestamp 1569543463
transform 1 0 1256 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2319
timestamp 1569543463
transform 1 0 1128 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2320
timestamp 1569543463
transform 1 0 1256 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2321
timestamp 1569543463
transform 1 0 1000 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2322
timestamp 1569543463
transform 1 0 1256 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2323
timestamp 1569543463
transform 1 0 1000 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2324
timestamp 1569543463
transform 1 0 1064 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2325
timestamp 1569543463
transform 1 0 1192 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2326
timestamp 1569543463
transform 1 0 1192 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2327
timestamp 1569543463
transform 1 0 1128 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2328
timestamp 1569543463
transform 1 0 1064 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2329
timestamp 1569543463
transform 1 0 1128 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2330
timestamp 1569543463
transform 1 0 1192 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2331
timestamp 1569543463
transform 1 0 1192 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2332
timestamp 1569543463
transform 1 0 1064 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2333
timestamp 1569543463
transform 1 0 1064 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2334
timestamp 1569543463
transform 1 0 1256 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2335
timestamp 1569543463
transform 1 0 1128 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2336
timestamp 1569543463
transform 1 0 488 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2337
timestamp 1569543463
transform 1 0 616 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2338
timestamp 1569543463
transform 1 0 552 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2339
timestamp 1569543463
transform 1 0 616 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2340
timestamp 1569543463
transform 1 0 616 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2341
timestamp 1569543463
transform 1 0 552 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2342
timestamp 1569543463
transform 1 0 488 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2343
timestamp 1569543463
transform 1 0 616 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2344
timestamp 1569543463
transform 1 0 552 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2345
timestamp 1569543463
transform 1 0 552 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2346
timestamp 1569543463
transform 1 0 488 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2347
timestamp 1569543463
transform 1 0 360 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2348
timestamp 1569543463
transform 1 0 424 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2349
timestamp 1569543463
transform 1 0 360 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2350
timestamp 1569543463
transform 1 0 488 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2351
timestamp 1569543463
transform 1 0 552 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2352
timestamp 1569543463
transform 1 0 424 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2353
timestamp 1569543463
transform 1 0 424 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2354
timestamp 1569543463
transform 1 0 360 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2355
timestamp 1569543463
transform 1 0 488 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2356
timestamp 1569543463
transform 1 0 424 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2357
timestamp 1569543463
transform 1 0 360 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2358
timestamp 1569543463
transform 1 0 616 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2359
timestamp 1569543463
transform 1 0 424 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2360
timestamp 1569543463
transform 1 0 360 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2361
timestamp 1569543463
transform 1 0 232 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2362
timestamp 1569543463
transform 1 0 232 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2363
timestamp 1569543463
transform 1 0 296 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2364
timestamp 1569543463
transform 1 0 296 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2365
timestamp 1569543463
transform 1 0 104 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2366
timestamp 1569543463
transform 1 0 232 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2367
timestamp 1569543463
transform 1 0 168 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2368
timestamp 1569543463
transform 1 0 104 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2369
timestamp 1569543463
transform 1 0 296 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2370
timestamp 1569543463
transform 1 0 104 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2371
timestamp 1569543463
transform 1 0 40 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2372
timestamp 1569543463
transform 1 0 232 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2373
timestamp 1569543463
transform 1 0 40 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2374
timestamp 1569543463
transform 1 0 104 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2375
timestamp 1569543463
transform 1 0 168 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2376
timestamp 1569543463
transform 1 0 168 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2377
timestamp 1569543463
transform 1 0 40 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2378
timestamp 1569543463
transform 1 0 296 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2379
timestamp 1569543463
transform 1 0 168 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2380
timestamp 1569543463
transform 1 0 40 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_2381
timestamp 1569543463
transform 1 0 296 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2382
timestamp 1569543463
transform 1 0 104 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_2383
timestamp 1569543463
transform 1 0 40 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_2384
timestamp 1569543463
transform 1 0 232 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_2385
timestamp 1569543463
transform 1 0 168 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_2386
timestamp 1569543463
transform 1 0 232 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2387
timestamp 1569543463
transform 1 0 168 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2388
timestamp 1569543463
transform 1 0 232 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2389
timestamp 1569543463
transform 1 0 232 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2390
timestamp 1569543463
transform 1 0 232 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2391
timestamp 1569543463
transform 1 0 168 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2392
timestamp 1569543463
transform 1 0 40 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2393
timestamp 1569543463
transform 1 0 40 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2394
timestamp 1569543463
transform 1 0 296 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2395
timestamp 1569543463
transform 1 0 232 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2396
timestamp 1569543463
transform 1 0 296 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2397
timestamp 1569543463
transform 1 0 40 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2398
timestamp 1569543463
transform 1 0 168 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2399
timestamp 1569543463
transform 1 0 104 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2400
timestamp 1569543463
transform 1 0 168 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2401
timestamp 1569543463
transform 1 0 104 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2402
timestamp 1569543463
transform 1 0 104 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2403
timestamp 1569543463
transform 1 0 40 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2404
timestamp 1569543463
transform 1 0 296 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2405
timestamp 1569543463
transform 1 0 296 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2406
timestamp 1569543463
transform 1 0 296 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2407
timestamp 1569543463
transform 1 0 104 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2408
timestamp 1569543463
transform 1 0 40 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2409
timestamp 1569543463
transform 1 0 104 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2410
timestamp 1569543463
transform 1 0 168 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2411
timestamp 1569543463
transform 1 0 616 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2412
timestamp 1569543463
transform 1 0 360 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2413
timestamp 1569543463
transform 1 0 616 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2414
timestamp 1569543463
transform 1 0 616 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2415
timestamp 1569543463
transform 1 0 488 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2416
timestamp 1569543463
transform 1 0 616 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2417
timestamp 1569543463
transform 1 0 360 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2418
timestamp 1569543463
transform 1 0 616 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2419
timestamp 1569543463
transform 1 0 488 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2420
timestamp 1569543463
transform 1 0 360 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2421
timestamp 1569543463
transform 1 0 424 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2422
timestamp 1569543463
transform 1 0 552 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2423
timestamp 1569543463
transform 1 0 488 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2424
timestamp 1569543463
transform 1 0 360 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2425
timestamp 1569543463
transform 1 0 424 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2426
timestamp 1569543463
transform 1 0 488 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2427
timestamp 1569543463
transform 1 0 552 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2428
timestamp 1569543463
transform 1 0 488 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2429
timestamp 1569543463
transform 1 0 424 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2430
timestamp 1569543463
transform 1 0 424 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2431
timestamp 1569543463
transform 1 0 552 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_2432
timestamp 1569543463
transform 1 0 552 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_2433
timestamp 1569543463
transform 1 0 552 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_2434
timestamp 1569543463
transform 1 0 360 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_2435
timestamp 1569543463
transform 1 0 424 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_2436
timestamp 1569543463
transform 1 0 616 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2437
timestamp 1569543463
transform 1 0 552 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2438
timestamp 1569543463
transform 1 0 616 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2439
timestamp 1569543463
transform 1 0 424 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2440
timestamp 1569543463
transform 1 0 360 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2441
timestamp 1569543463
transform 1 0 488 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2442
timestamp 1569543463
transform 1 0 552 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2443
timestamp 1569543463
transform 1 0 360 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2444
timestamp 1569543463
transform 1 0 424 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2445
timestamp 1569543463
transform 1 0 424 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2446
timestamp 1569543463
transform 1 0 488 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2447
timestamp 1569543463
transform 1 0 360 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2448
timestamp 1569543463
transform 1 0 488 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2449
timestamp 1569543463
transform 1 0 552 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2450
timestamp 1569543463
transform 1 0 616 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2451
timestamp 1569543463
transform 1 0 424 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2452
timestamp 1569543463
transform 1 0 616 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2453
timestamp 1569543463
transform 1 0 552 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2454
timestamp 1569543463
transform 1 0 488 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2455
timestamp 1569543463
transform 1 0 360 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2456
timestamp 1569543463
transform 1 0 232 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2457
timestamp 1569543463
transform 1 0 104 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2458
timestamp 1569543463
transform 1 0 168 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2459
timestamp 1569543463
transform 1 0 40 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2460
timestamp 1569543463
transform 1 0 168 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2461
timestamp 1569543463
transform 1 0 296 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2462
timestamp 1569543463
transform 1 0 40 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2463
timestamp 1569543463
transform 1 0 232 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2464
timestamp 1569543463
transform 1 0 40 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2465
timestamp 1569543463
transform 1 0 40 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2466
timestamp 1569543463
transform 1 0 104 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2467
timestamp 1569543463
transform 1 0 296 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2468
timestamp 1569543463
transform 1 0 232 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2469
timestamp 1569543463
transform 1 0 168 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2470
timestamp 1569543463
transform 1 0 296 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2471
timestamp 1569543463
transform 1 0 104 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2472
timestamp 1569543463
transform 1 0 296 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2473
timestamp 1569543463
transform 1 0 168 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2474
timestamp 1569543463
transform 1 0 232 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2475
timestamp 1569543463
transform 1 0 104 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2476
timestamp 1569543463
transform 1 0 296 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2477
timestamp 1569543463
transform 1 0 232 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2478
timestamp 1569543463
transform 1 0 40 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2479
timestamp 1569543463
transform 1 0 104 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2480
timestamp 1569543463
transform 1 0 232 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2481
timestamp 1569543463
transform 1 0 168 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2482
timestamp 1569543463
transform 1 0 104 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2483
timestamp 1569543463
transform 1 0 168 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2484
timestamp 1569543463
transform 1 0 232 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2485
timestamp 1569543463
transform 1 0 296 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2486
timestamp 1569543463
transform 1 0 168 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2487
timestamp 1569543463
transform 1 0 104 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2488
timestamp 1569543463
transform 1 0 296 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2489
timestamp 1569543463
transform 1 0 296 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2490
timestamp 1569543463
transform 1 0 40 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2491
timestamp 1569543463
transform 1 0 40 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2492
timestamp 1569543463
transform 1 0 40 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2493
timestamp 1569543463
transform 1 0 168 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2494
timestamp 1569543463
transform 1 0 232 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2495
timestamp 1569543463
transform 1 0 104 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2496
timestamp 1569543463
transform 1 0 552 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2497
timestamp 1569543463
transform 1 0 360 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2498
timestamp 1569543463
transform 1 0 552 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2499
timestamp 1569543463
transform 1 0 616 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2500
timestamp 1569543463
transform 1 0 424 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2501
timestamp 1569543463
transform 1 0 488 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2502
timestamp 1569543463
transform 1 0 424 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2503
timestamp 1569543463
transform 1 0 616 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2504
timestamp 1569543463
transform 1 0 488 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2505
timestamp 1569543463
transform 1 0 424 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2506
timestamp 1569543463
transform 1 0 616 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2507
timestamp 1569543463
transform 1 0 488 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2508
timestamp 1569543463
transform 1 0 616 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2509
timestamp 1569543463
transform 1 0 552 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2510
timestamp 1569543463
transform 1 0 360 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2511
timestamp 1569543463
transform 1 0 552 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2512
timestamp 1569543463
transform 1 0 360 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2513
timestamp 1569543463
transform 1 0 424 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2514
timestamp 1569543463
transform 1 0 488 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2515
timestamp 1569543463
transform 1 0 360 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2516
timestamp 1569543463
transform 1 0 424 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2517
timestamp 1569543463
transform 1 0 40 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2518
timestamp 1569543463
transform 1 0 296 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2519
timestamp 1569543463
transform 1 0 168 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2520
timestamp 1569543463
transform 1 0 616 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2521
timestamp 1569543463
transform 1 0 488 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2522
timestamp 1569543463
transform 1 0 360 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2523
timestamp 1569543463
transform 1 0 232 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2524
timestamp 1569543463
transform 1 0 104 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2525
timestamp 1569543463
transform 1 0 552 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2526
timestamp 1569543463
transform 1 0 1064 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2527
timestamp 1569543463
transform 1 0 1128 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2528
timestamp 1569543463
transform 1 0 1192 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2529
timestamp 1569543463
transform 1 0 1064 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2530
timestamp 1569543463
transform 1 0 1192 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2531
timestamp 1569543463
transform 1 0 1256 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2532
timestamp 1569543463
transform 1 0 1000 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2533
timestamp 1569543463
transform 1 0 1256 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2534
timestamp 1569543463
transform 1 0 1256 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2535
timestamp 1569543463
transform 1 0 1192 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2536
timestamp 1569543463
transform 1 0 1000 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2537
timestamp 1569543463
transform 1 0 1128 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2538
timestamp 1569543463
transform 1 0 1000 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2539
timestamp 1569543463
transform 1 0 1192 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2540
timestamp 1569543463
transform 1 0 1256 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2541
timestamp 1569543463
transform 1 0 1064 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2542
timestamp 1569543463
transform 1 0 1128 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2543
timestamp 1569543463
transform 1 0 1000 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2544
timestamp 1569543463
transform 1 0 1064 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2545
timestamp 1569543463
transform 1 0 1128 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2546
timestamp 1569543463
transform 1 0 872 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2547
timestamp 1569543463
transform 1 0 680 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2548
timestamp 1569543463
transform 1 0 808 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2549
timestamp 1569543463
transform 1 0 808 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2550
timestamp 1569543463
transform 1 0 936 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2551
timestamp 1569543463
transform 1 0 680 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2552
timestamp 1569543463
transform 1 0 872 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2553
timestamp 1569543463
transform 1 0 744 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2554
timestamp 1569543463
transform 1 0 744 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2555
timestamp 1569543463
transform 1 0 872 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2556
timestamp 1569543463
transform 1 0 872 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2557
timestamp 1569543463
transform 1 0 680 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2558
timestamp 1569543463
transform 1 0 808 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2559
timestamp 1569543463
transform 1 0 744 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_2560
timestamp 1569543463
transform 1 0 936 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_2561
timestamp 1569543463
transform 1 0 936 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2562
timestamp 1569543463
transform 1 0 808 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2563
timestamp 1569543463
transform 1 0 744 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_2564
timestamp 1569543463
transform 1 0 936 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2565
timestamp 1569543463
transform 1 0 680 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_2566
timestamp 1569543463
transform 1 0 680 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2567
timestamp 1569543463
transform 1 0 680 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2568
timestamp 1569543463
transform 1 0 744 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2569
timestamp 1569543463
transform 1 0 808 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2570
timestamp 1569543463
transform 1 0 744 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2571
timestamp 1569543463
transform 1 0 808 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2572
timestamp 1569543463
transform 1 0 936 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2573
timestamp 1569543463
transform 1 0 808 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2574
timestamp 1569543463
transform 1 0 872 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2575
timestamp 1569543463
transform 1 0 936 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2576
timestamp 1569543463
transform 1 0 808 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2577
timestamp 1569543463
transform 1 0 872 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2578
timestamp 1569543463
transform 1 0 936 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2579
timestamp 1569543463
transform 1 0 936 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2580
timestamp 1569543463
transform 1 0 680 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2581
timestamp 1569543463
transform 1 0 680 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2582
timestamp 1569543463
transform 1 0 872 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2583
timestamp 1569543463
transform 1 0 744 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2584
timestamp 1569543463
transform 1 0 872 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2585
timestamp 1569543463
transform 1 0 744 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2586
timestamp 1569543463
transform 1 0 1064 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2587
timestamp 1569543463
transform 1 0 1192 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2588
timestamp 1569543463
transform 1 0 1064 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2589
timestamp 1569543463
transform 1 0 1128 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2590
timestamp 1569543463
transform 1 0 1000 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2591
timestamp 1569543463
transform 1 0 1256 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2592
timestamp 1569543463
transform 1 0 1256 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2593
timestamp 1569543463
transform 1 0 1000 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2594
timestamp 1569543463
transform 1 0 1064 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2595
timestamp 1569543463
transform 1 0 1000 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2596
timestamp 1569543463
transform 1 0 1256 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2597
timestamp 1569543463
transform 1 0 1192 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2598
timestamp 1569543463
transform 1 0 1064 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2599
timestamp 1569543463
transform 1 0 1256 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2600
timestamp 1569543463
transform 1 0 1128 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2601
timestamp 1569543463
transform 1 0 1192 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2602
timestamp 1569543463
transform 1 0 1192 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_2603
timestamp 1569543463
transform 1 0 1128 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_2604
timestamp 1569543463
transform 1 0 1000 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_2605
timestamp 1569543463
transform 1 0 1128 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_2606
timestamp 1569543463
transform 1 0 872 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2607
timestamp 1569543463
transform 1 0 1256 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2608
timestamp 1569543463
transform 1 0 1000 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2609
timestamp 1569543463
transform 1 0 680 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2610
timestamp 1569543463
transform 1 0 1192 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2611
timestamp 1569543463
transform 1 0 744 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2612
timestamp 1569543463
transform 1 0 808 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2613
timestamp 1569543463
transform 1 0 1064 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2614
timestamp 1569543463
transform 1 0 1128 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2615
timestamp 1569543463
transform 1 0 936 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_2616
timestamp 1569543463
transform 1 0 1192 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2617
timestamp 1569543463
transform 1 0 1000 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2618
timestamp 1569543463
transform 1 0 1256 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2619
timestamp 1569543463
transform 1 0 1128 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2620
timestamp 1569543463
transform 1 0 1064 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2621
timestamp 1569543463
transform 1 0 1192 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2622
timestamp 1569543463
transform 1 0 1000 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2623
timestamp 1569543463
transform 1 0 1000 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2624
timestamp 1569543463
transform 1 0 1128 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2625
timestamp 1569543463
transform 1 0 1192 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2626
timestamp 1569543463
transform 1 0 1256 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2627
timestamp 1569543463
transform 1 0 1064 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2628
timestamp 1569543463
transform 1 0 1256 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2629
timestamp 1569543463
transform 1 0 1064 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2630
timestamp 1569543463
transform 1 0 1192 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2631
timestamp 1569543463
transform 1 0 1064 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2632
timestamp 1569543463
transform 1 0 1256 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2633
timestamp 1569543463
transform 1 0 1000 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2634
timestamp 1569543463
transform 1 0 1128 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2635
timestamp 1569543463
transform 1 0 1000 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2636
timestamp 1569543463
transform 1 0 1256 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2637
timestamp 1569543463
transform 1 0 1064 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2638
timestamp 1569543463
transform 1 0 1128 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2639
timestamp 1569543463
transform 1 0 1192 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2640
timestamp 1569543463
transform 1 0 1128 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2641
timestamp 1569543463
transform 1 0 744 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2642
timestamp 1569543463
transform 1 0 936 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2643
timestamp 1569543463
transform 1 0 936 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2644
timestamp 1569543463
transform 1 0 936 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2645
timestamp 1569543463
transform 1 0 872 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2646
timestamp 1569543463
transform 1 0 680 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2647
timestamp 1569543463
transform 1 0 936 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2648
timestamp 1569543463
transform 1 0 872 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2649
timestamp 1569543463
transform 1 0 744 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2650
timestamp 1569543463
transform 1 0 808 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2651
timestamp 1569543463
transform 1 0 744 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2652
timestamp 1569543463
transform 1 0 872 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2653
timestamp 1569543463
transform 1 0 808 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2654
timestamp 1569543463
transform 1 0 744 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2655
timestamp 1569543463
transform 1 0 680 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2656
timestamp 1569543463
transform 1 0 680 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2657
timestamp 1569543463
transform 1 0 808 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2658
timestamp 1569543463
transform 1 0 680 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2659
timestamp 1569543463
transform 1 0 936 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2660
timestamp 1569543463
transform 1 0 872 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2661
timestamp 1569543463
transform 1 0 808 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2662
timestamp 1569543463
transform 1 0 744 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2663
timestamp 1569543463
transform 1 0 808 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2664
timestamp 1569543463
transform 1 0 872 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2665
timestamp 1569543463
transform 1 0 680 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2666
timestamp 1569543463
transform 1 0 744 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2667
timestamp 1569543463
transform 1 0 936 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2668
timestamp 1569543463
transform 1 0 872 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2669
timestamp 1569543463
transform 1 0 936 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2670
timestamp 1569543463
transform 1 0 808 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2671
timestamp 1569543463
transform 1 0 808 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2672
timestamp 1569543463
transform 1 0 872 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2673
timestamp 1569543463
transform 1 0 872 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2674
timestamp 1569543463
transform 1 0 808 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2675
timestamp 1569543463
transform 1 0 936 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2676
timestamp 1569543463
transform 1 0 680 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2677
timestamp 1569543463
transform 1 0 872 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2678
timestamp 1569543463
transform 1 0 680 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2679
timestamp 1569543463
transform 1 0 744 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2680
timestamp 1569543463
transform 1 0 680 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2681
timestamp 1569543463
transform 1 0 872 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2682
timestamp 1569543463
transform 1 0 680 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2683
timestamp 1569543463
transform 1 0 744 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2684
timestamp 1569543463
transform 1 0 808 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2685
timestamp 1569543463
transform 1 0 936 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2686
timestamp 1569543463
transform 1 0 936 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2687
timestamp 1569543463
transform 1 0 744 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2688
timestamp 1569543463
transform 1 0 744 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2689
timestamp 1569543463
transform 1 0 808 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2690
timestamp 1569543463
transform 1 0 680 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2691
timestamp 1569543463
transform 1 0 1128 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2692
timestamp 1569543463
transform 1 0 1000 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2693
timestamp 1569543463
transform 1 0 1256 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2694
timestamp 1569543463
transform 1 0 1256 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2695
timestamp 1569543463
transform 1 0 1256 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2696
timestamp 1569543463
transform 1 0 1256 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2697
timestamp 1569543463
transform 1 0 1192 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2698
timestamp 1569543463
transform 1 0 1128 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2699
timestamp 1569543463
transform 1 0 1000 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2700
timestamp 1569543463
transform 1 0 1192 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2701
timestamp 1569543463
transform 1 0 1000 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2702
timestamp 1569543463
transform 1 0 1064 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2703
timestamp 1569543463
transform 1 0 1192 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2704
timestamp 1569543463
transform 1 0 1000 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2705
timestamp 1569543463
transform 1 0 1000 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2706
timestamp 1569543463
transform 1 0 1192 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2707
timestamp 1569543463
transform 1 0 1064 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2708
timestamp 1569543463
transform 1 0 1064 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2709
timestamp 1569543463
transform 1 0 1064 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2710
timestamp 1569543463
transform 1 0 1128 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2711
timestamp 1569543463
transform 1 0 1256 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2712
timestamp 1569543463
transform 1 0 1128 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2713
timestamp 1569543463
transform 1 0 1128 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2714
timestamp 1569543463
transform 1 0 1192 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2715
timestamp 1569543463
transform 1 0 1064 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2716
timestamp 1569543463
transform 1 0 424 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2717
timestamp 1569543463
transform 1 0 424 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2718
timestamp 1569543463
transform 1 0 488 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2719
timestamp 1569543463
transform 1 0 616 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2720
timestamp 1569543463
transform 1 0 552 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2721
timestamp 1569543463
transform 1 0 360 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2722
timestamp 1569543463
transform 1 0 488 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2723
timestamp 1569543463
transform 1 0 360 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2724
timestamp 1569543463
transform 1 0 424 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2725
timestamp 1569543463
transform 1 0 488 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2726
timestamp 1569543463
transform 1 0 424 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2727
timestamp 1569543463
transform 1 0 616 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2728
timestamp 1569543463
transform 1 0 488 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2729
timestamp 1569543463
transform 1 0 616 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2730
timestamp 1569543463
transform 1 0 552 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2731
timestamp 1569543463
transform 1 0 360 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2732
timestamp 1569543463
transform 1 0 360 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2733
timestamp 1569543463
transform 1 0 616 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2734
timestamp 1569543463
transform 1 0 552 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2735
timestamp 1569543463
transform 1 0 424 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2736
timestamp 1569543463
transform 1 0 552 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2737
timestamp 1569543463
transform 1 0 616 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2738
timestamp 1569543463
transform 1 0 552 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2739
timestamp 1569543463
transform 1 0 360 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2740
timestamp 1569543463
transform 1 0 488 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2741
timestamp 1569543463
transform 1 0 104 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2742
timestamp 1569543463
transform 1 0 104 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2743
timestamp 1569543463
transform 1 0 40 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2744
timestamp 1569543463
transform 1 0 232 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2745
timestamp 1569543463
transform 1 0 232 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2746
timestamp 1569543463
transform 1 0 40 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2747
timestamp 1569543463
transform 1 0 40 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2748
timestamp 1569543463
transform 1 0 40 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2749
timestamp 1569543463
transform 1 0 104 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2750
timestamp 1569543463
transform 1 0 168 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2751
timestamp 1569543463
transform 1 0 232 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2752
timestamp 1569543463
transform 1 0 296 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_2753
timestamp 1569543463
transform 1 0 232 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2754
timestamp 1569543463
transform 1 0 104 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2755
timestamp 1569543463
transform 1 0 40 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2756
timestamp 1569543463
transform 1 0 168 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2757
timestamp 1569543463
transform 1 0 296 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2758
timestamp 1569543463
transform 1 0 168 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2759
timestamp 1569543463
transform 1 0 232 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2760
timestamp 1569543463
transform 1 0 296 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2761
timestamp 1569543463
transform 1 0 168 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_2762
timestamp 1569543463
transform 1 0 168 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2763
timestamp 1569543463
transform 1 0 296 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2764
timestamp 1569543463
transform 1 0 104 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_2765
timestamp 1569543463
transform 1 0 296 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_2766
timestamp 1569543463
transform 1 0 232 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2767
timestamp 1569543463
transform 1 0 168 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2768
timestamp 1569543463
transform 1 0 168 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2769
timestamp 1569543463
transform 1 0 232 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2770
timestamp 1569543463
transform 1 0 104 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2771
timestamp 1569543463
transform 1 0 232 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2772
timestamp 1569543463
transform 1 0 168 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2773
timestamp 1569543463
transform 1 0 296 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2774
timestamp 1569543463
transform 1 0 104 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2775
timestamp 1569543463
transform 1 0 40 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2776
timestamp 1569543463
transform 1 0 296 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2777
timestamp 1569543463
transform 1 0 296 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2778
timestamp 1569543463
transform 1 0 296 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2779
timestamp 1569543463
transform 1 0 104 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2780
timestamp 1569543463
transform 1 0 232 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2781
timestamp 1569543463
transform 1 0 40 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2782
timestamp 1569543463
transform 1 0 40 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2783
timestamp 1569543463
transform 1 0 40 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2784
timestamp 1569543463
transform 1 0 168 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2785
timestamp 1569543463
transform 1 0 232 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2786
timestamp 1569543463
transform 1 0 104 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2787
timestamp 1569543463
transform 1 0 104 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2788
timestamp 1569543463
transform 1 0 296 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2789
timestamp 1569543463
transform 1 0 40 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2790
timestamp 1569543463
transform 1 0 168 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2791
timestamp 1569543463
transform 1 0 616 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2792
timestamp 1569543463
transform 1 0 616 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2793
timestamp 1569543463
transform 1 0 424 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2794
timestamp 1569543463
transform 1 0 488 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2795
timestamp 1569543463
transform 1 0 488 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2796
timestamp 1569543463
transform 1 0 424 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2797
timestamp 1569543463
transform 1 0 424 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2798
timestamp 1569543463
transform 1 0 552 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2799
timestamp 1569543463
transform 1 0 360 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2800
timestamp 1569543463
transform 1 0 424 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2801
timestamp 1569543463
transform 1 0 552 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2802
timestamp 1569543463
transform 1 0 360 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2803
timestamp 1569543463
transform 1 0 552 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2804
timestamp 1569543463
transform 1 0 360 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2805
timestamp 1569543463
transform 1 0 360 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2806
timestamp 1569543463
transform 1 0 552 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2807
timestamp 1569543463
transform 1 0 616 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2808
timestamp 1569543463
transform 1 0 616 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2809
timestamp 1569543463
transform 1 0 616 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_2810
timestamp 1569543463
transform 1 0 360 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2811
timestamp 1569543463
transform 1 0 424 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_2812
timestamp 1569543463
transform 1 0 488 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2813
timestamp 1569543463
transform 1 0 488 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2814
timestamp 1569543463
transform 1 0 552 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_2815
timestamp 1569543463
transform 1 0 488 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2816
timestamp 1569543463
transform 1 0 424 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2817
timestamp 1569543463
transform 1 0 424 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2818
timestamp 1569543463
transform 1 0 360 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2819
timestamp 1569543463
transform 1 0 616 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2820
timestamp 1569543463
transform 1 0 488 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2821
timestamp 1569543463
transform 1 0 488 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2822
timestamp 1569543463
transform 1 0 424 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2823
timestamp 1569543463
transform 1 0 360 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2824
timestamp 1569543463
transform 1 0 488 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2825
timestamp 1569543463
transform 1 0 552 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2826
timestamp 1569543463
transform 1 0 552 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2827
timestamp 1569543463
transform 1 0 360 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2828
timestamp 1569543463
transform 1 0 616 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2829
timestamp 1569543463
transform 1 0 616 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2830
timestamp 1569543463
transform 1 0 488 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2831
timestamp 1569543463
transform 1 0 360 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2832
timestamp 1569543463
transform 1 0 360 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2833
timestamp 1569543463
transform 1 0 424 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2834
timestamp 1569543463
transform 1 0 616 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2835
timestamp 1569543463
transform 1 0 552 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2836
timestamp 1569543463
transform 1 0 488 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2837
timestamp 1569543463
transform 1 0 552 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2838
timestamp 1569543463
transform 1 0 424 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2839
timestamp 1569543463
transform 1 0 616 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2840
timestamp 1569543463
transform 1 0 552 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2841
timestamp 1569543463
transform 1 0 40 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2842
timestamp 1569543463
transform 1 0 232 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2843
timestamp 1569543463
transform 1 0 104 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2844
timestamp 1569543463
transform 1 0 232 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2845
timestamp 1569543463
transform 1 0 232 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2846
timestamp 1569543463
transform 1 0 168 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2847
timestamp 1569543463
transform 1 0 296 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2848
timestamp 1569543463
transform 1 0 296 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2849
timestamp 1569543463
transform 1 0 232 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2850
timestamp 1569543463
transform 1 0 40 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2851
timestamp 1569543463
transform 1 0 296 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2852
timestamp 1569543463
transform 1 0 104 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2853
timestamp 1569543463
transform 1 0 296 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2854
timestamp 1569543463
transform 1 0 296 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2855
timestamp 1569543463
transform 1 0 104 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2856
timestamp 1569543463
transform 1 0 232 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2857
timestamp 1569543463
transform 1 0 104 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2858
timestamp 1569543463
transform 1 0 168 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2859
timestamp 1569543463
transform 1 0 104 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2860
timestamp 1569543463
transform 1 0 168 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2861
timestamp 1569543463
transform 1 0 40 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2862
timestamp 1569543463
transform 1 0 168 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2863
timestamp 1569543463
transform 1 0 40 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2864
timestamp 1569543463
transform 1 0 40 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2865
timestamp 1569543463
transform 1 0 168 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2866
timestamp 1569543463
transform 1 0 40 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2867
timestamp 1569543463
transform 1 0 232 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2868
timestamp 1569543463
transform 1 0 296 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2869
timestamp 1569543463
transform 1 0 232 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2870
timestamp 1569543463
transform 1 0 168 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2871
timestamp 1569543463
transform 1 0 168 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2872
timestamp 1569543463
transform 1 0 104 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2873
timestamp 1569543463
transform 1 0 232 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2874
timestamp 1569543463
transform 1 0 296 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2875
timestamp 1569543463
transform 1 0 296 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2876
timestamp 1569543463
transform 1 0 104 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2877
timestamp 1569543463
transform 1 0 296 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2878
timestamp 1569543463
transform 1 0 104 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2879
timestamp 1569543463
transform 1 0 232 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2880
timestamp 1569543463
transform 1 0 168 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2881
timestamp 1569543463
transform 1 0 168 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2882
timestamp 1569543463
transform 1 0 40 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2883
timestamp 1569543463
transform 1 0 40 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2884
timestamp 1569543463
transform 1 0 40 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2885
timestamp 1569543463
transform 1 0 104 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2886
timestamp 1569543463
transform 1 0 552 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2887
timestamp 1569543463
transform 1 0 424 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2888
timestamp 1569543463
transform 1 0 488 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2889
timestamp 1569543463
transform 1 0 424 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2890
timestamp 1569543463
transform 1 0 552 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2891
timestamp 1569543463
transform 1 0 360 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2892
timestamp 1569543463
transform 1 0 616 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2893
timestamp 1569543463
transform 1 0 616 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2894
timestamp 1569543463
transform 1 0 552 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2895
timestamp 1569543463
transform 1 0 616 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2896
timestamp 1569543463
transform 1 0 616 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2897
timestamp 1569543463
transform 1 0 488 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2898
timestamp 1569543463
transform 1 0 424 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2899
timestamp 1569543463
transform 1 0 488 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2900
timestamp 1569543463
transform 1 0 360 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2901
timestamp 1569543463
transform 1 0 360 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2902
timestamp 1569543463
transform 1 0 552 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2903
timestamp 1569543463
transform 1 0 424 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2904
timestamp 1569543463
transform 1 0 488 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2905
timestamp 1569543463
transform 1 0 360 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2906
timestamp 1569543463
transform 1 0 1128 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2907
timestamp 1569543463
transform 1 0 1000 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2908
timestamp 1569543463
transform 1 0 1256 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2909
timestamp 1569543463
transform 1 0 1064 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2910
timestamp 1569543463
transform 1 0 1192 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2911
timestamp 1569543463
transform 1 0 1192 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2912
timestamp 1569543463
transform 1 0 1192 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2913
timestamp 1569543463
transform 1 0 1256 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2914
timestamp 1569543463
transform 1 0 1256 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2915
timestamp 1569543463
transform 1 0 1256 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2916
timestamp 1569543463
transform 1 0 1256 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2917
timestamp 1569543463
transform 1 0 1064 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2918
timestamp 1569543463
transform 1 0 1064 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2919
timestamp 1569543463
transform 1 0 1192 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2920
timestamp 1569543463
transform 1 0 1000 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2921
timestamp 1569543463
transform 1 0 1064 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2922
timestamp 1569543463
transform 1 0 1128 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2923
timestamp 1569543463
transform 1 0 1000 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2924
timestamp 1569543463
transform 1 0 1000 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2925
timestamp 1569543463
transform 1 0 1128 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2926
timestamp 1569543463
transform 1 0 1128 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2927
timestamp 1569543463
transform 1 0 1128 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2928
timestamp 1569543463
transform 1 0 1064 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2929
timestamp 1569543463
transform 1 0 1000 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2930
timestamp 1569543463
transform 1 0 1192 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2931
timestamp 1569543463
transform 1 0 936 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2932
timestamp 1569543463
transform 1 0 808 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2933
timestamp 1569543463
transform 1 0 936 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2934
timestamp 1569543463
transform 1 0 808 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2935
timestamp 1569543463
transform 1 0 872 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2936
timestamp 1569543463
transform 1 0 936 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2937
timestamp 1569543463
transform 1 0 872 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2938
timestamp 1569543463
transform 1 0 872 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2939
timestamp 1569543463
transform 1 0 680 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2940
timestamp 1569543463
transform 1 0 680 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2941
timestamp 1569543463
transform 1 0 680 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2942
timestamp 1569543463
transform 1 0 872 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2943
timestamp 1569543463
transform 1 0 680 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2944
timestamp 1569543463
transform 1 0 680 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2945
timestamp 1569543463
transform 1 0 936 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2946
timestamp 1569543463
transform 1 0 744 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_2947
timestamp 1569543463
transform 1 0 808 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2948
timestamp 1569543463
transform 1 0 744 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2949
timestamp 1569543463
transform 1 0 808 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2950
timestamp 1569543463
transform 1 0 744 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_2951
timestamp 1569543463
transform 1 0 808 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2952
timestamp 1569543463
transform 1 0 744 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_2953
timestamp 1569543463
transform 1 0 744 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2954
timestamp 1569543463
transform 1 0 872 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_2955
timestamp 1569543463
transform 1 0 936 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_2956
timestamp 1569543463
transform 1 0 808 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2957
timestamp 1569543463
transform 1 0 872 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2958
timestamp 1569543463
transform 1 0 936 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2959
timestamp 1569543463
transform 1 0 808 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2960
timestamp 1569543463
transform 1 0 872 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2961
timestamp 1569543463
transform 1 0 872 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2962
timestamp 1569543463
transform 1 0 680 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2963
timestamp 1569543463
transform 1 0 680 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2964
timestamp 1569543463
transform 1 0 680 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2965
timestamp 1569543463
transform 1 0 680 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2966
timestamp 1569543463
transform 1 0 872 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2967
timestamp 1569543463
transform 1 0 808 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2968
timestamp 1569543463
transform 1 0 936 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2969
timestamp 1569543463
transform 1 0 744 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2970
timestamp 1569543463
transform 1 0 744 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2971
timestamp 1569543463
transform 1 0 744 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2972
timestamp 1569543463
transform 1 0 744 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2973
timestamp 1569543463
transform 1 0 936 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2974
timestamp 1569543463
transform 1 0 808 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2975
timestamp 1569543463
transform 1 0 936 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2976
timestamp 1569543463
transform 1 0 1192 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2977
timestamp 1569543463
transform 1 0 1064 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2978
timestamp 1569543463
transform 1 0 1256 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2979
timestamp 1569543463
transform 1 0 1256 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2980
timestamp 1569543463
transform 1 0 1256 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2981
timestamp 1569543463
transform 1 0 1256 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2982
timestamp 1569543463
transform 1 0 1192 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2983
timestamp 1569543463
transform 1 0 1128 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2984
timestamp 1569543463
transform 1 0 1064 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2985
timestamp 1569543463
transform 1 0 1000 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2986
timestamp 1569543463
transform 1 0 1000 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2987
timestamp 1569543463
transform 1 0 1128 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2988
timestamp 1569543463
transform 1 0 1192 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2989
timestamp 1569543463
transform 1 0 1064 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2990
timestamp 1569543463
transform 1 0 1192 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2991
timestamp 1569543463
transform 1 0 1000 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2992
timestamp 1569543463
transform 1 0 1128 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_2993
timestamp 1569543463
transform 1 0 1064 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_2994
timestamp 1569543463
transform 1 0 1000 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_2995
timestamp 1569543463
transform 1 0 1128 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_2996
timestamp 1569543463
transform 1 0 2344 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_2997
timestamp 1569543463
transform 1 0 2344 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_2998
timestamp 1569543463
transform 1 0 2344 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_2999
timestamp 1569543463
transform 1 0 2408 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3000
timestamp 1569543463
transform 1 0 2408 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3001
timestamp 1569543463
transform 1 0 2408 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3002
timestamp 1569543463
transform 1 0 2344 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3003
timestamp 1569543463
transform 1 0 2408 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3004
timestamp 1569543463
transform 1 0 2408 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3005
timestamp 1569543463
transform 1 0 2408 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3006
timestamp 1569543463
transform 1 0 2408 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3007
timestamp 1569543463
transform 1 0 2344 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3008
timestamp 1569543463
transform 1 0 2408 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3009
timestamp 1569543463
transform 1 0 2472 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3010
timestamp 1569543463
transform 1 0 2472 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3011
timestamp 1569543463
transform 1 0 2472 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3012
timestamp 1569543463
transform 1 0 2344 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3013
timestamp 1569543463
transform 1 0 2472 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3014
timestamp 1569543463
transform 1 0 2472 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3015
timestamp 1569543463
transform 1 0 2472 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3016
timestamp 1569543463
transform 1 0 2344 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3017
timestamp 1569543463
transform 1 0 2472 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3018
timestamp 1569543463
transform 1 0 2472 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3019
timestamp 1569543463
transform 1 0 2472 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3020
timestamp 1569543463
transform 1 0 2408 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3021
timestamp 1569543463
transform 1 0 2472 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3022
timestamp 1569543463
transform 1 0 2344 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3023
timestamp 1569543463
transform 1 0 2344 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3024
timestamp 1569543463
transform 1 0 2408 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3025
timestamp 1569543463
transform 1 0 2344 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3026
timestamp 1569543463
transform 1 0 1384 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3027
timestamp 1569543463
transform 1 0 1384 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3028
timestamp 1569543463
transform 1 0 1384 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3029
timestamp 1569543463
transform 1 0 1384 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3030
timestamp 1569543463
transform 1 0 1320 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3031
timestamp 1569543463
transform 1 0 1320 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3032
timestamp 1569543463
transform 1 0 1448 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3033
timestamp 1569543463
transform 1 0 1384 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3034
timestamp 1569543463
transform 1 0 1384 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3035
timestamp 1569543463
transform 1 0 1448 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3036
timestamp 1569543463
transform 1 0 1448 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3037
timestamp 1569543463
transform 1 0 1448 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3038
timestamp 1569543463
transform 1 0 1448 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3039
timestamp 1569543463
transform 1 0 1384 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3040
timestamp 1569543463
transform 1 0 1448 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3041
timestamp 1569543463
transform 1 0 1384 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3042
timestamp 1569543463
transform 1 0 1384 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3043
timestamp 1569543463
transform 1 0 1448 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3044
timestamp 1569543463
transform 1 0 1448 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3045
timestamp 1569543463
transform 1 0 1448 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3046
timestamp 1569543463
transform 1 0 1448 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3047
timestamp 1569543463
transform 1 0 1512 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3048
timestamp 1569543463
transform 1 0 1512 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3049
timestamp 1569543463
transform 1 0 1512 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3050
timestamp 1569543463
transform 1 0 1512 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3051
timestamp 1569543463
transform 1 0 1512 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3052
timestamp 1569543463
transform 1 0 1512 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3053
timestamp 1569543463
transform 1 0 1512 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3054
timestamp 1569543463
transform 1 0 1512 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3055
timestamp 1569543463
transform 1 0 1320 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3056
timestamp 1569543463
transform 1 0 1320 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3057
timestamp 1569543463
transform 1 0 1320 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3058
timestamp 1569543463
transform 1 0 1320 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3059
timestamp 1569543463
transform 1 0 1320 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3060
timestamp 1569543463
transform 1 0 1320 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3061
timestamp 1569543463
transform 1 0 1320 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3062
timestamp 1569543463
transform 1 0 1512 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3063
timestamp 1569543463
transform 1 0 1320 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3064
timestamp 1569543463
transform 1 0 1384 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3065
timestamp 1569543463
transform 1 0 1512 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3066
timestamp 1569543463
transform 1 0 1512 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3067
timestamp 1569543463
transform 1 0 1448 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3068
timestamp 1569543463
transform 1 0 1512 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3069
timestamp 1569543463
transform 1 0 1448 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3070
timestamp 1569543463
transform 1 0 1448 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3071
timestamp 1569543463
transform 1 0 1512 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3072
timestamp 1569543463
transform 1 0 1320 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3073
timestamp 1569543463
transform 1 0 1320 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3074
timestamp 1569543463
transform 1 0 1320 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3075
timestamp 1569543463
transform 1 0 1320 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3076
timestamp 1569543463
transform 1 0 1320 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3077
timestamp 1569543463
transform 1 0 1512 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3078
timestamp 1569543463
transform 1 0 1320 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3079
timestamp 1569543463
transform 1 0 1320 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3080
timestamp 1569543463
transform 1 0 1320 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3081
timestamp 1569543463
transform 1 0 1320 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3082
timestamp 1569543463
transform 1 0 1384 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3083
timestamp 1569543463
transform 1 0 1384 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3084
timestamp 1569543463
transform 1 0 1512 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3085
timestamp 1569543463
transform 1 0 1384 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3086
timestamp 1569543463
transform 1 0 1448 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3087
timestamp 1569543463
transform 1 0 1384 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3088
timestamp 1569543463
transform 1 0 1384 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3089
timestamp 1569543463
transform 1 0 1384 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3090
timestamp 1569543463
transform 1 0 1384 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3091
timestamp 1569543463
transform 1 0 1384 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3092
timestamp 1569543463
transform 1 0 1384 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3093
timestamp 1569543463
transform 1 0 1448 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3094
timestamp 1569543463
transform 1 0 1448 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3095
timestamp 1569543463
transform 1 0 1448 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3096
timestamp 1569543463
transform 1 0 1448 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3097
timestamp 1569543463
transform 1 0 1512 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3098
timestamp 1569543463
transform 1 0 1512 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3099
timestamp 1569543463
transform 1 0 1512 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3100
timestamp 1569543463
transform 1 0 1512 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3101
timestamp 1569543463
transform 1 0 1448 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3102
timestamp 1569543463
transform 1 0 2344 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3103
timestamp 1569543463
transform 1 0 2344 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3104
timestamp 1569543463
transform 1 0 2344 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3105
timestamp 1569543463
transform 1 0 2344 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3106
timestamp 1569543463
transform 1 0 2408 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3107
timestamp 1569543463
transform 1 0 2472 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3108
timestamp 1569543463
transform 1 0 2344 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_3109
timestamp 1569543463
transform 1 0 2344 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3110
timestamp 1569543463
transform 1 0 2472 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3111
timestamp 1569543463
transform 1 0 2472 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3112
timestamp 1569543463
transform 1 0 2344 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3113
timestamp 1569543463
transform 1 0 2344 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3114
timestamp 1569543463
transform 1 0 2344 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3115
timestamp 1569543463
transform 1 0 2472 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3116
timestamp 1569543463
transform 1 0 2472 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3117
timestamp 1569543463
transform 1 0 2408 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3118
timestamp 1569543463
transform 1 0 2408 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3119
timestamp 1569543463
transform 1 0 2408 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3120
timestamp 1569543463
transform 1 0 2408 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3121
timestamp 1569543463
transform 1 0 2408 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3122
timestamp 1569543463
transform 1 0 2408 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_3123
timestamp 1569543463
transform 1 0 2408 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3124
timestamp 1569543463
transform 1 0 2472 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_3125
timestamp 1569543463
transform 1 0 2408 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3126
timestamp 1569543463
transform 1 0 2472 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_3127
timestamp 1569543463
transform 1 0 2472 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3128
timestamp 1569543463
transform 1 0 2472 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3129
timestamp 1569543463
transform 1 0 4840 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3130
timestamp 1569543463
transform 1 0 4840 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3131
timestamp 1569543463
transform 1 0 4904 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3132
timestamp 1569543463
transform 1 0 4712 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3133
timestamp 1569543463
transform 1 0 4776 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3134
timestamp 1569543463
transform 1 0 4904 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3135
timestamp 1569543463
transform 1 0 4840 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3136
timestamp 1569543463
transform 1 0 4904 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3137
timestamp 1569543463
transform 1 0 4776 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3138
timestamp 1569543463
transform 1 0 4776 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3139
timestamp 1569543463
transform 1 0 4840 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3140
timestamp 1569543463
transform 1 0 4712 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3141
timestamp 1569543463
transform 1 0 4712 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3142
timestamp 1569543463
transform 1 0 4776 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3143
timestamp 1569543463
transform 1 0 4712 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3144
timestamp 1569543463
transform 1 0 4712 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3145
timestamp 1569543463
transform 1 0 4840 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3146
timestamp 1569543463
transform 1 0 4904 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3147
timestamp 1569543463
transform 1 0 4776 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3148
timestamp 1569543463
transform 1 0 4904 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3149
timestamp 1569543463
transform 1 0 4520 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3150
timestamp 1569543463
transform 1 0 4648 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3151
timestamp 1569543463
transform 1 0 4456 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3152
timestamp 1569543463
transform 1 0 4456 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3153
timestamp 1569543463
transform 1 0 4648 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3154
timestamp 1569543463
transform 1 0 4392 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3155
timestamp 1569543463
transform 1 0 4584 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3156
timestamp 1569543463
transform 1 0 4392 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3157
timestamp 1569543463
transform 1 0 4520 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3158
timestamp 1569543463
transform 1 0 4648 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3159
timestamp 1569543463
transform 1 0 4584 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3160
timestamp 1569543463
transform 1 0 4456 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3161
timestamp 1569543463
transform 1 0 4584 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3162
timestamp 1569543463
transform 1 0 4648 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3163
timestamp 1569543463
transform 1 0 4392 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3164
timestamp 1569543463
transform 1 0 4520 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3165
timestamp 1569543463
transform 1 0 4520 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3166
timestamp 1569543463
transform 1 0 4520 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3167
timestamp 1569543463
transform 1 0 4456 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3168
timestamp 1569543463
transform 1 0 4584 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3169
timestamp 1569543463
transform 1 0 4392 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3170
timestamp 1569543463
transform 1 0 4392 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3171
timestamp 1569543463
transform 1 0 4456 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3172
timestamp 1569543463
transform 1 0 4584 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3173
timestamp 1569543463
transform 1 0 4648 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3174
timestamp 1569543463
transform 1 0 4392 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3175
timestamp 1569543463
transform 1 0 4456 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3176
timestamp 1569543463
transform 1 0 4520 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3177
timestamp 1569543463
transform 1 0 4392 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3178
timestamp 1569543463
transform 1 0 4584 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3179
timestamp 1569543463
transform 1 0 4392 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3180
timestamp 1569543463
transform 1 0 4520 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3181
timestamp 1569543463
transform 1 0 4584 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3182
timestamp 1569543463
transform 1 0 4392 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3183
timestamp 1569543463
transform 1 0 4392 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3184
timestamp 1569543463
transform 1 0 4456 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3185
timestamp 1569543463
transform 1 0 4456 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3186
timestamp 1569543463
transform 1 0 4648 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3187
timestamp 1569543463
transform 1 0 4584 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3188
timestamp 1569543463
transform 1 0 4456 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3189
timestamp 1569543463
transform 1 0 4520 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3190
timestamp 1569543463
transform 1 0 4584 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3191
timestamp 1569543463
transform 1 0 4520 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3192
timestamp 1569543463
transform 1 0 4648 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3193
timestamp 1569543463
transform 1 0 4648 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3194
timestamp 1569543463
transform 1 0 4648 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3195
timestamp 1569543463
transform 1 0 4584 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3196
timestamp 1569543463
transform 1 0 4520 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3197
timestamp 1569543463
transform 1 0 4456 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3198
timestamp 1569543463
transform 1 0 4648 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3199
timestamp 1569543463
transform 1 0 4776 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3200
timestamp 1569543463
transform 1 0 4904 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3201
timestamp 1569543463
transform 1 0 4904 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3202
timestamp 1569543463
transform 1 0 4840 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3203
timestamp 1569543463
transform 1 0 4712 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3204
timestamp 1569543463
transform 1 0 4904 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3205
timestamp 1569543463
transform 1 0 4712 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3206
timestamp 1569543463
transform 1 0 4776 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3207
timestamp 1569543463
transform 1 0 4840 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3208
timestamp 1569543463
transform 1 0 4712 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3209
timestamp 1569543463
transform 1 0 4904 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3210
timestamp 1569543463
transform 1 0 4776 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3211
timestamp 1569543463
transform 1 0 4776 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3212
timestamp 1569543463
transform 1 0 4840 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3213
timestamp 1569543463
transform 1 0 4712 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3214
timestamp 1569543463
transform 1 0 4776 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3215
timestamp 1569543463
transform 1 0 4840 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3216
timestamp 1569543463
transform 1 0 4904 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3217
timestamp 1569543463
transform 1 0 4840 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3218
timestamp 1569543463
transform 1 0 4712 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3219
timestamp 1569543463
transform 1 0 4328 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3220
timestamp 1569543463
transform 1 0 4136 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3221
timestamp 1569543463
transform 1 0 4200 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3222
timestamp 1569543463
transform 1 0 4264 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3223
timestamp 1569543463
transform 1 0 4264 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3224
timestamp 1569543463
transform 1 0 4264 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3225
timestamp 1569543463
transform 1 0 4072 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3226
timestamp 1569543463
transform 1 0 4328 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3227
timestamp 1569543463
transform 1 0 4264 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3228
timestamp 1569543463
transform 1 0 4200 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3229
timestamp 1569543463
transform 1 0 4136 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3230
timestamp 1569543463
transform 1 0 4136 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3231
timestamp 1569543463
transform 1 0 4072 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3232
timestamp 1569543463
transform 1 0 4328 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3233
timestamp 1569543463
transform 1 0 4200 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3234
timestamp 1569543463
transform 1 0 4072 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3235
timestamp 1569543463
transform 1 0 4072 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3236
timestamp 1569543463
transform 1 0 4264 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3237
timestamp 1569543463
transform 1 0 4200 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3238
timestamp 1569543463
transform 1 0 4136 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3239
timestamp 1569543463
transform 1 0 4328 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3240
timestamp 1569543463
transform 1 0 4136 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3241
timestamp 1569543463
transform 1 0 4200 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3242
timestamp 1569543463
transform 1 0 4328 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3243
timestamp 1569543463
transform 1 0 4072 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3244
timestamp 1569543463
transform 1 0 3816 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3245
timestamp 1569543463
transform 1 0 3880 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3246
timestamp 1569543463
transform 1 0 3752 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3247
timestamp 1569543463
transform 1 0 4008 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3248
timestamp 1569543463
transform 1 0 3752 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3249
timestamp 1569543463
transform 1 0 3880 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3250
timestamp 1569543463
transform 1 0 3944 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3251
timestamp 1569543463
transform 1 0 3944 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3252
timestamp 1569543463
transform 1 0 3944 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3253
timestamp 1569543463
transform 1 0 4008 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3254
timestamp 1569543463
transform 1 0 3752 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3255
timestamp 1569543463
transform 1 0 3944 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3256
timestamp 1569543463
transform 1 0 3944 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3257
timestamp 1569543463
transform 1 0 3752 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3258
timestamp 1569543463
transform 1 0 4008 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3259
timestamp 1569543463
transform 1 0 3880 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3260
timestamp 1569543463
transform 1 0 3816 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3261
timestamp 1569543463
transform 1 0 4008 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3262
timestamp 1569543463
transform 1 0 3816 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3263
timestamp 1569543463
transform 1 0 3880 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3264
timestamp 1569543463
transform 1 0 4008 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3265
timestamp 1569543463
transform 1 0 3816 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3266
timestamp 1569543463
transform 1 0 3816 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3267
timestamp 1569543463
transform 1 0 3752 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3268
timestamp 1569543463
transform 1 0 3880 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3269
timestamp 1569543463
transform 1 0 3944 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3270
timestamp 1569543463
transform 1 0 3752 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3271
timestamp 1569543463
transform 1 0 4008 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3272
timestamp 1569543463
transform 1 0 3880 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3273
timestamp 1569543463
transform 1 0 3752 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3274
timestamp 1569543463
transform 1 0 3944 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3275
timestamp 1569543463
transform 1 0 3880 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3276
timestamp 1569543463
transform 1 0 3752 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3277
timestamp 1569543463
transform 1 0 3752 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3278
timestamp 1569543463
transform 1 0 3944 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3279
timestamp 1569543463
transform 1 0 3816 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3280
timestamp 1569543463
transform 1 0 3944 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3281
timestamp 1569543463
transform 1 0 4008 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3282
timestamp 1569543463
transform 1 0 3880 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3283
timestamp 1569543463
transform 1 0 3816 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3284
timestamp 1569543463
transform 1 0 3816 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3285
timestamp 1569543463
transform 1 0 3816 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3286
timestamp 1569543463
transform 1 0 3816 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3287
timestamp 1569543463
transform 1 0 4008 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3288
timestamp 1569543463
transform 1 0 3752 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3289
timestamp 1569543463
transform 1 0 4008 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3290
timestamp 1569543463
transform 1 0 4008 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3291
timestamp 1569543463
transform 1 0 3944 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3292
timestamp 1569543463
transform 1 0 3880 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3293
timestamp 1569543463
transform 1 0 3880 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3294
timestamp 1569543463
transform 1 0 4136 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3295
timestamp 1569543463
transform 1 0 4200 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3296
timestamp 1569543463
transform 1 0 4136 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3297
timestamp 1569543463
transform 1 0 4264 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3298
timestamp 1569543463
transform 1 0 4264 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3299
timestamp 1569543463
transform 1 0 4072 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3300
timestamp 1569543463
transform 1 0 4200 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3301
timestamp 1569543463
transform 1 0 4072 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3302
timestamp 1569543463
transform 1 0 4136 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3303
timestamp 1569543463
transform 1 0 4264 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3304
timestamp 1569543463
transform 1 0 4072 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3305
timestamp 1569543463
transform 1 0 4136 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3306
timestamp 1569543463
transform 1 0 4264 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3307
timestamp 1569543463
transform 1 0 4136 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3308
timestamp 1569543463
transform 1 0 4200 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3309
timestamp 1569543463
transform 1 0 4264 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3310
timestamp 1569543463
transform 1 0 4328 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3311
timestamp 1569543463
transform 1 0 4328 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3312
timestamp 1569543463
transform 1 0 4328 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3313
timestamp 1569543463
transform 1 0 4200 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3314
timestamp 1569543463
transform 1 0 4328 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3315
timestamp 1569543463
transform 1 0 4328 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3316
timestamp 1569543463
transform 1 0 4072 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3317
timestamp 1569543463
transform 1 0 4200 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3318
timestamp 1569543463
transform 1 0 4072 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3319
timestamp 1569543463
transform 1 0 4328 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3320
timestamp 1569543463
transform 1 0 4264 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3321
timestamp 1569543463
transform 1 0 4072 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3322
timestamp 1569543463
transform 1 0 4200 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3323
timestamp 1569543463
transform 1 0 4200 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3324
timestamp 1569543463
transform 1 0 4136 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3325
timestamp 1569543463
transform 1 0 4264 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3326
timestamp 1569543463
transform 1 0 4136 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3327
timestamp 1569543463
transform 1 0 4136 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3328
timestamp 1569543463
transform 1 0 4072 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3329
timestamp 1569543463
transform 1 0 4200 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3330
timestamp 1569543463
transform 1 0 4328 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3331
timestamp 1569543463
transform 1 0 4072 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3332
timestamp 1569543463
transform 1 0 4072 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3333
timestamp 1569543463
transform 1 0 4264 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3334
timestamp 1569543463
transform 1 0 4328 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3335
timestamp 1569543463
transform 1 0 4264 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3336
timestamp 1569543463
transform 1 0 4200 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3337
timestamp 1569543463
transform 1 0 4136 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3338
timestamp 1569543463
transform 1 0 4328 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3339
timestamp 1569543463
transform 1 0 3816 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3340
timestamp 1569543463
transform 1 0 3880 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3341
timestamp 1569543463
transform 1 0 3944 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3342
timestamp 1569543463
transform 1 0 3944 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3343
timestamp 1569543463
transform 1 0 3880 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3344
timestamp 1569543463
transform 1 0 3752 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3345
timestamp 1569543463
transform 1 0 3944 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3346
timestamp 1569543463
transform 1 0 3944 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3347
timestamp 1569543463
transform 1 0 4008 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3348
timestamp 1569543463
transform 1 0 3816 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3349
timestamp 1569543463
transform 1 0 3752 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3350
timestamp 1569543463
transform 1 0 4008 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3351
timestamp 1569543463
transform 1 0 4008 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3352
timestamp 1569543463
transform 1 0 3816 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3353
timestamp 1569543463
transform 1 0 3880 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3354
timestamp 1569543463
transform 1 0 3752 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3355
timestamp 1569543463
transform 1 0 3752 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3356
timestamp 1569543463
transform 1 0 4008 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3357
timestamp 1569543463
transform 1 0 3816 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3358
timestamp 1569543463
transform 1 0 3880 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3359
timestamp 1569543463
transform 1 0 3752 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3360
timestamp 1569543463
transform 1 0 4008 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3361
timestamp 1569543463
transform 1 0 3880 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3362
timestamp 1569543463
transform 1 0 4008 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3363
timestamp 1569543463
transform 1 0 3752 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3364
timestamp 1569543463
transform 1 0 3880 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3365
timestamp 1569543463
transform 1 0 3880 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3366
timestamp 1569543463
transform 1 0 3944 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3367
timestamp 1569543463
transform 1 0 3944 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3368
timestamp 1569543463
transform 1 0 4008 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3369
timestamp 1569543463
transform 1 0 3816 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3370
timestamp 1569543463
transform 1 0 4008 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3371
timestamp 1569543463
transform 1 0 3880 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3372
timestamp 1569543463
transform 1 0 3944 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3373
timestamp 1569543463
transform 1 0 3816 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3374
timestamp 1569543463
transform 1 0 3816 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3375
timestamp 1569543463
transform 1 0 3816 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3376
timestamp 1569543463
transform 1 0 3752 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3377
timestamp 1569543463
transform 1 0 3752 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3378
timestamp 1569543463
transform 1 0 3944 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3379
timestamp 1569543463
transform 1 0 4072 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3380
timestamp 1569543463
transform 1 0 4264 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3381
timestamp 1569543463
transform 1 0 4264 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3382
timestamp 1569543463
transform 1 0 4200 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3383
timestamp 1569543463
transform 1 0 4072 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3384
timestamp 1569543463
transform 1 0 4136 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3385
timestamp 1569543463
transform 1 0 4328 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3386
timestamp 1569543463
transform 1 0 4072 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3387
timestamp 1569543463
transform 1 0 4200 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3388
timestamp 1569543463
transform 1 0 4136 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3389
timestamp 1569543463
transform 1 0 4328 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3390
timestamp 1569543463
transform 1 0 4328 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3391
timestamp 1569543463
transform 1 0 4264 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3392
timestamp 1569543463
transform 1 0 4328 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3393
timestamp 1569543463
transform 1 0 4200 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3394
timestamp 1569543463
transform 1 0 4136 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3395
timestamp 1569543463
transform 1 0 4200 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3396
timestamp 1569543463
transform 1 0 4072 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3397
timestamp 1569543463
transform 1 0 4264 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3398
timestamp 1569543463
transform 1 0 4136 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3399
timestamp 1569543463
transform 1 0 4264 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3400
timestamp 1569543463
transform 1 0 4072 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3401
timestamp 1569543463
transform 1 0 4328 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3402
timestamp 1569543463
transform 1 0 3944 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3403
timestamp 1569543463
transform 1 0 4200 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3404
timestamp 1569543463
transform 1 0 4136 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3405
timestamp 1569543463
transform 1 0 3752 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3406
timestamp 1569543463
transform 1 0 4008 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3407
timestamp 1569543463
transform 1 0 3816 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3408
timestamp 1569543463
transform 1 0 3880 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3409
timestamp 1569543463
transform 1 0 4776 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3410
timestamp 1569543463
transform 1 0 4840 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3411
timestamp 1569543463
transform 1 0 4712 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3412
timestamp 1569543463
transform 1 0 4840 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3413
timestamp 1569543463
transform 1 0 4712 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3414
timestamp 1569543463
transform 1 0 4776 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3415
timestamp 1569543463
transform 1 0 4904 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3416
timestamp 1569543463
transform 1 0 4776 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3417
timestamp 1569543463
transform 1 0 4904 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3418
timestamp 1569543463
transform 1 0 4840 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3419
timestamp 1569543463
transform 1 0 4840 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3420
timestamp 1569543463
transform 1 0 4712 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3421
timestamp 1569543463
transform 1 0 4904 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3422
timestamp 1569543463
transform 1 0 4776 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3423
timestamp 1569543463
transform 1 0 4712 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3424
timestamp 1569543463
transform 1 0 4904 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3425
timestamp 1569543463
transform 1 0 4648 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3426
timestamp 1569543463
transform 1 0 4584 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3427
timestamp 1569543463
transform 1 0 4456 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3428
timestamp 1569543463
transform 1 0 4456 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3429
timestamp 1569543463
transform 1 0 4648 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3430
timestamp 1569543463
transform 1 0 4456 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3431
timestamp 1569543463
transform 1 0 4456 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3432
timestamp 1569543463
transform 1 0 4584 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3433
timestamp 1569543463
transform 1 0 4584 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3434
timestamp 1569543463
transform 1 0 4520 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3435
timestamp 1569543463
transform 1 0 4520 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3436
timestamp 1569543463
transform 1 0 4392 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3437
timestamp 1569543463
transform 1 0 4520 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3438
timestamp 1569543463
transform 1 0 4520 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3439
timestamp 1569543463
transform 1 0 4392 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3440
timestamp 1569543463
transform 1 0 4392 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3441
timestamp 1569543463
transform 1 0 4392 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3442
timestamp 1569543463
transform 1 0 4584 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3443
timestamp 1569543463
transform 1 0 4648 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3444
timestamp 1569543463
transform 1 0 4648 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3445
timestamp 1569543463
transform 1 0 4392 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3446
timestamp 1569543463
transform 1 0 4392 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3447
timestamp 1569543463
transform 1 0 4648 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3448
timestamp 1569543463
transform 1 0 4520 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3449
timestamp 1569543463
transform 1 0 4584 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3450
timestamp 1569543463
transform 1 0 4520 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3451
timestamp 1569543463
transform 1 0 4392 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3452
timestamp 1569543463
transform 1 0 4456 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3453
timestamp 1569543463
transform 1 0 4520 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3454
timestamp 1569543463
transform 1 0 4392 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3455
timestamp 1569543463
transform 1 0 4456 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3456
timestamp 1569543463
transform 1 0 4648 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3457
timestamp 1569543463
transform 1 0 4456 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3458
timestamp 1569543463
transform 1 0 4584 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3459
timestamp 1569543463
transform 1 0 4648 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3460
timestamp 1569543463
transform 1 0 4584 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3461
timestamp 1569543463
transform 1 0 4456 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3462
timestamp 1569543463
transform 1 0 4648 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3463
timestamp 1569543463
transform 1 0 4584 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3464
timestamp 1569543463
transform 1 0 4520 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3465
timestamp 1569543463
transform 1 0 4712 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3466
timestamp 1569543463
transform 1 0 4904 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3467
timestamp 1569543463
transform 1 0 4776 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3468
timestamp 1569543463
transform 1 0 4840 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3469
timestamp 1569543463
transform 1 0 4712 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3470
timestamp 1569543463
transform 1 0 4840 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3471
timestamp 1569543463
transform 1 0 4712 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3472
timestamp 1569543463
transform 1 0 4904 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3473
timestamp 1569543463
transform 1 0 4712 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3474
timestamp 1569543463
transform 1 0 4904 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3475
timestamp 1569543463
transform 1 0 4904 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3476
timestamp 1569543463
transform 1 0 4840 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3477
timestamp 1569543463
transform 1 0 4776 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3478
timestamp 1569543463
transform 1 0 4840 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3479
timestamp 1569543463
transform 1 0 4776 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3480
timestamp 1569543463
transform 1 0 4776 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3481
timestamp 1569543463
transform 1 0 4840 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3482
timestamp 1569543463
transform 1 0 4712 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3483
timestamp 1569543463
transform 1 0 4392 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3484
timestamp 1569543463
transform 1 0 4776 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3485
timestamp 1569543463
transform 1 0 4456 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3486
timestamp 1569543463
transform 1 0 4520 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3487
timestamp 1569543463
transform 1 0 4904 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3488
timestamp 1569543463
transform 1 0 4584 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3489
timestamp 1569543463
transform 1 0 4648 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3490
timestamp 1569543463
transform 1 0 3624 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3491
timestamp 1569543463
transform 1 0 3496 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3492
timestamp 1569543463
transform 1 0 3496 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3493
timestamp 1569543463
transform 1 0 3496 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3494
timestamp 1569543463
transform 1 0 3624 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3495
timestamp 1569543463
transform 1 0 3560 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3496
timestamp 1569543463
transform 1 0 3560 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3497
timestamp 1569543463
transform 1 0 3624 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3498
timestamp 1569543463
transform 1 0 3624 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3499
timestamp 1569543463
transform 1 0 3560 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3500
timestamp 1569543463
transform 1 0 3688 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3501
timestamp 1569543463
transform 1 0 3688 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3502
timestamp 1569543463
transform 1 0 3688 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3503
timestamp 1569543463
transform 1 0 3560 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3504
timestamp 1569543463
transform 1 0 3688 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3505
timestamp 1569543463
transform 1 0 3688 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3506
timestamp 1569543463
transform 1 0 3560 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3507
timestamp 1569543463
transform 1 0 3496 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3508
timestamp 1569543463
transform 1 0 3624 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3509
timestamp 1569543463
transform 1 0 3496 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3510
timestamp 1569543463
transform 1 0 3368 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3511
timestamp 1569543463
transform 1 0 3368 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3512
timestamp 1569543463
transform 1 0 3304 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3513
timestamp 1569543463
transform 1 0 3176 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3514
timestamp 1569543463
transform 1 0 3176 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3515
timestamp 1569543463
transform 1 0 3176 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3516
timestamp 1569543463
transform 1 0 3176 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3517
timestamp 1569543463
transform 1 0 3176 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3518
timestamp 1569543463
transform 1 0 3304 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3519
timestamp 1569543463
transform 1 0 3240 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3520
timestamp 1569543463
transform 1 0 3240 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3521
timestamp 1569543463
transform 1 0 3240 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3522
timestamp 1569543463
transform 1 0 3240 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3523
timestamp 1569543463
transform 1 0 3240 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3524
timestamp 1569543463
transform 1 0 3304 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3525
timestamp 1569543463
transform 1 0 3304 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3526
timestamp 1569543463
transform 1 0 3304 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3527
timestamp 1569543463
transform 1 0 3368 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3528
timestamp 1569543463
transform 1 0 3368 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3529
timestamp 1569543463
transform 1 0 3368 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3530
timestamp 1569543463
transform 1 0 3176 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3531
timestamp 1569543463
transform 1 0 3240 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3532
timestamp 1569543463
transform 1 0 3304 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3533
timestamp 1569543463
transform 1 0 3368 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3534
timestamp 1569543463
transform 1 0 3304 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3535
timestamp 1569543463
transform 1 0 3304 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3536
timestamp 1569543463
transform 1 0 3176 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3537
timestamp 1569543463
transform 1 0 3368 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3538
timestamp 1569543463
transform 1 0 3368 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3539
timestamp 1569543463
transform 1 0 3368 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3540
timestamp 1569543463
transform 1 0 3176 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3541
timestamp 1569543463
transform 1 0 3368 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3542
timestamp 1569543463
transform 1 0 3304 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3543
timestamp 1569543463
transform 1 0 3240 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3544
timestamp 1569543463
transform 1 0 3240 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3545
timestamp 1569543463
transform 1 0 3240 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3546
timestamp 1569543463
transform 1 0 3240 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3547
timestamp 1569543463
transform 1 0 3304 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3548
timestamp 1569543463
transform 1 0 3176 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3549
timestamp 1569543463
transform 1 0 3176 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3550
timestamp 1569543463
transform 1 0 3688 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3551
timestamp 1569543463
transform 1 0 3624 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3552
timestamp 1569543463
transform 1 0 3688 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3553
timestamp 1569543463
transform 1 0 3496 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3554
timestamp 1569543463
transform 1 0 3496 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3555
timestamp 1569543463
transform 1 0 3688 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3556
timestamp 1569543463
transform 1 0 3496 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3557
timestamp 1569543463
transform 1 0 3496 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3558
timestamp 1569543463
transform 1 0 3688 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3559
timestamp 1569543463
transform 1 0 3688 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3560
timestamp 1569543463
transform 1 0 3560 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3561
timestamp 1569543463
transform 1 0 3496 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3562
timestamp 1569543463
transform 1 0 3560 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3563
timestamp 1569543463
transform 1 0 3560 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3564
timestamp 1569543463
transform 1 0 3560 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3565
timestamp 1569543463
transform 1 0 3560 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3566
timestamp 1569543463
transform 1 0 3624 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3567
timestamp 1569543463
transform 1 0 3624 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3568
timestamp 1569543463
transform 1 0 3624 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3569
timestamp 1569543463
transform 1 0 3624 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3570
timestamp 1569543463
transform 1 0 3432 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3571
timestamp 1569543463
transform 1 0 3432 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3572
timestamp 1569543463
transform 1 0 3432 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3573
timestamp 1569543463
transform 1 0 3432 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3574
timestamp 1569543463
transform 1 0 3432 0 1 2536
box -8 -8 8 8
use VIA2$5  VIA2$5_3575
timestamp 1569543463
transform 1 0 3432 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3576
timestamp 1569543463
transform 1 0 3432 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3577
timestamp 1569543463
transform 1 0 3432 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3578
timestamp 1569543463
transform 1 0 3432 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3579
timestamp 1569543463
transform 1 0 3432 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3580
timestamp 1569543463
transform 1 0 3048 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3581
timestamp 1569543463
transform 1 0 3048 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3582
timestamp 1569543463
transform 1 0 3112 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3583
timestamp 1569543463
transform 1 0 2600 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3584
timestamp 1569543463
transform 1 0 2856 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3585
timestamp 1569543463
transform 1 0 2856 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3586
timestamp 1569543463
transform 1 0 2856 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3587
timestamp 1569543463
transform 1 0 2856 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3588
timestamp 1569543463
transform 1 0 2792 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3589
timestamp 1569543463
transform 1 0 2792 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3590
timestamp 1569543463
transform 1 0 2792 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3591
timestamp 1569543463
transform 1 0 2792 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3592
timestamp 1569543463
transform 1 0 3112 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3593
timestamp 1569543463
transform 1 0 3112 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3594
timestamp 1569543463
transform 1 0 2920 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3595
timestamp 1569543463
transform 1 0 2920 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3596
timestamp 1569543463
transform 1 0 2920 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3597
timestamp 1569543463
transform 1 0 2920 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3598
timestamp 1569543463
transform 1 0 3112 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3599
timestamp 1569543463
transform 1 0 3048 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3600
timestamp 1569543463
transform 1 0 3048 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3601
timestamp 1569543463
transform 1 0 3048 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3602
timestamp 1569543463
transform 1 0 3048 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3603
timestamp 1569543463
transform 1 0 3112 0 1 2600
box -8 -8 8 8
use VIA2$5  VIA2$5_3604
timestamp 1569543463
transform 1 0 2664 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3605
timestamp 1569543463
transform 1 0 2664 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3606
timestamp 1569543463
transform 1 0 3112 0 1 2664
box -8 -8 8 8
use VIA2$5  VIA2$5_3607
timestamp 1569543463
transform 1 0 3112 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3608
timestamp 1569543463
transform 1 0 3112 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3609
timestamp 1569543463
transform 1 0 3112 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3610
timestamp 1569543463
transform 1 0 2856 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3611
timestamp 1569543463
transform 1 0 2920 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3612
timestamp 1569543463
transform 1 0 2920 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3613
timestamp 1569543463
transform 1 0 2984 0 1 2728
box -8 -8 8 8
use VIA2$5  VIA2$5_3614
timestamp 1569543463
transform 1 0 2984 0 1 2792
box -8 -8 8 8
use VIA2$5  VIA2$5_3615
timestamp 1569543463
transform 1 0 2984 0 1 2856
box -8 -8 8 8
use VIA2$5  VIA2$5_3616
timestamp 1569543463
transform 1 0 2728 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3617
timestamp 1569543463
transform 1 0 2728 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3618
timestamp 1569543463
transform 1 0 2984 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3619
timestamp 1569543463
transform 1 0 2984 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3620
timestamp 1569543463
transform 1 0 2984 0 1 3048
box -8 -8 8 8
use VIA2$5  VIA2$5_3621
timestamp 1569543463
transform 1 0 2984 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3622
timestamp 1569543463
transform 1 0 2728 0 1 3112
box -8 -8 8 8
use VIA2$5  VIA2$5_3623
timestamp 1569543463
transform 1 0 3048 0 1 2920
box -8 -8 8 8
use VIA2$5  VIA2$5_3624
timestamp 1569543463
transform 1 0 3048 0 1 2984
box -8 -8 8 8
use VIA2$5  VIA2$5_3625
timestamp 1569543463
transform 1 0 2984 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3626
timestamp 1569543463
transform 1 0 2984 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3627
timestamp 1569543463
transform 1 0 2920 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3628
timestamp 1569543463
transform 1 0 3112 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3629
timestamp 1569543463
transform 1 0 3048 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3630
timestamp 1569543463
transform 1 0 3112 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3631
timestamp 1569543463
transform 1 0 2920 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3632
timestamp 1569543463
transform 1 0 2920 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3633
timestamp 1569543463
transform 1 0 3048 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3634
timestamp 1569543463
transform 1 0 2856 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3635
timestamp 1569543463
transform 1 0 3112 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3636
timestamp 1569543463
transform 1 0 2920 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3637
timestamp 1569543463
transform 1 0 3048 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3638
timestamp 1569543463
transform 1 0 2856 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3639
timestamp 1569543463
transform 1 0 2856 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3640
timestamp 1569543463
transform 1 0 2856 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3641
timestamp 1569543463
transform 1 0 2984 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3642
timestamp 1569543463
transform 1 0 3048 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3643
timestamp 1569543463
transform 1 0 3112 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3644
timestamp 1569543463
transform 1 0 2984 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3645
timestamp 1569543463
transform 1 0 2600 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3646
timestamp 1569543463
transform 1 0 2600 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3647
timestamp 1569543463
transform 1 0 2792 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3648
timestamp 1569543463
transform 1 0 2600 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3649
timestamp 1569543463
transform 1 0 2536 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3650
timestamp 1569543463
transform 1 0 2536 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3651
timestamp 1569543463
transform 1 0 2728 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3652
timestamp 1569543463
transform 1 0 2792 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3653
timestamp 1569543463
transform 1 0 2728 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3654
timestamp 1569543463
transform 1 0 2600 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3655
timestamp 1569543463
transform 1 0 2536 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3656
timestamp 1569543463
transform 1 0 2728 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3657
timestamp 1569543463
transform 1 0 2664 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3658
timestamp 1569543463
transform 1 0 2792 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3659
timestamp 1569543463
transform 1 0 2664 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3660
timestamp 1569543463
transform 1 0 2536 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3661
timestamp 1569543463
transform 1 0 2728 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3662
timestamp 1569543463
transform 1 0 2664 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3663
timestamp 1569543463
transform 1 0 2792 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3664
timestamp 1569543463
transform 1 0 2664 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3665
timestamp 1569543463
transform 1 0 2600 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3666
timestamp 1569543463
transform 1 0 2536 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3667
timestamp 1569543463
transform 1 0 2728 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3668
timestamp 1569543463
transform 1 0 2728 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3669
timestamp 1569543463
transform 1 0 2792 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3670
timestamp 1569543463
transform 1 0 2536 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3671
timestamp 1569543463
transform 1 0 2728 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3672
timestamp 1569543463
transform 1 0 2792 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3673
timestamp 1569543463
transform 1 0 2728 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3674
timestamp 1569543463
transform 1 0 2792 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3675
timestamp 1569543463
transform 1 0 2792 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3676
timestamp 1569543463
transform 1 0 2600 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3677
timestamp 1569543463
transform 1 0 2664 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3678
timestamp 1569543463
transform 1 0 2664 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3679
timestamp 1569543463
transform 1 0 2664 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3680
timestamp 1569543463
transform 1 0 2536 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3681
timestamp 1569543463
transform 1 0 2600 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3682
timestamp 1569543463
transform 1 0 2664 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3683
timestamp 1569543463
transform 1 0 2536 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3684
timestamp 1569543463
transform 1 0 2600 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3685
timestamp 1569543463
transform 1 0 2856 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3686
timestamp 1569543463
transform 1 0 2984 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3687
timestamp 1569543463
transform 1 0 2984 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3688
timestamp 1569543463
transform 1 0 2984 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3689
timestamp 1569543463
transform 1 0 2856 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3690
timestamp 1569543463
transform 1 0 2856 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3691
timestamp 1569543463
transform 1 0 3048 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3692
timestamp 1569543463
transform 1 0 2984 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3693
timestamp 1569543463
transform 1 0 3048 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3694
timestamp 1569543463
transform 1 0 2920 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3695
timestamp 1569543463
transform 1 0 2920 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3696
timestamp 1569543463
transform 1 0 3112 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3697
timestamp 1569543463
transform 1 0 2920 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3698
timestamp 1569543463
transform 1 0 3048 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3699
timestamp 1569543463
transform 1 0 3048 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3700
timestamp 1569543463
transform 1 0 3112 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3701
timestamp 1569543463
transform 1 0 3112 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3702
timestamp 1569543463
transform 1 0 2920 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3703
timestamp 1569543463
transform 1 0 3112 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3704
timestamp 1569543463
transform 1 0 2856 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3705
timestamp 1569543463
transform 1 0 2984 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3706
timestamp 1569543463
transform 1 0 3048 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3707
timestamp 1569543463
transform 1 0 2728 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3708
timestamp 1569543463
transform 1 0 2600 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3709
timestamp 1569543463
transform 1 0 2792 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3710
timestamp 1569543463
transform 1 0 2664 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3711
timestamp 1569543463
transform 1 0 3112 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3712
timestamp 1569543463
transform 1 0 2856 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3713
timestamp 1569543463
transform 1 0 2920 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3714
timestamp 1569543463
transform 1 0 2536 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3715
timestamp 1569543463
transform 1 0 3688 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3716
timestamp 1569543463
transform 1 0 3496 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3717
timestamp 1569543463
transform 1 0 3496 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3718
timestamp 1569543463
transform 1 0 3496 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3719
timestamp 1569543463
transform 1 0 3496 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3720
timestamp 1569543463
transform 1 0 3688 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3721
timestamp 1569543463
transform 1 0 3560 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3722
timestamp 1569543463
transform 1 0 3560 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3723
timestamp 1569543463
transform 1 0 3560 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3724
timestamp 1569543463
transform 1 0 3560 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3725
timestamp 1569543463
transform 1 0 3688 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3726
timestamp 1569543463
transform 1 0 3624 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3727
timestamp 1569543463
transform 1 0 3624 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3728
timestamp 1569543463
transform 1 0 3688 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3729
timestamp 1569543463
transform 1 0 3624 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3730
timestamp 1569543463
transform 1 0 3624 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3731
timestamp 1569543463
transform 1 0 3304 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3732
timestamp 1569543463
transform 1 0 3176 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3733
timestamp 1569543463
transform 1 0 3176 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3734
timestamp 1569543463
transform 1 0 3304 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3735
timestamp 1569543463
transform 1 0 3304 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3736
timestamp 1569543463
transform 1 0 3304 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3737
timestamp 1569543463
transform 1 0 3176 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3738
timestamp 1569543463
transform 1 0 3176 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3739
timestamp 1569543463
transform 1 0 3240 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3740
timestamp 1569543463
transform 1 0 3240 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3741
timestamp 1569543463
transform 1 0 3240 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3742
timestamp 1569543463
transform 1 0 3240 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3743
timestamp 1569543463
transform 1 0 3368 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3744
timestamp 1569543463
transform 1 0 3368 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3745
timestamp 1569543463
transform 1 0 3368 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3746
timestamp 1569543463
transform 1 0 3368 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3747
timestamp 1569543463
transform 1 0 3176 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3748
timestamp 1569543463
transform 1 0 3176 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3749
timestamp 1569543463
transform 1 0 3368 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3750
timestamp 1569543463
transform 1 0 3240 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3751
timestamp 1569543463
transform 1 0 3240 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3752
timestamp 1569543463
transform 1 0 3240 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3753
timestamp 1569543463
transform 1 0 3240 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3754
timestamp 1569543463
transform 1 0 3368 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3755
timestamp 1569543463
transform 1 0 3368 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3756
timestamp 1569543463
transform 1 0 3176 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3757
timestamp 1569543463
transform 1 0 3176 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3758
timestamp 1569543463
transform 1 0 3304 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3759
timestamp 1569543463
transform 1 0 3304 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3760
timestamp 1569543463
transform 1 0 3304 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3761
timestamp 1569543463
transform 1 0 3304 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3762
timestamp 1569543463
transform 1 0 3368 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3763
timestamp 1569543463
transform 1 0 3688 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3764
timestamp 1569543463
transform 1 0 3688 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3765
timestamp 1569543463
transform 1 0 3688 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3766
timestamp 1569543463
transform 1 0 3688 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3767
timestamp 1569543463
transform 1 0 3496 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3768
timestamp 1569543463
transform 1 0 3496 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3769
timestamp 1569543463
transform 1 0 3560 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3770
timestamp 1569543463
transform 1 0 3560 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3771
timestamp 1569543463
transform 1 0 3624 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3772
timestamp 1569543463
transform 1 0 3624 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3773
timestamp 1569543463
transform 1 0 3496 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3774
timestamp 1569543463
transform 1 0 3496 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3775
timestamp 1569543463
transform 1 0 3624 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3776
timestamp 1569543463
transform 1 0 3624 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3777
timestamp 1569543463
transform 1 0 3560 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3778
timestamp 1569543463
transform 1 0 3560 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3779
timestamp 1569543463
transform 1 0 3240 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3780
timestamp 1569543463
transform 1 0 3304 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3781
timestamp 1569543463
transform 1 0 3432 0 1 3560
box -8 -8 8 8
use VIA2$5  VIA2$5_3782
timestamp 1569543463
transform 1 0 3496 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3783
timestamp 1569543463
transform 1 0 3560 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3784
timestamp 1569543463
transform 1 0 3624 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3785
timestamp 1569543463
transform 1 0 3432 0 1 3624
box -8 -8 8 8
use VIA2$5  VIA2$5_3786
timestamp 1569543463
transform 1 0 3432 0 1 3688
box -8 -8 8 8
use VIA2$5  VIA2$5_3787
timestamp 1569543463
transform 1 0 3368 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3788
timestamp 1569543463
transform 1 0 3432 0 1 3176
box -8 -8 8 8
use VIA2$5  VIA2$5_3789
timestamp 1569543463
transform 1 0 3432 0 1 3240
box -8 -8 8 8
use VIA2$5  VIA2$5_3790
timestamp 1569543463
transform 1 0 3432 0 1 3304
box -8 -8 8 8
use VIA2$5  VIA2$5_3791
timestamp 1569543463
transform 1 0 3432 0 1 3368
box -8 -8 8 8
use VIA2$5  VIA2$5_3792
timestamp 1569543463
transform 1 0 3432 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3793
timestamp 1569543463
transform 1 0 3432 0 1 3496
box -8 -8 8 8
use VIA2$5  VIA2$5_3794
timestamp 1569543463
transform 1 0 3688 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3795
timestamp 1569543463
transform 1 0 3176 0 1 3432
box -8 -8 8 8
use VIA2$5  VIA2$5_3796
timestamp 1569543463
transform 1 0 3688 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3797
timestamp 1569543463
transform 1 0 3624 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3798
timestamp 1569543463
transform 1 0 3560 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3799
timestamp 1569543463
transform 1 0 3496 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3800
timestamp 1569543463
transform 1 0 3688 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3801
timestamp 1569543463
transform 1 0 3624 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3802
timestamp 1569543463
transform 1 0 3688 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3803
timestamp 1569543463
transform 1 0 3624 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3804
timestamp 1569543463
transform 1 0 3496 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3805
timestamp 1569543463
transform 1 0 3560 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3806
timestamp 1569543463
transform 1 0 3496 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3807
timestamp 1569543463
transform 1 0 3560 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3808
timestamp 1569543463
transform 1 0 3624 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3809
timestamp 1569543463
transform 1 0 3560 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3810
timestamp 1569543463
transform 1 0 3688 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3811
timestamp 1569543463
transform 1 0 3560 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3812
timestamp 1569543463
transform 1 0 3688 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3813
timestamp 1569543463
transform 1 0 3624 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3814
timestamp 1569543463
transform 1 0 3496 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3815
timestamp 1569543463
transform 1 0 3496 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3816
timestamp 1569543463
transform 1 0 3368 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3817
timestamp 1569543463
transform 1 0 3368 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3818
timestamp 1569543463
transform 1 0 3240 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3819
timestamp 1569543463
transform 1 0 3176 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3820
timestamp 1569543463
transform 1 0 3240 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3821
timestamp 1569543463
transform 1 0 3240 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3822
timestamp 1569543463
transform 1 0 3304 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3823
timestamp 1569543463
transform 1 0 3176 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3824
timestamp 1569543463
transform 1 0 3368 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3825
timestamp 1569543463
transform 1 0 3304 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3826
timestamp 1569543463
transform 1 0 3304 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3827
timestamp 1569543463
transform 1 0 3304 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3828
timestamp 1569543463
transform 1 0 3240 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3829
timestamp 1569543463
transform 1 0 3176 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3830
timestamp 1569543463
transform 1 0 3176 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3831
timestamp 1569543463
transform 1 0 3368 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3832
timestamp 1569543463
transform 1 0 3304 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3833
timestamp 1569543463
transform 1 0 3368 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3834
timestamp 1569543463
transform 1 0 3176 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3835
timestamp 1569543463
transform 1 0 3240 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3836
timestamp 1569543463
transform 1 0 3304 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3837
timestamp 1569543463
transform 1 0 3240 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3838
timestamp 1569543463
transform 1 0 3176 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3839
timestamp 1569543463
transform 1 0 3240 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3840
timestamp 1569543463
transform 1 0 3176 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3841
timestamp 1569543463
transform 1 0 3176 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3842
timestamp 1569543463
transform 1 0 3368 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3843
timestamp 1569543463
transform 1 0 3304 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3844
timestamp 1569543463
transform 1 0 3240 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3845
timestamp 1569543463
transform 1 0 3240 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3846
timestamp 1569543463
transform 1 0 3368 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3847
timestamp 1569543463
transform 1 0 3176 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3848
timestamp 1569543463
transform 1 0 3304 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3849
timestamp 1569543463
transform 1 0 3368 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3850
timestamp 1569543463
transform 1 0 3304 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3851
timestamp 1569543463
transform 1 0 3304 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3852
timestamp 1569543463
transform 1 0 3240 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3853
timestamp 1569543463
transform 1 0 3368 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3854
timestamp 1569543463
transform 1 0 3176 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3855
timestamp 1569543463
transform 1 0 3368 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3856
timestamp 1569543463
transform 1 0 3624 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3857
timestamp 1569543463
transform 1 0 3624 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3858
timestamp 1569543463
transform 1 0 3688 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3859
timestamp 1569543463
transform 1 0 3496 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3860
timestamp 1569543463
transform 1 0 3624 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3861
timestamp 1569543463
transform 1 0 3688 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3862
timestamp 1569543463
transform 1 0 3560 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3863
timestamp 1569543463
transform 1 0 3688 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3864
timestamp 1569543463
transform 1 0 3688 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3865
timestamp 1569543463
transform 1 0 3496 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3866
timestamp 1569543463
transform 1 0 3688 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3867
timestamp 1569543463
transform 1 0 3624 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3868
timestamp 1569543463
transform 1 0 3496 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3869
timestamp 1569543463
transform 1 0 3496 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3870
timestamp 1569543463
transform 1 0 3560 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3871
timestamp 1569543463
transform 1 0 3560 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3872
timestamp 1569543463
transform 1 0 3496 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3873
timestamp 1569543463
transform 1 0 3560 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3874
timestamp 1569543463
transform 1 0 3560 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3875
timestamp 1569543463
transform 1 0 3624 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3876
timestamp 1569543463
transform 1 0 3432 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3877
timestamp 1569543463
transform 1 0 3432 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3878
timestamp 1569543463
transform 1 0 3432 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3879
timestamp 1569543463
transform 1 0 3432 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3880
timestamp 1569543463
transform 1 0 3432 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3881
timestamp 1569543463
transform 1 0 3432 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3882
timestamp 1569543463
transform 1 0 3432 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3883
timestamp 1569543463
transform 1 0 3432 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3884
timestamp 1569543463
transform 1 0 3432 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3885
timestamp 1569543463
transform 1 0 3432 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3886
timestamp 1569543463
transform 1 0 2984 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3887
timestamp 1569543463
transform 1 0 3112 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3888
timestamp 1569543463
transform 1 0 2984 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3889
timestamp 1569543463
transform 1 0 2920 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3890
timestamp 1569543463
transform 1 0 3112 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3891
timestamp 1569543463
transform 1 0 2920 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3892
timestamp 1569543463
transform 1 0 2856 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3893
timestamp 1569543463
transform 1 0 2984 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3894
timestamp 1569543463
transform 1 0 2984 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3895
timestamp 1569543463
transform 1 0 2984 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3896
timestamp 1569543463
transform 1 0 3112 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3897
timestamp 1569543463
transform 1 0 2856 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3898
timestamp 1569543463
transform 1 0 3048 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3899
timestamp 1569543463
transform 1 0 2856 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3900
timestamp 1569543463
transform 1 0 2920 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3901
timestamp 1569543463
transform 1 0 2920 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3902
timestamp 1569543463
transform 1 0 3048 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3903
timestamp 1569543463
transform 1 0 3112 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3904
timestamp 1569543463
transform 1 0 2856 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3905
timestamp 1569543463
transform 1 0 3048 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3906
timestamp 1569543463
transform 1 0 3048 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3907
timestamp 1569543463
transform 1 0 3112 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3908
timestamp 1569543463
transform 1 0 3048 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3909
timestamp 1569543463
transform 1 0 2920 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3910
timestamp 1569543463
transform 1 0 2856 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3911
timestamp 1569543463
transform 1 0 2664 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3912
timestamp 1569543463
transform 1 0 2536 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3913
timestamp 1569543463
transform 1 0 2728 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3914
timestamp 1569543463
transform 1 0 2536 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3915
timestamp 1569543463
transform 1 0 2728 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3916
timestamp 1569543463
transform 1 0 2536 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3917
timestamp 1569543463
transform 1 0 2728 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3918
timestamp 1569543463
transform 1 0 2600 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3919
timestamp 1569543463
transform 1 0 2600 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3920
timestamp 1569543463
transform 1 0 2664 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3921
timestamp 1569543463
transform 1 0 2600 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3922
timestamp 1569543463
transform 1 0 2664 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3923
timestamp 1569543463
transform 1 0 2728 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3924
timestamp 1569543463
transform 1 0 2728 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3925
timestamp 1569543463
transform 1 0 2600 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3926
timestamp 1569543463
transform 1 0 2664 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3927
timestamp 1569543463
transform 1 0 2792 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3928
timestamp 1569543463
transform 1 0 2600 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3929
timestamp 1569543463
transform 1 0 2792 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3930
timestamp 1569543463
transform 1 0 2536 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3931
timestamp 1569543463
transform 1 0 2792 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_3932
timestamp 1569543463
transform 1 0 2664 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_3933
timestamp 1569543463
transform 1 0 2536 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_3934
timestamp 1569543463
transform 1 0 2792 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_3935
timestamp 1569543463
transform 1 0 2792 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_3936
timestamp 1569543463
transform 1 0 2792 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3937
timestamp 1569543463
transform 1 0 2664 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3938
timestamp 1569543463
transform 1 0 2536 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3939
timestamp 1569543463
transform 1 0 2536 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3940
timestamp 1569543463
transform 1 0 2600 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3941
timestamp 1569543463
transform 1 0 2600 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3942
timestamp 1569543463
transform 1 0 2728 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3943
timestamp 1569543463
transform 1 0 2600 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3944
timestamp 1569543463
transform 1 0 2664 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3945
timestamp 1569543463
transform 1 0 2728 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3946
timestamp 1569543463
transform 1 0 2792 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3947
timestamp 1569543463
transform 1 0 2792 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3948
timestamp 1569543463
transform 1 0 2728 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3949
timestamp 1569543463
transform 1 0 2664 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3950
timestamp 1569543463
transform 1 0 2792 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3951
timestamp 1569543463
transform 1 0 2536 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3952
timestamp 1569543463
transform 1 0 2792 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3953
timestamp 1569543463
transform 1 0 2536 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3954
timestamp 1569543463
transform 1 0 2536 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3955
timestamp 1569543463
transform 1 0 2728 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3956
timestamp 1569543463
transform 1 0 2600 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3957
timestamp 1569543463
transform 1 0 2664 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3958
timestamp 1569543463
transform 1 0 2664 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3959
timestamp 1569543463
transform 1 0 2728 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3960
timestamp 1569543463
transform 1 0 2600 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3961
timestamp 1569543463
transform 1 0 2856 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3962
timestamp 1569543463
transform 1 0 2984 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3963
timestamp 1569543463
transform 1 0 2984 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3964
timestamp 1569543463
transform 1 0 3112 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3965
timestamp 1569543463
transform 1 0 3112 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3966
timestamp 1569543463
transform 1 0 2984 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3967
timestamp 1569543463
transform 1 0 2920 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3968
timestamp 1569543463
transform 1 0 2920 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3969
timestamp 1569543463
transform 1 0 3048 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3970
timestamp 1569543463
transform 1 0 3048 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3971
timestamp 1569543463
transform 1 0 2920 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3972
timestamp 1569543463
transform 1 0 2920 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3973
timestamp 1569543463
transform 1 0 2920 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3974
timestamp 1569543463
transform 1 0 2984 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3975
timestamp 1569543463
transform 1 0 2984 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_3976
timestamp 1569543463
transform 1 0 3048 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3977
timestamp 1569543463
transform 1 0 3048 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3978
timestamp 1569543463
transform 1 0 3048 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3979
timestamp 1569543463
transform 1 0 3112 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3980
timestamp 1569543463
transform 1 0 3112 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3981
timestamp 1569543463
transform 1 0 3112 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3982
timestamp 1569543463
transform 1 0 2856 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_3983
timestamp 1569543463
transform 1 0 2856 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_3984
timestamp 1569543463
transform 1 0 2856 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_3985
timestamp 1569543463
transform 1 0 2856 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_3986
timestamp 1569543463
transform 1 0 2856 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3987
timestamp 1569543463
transform 1 0 3112 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3988
timestamp 1569543463
transform 1 0 2920 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3989
timestamp 1569543463
transform 1 0 3048 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3990
timestamp 1569543463
transform 1 0 2920 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_3991
timestamp 1569543463
transform 1 0 3048 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3992
timestamp 1569543463
transform 1 0 3112 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3993
timestamp 1569543463
transform 1 0 3048 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_3994
timestamp 1569543463
transform 1 0 2856 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_3995
timestamp 1569543463
transform 1 0 2920 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3996
timestamp 1569543463
transform 1 0 2984 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_3997
timestamp 1569543463
transform 1 0 2856 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3998
timestamp 1569543463
transform 1 0 3112 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_3999
timestamp 1569543463
transform 1 0 2984 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4000
timestamp 1569543463
transform 1 0 2920 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4001
timestamp 1569543463
transform 1 0 3048 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4002
timestamp 1569543463
transform 1 0 2920 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4003
timestamp 1569543463
transform 1 0 2984 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4004
timestamp 1569543463
transform 1 0 2856 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4005
timestamp 1569543463
transform 1 0 3048 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4006
timestamp 1569543463
transform 1 0 2984 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4007
timestamp 1569543463
transform 1 0 2856 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4008
timestamp 1569543463
transform 1 0 3112 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4009
timestamp 1569543463
transform 1 0 2984 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4010
timestamp 1569543463
transform 1 0 3112 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4011
timestamp 1569543463
transform 1 0 2536 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4012
timestamp 1569543463
transform 1 0 2600 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4013
timestamp 1569543463
transform 1 0 2664 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4014
timestamp 1569543463
transform 1 0 2664 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4015
timestamp 1569543463
transform 1 0 2536 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4016
timestamp 1569543463
transform 1 0 2728 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4017
timestamp 1569543463
transform 1 0 2664 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4018
timestamp 1569543463
transform 1 0 2536 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4019
timestamp 1569543463
transform 1 0 2728 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4020
timestamp 1569543463
transform 1 0 2664 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4021
timestamp 1569543463
transform 1 0 2536 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4022
timestamp 1569543463
transform 1 0 2664 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4023
timestamp 1569543463
transform 1 0 2536 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4024
timestamp 1569543463
transform 1 0 2792 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4025
timestamp 1569543463
transform 1 0 2600 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4026
timestamp 1569543463
transform 1 0 2728 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4027
timestamp 1569543463
transform 1 0 2728 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4028
timestamp 1569543463
transform 1 0 2600 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4029
timestamp 1569543463
transform 1 0 2792 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4030
timestamp 1569543463
transform 1 0 2792 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4031
timestamp 1569543463
transform 1 0 2728 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4032
timestamp 1569543463
transform 1 0 2600 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4033
timestamp 1569543463
transform 1 0 2792 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4034
timestamp 1569543463
transform 1 0 2600 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4035
timestamp 1569543463
transform 1 0 2792 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4036
timestamp 1569543463
transform 1 0 2536 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4037
timestamp 1569543463
transform 1 0 2792 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4038
timestamp 1569543463
transform 1 0 2664 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4039
timestamp 1569543463
transform 1 0 2664 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4040
timestamp 1569543463
transform 1 0 2728 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4041
timestamp 1569543463
transform 1 0 2664 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4042
timestamp 1569543463
transform 1 0 2728 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4043
timestamp 1569543463
transform 1 0 2600 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4044
timestamp 1569543463
transform 1 0 2536 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4045
timestamp 1569543463
transform 1 0 2600 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4046
timestamp 1569543463
transform 1 0 2664 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4047
timestamp 1569543463
transform 1 0 2792 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4048
timestamp 1569543463
transform 1 0 2536 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4049
timestamp 1569543463
transform 1 0 2728 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4050
timestamp 1569543463
transform 1 0 2536 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4051
timestamp 1569543463
transform 1 0 2728 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4052
timestamp 1569543463
transform 1 0 2792 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4053
timestamp 1569543463
transform 1 0 2600 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4054
timestamp 1569543463
transform 1 0 2600 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4055
timestamp 1569543463
transform 1 0 2792 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4056
timestamp 1569543463
transform 1 0 3112 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4057
timestamp 1569543463
transform 1 0 2920 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4058
timestamp 1569543463
transform 1 0 2920 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4059
timestamp 1569543463
transform 1 0 2984 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4060
timestamp 1569543463
transform 1 0 2984 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4061
timestamp 1569543463
transform 1 0 2984 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4062
timestamp 1569543463
transform 1 0 3048 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4063
timestamp 1569543463
transform 1 0 3112 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4064
timestamp 1569543463
transform 1 0 3112 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4065
timestamp 1569543463
transform 1 0 3048 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4066
timestamp 1569543463
transform 1 0 2856 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4067
timestamp 1569543463
transform 1 0 2920 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4068
timestamp 1569543463
transform 1 0 3048 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4069
timestamp 1569543463
transform 1 0 2984 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4070
timestamp 1569543463
transform 1 0 3112 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4071
timestamp 1569543463
transform 1 0 3048 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4072
timestamp 1569543463
transform 1 0 2856 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4073
timestamp 1569543463
transform 1 0 2856 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4074
timestamp 1569543463
transform 1 0 2856 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4075
timestamp 1569543463
transform 1 0 2920 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4076
timestamp 1569543463
transform 1 0 3496 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4077
timestamp 1569543463
transform 1 0 3496 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4078
timestamp 1569543463
transform 1 0 3496 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4079
timestamp 1569543463
transform 1 0 3688 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4080
timestamp 1569543463
transform 1 0 3688 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4081
timestamp 1569543463
transform 1 0 3688 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4082
timestamp 1569543463
transform 1 0 3560 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4083
timestamp 1569543463
transform 1 0 3560 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4084
timestamp 1569543463
transform 1 0 3560 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4085
timestamp 1569543463
transform 1 0 3560 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4086
timestamp 1569543463
transform 1 0 3560 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4087
timestamp 1569543463
transform 1 0 3688 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4088
timestamp 1569543463
transform 1 0 3688 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4089
timestamp 1569543463
transform 1 0 3624 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4090
timestamp 1569543463
transform 1 0 3624 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4091
timestamp 1569543463
transform 1 0 3624 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4092
timestamp 1569543463
transform 1 0 3624 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4093
timestamp 1569543463
transform 1 0 3496 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4094
timestamp 1569543463
transform 1 0 3624 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4095
timestamp 1569543463
transform 1 0 3496 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4096
timestamp 1569543463
transform 1 0 3304 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4097
timestamp 1569543463
transform 1 0 3240 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4098
timestamp 1569543463
transform 1 0 3176 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4099
timestamp 1569543463
transform 1 0 3304 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4100
timestamp 1569543463
transform 1 0 3176 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4101
timestamp 1569543463
transform 1 0 3240 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4102
timestamp 1569543463
transform 1 0 3176 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4103
timestamp 1569543463
transform 1 0 3176 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4104
timestamp 1569543463
transform 1 0 3176 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4105
timestamp 1569543463
transform 1 0 3240 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4106
timestamp 1569543463
transform 1 0 3368 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4107
timestamp 1569543463
transform 1 0 3368 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4108
timestamp 1569543463
transform 1 0 3368 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4109
timestamp 1569543463
transform 1 0 3304 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4110
timestamp 1569543463
transform 1 0 3240 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4111
timestamp 1569543463
transform 1 0 3304 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4112
timestamp 1569543463
transform 1 0 3240 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4113
timestamp 1569543463
transform 1 0 3368 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4114
timestamp 1569543463
transform 1 0 3368 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4115
timestamp 1569543463
transform 1 0 3304 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4116
timestamp 1569543463
transform 1 0 3368 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4117
timestamp 1569543463
transform 1 0 3240 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4118
timestamp 1569543463
transform 1 0 3240 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4119
timestamp 1569543463
transform 1 0 3368 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4120
timestamp 1569543463
transform 1 0 3240 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4121
timestamp 1569543463
transform 1 0 3176 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4122
timestamp 1569543463
transform 1 0 3304 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4123
timestamp 1569543463
transform 1 0 3304 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4124
timestamp 1569543463
transform 1 0 3176 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4125
timestamp 1569543463
transform 1 0 3304 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4126
timestamp 1569543463
transform 1 0 3176 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4127
timestamp 1569543463
transform 1 0 3176 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4128
timestamp 1569543463
transform 1 0 3240 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4129
timestamp 1569543463
transform 1 0 3304 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4130
timestamp 1569543463
transform 1 0 3368 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4131
timestamp 1569543463
transform 1 0 3368 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4132
timestamp 1569543463
transform 1 0 3624 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4133
timestamp 1569543463
transform 1 0 3624 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4134
timestamp 1569543463
transform 1 0 3496 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4135
timestamp 1569543463
transform 1 0 3560 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4136
timestamp 1569543463
transform 1 0 3624 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4137
timestamp 1569543463
transform 1 0 3624 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4138
timestamp 1569543463
transform 1 0 3496 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4139
timestamp 1569543463
transform 1 0 3496 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4140
timestamp 1569543463
transform 1 0 3496 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4141
timestamp 1569543463
transform 1 0 3560 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4142
timestamp 1569543463
transform 1 0 3560 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4143
timestamp 1569543463
transform 1 0 3560 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4144
timestamp 1569543463
transform 1 0 3688 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4145
timestamp 1569543463
transform 1 0 3688 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4146
timestamp 1569543463
transform 1 0 3688 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4147
timestamp 1569543463
transform 1 0 3688 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4148
timestamp 1569543463
transform 1 0 3432 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4149
timestamp 1569543463
transform 1 0 3432 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4150
timestamp 1569543463
transform 1 0 3432 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4151
timestamp 1569543463
transform 1 0 3432 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4152
timestamp 1569543463
transform 1 0 3432 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4153
timestamp 1569543463
transform 1 0 3432 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4154
timestamp 1569543463
transform 1 0 3432 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4155
timestamp 1569543463
transform 1 0 3432 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4156
timestamp 1569543463
transform 1 0 3432 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4157
timestamp 1569543463
transform 1 0 4712 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4158
timestamp 1569543463
transform 1 0 4520 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4159
timestamp 1569543463
transform 1 0 4520 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4160
timestamp 1569543463
transform 1 0 4712 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4161
timestamp 1569543463
transform 1 0 4904 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4162
timestamp 1569543463
transform 1 0 4584 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4163
timestamp 1569543463
transform 1 0 4840 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4164
timestamp 1569543463
transform 1 0 4840 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4165
timestamp 1569543463
transform 1 0 4648 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4166
timestamp 1569543463
transform 1 0 4456 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4167
timestamp 1569543463
transform 1 0 4456 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4168
timestamp 1569543463
transform 1 0 4648 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4169
timestamp 1569543463
transform 1 0 4584 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4170
timestamp 1569543463
transform 1 0 4584 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4171
timestamp 1569543463
transform 1 0 4904 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4172
timestamp 1569543463
transform 1 0 4776 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4173
timestamp 1569543463
transform 1 0 4904 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4174
timestamp 1569543463
transform 1 0 4648 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4175
timestamp 1569543463
transform 1 0 4712 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4176
timestamp 1569543463
transform 1 0 4520 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4177
timestamp 1569543463
transform 1 0 4392 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4178
timestamp 1569543463
transform 1 0 4840 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4179
timestamp 1569543463
transform 1 0 4776 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4180
timestamp 1569543463
transform 1 0 4776 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4181
timestamp 1569543463
transform 1 0 4328 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4182
timestamp 1569543463
transform 1 0 3752 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4183
timestamp 1569543463
transform 1 0 3752 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4184
timestamp 1569543463
transform 1 0 3752 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4185
timestamp 1569543463
transform 1 0 3752 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_4186
timestamp 1569543463
transform 1 0 3752 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_4187
timestamp 1569543463
transform 1 0 3752 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_4188
timestamp 1569543463
transform 1 0 3752 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_4189
timestamp 1569543463
transform 1 0 3752 0 1 4200
box -8 -8 8 8
use VIA2$5  VIA2$5_4190
timestamp 1569543463
transform 1 0 3816 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4191
timestamp 1569543463
transform 1 0 3816 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4192
timestamp 1569543463
transform 1 0 3816 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4193
timestamp 1569543463
transform 1 0 3816 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_4194
timestamp 1569543463
transform 1 0 3816 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_4195
timestamp 1569543463
transform 1 0 3816 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_4196
timestamp 1569543463
transform 1 0 3816 0 1 4136
box -8 -8 8 8
use VIA2$5  VIA2$5_4197
timestamp 1569543463
transform 1 0 3880 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4198
timestamp 1569543463
transform 1 0 3880 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4199
timestamp 1569543463
transform 1 0 3880 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4200
timestamp 1569543463
transform 1 0 3880 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_4201
timestamp 1569543463
transform 1 0 3880 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_4202
timestamp 1569543463
transform 1 0 3880 0 1 4072
box -8 -8 8 8
use VIA2$5  VIA2$5_4203
timestamp 1569543463
transform 1 0 3944 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4204
timestamp 1569543463
transform 1 0 3944 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4205
timestamp 1569543463
transform 1 0 3944 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4206
timestamp 1569543463
transform 1 0 3944 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_4207
timestamp 1569543463
transform 1 0 3944 0 1 4008
box -8 -8 8 8
use VIA2$5  VIA2$5_4208
timestamp 1569543463
transform 1 0 4008 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4209
timestamp 1569543463
transform 1 0 4008 0 1 3944
box -8 -8 8 8
use VIA2$5  VIA2$5_4210
timestamp 1569543463
transform 1 0 4072 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4211
timestamp 1569543463
transform 1 0 4072 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4212
timestamp 1569543463
transform 1 0 4072 0 1 3880
box -8 -8 8 8
use VIA2$5  VIA2$5_4213
timestamp 1569543463
transform 1 0 4136 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4214
timestamp 1569543463
transform 1 0 4136 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4215
timestamp 1569543463
transform 1 0 3752 0 1 4264
box -8 -8 8 8
use VIA2$5  VIA2$5_4216
timestamp 1569543463
transform 1 0 3752 0 1 4328
box -8 -8 8 8
use VIA2$5  VIA2$5_4217
timestamp 1569543463
transform 1 0 4200 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4218
timestamp 1569543463
transform 1 0 4264 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4219
timestamp 1569543463
transform 1 0 4008 0 1 3752
box -8 -8 8 8
use VIA2$5  VIA2$5_4220
timestamp 1569543463
transform 1 0 4008 0 1 3816
box -8 -8 8 8
use VIA2$5  VIA2$5_4221
timestamp 1569543463
transform 1 0 4264 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4222
timestamp 1569543463
transform 1 0 4328 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4223
timestamp 1569543463
transform 1 0 4264 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4224
timestamp 1569543463
transform 1 0 3752 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4225
timestamp 1569543463
transform 1 0 3752 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4226
timestamp 1569543463
transform 1 0 3752 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4227
timestamp 1569543463
transform 1 0 3752 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4228
timestamp 1569543463
transform 1 0 3752 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4229
timestamp 1569543463
transform 1 0 4264 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4230
timestamp 1569543463
transform 1 0 3752 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4231
timestamp 1569543463
transform 1 0 4328 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4232
timestamp 1569543463
transform 1 0 4328 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4233
timestamp 1569543463
transform 1 0 4328 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4234
timestamp 1569543463
transform 1 0 4328 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4235
timestamp 1569543463
transform 1 0 4328 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4236
timestamp 1569543463
transform 1 0 4328 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4237
timestamp 1569543463
transform 1 0 4328 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4238
timestamp 1569543463
transform 1 0 3752 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4239
timestamp 1569543463
transform 1 0 4264 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4240
timestamp 1569543463
transform 1 0 4264 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4241
timestamp 1569543463
transform 1 0 3752 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4242
timestamp 1569543463
transform 1 0 4264 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4243
timestamp 1569543463
transform 1 0 3752 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4244
timestamp 1569543463
transform 1 0 4264 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4245
timestamp 1569543463
transform 1 0 4456 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4246
timestamp 1569543463
transform 1 0 4520 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4247
timestamp 1569543463
transform 1 0 4520 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4248
timestamp 1569543463
transform 1 0 4520 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4249
timestamp 1569543463
transform 1 0 4520 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4250
timestamp 1569543463
transform 1 0 4584 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4251
timestamp 1569543463
transform 1 0 4584 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4252
timestamp 1569543463
transform 1 0 4584 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4253
timestamp 1569543463
transform 1 0 4392 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4254
timestamp 1569543463
transform 1 0 4456 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4255
timestamp 1569543463
transform 1 0 4648 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4256
timestamp 1569543463
transform 1 0 4776 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4257
timestamp 1569543463
transform 1 0 4776 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4258
timestamp 1569543463
transform 1 0 4648 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4259
timestamp 1569543463
transform 1 0 4776 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4260
timestamp 1569543463
transform 1 0 4776 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4261
timestamp 1569543463
transform 1 0 4776 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4262
timestamp 1569543463
transform 1 0 4840 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4263
timestamp 1569543463
transform 1 0 4840 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4264
timestamp 1569543463
transform 1 0 4840 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4265
timestamp 1569543463
transform 1 0 4840 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4266
timestamp 1569543463
transform 1 0 4840 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4267
timestamp 1569543463
transform 1 0 4840 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4268
timestamp 1569543463
transform 1 0 4904 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4269
timestamp 1569543463
transform 1 0 4904 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4270
timestamp 1569543463
transform 1 0 4904 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4271
timestamp 1569543463
transform 1 0 4904 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4272
timestamp 1569543463
transform 1 0 4712 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4273
timestamp 1569543463
transform 1 0 4904 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4274
timestamp 1569543463
transform 1 0 4904 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4275
timestamp 1569543463
transform 1 0 4712 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4276
timestamp 1569543463
transform 1 0 4712 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4277
timestamp 1569543463
transform 1 0 4712 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4278
timestamp 1569543463
transform 1 0 4968 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4279
timestamp 1569543463
transform 1 0 4968 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4280
timestamp 1569543463
transform 1 0 4968 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4281
timestamp 1569543463
transform 1 0 4968 0 1 4904
box -8 -8 8 8
use VIA2$5  VIA2$5_4282
timestamp 1569543463
transform 1 0 4712 0 1 4968
box -8 -8 8 8
use VIA2$5  VIA2$5_4283
timestamp 1569543463
transform 1 0 4776 0 1 4968
box -8 -8 8 8
use VIA2$5  VIA2$5_4284
timestamp 1569543463
transform 1 0 4840 0 1 4968
box -8 -8 8 8
use VIA2$5  VIA2$5_4285
timestamp 1569543463
transform 1 0 4904 0 1 4968
box -8 -8 8 8
use VIA2$5  VIA2$5_4286
timestamp 1569543463
transform 1 0 4968 0 1 4968
box -8 -8 8 8
use VIA2$5  VIA2$5_4287
timestamp 1569543463
transform 1 0 4392 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4288
timestamp 1569543463
transform 1 0 4392 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4289
timestamp 1569543463
transform 1 0 4392 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4290
timestamp 1569543463
transform 1 0 4392 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4291
timestamp 1569543463
transform 1 0 4392 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4292
timestamp 1569543463
transform 1 0 4392 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4293
timestamp 1569543463
transform 1 0 4392 0 1 4776
box -8 -8 8 8
use VIA2$5  VIA2$5_4294
timestamp 1569543463
transform 1 0 4392 0 1 4840
box -8 -8 8 8
use VIA2$5  VIA2$5_4295
timestamp 1569543463
transform 1 0 4456 0 1 4392
box -8 -8 8 8
use VIA2$5  VIA2$5_4296
timestamp 1569543463
transform 1 0 4456 0 1 4456
box -8 -8 8 8
use VIA2$5  VIA2$5_4297
timestamp 1569543463
transform 1 0 4456 0 1 4520
box -8 -8 8 8
use VIA2$5  VIA2$5_4298
timestamp 1569543463
transform 1 0 4456 0 1 4584
box -8 -8 8 8
use VIA2$5  VIA2$5_4299
timestamp 1569543463
transform 1 0 4456 0 1 4648
box -8 -8 8 8
use VIA2$5  VIA2$5_4300
timestamp 1569543463
transform 1 0 4456 0 1 4712
box -8 -8 8 8
use VIA2$5  VIA2$5_4301
timestamp 1569543463
transform 1 0 4456 0 1 4776
box -8 -8 8 8
<< end >>
