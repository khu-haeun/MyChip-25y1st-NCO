magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect 8680 8700 29300 29300
<< metal1 >>
rect 11740 28979 28180 28980
rect 10061 28966 28180 28979
rect 10061 28950 10076 28966
rect 10092 28950 10108 28966
rect 10124 28950 10140 28966
rect 10156 28950 10172 28966
rect 10188 28950 10204 28966
rect 10220 28950 10236 28966
rect 10252 28950 10268 28966
rect 10284 28950 10300 28966
rect 10316 28950 10332 28966
rect 10348 28950 10364 28966
rect 10380 28950 10396 28966
rect 10412 28950 10428 28966
rect 10444 28950 10460 28966
rect 10476 28950 10492 28966
rect 10508 28950 10524 28966
rect 10540 28950 10556 28966
rect 10572 28950 10588 28966
rect 10604 28950 10620 28966
rect 10636 28950 10652 28966
rect 10668 28950 10684 28966
rect 10700 28950 10716 28966
rect 10732 28950 10748 28966
rect 10764 28950 10780 28966
rect 10796 28950 10812 28966
rect 10828 28950 10844 28966
rect 10860 28950 10876 28966
rect 10892 28950 10908 28966
rect 10924 28950 10940 28966
rect 10956 28950 10972 28966
rect 10988 28950 11004 28966
rect 11020 28950 11036 28966
rect 11052 28950 11068 28966
rect 11084 28950 11100 28966
rect 11116 28950 11132 28966
rect 11148 28950 11164 28966
rect 11180 28950 11196 28966
rect 11212 28950 11228 28966
rect 11244 28950 11260 28966
rect 11276 28950 11292 28966
rect 11308 28950 11324 28966
rect 11340 28950 11356 28966
rect 11372 28950 11388 28966
rect 11404 28950 11420 28966
rect 11436 28950 11452 28966
rect 11468 28950 11484 28966
rect 11500 28950 11516 28966
rect 11532 28950 11548 28966
rect 11564 28950 11580 28966
rect 11596 28950 11612 28966
rect 11628 28950 11644 28966
rect 11660 28950 11676 28966
rect 11692 28950 11708 28966
rect 11724 28950 28180 28966
rect 10061 28934 28180 28950
rect 10061 28918 10076 28934
rect 10092 28918 10108 28934
rect 10124 28918 10140 28934
rect 10156 28918 10172 28934
rect 10188 28918 10204 28934
rect 10220 28918 10236 28934
rect 10252 28918 10268 28934
rect 10284 28918 10300 28934
rect 10316 28918 10332 28934
rect 10348 28918 10364 28934
rect 10380 28918 10396 28934
rect 10412 28918 10428 28934
rect 10444 28918 10460 28934
rect 10476 28918 10492 28934
rect 10508 28918 10524 28934
rect 10540 28918 10556 28934
rect 10572 28918 10588 28934
rect 10604 28918 10620 28934
rect 10636 28918 10652 28934
rect 10668 28918 10684 28934
rect 10700 28918 10716 28934
rect 10732 28918 10748 28934
rect 10764 28918 10780 28934
rect 10796 28918 10812 28934
rect 10828 28918 10844 28934
rect 10860 28918 10876 28934
rect 10892 28918 10908 28934
rect 10924 28918 10940 28934
rect 10956 28918 10972 28934
rect 10988 28918 11004 28934
rect 11020 28918 11036 28934
rect 11052 28918 11068 28934
rect 11084 28918 11100 28934
rect 11116 28918 11132 28934
rect 11148 28918 11164 28934
rect 11180 28918 11196 28934
rect 11212 28918 11228 28934
rect 11244 28918 11260 28934
rect 11276 28918 11292 28934
rect 11308 28918 11324 28934
rect 11340 28918 11356 28934
rect 11372 28918 11388 28934
rect 11404 28918 11420 28934
rect 11436 28918 11452 28934
rect 11468 28918 11484 28934
rect 11500 28918 11516 28934
rect 11532 28918 11548 28934
rect 11564 28918 11580 28934
rect 11596 28918 11612 28934
rect 11628 28918 11644 28934
rect 11660 28918 11676 28934
rect 11692 28918 11708 28934
rect 11724 28918 28180 28934
rect 10061 28902 28180 28918
rect 10061 28886 10076 28902
rect 10092 28886 10108 28902
rect 10124 28886 10140 28902
rect 10156 28886 10172 28902
rect 10188 28886 10204 28902
rect 10220 28886 10236 28902
rect 10252 28886 10268 28902
rect 10284 28886 10300 28902
rect 10316 28886 10332 28902
rect 10348 28886 10364 28902
rect 10380 28886 10396 28902
rect 10412 28886 10428 28902
rect 10444 28886 10460 28902
rect 10476 28886 10492 28902
rect 10508 28886 10524 28902
rect 10540 28886 10556 28902
rect 10572 28886 10588 28902
rect 10604 28886 10620 28902
rect 10636 28886 10652 28902
rect 10668 28886 10684 28902
rect 10700 28886 10716 28902
rect 10732 28886 10748 28902
rect 10764 28886 10780 28902
rect 10796 28886 10812 28902
rect 10828 28886 10844 28902
rect 10860 28886 10876 28902
rect 10892 28886 10908 28902
rect 10924 28886 10940 28902
rect 10956 28886 10972 28902
rect 10988 28886 11004 28902
rect 11020 28886 11036 28902
rect 11052 28886 11068 28902
rect 11084 28886 11100 28902
rect 11116 28886 11132 28902
rect 11148 28886 11164 28902
rect 11180 28886 11196 28902
rect 11212 28886 11228 28902
rect 11244 28886 11260 28902
rect 11276 28886 11292 28902
rect 11308 28886 11324 28902
rect 11340 28886 11356 28902
rect 11372 28886 11388 28902
rect 11404 28886 11420 28902
rect 11436 28886 11452 28902
rect 11468 28886 11484 28902
rect 11500 28886 11516 28902
rect 11532 28886 11548 28902
rect 11564 28886 11580 28902
rect 11596 28886 11612 28902
rect 11628 28886 11644 28902
rect 11660 28886 11676 28902
rect 11692 28886 11708 28902
rect 11724 28886 28180 28902
rect 10061 28870 28180 28886
rect 10061 28854 10076 28870
rect 10092 28854 10108 28870
rect 10124 28854 10140 28870
rect 10156 28854 10172 28870
rect 10188 28854 10204 28870
rect 10220 28854 10236 28870
rect 10252 28854 10268 28870
rect 10284 28854 10300 28870
rect 10316 28854 10332 28870
rect 10348 28854 10364 28870
rect 10380 28854 10396 28870
rect 10412 28854 10428 28870
rect 10444 28854 10460 28870
rect 10476 28854 10492 28870
rect 10508 28854 10524 28870
rect 10540 28854 10556 28870
rect 10572 28854 10588 28870
rect 10604 28854 10620 28870
rect 10636 28854 10652 28870
rect 10668 28854 10684 28870
rect 10700 28854 10716 28870
rect 10732 28854 10748 28870
rect 10764 28854 10780 28870
rect 10796 28854 10812 28870
rect 10828 28854 10844 28870
rect 10860 28854 10876 28870
rect 10892 28854 10908 28870
rect 10924 28854 10940 28870
rect 10956 28854 10972 28870
rect 10988 28854 11004 28870
rect 11020 28854 11036 28870
rect 11052 28854 11068 28870
rect 11084 28854 11100 28870
rect 11116 28854 11132 28870
rect 11148 28854 11164 28870
rect 11180 28854 11196 28870
rect 11212 28854 11228 28870
rect 11244 28854 11260 28870
rect 11276 28854 11292 28870
rect 11308 28854 11324 28870
rect 11340 28854 11356 28870
rect 11372 28854 11388 28870
rect 11404 28854 11420 28870
rect 11436 28854 11452 28870
rect 11468 28854 11484 28870
rect 11500 28854 11516 28870
rect 11532 28854 11548 28870
rect 11564 28854 11580 28870
rect 11596 28854 11612 28870
rect 11628 28854 11644 28870
rect 11660 28854 11676 28870
rect 11692 28854 11708 28870
rect 11724 28854 28180 28870
rect 10061 28838 28180 28854
rect 10061 28822 10076 28838
rect 10092 28822 10108 28838
rect 10124 28822 10140 28838
rect 10156 28822 10172 28838
rect 10188 28822 10204 28838
rect 10220 28822 10236 28838
rect 10252 28822 10268 28838
rect 10284 28822 10300 28838
rect 10316 28822 10332 28838
rect 10348 28822 10364 28838
rect 10380 28822 10396 28838
rect 10412 28822 10428 28838
rect 10444 28822 10460 28838
rect 10476 28822 10492 28838
rect 10508 28822 10524 28838
rect 10540 28822 10556 28838
rect 10572 28822 10588 28838
rect 10604 28822 10620 28838
rect 10636 28822 10652 28838
rect 10668 28822 10684 28838
rect 10700 28822 10716 28838
rect 10732 28822 10748 28838
rect 10764 28822 10780 28838
rect 10796 28822 10812 28838
rect 10828 28822 10844 28838
rect 10860 28822 10876 28838
rect 10892 28822 10908 28838
rect 10924 28822 10940 28838
rect 10956 28822 10972 28838
rect 10988 28822 11004 28838
rect 11020 28822 11036 28838
rect 11052 28822 11068 28838
rect 11084 28822 11100 28838
rect 11116 28822 11132 28838
rect 11148 28822 11164 28838
rect 11180 28822 11196 28838
rect 11212 28822 11228 28838
rect 11244 28822 11260 28838
rect 11276 28822 11292 28838
rect 11308 28822 11324 28838
rect 11340 28822 11356 28838
rect 11372 28822 11388 28838
rect 11404 28822 11420 28838
rect 11436 28822 11452 28838
rect 11468 28822 11484 28838
rect 11500 28822 11516 28838
rect 11532 28822 11548 28838
rect 11564 28822 11580 28838
rect 11596 28822 11612 28838
rect 11628 28822 11644 28838
rect 11660 28822 11676 28838
rect 11692 28822 11708 28838
rect 11724 28822 28180 28838
rect 10061 28806 28180 28822
rect 10061 28790 10076 28806
rect 10092 28790 10108 28806
rect 10124 28790 10140 28806
rect 10156 28790 10172 28806
rect 10188 28790 10204 28806
rect 10220 28790 10236 28806
rect 10252 28790 10268 28806
rect 10284 28790 10300 28806
rect 10316 28790 10332 28806
rect 10348 28790 10364 28806
rect 10380 28790 10396 28806
rect 10412 28790 10428 28806
rect 10444 28790 10460 28806
rect 10476 28790 10492 28806
rect 10508 28790 10524 28806
rect 10540 28790 10556 28806
rect 10572 28790 10588 28806
rect 10604 28790 10620 28806
rect 10636 28790 10652 28806
rect 10668 28790 10684 28806
rect 10700 28790 10716 28806
rect 10732 28790 10748 28806
rect 10764 28790 10780 28806
rect 10796 28790 10812 28806
rect 10828 28790 10844 28806
rect 10860 28790 10876 28806
rect 10892 28790 10908 28806
rect 10924 28790 10940 28806
rect 10956 28790 10972 28806
rect 10988 28790 11004 28806
rect 11020 28790 11036 28806
rect 11052 28790 11068 28806
rect 11084 28790 11100 28806
rect 11116 28790 11132 28806
rect 11148 28790 11164 28806
rect 11180 28790 11196 28806
rect 11212 28790 11228 28806
rect 11244 28790 11260 28806
rect 11276 28790 11292 28806
rect 11308 28790 11324 28806
rect 11340 28790 11356 28806
rect 11372 28790 11388 28806
rect 11404 28790 11420 28806
rect 11436 28790 11452 28806
rect 11468 28790 11484 28806
rect 11500 28790 11516 28806
rect 11532 28790 11548 28806
rect 11564 28790 11580 28806
rect 11596 28790 11612 28806
rect 11628 28790 11644 28806
rect 11660 28790 11676 28806
rect 11692 28790 11708 28806
rect 11724 28790 28180 28806
rect 10061 28774 28180 28790
rect 10061 28758 10076 28774
rect 10092 28758 10108 28774
rect 10124 28758 10140 28774
rect 10156 28758 10172 28774
rect 10188 28758 10204 28774
rect 10220 28758 10236 28774
rect 10252 28758 10268 28774
rect 10284 28758 10300 28774
rect 10316 28758 10332 28774
rect 10348 28758 10364 28774
rect 10380 28758 10396 28774
rect 10412 28758 10428 28774
rect 10444 28758 10460 28774
rect 10476 28758 10492 28774
rect 10508 28758 10524 28774
rect 10540 28758 10556 28774
rect 10572 28758 10588 28774
rect 10604 28758 10620 28774
rect 10636 28758 10652 28774
rect 10668 28758 10684 28774
rect 10700 28758 10716 28774
rect 10732 28758 10748 28774
rect 10764 28758 10780 28774
rect 10796 28758 10812 28774
rect 10828 28758 10844 28774
rect 10860 28758 10876 28774
rect 10892 28758 10908 28774
rect 10924 28758 10940 28774
rect 10956 28758 10972 28774
rect 10988 28758 11004 28774
rect 11020 28758 11036 28774
rect 11052 28758 11068 28774
rect 11084 28758 11100 28774
rect 11116 28758 11132 28774
rect 11148 28758 11164 28774
rect 11180 28758 11196 28774
rect 11212 28758 11228 28774
rect 11244 28758 11260 28774
rect 11276 28758 11292 28774
rect 11308 28758 11324 28774
rect 11340 28758 11356 28774
rect 11372 28758 11388 28774
rect 11404 28758 11420 28774
rect 11436 28758 11452 28774
rect 11468 28758 11484 28774
rect 11500 28758 11516 28774
rect 11532 28758 11548 28774
rect 11564 28758 11580 28774
rect 11596 28758 11612 28774
rect 11628 28758 11644 28774
rect 11660 28758 11676 28774
rect 11692 28758 11708 28774
rect 11724 28758 28180 28774
rect 10061 28742 28180 28758
rect 10061 28726 10076 28742
rect 10092 28726 10108 28742
rect 10124 28726 10140 28742
rect 10156 28726 10172 28742
rect 10188 28726 10204 28742
rect 10220 28726 10236 28742
rect 10252 28726 10268 28742
rect 10284 28726 10300 28742
rect 10316 28726 10332 28742
rect 10348 28726 10364 28742
rect 10380 28726 10396 28742
rect 10412 28726 10428 28742
rect 10444 28726 10460 28742
rect 10476 28726 10492 28742
rect 10508 28726 10524 28742
rect 10540 28726 10556 28742
rect 10572 28726 10588 28742
rect 10604 28726 10620 28742
rect 10636 28726 10652 28742
rect 10668 28726 10684 28742
rect 10700 28726 10716 28742
rect 10732 28726 10748 28742
rect 10764 28726 10780 28742
rect 10796 28726 10812 28742
rect 10828 28726 10844 28742
rect 10860 28726 10876 28742
rect 10892 28726 10908 28742
rect 10924 28726 10940 28742
rect 10956 28726 10972 28742
rect 10988 28726 11004 28742
rect 11020 28726 11036 28742
rect 11052 28726 11068 28742
rect 11084 28726 11100 28742
rect 11116 28726 11132 28742
rect 11148 28726 11164 28742
rect 11180 28726 11196 28742
rect 11212 28726 11228 28742
rect 11244 28726 11260 28742
rect 11276 28726 11292 28742
rect 11308 28726 11324 28742
rect 11340 28726 11356 28742
rect 11372 28726 11388 28742
rect 11404 28726 11420 28742
rect 11436 28726 11452 28742
rect 11468 28726 11484 28742
rect 11500 28726 11516 28742
rect 11532 28726 11548 28742
rect 11564 28726 11580 28742
rect 11596 28726 11612 28742
rect 11628 28726 11644 28742
rect 11660 28726 11676 28742
rect 11692 28726 11708 28742
rect 11724 28726 28180 28742
rect 10061 28710 28180 28726
rect 10061 28694 10076 28710
rect 10092 28694 10108 28710
rect 10124 28694 10140 28710
rect 10156 28694 10172 28710
rect 10188 28694 10204 28710
rect 10220 28694 10236 28710
rect 10252 28694 10268 28710
rect 10284 28694 10300 28710
rect 10316 28694 10332 28710
rect 10348 28694 10364 28710
rect 10380 28694 10396 28710
rect 10412 28694 10428 28710
rect 10444 28694 10460 28710
rect 10476 28694 10492 28710
rect 10508 28694 10524 28710
rect 10540 28694 10556 28710
rect 10572 28694 10588 28710
rect 10604 28694 10620 28710
rect 10636 28694 10652 28710
rect 10668 28694 10684 28710
rect 10700 28694 10716 28710
rect 10732 28694 10748 28710
rect 10764 28694 10780 28710
rect 10796 28694 10812 28710
rect 10828 28694 10844 28710
rect 10860 28694 10876 28710
rect 10892 28694 10908 28710
rect 10924 28694 10940 28710
rect 10956 28694 10972 28710
rect 10988 28694 11004 28710
rect 11020 28694 11036 28710
rect 11052 28694 11068 28710
rect 11084 28694 11100 28710
rect 11116 28694 11132 28710
rect 11148 28694 11164 28710
rect 11180 28694 11196 28710
rect 11212 28694 11228 28710
rect 11244 28694 11260 28710
rect 11276 28694 11292 28710
rect 11308 28694 11324 28710
rect 11340 28694 11356 28710
rect 11372 28694 11388 28710
rect 11404 28694 11420 28710
rect 11436 28694 11452 28710
rect 11468 28694 11484 28710
rect 11500 28694 11516 28710
rect 11532 28694 11548 28710
rect 11564 28694 11580 28710
rect 11596 28694 11612 28710
rect 11628 28694 11644 28710
rect 11660 28694 11676 28710
rect 11692 28694 11708 28710
rect 11724 28694 28180 28710
rect 10061 28681 28180 28694
rect 11740 28680 28180 28681
rect 27960 27820 28180 28680
rect 9660 27679 10100 27680
rect 9081 27668 10100 27679
rect 9081 27652 9106 27668
rect 9122 27652 9138 27668
rect 9154 27652 9170 27668
rect 9186 27652 9202 27668
rect 9218 27652 9234 27668
rect 9250 27652 9266 27668
rect 9282 27652 9298 27668
rect 9314 27652 9330 27668
rect 9346 27652 9362 27668
rect 9378 27652 9394 27668
rect 9410 27652 9426 27668
rect 9442 27652 9458 27668
rect 9474 27652 9490 27668
rect 9506 27652 9522 27668
rect 9538 27652 9554 27668
rect 9570 27652 9586 27668
rect 9602 27652 9618 27668
rect 9634 27652 10100 27668
rect 9081 27636 10100 27652
rect 9081 27620 9106 27636
rect 9122 27620 9138 27636
rect 9154 27620 9170 27636
rect 9186 27620 9202 27636
rect 9218 27620 9234 27636
rect 9250 27620 9266 27636
rect 9282 27620 9298 27636
rect 9314 27620 9330 27636
rect 9346 27620 9362 27636
rect 9378 27620 9394 27636
rect 9410 27620 9426 27636
rect 9442 27620 9458 27636
rect 9474 27620 9490 27636
rect 9506 27620 9522 27636
rect 9538 27620 9554 27636
rect 9570 27620 9586 27636
rect 9602 27620 9618 27636
rect 9634 27620 10100 27636
rect 9081 27604 10100 27620
rect 9081 27588 9106 27604
rect 9122 27588 9138 27604
rect 9154 27588 9170 27604
rect 9186 27588 9202 27604
rect 9218 27588 9234 27604
rect 9250 27588 9266 27604
rect 9282 27588 9298 27604
rect 9314 27588 9330 27604
rect 9346 27588 9362 27604
rect 9378 27588 9394 27604
rect 9410 27588 9426 27604
rect 9442 27588 9458 27604
rect 9474 27588 9490 27604
rect 9506 27588 9522 27604
rect 9538 27588 9554 27604
rect 9570 27588 9586 27604
rect 9602 27588 9618 27604
rect 9634 27588 10100 27604
rect 9081 27572 10100 27588
rect 9081 27556 9106 27572
rect 9122 27556 9138 27572
rect 9154 27556 9170 27572
rect 9186 27556 9202 27572
rect 9218 27556 9234 27572
rect 9250 27556 9266 27572
rect 9282 27556 9298 27572
rect 9314 27556 9330 27572
rect 9346 27556 9362 27572
rect 9378 27556 9394 27572
rect 9410 27556 9426 27572
rect 9442 27556 9458 27572
rect 9474 27556 9490 27572
rect 9506 27556 9522 27572
rect 9538 27556 9554 27572
rect 9570 27556 9586 27572
rect 9602 27556 9618 27572
rect 9634 27556 10100 27572
rect 9081 27540 10100 27556
rect 9081 27524 9106 27540
rect 9122 27524 9138 27540
rect 9154 27524 9170 27540
rect 9186 27524 9202 27540
rect 9218 27524 9234 27540
rect 9250 27524 9266 27540
rect 9282 27524 9298 27540
rect 9314 27524 9330 27540
rect 9346 27524 9362 27540
rect 9378 27524 9394 27540
rect 9410 27524 9426 27540
rect 9442 27524 9458 27540
rect 9474 27524 9490 27540
rect 9506 27524 9522 27540
rect 9538 27524 9554 27540
rect 9570 27524 9586 27540
rect 9602 27524 9618 27540
rect 9634 27524 10100 27540
rect 9081 27508 10100 27524
rect 9081 27492 9106 27508
rect 9122 27492 9138 27508
rect 9154 27492 9170 27508
rect 9186 27492 9202 27508
rect 9218 27492 9234 27508
rect 9250 27492 9266 27508
rect 9282 27492 9298 27508
rect 9314 27492 9330 27508
rect 9346 27492 9362 27508
rect 9378 27492 9394 27508
rect 9410 27492 9426 27508
rect 9442 27492 9458 27508
rect 9474 27492 9490 27508
rect 9506 27492 9522 27508
rect 9538 27492 9554 27508
rect 9570 27492 9586 27508
rect 9602 27492 9618 27508
rect 9634 27492 10100 27508
rect 9081 27476 10100 27492
rect 9081 27460 9106 27476
rect 9122 27460 9138 27476
rect 9154 27460 9170 27476
rect 9186 27460 9202 27476
rect 9218 27460 9234 27476
rect 9250 27460 9266 27476
rect 9282 27460 9298 27476
rect 9314 27460 9330 27476
rect 9346 27460 9362 27476
rect 9378 27460 9394 27476
rect 9410 27460 9426 27476
rect 9442 27460 9458 27476
rect 9474 27460 9490 27476
rect 9506 27460 9522 27476
rect 9538 27460 9554 27476
rect 9570 27460 9586 27476
rect 9602 27460 9618 27476
rect 9634 27460 10100 27476
rect 9081 27444 10100 27460
rect 9081 27428 9106 27444
rect 9122 27428 9138 27444
rect 9154 27428 9170 27444
rect 9186 27428 9202 27444
rect 9218 27428 9234 27444
rect 9250 27428 9266 27444
rect 9282 27428 9298 27444
rect 9314 27428 9330 27444
rect 9346 27428 9362 27444
rect 9378 27428 9394 27444
rect 9410 27428 9426 27444
rect 9442 27428 9458 27444
rect 9474 27428 9490 27444
rect 9506 27428 9522 27444
rect 9538 27428 9554 27444
rect 9570 27428 9586 27444
rect 9602 27428 9618 27444
rect 9634 27428 10100 27444
rect 9081 27412 10100 27428
rect 9081 27396 9106 27412
rect 9122 27396 9138 27412
rect 9154 27396 9170 27412
rect 9186 27396 9202 27412
rect 9218 27396 9234 27412
rect 9250 27396 9266 27412
rect 9282 27396 9298 27412
rect 9314 27396 9330 27412
rect 9346 27396 9362 27412
rect 9378 27396 9394 27412
rect 9410 27396 9426 27412
rect 9442 27396 9458 27412
rect 9474 27396 9490 27412
rect 9506 27396 9522 27412
rect 9538 27396 9554 27412
rect 9570 27396 9586 27412
rect 9602 27396 9618 27412
rect 9634 27396 10100 27412
rect 9081 27380 10100 27396
rect 9081 27364 9106 27380
rect 9122 27364 9138 27380
rect 9154 27364 9170 27380
rect 9186 27364 9202 27380
rect 9218 27364 9234 27380
rect 9250 27364 9266 27380
rect 9282 27364 9298 27380
rect 9314 27364 9330 27380
rect 9346 27364 9362 27380
rect 9378 27364 9394 27380
rect 9410 27364 9426 27380
rect 9442 27364 9458 27380
rect 9474 27364 9490 27380
rect 9506 27364 9522 27380
rect 9538 27364 9554 27380
rect 9570 27364 9586 27380
rect 9602 27364 9618 27380
rect 9634 27364 10100 27380
rect 9081 27348 10100 27364
rect 9081 27332 9106 27348
rect 9122 27332 9138 27348
rect 9154 27332 9170 27348
rect 9186 27332 9202 27348
rect 9218 27332 9234 27348
rect 9250 27332 9266 27348
rect 9282 27332 9298 27348
rect 9314 27332 9330 27348
rect 9346 27332 9362 27348
rect 9378 27332 9394 27348
rect 9410 27332 9426 27348
rect 9442 27332 9458 27348
rect 9474 27332 9490 27348
rect 9506 27332 9522 27348
rect 9538 27332 9554 27348
rect 9570 27332 9586 27348
rect 9602 27332 9618 27348
rect 9634 27332 10100 27348
rect 9081 27316 10100 27332
rect 9081 27300 9106 27316
rect 9122 27300 9138 27316
rect 9154 27300 9170 27316
rect 9186 27300 9202 27316
rect 9218 27300 9234 27316
rect 9250 27300 9266 27316
rect 9282 27300 9298 27316
rect 9314 27300 9330 27316
rect 9346 27300 9362 27316
rect 9378 27300 9394 27316
rect 9410 27300 9426 27316
rect 9442 27300 9458 27316
rect 9474 27300 9490 27316
rect 9506 27300 9522 27316
rect 9538 27300 9554 27316
rect 9570 27300 9586 27316
rect 9602 27300 9618 27316
rect 9634 27300 10100 27316
rect 9081 27284 10100 27300
rect 9081 27268 9106 27284
rect 9122 27268 9138 27284
rect 9154 27268 9170 27284
rect 9186 27268 9202 27284
rect 9218 27268 9234 27284
rect 9250 27268 9266 27284
rect 9282 27268 9298 27284
rect 9314 27268 9330 27284
rect 9346 27268 9362 27284
rect 9378 27268 9394 27284
rect 9410 27268 9426 27284
rect 9442 27268 9458 27284
rect 9474 27268 9490 27284
rect 9506 27268 9522 27284
rect 9538 27268 9554 27284
rect 9570 27268 9586 27284
rect 9602 27268 9618 27284
rect 9634 27268 10100 27284
rect 9081 27252 10100 27268
rect 9081 27236 9106 27252
rect 9122 27236 9138 27252
rect 9154 27236 9170 27252
rect 9186 27236 9202 27252
rect 9218 27236 9234 27252
rect 9250 27236 9266 27252
rect 9282 27236 9298 27252
rect 9314 27236 9330 27252
rect 9346 27236 9362 27252
rect 9378 27236 9394 27252
rect 9410 27236 9426 27252
rect 9442 27236 9458 27252
rect 9474 27236 9490 27252
rect 9506 27236 9522 27252
rect 9538 27236 9554 27252
rect 9570 27236 9586 27252
rect 9602 27236 9618 27252
rect 9634 27236 10100 27252
rect 9081 27220 10100 27236
rect 9081 27204 9106 27220
rect 9122 27204 9138 27220
rect 9154 27204 9170 27220
rect 9186 27204 9202 27220
rect 9218 27204 9234 27220
rect 9250 27204 9266 27220
rect 9282 27204 9298 27220
rect 9314 27204 9330 27220
rect 9346 27204 9362 27220
rect 9378 27204 9394 27220
rect 9410 27204 9426 27220
rect 9442 27204 9458 27220
rect 9474 27204 9490 27220
rect 9506 27204 9522 27220
rect 9538 27204 9554 27220
rect 9570 27204 9586 27220
rect 9602 27204 9618 27220
rect 9634 27204 10100 27220
rect 9081 27188 10100 27204
rect 9081 27172 9106 27188
rect 9122 27172 9138 27188
rect 9154 27172 9170 27188
rect 9186 27172 9202 27188
rect 9218 27172 9234 27188
rect 9250 27172 9266 27188
rect 9282 27172 9298 27188
rect 9314 27172 9330 27188
rect 9346 27172 9362 27188
rect 9378 27172 9394 27188
rect 9410 27172 9426 27188
rect 9442 27172 9458 27188
rect 9474 27172 9490 27188
rect 9506 27172 9522 27188
rect 9538 27172 9554 27188
rect 9570 27172 9586 27188
rect 9602 27172 9618 27188
rect 9634 27172 10100 27188
rect 9081 27156 10100 27172
rect 9081 27140 9106 27156
rect 9122 27140 9138 27156
rect 9154 27140 9170 27156
rect 9186 27140 9202 27156
rect 9218 27140 9234 27156
rect 9250 27140 9266 27156
rect 9282 27140 9298 27156
rect 9314 27140 9330 27156
rect 9346 27140 9362 27156
rect 9378 27140 9394 27156
rect 9410 27140 9426 27156
rect 9442 27140 9458 27156
rect 9474 27140 9490 27156
rect 9506 27140 9522 27156
rect 9538 27140 9554 27156
rect 9570 27140 9586 27156
rect 9602 27140 9618 27156
rect 9634 27140 10100 27156
rect 9081 27124 10100 27140
rect 9081 27108 9106 27124
rect 9122 27108 9138 27124
rect 9154 27108 9170 27124
rect 9186 27108 9202 27124
rect 9218 27108 9234 27124
rect 9250 27108 9266 27124
rect 9282 27108 9298 27124
rect 9314 27108 9330 27124
rect 9346 27108 9362 27124
rect 9378 27108 9394 27124
rect 9410 27108 9426 27124
rect 9442 27108 9458 27124
rect 9474 27108 9490 27124
rect 9506 27108 9522 27124
rect 9538 27108 9554 27124
rect 9570 27108 9586 27124
rect 9602 27108 9618 27124
rect 9634 27108 10100 27124
rect 9081 27092 10100 27108
rect 9081 27076 9106 27092
rect 9122 27076 9138 27092
rect 9154 27076 9170 27092
rect 9186 27076 9202 27092
rect 9218 27076 9234 27092
rect 9250 27076 9266 27092
rect 9282 27076 9298 27092
rect 9314 27076 9330 27092
rect 9346 27076 9362 27092
rect 9378 27076 9394 27092
rect 9410 27076 9426 27092
rect 9442 27076 9458 27092
rect 9474 27076 9490 27092
rect 9506 27076 9522 27092
rect 9538 27076 9554 27092
rect 9570 27076 9586 27092
rect 9602 27076 9618 27092
rect 9634 27076 10100 27092
rect 9081 27060 10100 27076
rect 9081 27044 9106 27060
rect 9122 27044 9138 27060
rect 9154 27044 9170 27060
rect 9186 27044 9202 27060
rect 9218 27044 9234 27060
rect 9250 27044 9266 27060
rect 9282 27044 9298 27060
rect 9314 27044 9330 27060
rect 9346 27044 9362 27060
rect 9378 27044 9394 27060
rect 9410 27044 9426 27060
rect 9442 27044 9458 27060
rect 9474 27044 9490 27060
rect 9506 27044 9522 27060
rect 9538 27044 9554 27060
rect 9570 27044 9586 27060
rect 9602 27044 9618 27060
rect 9634 27044 10100 27060
rect 9081 27028 10100 27044
rect 9081 27012 9106 27028
rect 9122 27012 9138 27028
rect 9154 27012 9170 27028
rect 9186 27012 9202 27028
rect 9218 27012 9234 27028
rect 9250 27012 9266 27028
rect 9282 27012 9298 27028
rect 9314 27012 9330 27028
rect 9346 27012 9362 27028
rect 9378 27012 9394 27028
rect 9410 27012 9426 27028
rect 9442 27012 9458 27028
rect 9474 27012 9490 27028
rect 9506 27012 9522 27028
rect 9538 27012 9554 27028
rect 9570 27012 9586 27028
rect 9602 27012 9618 27028
rect 9634 27012 10100 27028
rect 9081 26996 10100 27012
rect 9081 26980 9106 26996
rect 9122 26980 9138 26996
rect 9154 26980 9170 26996
rect 9186 26980 9202 26996
rect 9218 26980 9234 26996
rect 9250 26980 9266 26996
rect 9282 26980 9298 26996
rect 9314 26980 9330 26996
rect 9346 26980 9362 26996
rect 9378 26980 9394 26996
rect 9410 26980 9426 26996
rect 9442 26980 9458 26996
rect 9474 26980 9490 26996
rect 9506 26980 9522 26996
rect 9538 26980 9554 26996
rect 9570 26980 9586 26996
rect 9602 26980 9618 26996
rect 9634 26980 10100 26996
rect 9081 26964 10100 26980
rect 9081 26948 9106 26964
rect 9122 26948 9138 26964
rect 9154 26948 9170 26964
rect 9186 26948 9202 26964
rect 9218 26948 9234 26964
rect 9250 26948 9266 26964
rect 9282 26948 9298 26964
rect 9314 26948 9330 26964
rect 9346 26948 9362 26964
rect 9378 26948 9394 26964
rect 9410 26948 9426 26964
rect 9442 26948 9458 26964
rect 9474 26948 9490 26964
rect 9506 26948 9522 26964
rect 9538 26948 9554 26964
rect 9570 26948 9586 26964
rect 9602 26948 9618 26964
rect 9634 26948 10100 26964
rect 9081 26932 10100 26948
rect 9081 26916 9106 26932
rect 9122 26916 9138 26932
rect 9154 26916 9170 26932
rect 9186 26916 9202 26932
rect 9218 26916 9234 26932
rect 9250 26916 9266 26932
rect 9282 26916 9298 26932
rect 9314 26916 9330 26932
rect 9346 26916 9362 26932
rect 9378 26916 9394 26932
rect 9410 26916 9426 26932
rect 9442 26916 9458 26932
rect 9474 26916 9490 26932
rect 9506 26916 9522 26932
rect 9538 26916 9554 26932
rect 9570 26916 9586 26932
rect 9602 26916 9618 26932
rect 9634 26916 10100 26932
rect 9081 26900 10100 26916
rect 9081 26884 9106 26900
rect 9122 26884 9138 26900
rect 9154 26884 9170 26900
rect 9186 26884 9202 26900
rect 9218 26884 9234 26900
rect 9250 26884 9266 26900
rect 9282 26884 9298 26900
rect 9314 26884 9330 26900
rect 9346 26884 9362 26900
rect 9378 26884 9394 26900
rect 9410 26884 9426 26900
rect 9442 26884 9458 26900
rect 9474 26884 9490 26900
rect 9506 26884 9522 26900
rect 9538 26884 9554 26900
rect 9570 26884 9586 26900
rect 9602 26884 9618 26900
rect 9634 26884 10100 26900
rect 9081 26868 10100 26884
rect 9081 26852 9106 26868
rect 9122 26852 9138 26868
rect 9154 26852 9170 26868
rect 9186 26852 9202 26868
rect 9218 26852 9234 26868
rect 9250 26852 9266 26868
rect 9282 26852 9298 26868
rect 9314 26852 9330 26868
rect 9346 26852 9362 26868
rect 9378 26852 9394 26868
rect 9410 26852 9426 26868
rect 9442 26852 9458 26868
rect 9474 26852 9490 26868
rect 9506 26852 9522 26868
rect 9538 26852 9554 26868
rect 9570 26852 9586 26868
rect 9602 26852 9618 26868
rect 9634 26852 10100 26868
rect 9081 26836 10100 26852
rect 9081 26820 9106 26836
rect 9122 26820 9138 26836
rect 9154 26820 9170 26836
rect 9186 26820 9202 26836
rect 9218 26820 9234 26836
rect 9250 26820 9266 26836
rect 9282 26820 9298 26836
rect 9314 26820 9330 26836
rect 9346 26820 9362 26836
rect 9378 26820 9394 26836
rect 9410 26820 9426 26836
rect 9442 26820 9458 26836
rect 9474 26820 9490 26836
rect 9506 26820 9522 26836
rect 9538 26820 9554 26836
rect 9570 26820 9586 26836
rect 9602 26820 9618 26836
rect 9634 26820 10100 26836
rect 9081 26804 10100 26820
rect 9081 26788 9106 26804
rect 9122 26788 9138 26804
rect 9154 26788 9170 26804
rect 9186 26788 9202 26804
rect 9218 26788 9234 26804
rect 9250 26788 9266 26804
rect 9282 26788 9298 26804
rect 9314 26788 9330 26804
rect 9346 26788 9362 26804
rect 9378 26788 9394 26804
rect 9410 26788 9426 26804
rect 9442 26788 9458 26804
rect 9474 26788 9490 26804
rect 9506 26788 9522 26804
rect 9538 26788 9554 26804
rect 9570 26788 9586 26804
rect 9602 26788 9618 26804
rect 9634 26788 10100 26804
rect 9081 26772 10100 26788
rect 9081 26756 9106 26772
rect 9122 26756 9138 26772
rect 9154 26756 9170 26772
rect 9186 26756 9202 26772
rect 9218 26756 9234 26772
rect 9250 26756 9266 26772
rect 9282 26756 9298 26772
rect 9314 26756 9330 26772
rect 9346 26756 9362 26772
rect 9378 26756 9394 26772
rect 9410 26756 9426 26772
rect 9442 26756 9458 26772
rect 9474 26756 9490 26772
rect 9506 26756 9522 26772
rect 9538 26756 9554 26772
rect 9570 26756 9586 26772
rect 9602 26756 9618 26772
rect 9634 26756 10100 26772
rect 9081 26740 10100 26756
rect 9081 26724 9106 26740
rect 9122 26724 9138 26740
rect 9154 26724 9170 26740
rect 9186 26724 9202 26740
rect 9218 26724 9234 26740
rect 9250 26724 9266 26740
rect 9282 26724 9298 26740
rect 9314 26724 9330 26740
rect 9346 26724 9362 26740
rect 9378 26724 9394 26740
rect 9410 26724 9426 26740
rect 9442 26724 9458 26740
rect 9474 26724 9490 26740
rect 9506 26724 9522 26740
rect 9538 26724 9554 26740
rect 9570 26724 9586 26740
rect 9602 26724 9618 26740
rect 9634 26724 10100 26740
rect 9081 26708 10100 26724
rect 9081 26692 9106 26708
rect 9122 26692 9138 26708
rect 9154 26692 9170 26708
rect 9186 26692 9202 26708
rect 9218 26692 9234 26708
rect 9250 26692 9266 26708
rect 9282 26692 9298 26708
rect 9314 26692 9330 26708
rect 9346 26692 9362 26708
rect 9378 26692 9394 26708
rect 9410 26692 9426 26708
rect 9442 26692 9458 26708
rect 9474 26692 9490 26708
rect 9506 26692 9522 26708
rect 9538 26692 9554 26708
rect 9570 26692 9586 26708
rect 9602 26692 9618 26708
rect 9634 26692 10100 26708
rect 9081 26676 10100 26692
rect 9081 26660 9106 26676
rect 9122 26660 9138 26676
rect 9154 26660 9170 26676
rect 9186 26660 9202 26676
rect 9218 26660 9234 26676
rect 9250 26660 9266 26676
rect 9282 26660 9298 26676
rect 9314 26660 9330 26676
rect 9346 26660 9362 26676
rect 9378 26660 9394 26676
rect 9410 26660 9426 26676
rect 9442 26660 9458 26676
rect 9474 26660 9490 26676
rect 9506 26660 9522 26676
rect 9538 26660 9554 26676
rect 9570 26660 9586 26676
rect 9602 26660 9618 26676
rect 9634 26660 10100 26676
rect 9081 26644 10100 26660
rect 9081 26628 9106 26644
rect 9122 26628 9138 26644
rect 9154 26628 9170 26644
rect 9186 26628 9202 26644
rect 9218 26628 9234 26644
rect 9250 26628 9266 26644
rect 9282 26628 9298 26644
rect 9314 26628 9330 26644
rect 9346 26628 9362 26644
rect 9378 26628 9394 26644
rect 9410 26628 9426 26644
rect 9442 26628 9458 26644
rect 9474 26628 9490 26644
rect 9506 26628 9522 26644
rect 9538 26628 9554 26644
rect 9570 26628 9586 26644
rect 9602 26628 9618 26644
rect 9634 26628 10100 26644
rect 9081 26612 10100 26628
rect 9081 26596 9106 26612
rect 9122 26596 9138 26612
rect 9154 26596 9170 26612
rect 9186 26596 9202 26612
rect 9218 26596 9234 26612
rect 9250 26596 9266 26612
rect 9282 26596 9298 26612
rect 9314 26596 9330 26612
rect 9346 26596 9362 26612
rect 9378 26596 9394 26612
rect 9410 26596 9426 26612
rect 9442 26596 9458 26612
rect 9474 26596 9490 26612
rect 9506 26596 9522 26612
rect 9538 26596 9554 26612
rect 9570 26596 9586 26612
rect 9602 26596 9618 26612
rect 9634 26596 10100 26612
rect 9081 26580 10100 26596
rect 9081 26564 9106 26580
rect 9122 26564 9138 26580
rect 9154 26564 9170 26580
rect 9186 26564 9202 26580
rect 9218 26564 9234 26580
rect 9250 26564 9266 26580
rect 9282 26564 9298 26580
rect 9314 26564 9330 26580
rect 9346 26564 9362 26580
rect 9378 26564 9394 26580
rect 9410 26564 9426 26580
rect 9442 26564 9458 26580
rect 9474 26564 9490 26580
rect 9506 26564 9522 26580
rect 9538 26564 9554 26580
rect 9570 26564 9586 26580
rect 9602 26564 9618 26580
rect 9634 26564 10100 26580
rect 9081 26548 10100 26564
rect 9081 26532 9106 26548
rect 9122 26532 9138 26548
rect 9154 26532 9170 26548
rect 9186 26532 9202 26548
rect 9218 26532 9234 26548
rect 9250 26532 9266 26548
rect 9282 26532 9298 26548
rect 9314 26532 9330 26548
rect 9346 26532 9362 26548
rect 9378 26532 9394 26548
rect 9410 26532 9426 26548
rect 9442 26532 9458 26548
rect 9474 26532 9490 26548
rect 9506 26532 9522 26548
rect 9538 26532 9554 26548
rect 9570 26532 9586 26548
rect 9602 26532 9618 26548
rect 9634 26532 10100 26548
rect 9081 26521 10100 26532
rect 9660 26520 10100 26521
rect 14740 9419 23940 9420
rect 14661 9404 24019 9419
rect 14661 9388 14676 9404
rect 14692 9388 14708 9404
rect 14724 9388 23956 9404
rect 23972 9388 23988 9404
rect 24004 9388 24019 9404
rect 14661 9372 24019 9388
rect 14661 9356 14676 9372
rect 14692 9356 14708 9372
rect 14724 9356 23956 9372
rect 23972 9356 23988 9372
rect 24004 9356 24019 9372
rect 14661 9341 24019 9356
rect 14740 9340 23940 9341
rect 12040 9259 24100 9260
rect 11961 9244 24179 9259
rect 11961 9228 11976 9244
rect 11992 9228 12008 9244
rect 12024 9228 24116 9244
rect 24132 9228 24148 9244
rect 24164 9228 24179 9244
rect 11961 9212 24179 9228
rect 11961 9196 11976 9212
rect 11992 9196 12008 9212
rect 12024 9196 24116 9212
rect 24132 9196 24148 9212
rect 24164 9196 24179 9212
rect 11961 9181 24179 9196
rect 12040 9180 24100 9181
<< m2contact >>
rect 10076 28950 10092 28966
rect 10108 28950 10124 28966
rect 10140 28950 10156 28966
rect 10172 28950 10188 28966
rect 10204 28950 10220 28966
rect 10236 28950 10252 28966
rect 10268 28950 10284 28966
rect 10300 28950 10316 28966
rect 10332 28950 10348 28966
rect 10364 28950 10380 28966
rect 10396 28950 10412 28966
rect 10428 28950 10444 28966
rect 10460 28950 10476 28966
rect 10492 28950 10508 28966
rect 10524 28950 10540 28966
rect 10556 28950 10572 28966
rect 10588 28950 10604 28966
rect 10620 28950 10636 28966
rect 10652 28950 10668 28966
rect 10684 28950 10700 28966
rect 10716 28950 10732 28966
rect 10748 28950 10764 28966
rect 10780 28950 10796 28966
rect 10812 28950 10828 28966
rect 10844 28950 10860 28966
rect 10876 28950 10892 28966
rect 10908 28950 10924 28966
rect 10940 28950 10956 28966
rect 10972 28950 10988 28966
rect 11004 28950 11020 28966
rect 11036 28950 11052 28966
rect 11068 28950 11084 28966
rect 11100 28950 11116 28966
rect 11132 28950 11148 28966
rect 11164 28950 11180 28966
rect 11196 28950 11212 28966
rect 11228 28950 11244 28966
rect 11260 28950 11276 28966
rect 11292 28950 11308 28966
rect 11324 28950 11340 28966
rect 11356 28950 11372 28966
rect 11388 28950 11404 28966
rect 11420 28950 11436 28966
rect 11452 28950 11468 28966
rect 11484 28950 11500 28966
rect 11516 28950 11532 28966
rect 11548 28950 11564 28966
rect 11580 28950 11596 28966
rect 11612 28950 11628 28966
rect 11644 28950 11660 28966
rect 11676 28950 11692 28966
rect 11708 28950 11724 28966
rect 10076 28918 10092 28934
rect 10108 28918 10124 28934
rect 10140 28918 10156 28934
rect 10172 28918 10188 28934
rect 10204 28918 10220 28934
rect 10236 28918 10252 28934
rect 10268 28918 10284 28934
rect 10300 28918 10316 28934
rect 10332 28918 10348 28934
rect 10364 28918 10380 28934
rect 10396 28918 10412 28934
rect 10428 28918 10444 28934
rect 10460 28918 10476 28934
rect 10492 28918 10508 28934
rect 10524 28918 10540 28934
rect 10556 28918 10572 28934
rect 10588 28918 10604 28934
rect 10620 28918 10636 28934
rect 10652 28918 10668 28934
rect 10684 28918 10700 28934
rect 10716 28918 10732 28934
rect 10748 28918 10764 28934
rect 10780 28918 10796 28934
rect 10812 28918 10828 28934
rect 10844 28918 10860 28934
rect 10876 28918 10892 28934
rect 10908 28918 10924 28934
rect 10940 28918 10956 28934
rect 10972 28918 10988 28934
rect 11004 28918 11020 28934
rect 11036 28918 11052 28934
rect 11068 28918 11084 28934
rect 11100 28918 11116 28934
rect 11132 28918 11148 28934
rect 11164 28918 11180 28934
rect 11196 28918 11212 28934
rect 11228 28918 11244 28934
rect 11260 28918 11276 28934
rect 11292 28918 11308 28934
rect 11324 28918 11340 28934
rect 11356 28918 11372 28934
rect 11388 28918 11404 28934
rect 11420 28918 11436 28934
rect 11452 28918 11468 28934
rect 11484 28918 11500 28934
rect 11516 28918 11532 28934
rect 11548 28918 11564 28934
rect 11580 28918 11596 28934
rect 11612 28918 11628 28934
rect 11644 28918 11660 28934
rect 11676 28918 11692 28934
rect 11708 28918 11724 28934
rect 10076 28886 10092 28902
rect 10108 28886 10124 28902
rect 10140 28886 10156 28902
rect 10172 28886 10188 28902
rect 10204 28886 10220 28902
rect 10236 28886 10252 28902
rect 10268 28886 10284 28902
rect 10300 28886 10316 28902
rect 10332 28886 10348 28902
rect 10364 28886 10380 28902
rect 10396 28886 10412 28902
rect 10428 28886 10444 28902
rect 10460 28886 10476 28902
rect 10492 28886 10508 28902
rect 10524 28886 10540 28902
rect 10556 28886 10572 28902
rect 10588 28886 10604 28902
rect 10620 28886 10636 28902
rect 10652 28886 10668 28902
rect 10684 28886 10700 28902
rect 10716 28886 10732 28902
rect 10748 28886 10764 28902
rect 10780 28886 10796 28902
rect 10812 28886 10828 28902
rect 10844 28886 10860 28902
rect 10876 28886 10892 28902
rect 10908 28886 10924 28902
rect 10940 28886 10956 28902
rect 10972 28886 10988 28902
rect 11004 28886 11020 28902
rect 11036 28886 11052 28902
rect 11068 28886 11084 28902
rect 11100 28886 11116 28902
rect 11132 28886 11148 28902
rect 11164 28886 11180 28902
rect 11196 28886 11212 28902
rect 11228 28886 11244 28902
rect 11260 28886 11276 28902
rect 11292 28886 11308 28902
rect 11324 28886 11340 28902
rect 11356 28886 11372 28902
rect 11388 28886 11404 28902
rect 11420 28886 11436 28902
rect 11452 28886 11468 28902
rect 11484 28886 11500 28902
rect 11516 28886 11532 28902
rect 11548 28886 11564 28902
rect 11580 28886 11596 28902
rect 11612 28886 11628 28902
rect 11644 28886 11660 28902
rect 11676 28886 11692 28902
rect 11708 28886 11724 28902
rect 10076 28854 10092 28870
rect 10108 28854 10124 28870
rect 10140 28854 10156 28870
rect 10172 28854 10188 28870
rect 10204 28854 10220 28870
rect 10236 28854 10252 28870
rect 10268 28854 10284 28870
rect 10300 28854 10316 28870
rect 10332 28854 10348 28870
rect 10364 28854 10380 28870
rect 10396 28854 10412 28870
rect 10428 28854 10444 28870
rect 10460 28854 10476 28870
rect 10492 28854 10508 28870
rect 10524 28854 10540 28870
rect 10556 28854 10572 28870
rect 10588 28854 10604 28870
rect 10620 28854 10636 28870
rect 10652 28854 10668 28870
rect 10684 28854 10700 28870
rect 10716 28854 10732 28870
rect 10748 28854 10764 28870
rect 10780 28854 10796 28870
rect 10812 28854 10828 28870
rect 10844 28854 10860 28870
rect 10876 28854 10892 28870
rect 10908 28854 10924 28870
rect 10940 28854 10956 28870
rect 10972 28854 10988 28870
rect 11004 28854 11020 28870
rect 11036 28854 11052 28870
rect 11068 28854 11084 28870
rect 11100 28854 11116 28870
rect 11132 28854 11148 28870
rect 11164 28854 11180 28870
rect 11196 28854 11212 28870
rect 11228 28854 11244 28870
rect 11260 28854 11276 28870
rect 11292 28854 11308 28870
rect 11324 28854 11340 28870
rect 11356 28854 11372 28870
rect 11388 28854 11404 28870
rect 11420 28854 11436 28870
rect 11452 28854 11468 28870
rect 11484 28854 11500 28870
rect 11516 28854 11532 28870
rect 11548 28854 11564 28870
rect 11580 28854 11596 28870
rect 11612 28854 11628 28870
rect 11644 28854 11660 28870
rect 11676 28854 11692 28870
rect 11708 28854 11724 28870
rect 10076 28822 10092 28838
rect 10108 28822 10124 28838
rect 10140 28822 10156 28838
rect 10172 28822 10188 28838
rect 10204 28822 10220 28838
rect 10236 28822 10252 28838
rect 10268 28822 10284 28838
rect 10300 28822 10316 28838
rect 10332 28822 10348 28838
rect 10364 28822 10380 28838
rect 10396 28822 10412 28838
rect 10428 28822 10444 28838
rect 10460 28822 10476 28838
rect 10492 28822 10508 28838
rect 10524 28822 10540 28838
rect 10556 28822 10572 28838
rect 10588 28822 10604 28838
rect 10620 28822 10636 28838
rect 10652 28822 10668 28838
rect 10684 28822 10700 28838
rect 10716 28822 10732 28838
rect 10748 28822 10764 28838
rect 10780 28822 10796 28838
rect 10812 28822 10828 28838
rect 10844 28822 10860 28838
rect 10876 28822 10892 28838
rect 10908 28822 10924 28838
rect 10940 28822 10956 28838
rect 10972 28822 10988 28838
rect 11004 28822 11020 28838
rect 11036 28822 11052 28838
rect 11068 28822 11084 28838
rect 11100 28822 11116 28838
rect 11132 28822 11148 28838
rect 11164 28822 11180 28838
rect 11196 28822 11212 28838
rect 11228 28822 11244 28838
rect 11260 28822 11276 28838
rect 11292 28822 11308 28838
rect 11324 28822 11340 28838
rect 11356 28822 11372 28838
rect 11388 28822 11404 28838
rect 11420 28822 11436 28838
rect 11452 28822 11468 28838
rect 11484 28822 11500 28838
rect 11516 28822 11532 28838
rect 11548 28822 11564 28838
rect 11580 28822 11596 28838
rect 11612 28822 11628 28838
rect 11644 28822 11660 28838
rect 11676 28822 11692 28838
rect 11708 28822 11724 28838
rect 10076 28790 10092 28806
rect 10108 28790 10124 28806
rect 10140 28790 10156 28806
rect 10172 28790 10188 28806
rect 10204 28790 10220 28806
rect 10236 28790 10252 28806
rect 10268 28790 10284 28806
rect 10300 28790 10316 28806
rect 10332 28790 10348 28806
rect 10364 28790 10380 28806
rect 10396 28790 10412 28806
rect 10428 28790 10444 28806
rect 10460 28790 10476 28806
rect 10492 28790 10508 28806
rect 10524 28790 10540 28806
rect 10556 28790 10572 28806
rect 10588 28790 10604 28806
rect 10620 28790 10636 28806
rect 10652 28790 10668 28806
rect 10684 28790 10700 28806
rect 10716 28790 10732 28806
rect 10748 28790 10764 28806
rect 10780 28790 10796 28806
rect 10812 28790 10828 28806
rect 10844 28790 10860 28806
rect 10876 28790 10892 28806
rect 10908 28790 10924 28806
rect 10940 28790 10956 28806
rect 10972 28790 10988 28806
rect 11004 28790 11020 28806
rect 11036 28790 11052 28806
rect 11068 28790 11084 28806
rect 11100 28790 11116 28806
rect 11132 28790 11148 28806
rect 11164 28790 11180 28806
rect 11196 28790 11212 28806
rect 11228 28790 11244 28806
rect 11260 28790 11276 28806
rect 11292 28790 11308 28806
rect 11324 28790 11340 28806
rect 11356 28790 11372 28806
rect 11388 28790 11404 28806
rect 11420 28790 11436 28806
rect 11452 28790 11468 28806
rect 11484 28790 11500 28806
rect 11516 28790 11532 28806
rect 11548 28790 11564 28806
rect 11580 28790 11596 28806
rect 11612 28790 11628 28806
rect 11644 28790 11660 28806
rect 11676 28790 11692 28806
rect 11708 28790 11724 28806
rect 10076 28758 10092 28774
rect 10108 28758 10124 28774
rect 10140 28758 10156 28774
rect 10172 28758 10188 28774
rect 10204 28758 10220 28774
rect 10236 28758 10252 28774
rect 10268 28758 10284 28774
rect 10300 28758 10316 28774
rect 10332 28758 10348 28774
rect 10364 28758 10380 28774
rect 10396 28758 10412 28774
rect 10428 28758 10444 28774
rect 10460 28758 10476 28774
rect 10492 28758 10508 28774
rect 10524 28758 10540 28774
rect 10556 28758 10572 28774
rect 10588 28758 10604 28774
rect 10620 28758 10636 28774
rect 10652 28758 10668 28774
rect 10684 28758 10700 28774
rect 10716 28758 10732 28774
rect 10748 28758 10764 28774
rect 10780 28758 10796 28774
rect 10812 28758 10828 28774
rect 10844 28758 10860 28774
rect 10876 28758 10892 28774
rect 10908 28758 10924 28774
rect 10940 28758 10956 28774
rect 10972 28758 10988 28774
rect 11004 28758 11020 28774
rect 11036 28758 11052 28774
rect 11068 28758 11084 28774
rect 11100 28758 11116 28774
rect 11132 28758 11148 28774
rect 11164 28758 11180 28774
rect 11196 28758 11212 28774
rect 11228 28758 11244 28774
rect 11260 28758 11276 28774
rect 11292 28758 11308 28774
rect 11324 28758 11340 28774
rect 11356 28758 11372 28774
rect 11388 28758 11404 28774
rect 11420 28758 11436 28774
rect 11452 28758 11468 28774
rect 11484 28758 11500 28774
rect 11516 28758 11532 28774
rect 11548 28758 11564 28774
rect 11580 28758 11596 28774
rect 11612 28758 11628 28774
rect 11644 28758 11660 28774
rect 11676 28758 11692 28774
rect 11708 28758 11724 28774
rect 10076 28726 10092 28742
rect 10108 28726 10124 28742
rect 10140 28726 10156 28742
rect 10172 28726 10188 28742
rect 10204 28726 10220 28742
rect 10236 28726 10252 28742
rect 10268 28726 10284 28742
rect 10300 28726 10316 28742
rect 10332 28726 10348 28742
rect 10364 28726 10380 28742
rect 10396 28726 10412 28742
rect 10428 28726 10444 28742
rect 10460 28726 10476 28742
rect 10492 28726 10508 28742
rect 10524 28726 10540 28742
rect 10556 28726 10572 28742
rect 10588 28726 10604 28742
rect 10620 28726 10636 28742
rect 10652 28726 10668 28742
rect 10684 28726 10700 28742
rect 10716 28726 10732 28742
rect 10748 28726 10764 28742
rect 10780 28726 10796 28742
rect 10812 28726 10828 28742
rect 10844 28726 10860 28742
rect 10876 28726 10892 28742
rect 10908 28726 10924 28742
rect 10940 28726 10956 28742
rect 10972 28726 10988 28742
rect 11004 28726 11020 28742
rect 11036 28726 11052 28742
rect 11068 28726 11084 28742
rect 11100 28726 11116 28742
rect 11132 28726 11148 28742
rect 11164 28726 11180 28742
rect 11196 28726 11212 28742
rect 11228 28726 11244 28742
rect 11260 28726 11276 28742
rect 11292 28726 11308 28742
rect 11324 28726 11340 28742
rect 11356 28726 11372 28742
rect 11388 28726 11404 28742
rect 11420 28726 11436 28742
rect 11452 28726 11468 28742
rect 11484 28726 11500 28742
rect 11516 28726 11532 28742
rect 11548 28726 11564 28742
rect 11580 28726 11596 28742
rect 11612 28726 11628 28742
rect 11644 28726 11660 28742
rect 11676 28726 11692 28742
rect 11708 28726 11724 28742
rect 10076 28694 10092 28710
rect 10108 28694 10124 28710
rect 10140 28694 10156 28710
rect 10172 28694 10188 28710
rect 10204 28694 10220 28710
rect 10236 28694 10252 28710
rect 10268 28694 10284 28710
rect 10300 28694 10316 28710
rect 10332 28694 10348 28710
rect 10364 28694 10380 28710
rect 10396 28694 10412 28710
rect 10428 28694 10444 28710
rect 10460 28694 10476 28710
rect 10492 28694 10508 28710
rect 10524 28694 10540 28710
rect 10556 28694 10572 28710
rect 10588 28694 10604 28710
rect 10620 28694 10636 28710
rect 10652 28694 10668 28710
rect 10684 28694 10700 28710
rect 10716 28694 10732 28710
rect 10748 28694 10764 28710
rect 10780 28694 10796 28710
rect 10812 28694 10828 28710
rect 10844 28694 10860 28710
rect 10876 28694 10892 28710
rect 10908 28694 10924 28710
rect 10940 28694 10956 28710
rect 10972 28694 10988 28710
rect 11004 28694 11020 28710
rect 11036 28694 11052 28710
rect 11068 28694 11084 28710
rect 11100 28694 11116 28710
rect 11132 28694 11148 28710
rect 11164 28694 11180 28710
rect 11196 28694 11212 28710
rect 11228 28694 11244 28710
rect 11260 28694 11276 28710
rect 11292 28694 11308 28710
rect 11324 28694 11340 28710
rect 11356 28694 11372 28710
rect 11388 28694 11404 28710
rect 11420 28694 11436 28710
rect 11452 28694 11468 28710
rect 11484 28694 11500 28710
rect 11516 28694 11532 28710
rect 11548 28694 11564 28710
rect 11580 28694 11596 28710
rect 11612 28694 11628 28710
rect 11644 28694 11660 28710
rect 11676 28694 11692 28710
rect 11708 28694 11724 28710
rect 9106 27652 9122 27668
rect 9138 27652 9154 27668
rect 9170 27652 9186 27668
rect 9202 27652 9218 27668
rect 9234 27652 9250 27668
rect 9266 27652 9282 27668
rect 9298 27652 9314 27668
rect 9330 27652 9346 27668
rect 9362 27652 9378 27668
rect 9394 27652 9410 27668
rect 9426 27652 9442 27668
rect 9458 27652 9474 27668
rect 9490 27652 9506 27668
rect 9522 27652 9538 27668
rect 9554 27652 9570 27668
rect 9586 27652 9602 27668
rect 9618 27652 9634 27668
rect 9106 27620 9122 27636
rect 9138 27620 9154 27636
rect 9170 27620 9186 27636
rect 9202 27620 9218 27636
rect 9234 27620 9250 27636
rect 9266 27620 9282 27636
rect 9298 27620 9314 27636
rect 9330 27620 9346 27636
rect 9362 27620 9378 27636
rect 9394 27620 9410 27636
rect 9426 27620 9442 27636
rect 9458 27620 9474 27636
rect 9490 27620 9506 27636
rect 9522 27620 9538 27636
rect 9554 27620 9570 27636
rect 9586 27620 9602 27636
rect 9618 27620 9634 27636
rect 9106 27588 9122 27604
rect 9138 27588 9154 27604
rect 9170 27588 9186 27604
rect 9202 27588 9218 27604
rect 9234 27588 9250 27604
rect 9266 27588 9282 27604
rect 9298 27588 9314 27604
rect 9330 27588 9346 27604
rect 9362 27588 9378 27604
rect 9394 27588 9410 27604
rect 9426 27588 9442 27604
rect 9458 27588 9474 27604
rect 9490 27588 9506 27604
rect 9522 27588 9538 27604
rect 9554 27588 9570 27604
rect 9586 27588 9602 27604
rect 9618 27588 9634 27604
rect 9106 27556 9122 27572
rect 9138 27556 9154 27572
rect 9170 27556 9186 27572
rect 9202 27556 9218 27572
rect 9234 27556 9250 27572
rect 9266 27556 9282 27572
rect 9298 27556 9314 27572
rect 9330 27556 9346 27572
rect 9362 27556 9378 27572
rect 9394 27556 9410 27572
rect 9426 27556 9442 27572
rect 9458 27556 9474 27572
rect 9490 27556 9506 27572
rect 9522 27556 9538 27572
rect 9554 27556 9570 27572
rect 9586 27556 9602 27572
rect 9618 27556 9634 27572
rect 9106 27524 9122 27540
rect 9138 27524 9154 27540
rect 9170 27524 9186 27540
rect 9202 27524 9218 27540
rect 9234 27524 9250 27540
rect 9266 27524 9282 27540
rect 9298 27524 9314 27540
rect 9330 27524 9346 27540
rect 9362 27524 9378 27540
rect 9394 27524 9410 27540
rect 9426 27524 9442 27540
rect 9458 27524 9474 27540
rect 9490 27524 9506 27540
rect 9522 27524 9538 27540
rect 9554 27524 9570 27540
rect 9586 27524 9602 27540
rect 9618 27524 9634 27540
rect 9106 27492 9122 27508
rect 9138 27492 9154 27508
rect 9170 27492 9186 27508
rect 9202 27492 9218 27508
rect 9234 27492 9250 27508
rect 9266 27492 9282 27508
rect 9298 27492 9314 27508
rect 9330 27492 9346 27508
rect 9362 27492 9378 27508
rect 9394 27492 9410 27508
rect 9426 27492 9442 27508
rect 9458 27492 9474 27508
rect 9490 27492 9506 27508
rect 9522 27492 9538 27508
rect 9554 27492 9570 27508
rect 9586 27492 9602 27508
rect 9618 27492 9634 27508
rect 9106 27460 9122 27476
rect 9138 27460 9154 27476
rect 9170 27460 9186 27476
rect 9202 27460 9218 27476
rect 9234 27460 9250 27476
rect 9266 27460 9282 27476
rect 9298 27460 9314 27476
rect 9330 27460 9346 27476
rect 9362 27460 9378 27476
rect 9394 27460 9410 27476
rect 9426 27460 9442 27476
rect 9458 27460 9474 27476
rect 9490 27460 9506 27476
rect 9522 27460 9538 27476
rect 9554 27460 9570 27476
rect 9586 27460 9602 27476
rect 9618 27460 9634 27476
rect 9106 27428 9122 27444
rect 9138 27428 9154 27444
rect 9170 27428 9186 27444
rect 9202 27428 9218 27444
rect 9234 27428 9250 27444
rect 9266 27428 9282 27444
rect 9298 27428 9314 27444
rect 9330 27428 9346 27444
rect 9362 27428 9378 27444
rect 9394 27428 9410 27444
rect 9426 27428 9442 27444
rect 9458 27428 9474 27444
rect 9490 27428 9506 27444
rect 9522 27428 9538 27444
rect 9554 27428 9570 27444
rect 9586 27428 9602 27444
rect 9618 27428 9634 27444
rect 9106 27396 9122 27412
rect 9138 27396 9154 27412
rect 9170 27396 9186 27412
rect 9202 27396 9218 27412
rect 9234 27396 9250 27412
rect 9266 27396 9282 27412
rect 9298 27396 9314 27412
rect 9330 27396 9346 27412
rect 9362 27396 9378 27412
rect 9394 27396 9410 27412
rect 9426 27396 9442 27412
rect 9458 27396 9474 27412
rect 9490 27396 9506 27412
rect 9522 27396 9538 27412
rect 9554 27396 9570 27412
rect 9586 27396 9602 27412
rect 9618 27396 9634 27412
rect 9106 27364 9122 27380
rect 9138 27364 9154 27380
rect 9170 27364 9186 27380
rect 9202 27364 9218 27380
rect 9234 27364 9250 27380
rect 9266 27364 9282 27380
rect 9298 27364 9314 27380
rect 9330 27364 9346 27380
rect 9362 27364 9378 27380
rect 9394 27364 9410 27380
rect 9426 27364 9442 27380
rect 9458 27364 9474 27380
rect 9490 27364 9506 27380
rect 9522 27364 9538 27380
rect 9554 27364 9570 27380
rect 9586 27364 9602 27380
rect 9618 27364 9634 27380
rect 9106 27332 9122 27348
rect 9138 27332 9154 27348
rect 9170 27332 9186 27348
rect 9202 27332 9218 27348
rect 9234 27332 9250 27348
rect 9266 27332 9282 27348
rect 9298 27332 9314 27348
rect 9330 27332 9346 27348
rect 9362 27332 9378 27348
rect 9394 27332 9410 27348
rect 9426 27332 9442 27348
rect 9458 27332 9474 27348
rect 9490 27332 9506 27348
rect 9522 27332 9538 27348
rect 9554 27332 9570 27348
rect 9586 27332 9602 27348
rect 9618 27332 9634 27348
rect 9106 27300 9122 27316
rect 9138 27300 9154 27316
rect 9170 27300 9186 27316
rect 9202 27300 9218 27316
rect 9234 27300 9250 27316
rect 9266 27300 9282 27316
rect 9298 27300 9314 27316
rect 9330 27300 9346 27316
rect 9362 27300 9378 27316
rect 9394 27300 9410 27316
rect 9426 27300 9442 27316
rect 9458 27300 9474 27316
rect 9490 27300 9506 27316
rect 9522 27300 9538 27316
rect 9554 27300 9570 27316
rect 9586 27300 9602 27316
rect 9618 27300 9634 27316
rect 9106 27268 9122 27284
rect 9138 27268 9154 27284
rect 9170 27268 9186 27284
rect 9202 27268 9218 27284
rect 9234 27268 9250 27284
rect 9266 27268 9282 27284
rect 9298 27268 9314 27284
rect 9330 27268 9346 27284
rect 9362 27268 9378 27284
rect 9394 27268 9410 27284
rect 9426 27268 9442 27284
rect 9458 27268 9474 27284
rect 9490 27268 9506 27284
rect 9522 27268 9538 27284
rect 9554 27268 9570 27284
rect 9586 27268 9602 27284
rect 9618 27268 9634 27284
rect 9106 27236 9122 27252
rect 9138 27236 9154 27252
rect 9170 27236 9186 27252
rect 9202 27236 9218 27252
rect 9234 27236 9250 27252
rect 9266 27236 9282 27252
rect 9298 27236 9314 27252
rect 9330 27236 9346 27252
rect 9362 27236 9378 27252
rect 9394 27236 9410 27252
rect 9426 27236 9442 27252
rect 9458 27236 9474 27252
rect 9490 27236 9506 27252
rect 9522 27236 9538 27252
rect 9554 27236 9570 27252
rect 9586 27236 9602 27252
rect 9618 27236 9634 27252
rect 9106 27204 9122 27220
rect 9138 27204 9154 27220
rect 9170 27204 9186 27220
rect 9202 27204 9218 27220
rect 9234 27204 9250 27220
rect 9266 27204 9282 27220
rect 9298 27204 9314 27220
rect 9330 27204 9346 27220
rect 9362 27204 9378 27220
rect 9394 27204 9410 27220
rect 9426 27204 9442 27220
rect 9458 27204 9474 27220
rect 9490 27204 9506 27220
rect 9522 27204 9538 27220
rect 9554 27204 9570 27220
rect 9586 27204 9602 27220
rect 9618 27204 9634 27220
rect 9106 27172 9122 27188
rect 9138 27172 9154 27188
rect 9170 27172 9186 27188
rect 9202 27172 9218 27188
rect 9234 27172 9250 27188
rect 9266 27172 9282 27188
rect 9298 27172 9314 27188
rect 9330 27172 9346 27188
rect 9362 27172 9378 27188
rect 9394 27172 9410 27188
rect 9426 27172 9442 27188
rect 9458 27172 9474 27188
rect 9490 27172 9506 27188
rect 9522 27172 9538 27188
rect 9554 27172 9570 27188
rect 9586 27172 9602 27188
rect 9618 27172 9634 27188
rect 9106 27140 9122 27156
rect 9138 27140 9154 27156
rect 9170 27140 9186 27156
rect 9202 27140 9218 27156
rect 9234 27140 9250 27156
rect 9266 27140 9282 27156
rect 9298 27140 9314 27156
rect 9330 27140 9346 27156
rect 9362 27140 9378 27156
rect 9394 27140 9410 27156
rect 9426 27140 9442 27156
rect 9458 27140 9474 27156
rect 9490 27140 9506 27156
rect 9522 27140 9538 27156
rect 9554 27140 9570 27156
rect 9586 27140 9602 27156
rect 9618 27140 9634 27156
rect 9106 27108 9122 27124
rect 9138 27108 9154 27124
rect 9170 27108 9186 27124
rect 9202 27108 9218 27124
rect 9234 27108 9250 27124
rect 9266 27108 9282 27124
rect 9298 27108 9314 27124
rect 9330 27108 9346 27124
rect 9362 27108 9378 27124
rect 9394 27108 9410 27124
rect 9426 27108 9442 27124
rect 9458 27108 9474 27124
rect 9490 27108 9506 27124
rect 9522 27108 9538 27124
rect 9554 27108 9570 27124
rect 9586 27108 9602 27124
rect 9618 27108 9634 27124
rect 9106 27076 9122 27092
rect 9138 27076 9154 27092
rect 9170 27076 9186 27092
rect 9202 27076 9218 27092
rect 9234 27076 9250 27092
rect 9266 27076 9282 27092
rect 9298 27076 9314 27092
rect 9330 27076 9346 27092
rect 9362 27076 9378 27092
rect 9394 27076 9410 27092
rect 9426 27076 9442 27092
rect 9458 27076 9474 27092
rect 9490 27076 9506 27092
rect 9522 27076 9538 27092
rect 9554 27076 9570 27092
rect 9586 27076 9602 27092
rect 9618 27076 9634 27092
rect 9106 27044 9122 27060
rect 9138 27044 9154 27060
rect 9170 27044 9186 27060
rect 9202 27044 9218 27060
rect 9234 27044 9250 27060
rect 9266 27044 9282 27060
rect 9298 27044 9314 27060
rect 9330 27044 9346 27060
rect 9362 27044 9378 27060
rect 9394 27044 9410 27060
rect 9426 27044 9442 27060
rect 9458 27044 9474 27060
rect 9490 27044 9506 27060
rect 9522 27044 9538 27060
rect 9554 27044 9570 27060
rect 9586 27044 9602 27060
rect 9618 27044 9634 27060
rect 9106 27012 9122 27028
rect 9138 27012 9154 27028
rect 9170 27012 9186 27028
rect 9202 27012 9218 27028
rect 9234 27012 9250 27028
rect 9266 27012 9282 27028
rect 9298 27012 9314 27028
rect 9330 27012 9346 27028
rect 9362 27012 9378 27028
rect 9394 27012 9410 27028
rect 9426 27012 9442 27028
rect 9458 27012 9474 27028
rect 9490 27012 9506 27028
rect 9522 27012 9538 27028
rect 9554 27012 9570 27028
rect 9586 27012 9602 27028
rect 9618 27012 9634 27028
rect 9106 26980 9122 26996
rect 9138 26980 9154 26996
rect 9170 26980 9186 26996
rect 9202 26980 9218 26996
rect 9234 26980 9250 26996
rect 9266 26980 9282 26996
rect 9298 26980 9314 26996
rect 9330 26980 9346 26996
rect 9362 26980 9378 26996
rect 9394 26980 9410 26996
rect 9426 26980 9442 26996
rect 9458 26980 9474 26996
rect 9490 26980 9506 26996
rect 9522 26980 9538 26996
rect 9554 26980 9570 26996
rect 9586 26980 9602 26996
rect 9618 26980 9634 26996
rect 9106 26948 9122 26964
rect 9138 26948 9154 26964
rect 9170 26948 9186 26964
rect 9202 26948 9218 26964
rect 9234 26948 9250 26964
rect 9266 26948 9282 26964
rect 9298 26948 9314 26964
rect 9330 26948 9346 26964
rect 9362 26948 9378 26964
rect 9394 26948 9410 26964
rect 9426 26948 9442 26964
rect 9458 26948 9474 26964
rect 9490 26948 9506 26964
rect 9522 26948 9538 26964
rect 9554 26948 9570 26964
rect 9586 26948 9602 26964
rect 9618 26948 9634 26964
rect 9106 26916 9122 26932
rect 9138 26916 9154 26932
rect 9170 26916 9186 26932
rect 9202 26916 9218 26932
rect 9234 26916 9250 26932
rect 9266 26916 9282 26932
rect 9298 26916 9314 26932
rect 9330 26916 9346 26932
rect 9362 26916 9378 26932
rect 9394 26916 9410 26932
rect 9426 26916 9442 26932
rect 9458 26916 9474 26932
rect 9490 26916 9506 26932
rect 9522 26916 9538 26932
rect 9554 26916 9570 26932
rect 9586 26916 9602 26932
rect 9618 26916 9634 26932
rect 9106 26884 9122 26900
rect 9138 26884 9154 26900
rect 9170 26884 9186 26900
rect 9202 26884 9218 26900
rect 9234 26884 9250 26900
rect 9266 26884 9282 26900
rect 9298 26884 9314 26900
rect 9330 26884 9346 26900
rect 9362 26884 9378 26900
rect 9394 26884 9410 26900
rect 9426 26884 9442 26900
rect 9458 26884 9474 26900
rect 9490 26884 9506 26900
rect 9522 26884 9538 26900
rect 9554 26884 9570 26900
rect 9586 26884 9602 26900
rect 9618 26884 9634 26900
rect 9106 26852 9122 26868
rect 9138 26852 9154 26868
rect 9170 26852 9186 26868
rect 9202 26852 9218 26868
rect 9234 26852 9250 26868
rect 9266 26852 9282 26868
rect 9298 26852 9314 26868
rect 9330 26852 9346 26868
rect 9362 26852 9378 26868
rect 9394 26852 9410 26868
rect 9426 26852 9442 26868
rect 9458 26852 9474 26868
rect 9490 26852 9506 26868
rect 9522 26852 9538 26868
rect 9554 26852 9570 26868
rect 9586 26852 9602 26868
rect 9618 26852 9634 26868
rect 9106 26820 9122 26836
rect 9138 26820 9154 26836
rect 9170 26820 9186 26836
rect 9202 26820 9218 26836
rect 9234 26820 9250 26836
rect 9266 26820 9282 26836
rect 9298 26820 9314 26836
rect 9330 26820 9346 26836
rect 9362 26820 9378 26836
rect 9394 26820 9410 26836
rect 9426 26820 9442 26836
rect 9458 26820 9474 26836
rect 9490 26820 9506 26836
rect 9522 26820 9538 26836
rect 9554 26820 9570 26836
rect 9586 26820 9602 26836
rect 9618 26820 9634 26836
rect 9106 26788 9122 26804
rect 9138 26788 9154 26804
rect 9170 26788 9186 26804
rect 9202 26788 9218 26804
rect 9234 26788 9250 26804
rect 9266 26788 9282 26804
rect 9298 26788 9314 26804
rect 9330 26788 9346 26804
rect 9362 26788 9378 26804
rect 9394 26788 9410 26804
rect 9426 26788 9442 26804
rect 9458 26788 9474 26804
rect 9490 26788 9506 26804
rect 9522 26788 9538 26804
rect 9554 26788 9570 26804
rect 9586 26788 9602 26804
rect 9618 26788 9634 26804
rect 9106 26756 9122 26772
rect 9138 26756 9154 26772
rect 9170 26756 9186 26772
rect 9202 26756 9218 26772
rect 9234 26756 9250 26772
rect 9266 26756 9282 26772
rect 9298 26756 9314 26772
rect 9330 26756 9346 26772
rect 9362 26756 9378 26772
rect 9394 26756 9410 26772
rect 9426 26756 9442 26772
rect 9458 26756 9474 26772
rect 9490 26756 9506 26772
rect 9522 26756 9538 26772
rect 9554 26756 9570 26772
rect 9586 26756 9602 26772
rect 9618 26756 9634 26772
rect 9106 26724 9122 26740
rect 9138 26724 9154 26740
rect 9170 26724 9186 26740
rect 9202 26724 9218 26740
rect 9234 26724 9250 26740
rect 9266 26724 9282 26740
rect 9298 26724 9314 26740
rect 9330 26724 9346 26740
rect 9362 26724 9378 26740
rect 9394 26724 9410 26740
rect 9426 26724 9442 26740
rect 9458 26724 9474 26740
rect 9490 26724 9506 26740
rect 9522 26724 9538 26740
rect 9554 26724 9570 26740
rect 9586 26724 9602 26740
rect 9618 26724 9634 26740
rect 9106 26692 9122 26708
rect 9138 26692 9154 26708
rect 9170 26692 9186 26708
rect 9202 26692 9218 26708
rect 9234 26692 9250 26708
rect 9266 26692 9282 26708
rect 9298 26692 9314 26708
rect 9330 26692 9346 26708
rect 9362 26692 9378 26708
rect 9394 26692 9410 26708
rect 9426 26692 9442 26708
rect 9458 26692 9474 26708
rect 9490 26692 9506 26708
rect 9522 26692 9538 26708
rect 9554 26692 9570 26708
rect 9586 26692 9602 26708
rect 9618 26692 9634 26708
rect 9106 26660 9122 26676
rect 9138 26660 9154 26676
rect 9170 26660 9186 26676
rect 9202 26660 9218 26676
rect 9234 26660 9250 26676
rect 9266 26660 9282 26676
rect 9298 26660 9314 26676
rect 9330 26660 9346 26676
rect 9362 26660 9378 26676
rect 9394 26660 9410 26676
rect 9426 26660 9442 26676
rect 9458 26660 9474 26676
rect 9490 26660 9506 26676
rect 9522 26660 9538 26676
rect 9554 26660 9570 26676
rect 9586 26660 9602 26676
rect 9618 26660 9634 26676
rect 9106 26628 9122 26644
rect 9138 26628 9154 26644
rect 9170 26628 9186 26644
rect 9202 26628 9218 26644
rect 9234 26628 9250 26644
rect 9266 26628 9282 26644
rect 9298 26628 9314 26644
rect 9330 26628 9346 26644
rect 9362 26628 9378 26644
rect 9394 26628 9410 26644
rect 9426 26628 9442 26644
rect 9458 26628 9474 26644
rect 9490 26628 9506 26644
rect 9522 26628 9538 26644
rect 9554 26628 9570 26644
rect 9586 26628 9602 26644
rect 9618 26628 9634 26644
rect 9106 26596 9122 26612
rect 9138 26596 9154 26612
rect 9170 26596 9186 26612
rect 9202 26596 9218 26612
rect 9234 26596 9250 26612
rect 9266 26596 9282 26612
rect 9298 26596 9314 26612
rect 9330 26596 9346 26612
rect 9362 26596 9378 26612
rect 9394 26596 9410 26612
rect 9426 26596 9442 26612
rect 9458 26596 9474 26612
rect 9490 26596 9506 26612
rect 9522 26596 9538 26612
rect 9554 26596 9570 26612
rect 9586 26596 9602 26612
rect 9618 26596 9634 26612
rect 9106 26564 9122 26580
rect 9138 26564 9154 26580
rect 9170 26564 9186 26580
rect 9202 26564 9218 26580
rect 9234 26564 9250 26580
rect 9266 26564 9282 26580
rect 9298 26564 9314 26580
rect 9330 26564 9346 26580
rect 9362 26564 9378 26580
rect 9394 26564 9410 26580
rect 9426 26564 9442 26580
rect 9458 26564 9474 26580
rect 9490 26564 9506 26580
rect 9522 26564 9538 26580
rect 9554 26564 9570 26580
rect 9586 26564 9602 26580
rect 9618 26564 9634 26580
rect 9106 26532 9122 26548
rect 9138 26532 9154 26548
rect 9170 26532 9186 26548
rect 9202 26532 9218 26548
rect 9234 26532 9250 26548
rect 9266 26532 9282 26548
rect 9298 26532 9314 26548
rect 9330 26532 9346 26548
rect 9362 26532 9378 26548
rect 9394 26532 9410 26548
rect 9426 26532 9442 26548
rect 9458 26532 9474 26548
rect 9490 26532 9506 26548
rect 9522 26532 9538 26548
rect 9554 26532 9570 26548
rect 9586 26532 9602 26548
rect 9618 26532 9634 26548
rect 14676 9388 14692 9404
rect 14708 9388 14724 9404
rect 23956 9388 23972 9404
rect 23988 9388 24004 9404
rect 14676 9356 14692 9372
rect 14708 9356 14724 9372
rect 23956 9356 23972 9372
rect 23988 9356 24004 9372
rect 11976 9228 11992 9244
rect 12008 9228 12024 9244
rect 24116 9228 24132 9244
rect 24148 9228 24164 9244
rect 11976 9196 11992 9212
rect 12008 9196 12024 9212
rect 24116 9196 24132 9212
rect 24148 9196 24164 9212
<< metal2 >>
rect 10060 28980 11740 29180
rect 10061 28966 11739 28980
rect 10061 28950 10076 28966
rect 10092 28950 10108 28966
rect 10124 28950 10140 28966
rect 10156 28950 10172 28966
rect 10188 28950 10204 28966
rect 10220 28950 10236 28966
rect 10252 28950 10268 28966
rect 10284 28950 10300 28966
rect 10316 28950 10332 28966
rect 10348 28950 10364 28966
rect 10380 28950 10396 28966
rect 10412 28950 10428 28966
rect 10444 28950 10460 28966
rect 10476 28950 10492 28966
rect 10508 28950 10524 28966
rect 10540 28950 10556 28966
rect 10572 28950 10588 28966
rect 10604 28950 10620 28966
rect 10636 28950 10652 28966
rect 10668 28950 10684 28966
rect 10700 28950 10716 28966
rect 10732 28950 10748 28966
rect 10764 28950 10780 28966
rect 10796 28950 10812 28966
rect 10828 28950 10844 28966
rect 10860 28950 10876 28966
rect 10892 28950 10908 28966
rect 10924 28950 10940 28966
rect 10956 28950 10972 28966
rect 10988 28950 11004 28966
rect 11020 28950 11036 28966
rect 11052 28950 11068 28966
rect 11084 28950 11100 28966
rect 11116 28950 11132 28966
rect 11148 28950 11164 28966
rect 11180 28950 11196 28966
rect 11212 28950 11228 28966
rect 11244 28950 11260 28966
rect 11276 28950 11292 28966
rect 11308 28950 11324 28966
rect 11340 28950 11356 28966
rect 11372 28950 11388 28966
rect 11404 28950 11420 28966
rect 11436 28950 11452 28966
rect 11468 28950 11484 28966
rect 11500 28950 11516 28966
rect 11532 28950 11548 28966
rect 11564 28950 11580 28966
rect 11596 28950 11612 28966
rect 11628 28950 11644 28966
rect 11660 28950 11676 28966
rect 11692 28950 11708 28966
rect 11724 28950 11739 28966
rect 10061 28934 11739 28950
rect 10061 28918 10076 28934
rect 10092 28918 10108 28934
rect 10124 28918 10140 28934
rect 10156 28918 10172 28934
rect 10188 28918 10204 28934
rect 10220 28918 10236 28934
rect 10252 28918 10268 28934
rect 10284 28918 10300 28934
rect 10316 28918 10332 28934
rect 10348 28918 10364 28934
rect 10380 28918 10396 28934
rect 10412 28918 10428 28934
rect 10444 28918 10460 28934
rect 10476 28918 10492 28934
rect 10508 28918 10524 28934
rect 10540 28918 10556 28934
rect 10572 28918 10588 28934
rect 10604 28918 10620 28934
rect 10636 28918 10652 28934
rect 10668 28918 10684 28934
rect 10700 28918 10716 28934
rect 10732 28918 10748 28934
rect 10764 28918 10780 28934
rect 10796 28918 10812 28934
rect 10828 28918 10844 28934
rect 10860 28918 10876 28934
rect 10892 28918 10908 28934
rect 10924 28918 10940 28934
rect 10956 28918 10972 28934
rect 10988 28918 11004 28934
rect 11020 28918 11036 28934
rect 11052 28918 11068 28934
rect 11084 28918 11100 28934
rect 11116 28918 11132 28934
rect 11148 28918 11164 28934
rect 11180 28918 11196 28934
rect 11212 28918 11228 28934
rect 11244 28918 11260 28934
rect 11276 28918 11292 28934
rect 11308 28918 11324 28934
rect 11340 28918 11356 28934
rect 11372 28918 11388 28934
rect 11404 28918 11420 28934
rect 11436 28918 11452 28934
rect 11468 28918 11484 28934
rect 11500 28918 11516 28934
rect 11532 28918 11548 28934
rect 11564 28918 11580 28934
rect 11596 28918 11612 28934
rect 11628 28918 11644 28934
rect 11660 28918 11676 28934
rect 11692 28918 11708 28934
rect 11724 28918 11739 28934
rect 10061 28902 11739 28918
rect 10061 28886 10076 28902
rect 10092 28886 10108 28902
rect 10124 28886 10140 28902
rect 10156 28886 10172 28902
rect 10188 28886 10204 28902
rect 10220 28886 10236 28902
rect 10252 28886 10268 28902
rect 10284 28886 10300 28902
rect 10316 28886 10332 28902
rect 10348 28886 10364 28902
rect 10380 28886 10396 28902
rect 10412 28886 10428 28902
rect 10444 28886 10460 28902
rect 10476 28886 10492 28902
rect 10508 28886 10524 28902
rect 10540 28886 10556 28902
rect 10572 28886 10588 28902
rect 10604 28886 10620 28902
rect 10636 28886 10652 28902
rect 10668 28886 10684 28902
rect 10700 28886 10716 28902
rect 10732 28886 10748 28902
rect 10764 28886 10780 28902
rect 10796 28886 10812 28902
rect 10828 28886 10844 28902
rect 10860 28886 10876 28902
rect 10892 28886 10908 28902
rect 10924 28886 10940 28902
rect 10956 28886 10972 28902
rect 10988 28886 11004 28902
rect 11020 28886 11036 28902
rect 11052 28886 11068 28902
rect 11084 28886 11100 28902
rect 11116 28886 11132 28902
rect 11148 28886 11164 28902
rect 11180 28886 11196 28902
rect 11212 28886 11228 28902
rect 11244 28886 11260 28902
rect 11276 28886 11292 28902
rect 11308 28886 11324 28902
rect 11340 28886 11356 28902
rect 11372 28886 11388 28902
rect 11404 28886 11420 28902
rect 11436 28886 11452 28902
rect 11468 28886 11484 28902
rect 11500 28886 11516 28902
rect 11532 28886 11548 28902
rect 11564 28886 11580 28902
rect 11596 28886 11612 28902
rect 11628 28886 11644 28902
rect 11660 28886 11676 28902
rect 11692 28886 11708 28902
rect 11724 28886 11739 28902
rect 10061 28870 11739 28886
rect 10061 28854 10076 28870
rect 10092 28854 10108 28870
rect 10124 28854 10140 28870
rect 10156 28854 10172 28870
rect 10188 28854 10204 28870
rect 10220 28854 10236 28870
rect 10252 28854 10268 28870
rect 10284 28854 10300 28870
rect 10316 28854 10332 28870
rect 10348 28854 10364 28870
rect 10380 28854 10396 28870
rect 10412 28854 10428 28870
rect 10444 28854 10460 28870
rect 10476 28854 10492 28870
rect 10508 28854 10524 28870
rect 10540 28854 10556 28870
rect 10572 28854 10588 28870
rect 10604 28854 10620 28870
rect 10636 28854 10652 28870
rect 10668 28854 10684 28870
rect 10700 28854 10716 28870
rect 10732 28854 10748 28870
rect 10764 28854 10780 28870
rect 10796 28854 10812 28870
rect 10828 28854 10844 28870
rect 10860 28854 10876 28870
rect 10892 28854 10908 28870
rect 10924 28854 10940 28870
rect 10956 28854 10972 28870
rect 10988 28854 11004 28870
rect 11020 28854 11036 28870
rect 11052 28854 11068 28870
rect 11084 28854 11100 28870
rect 11116 28854 11132 28870
rect 11148 28854 11164 28870
rect 11180 28854 11196 28870
rect 11212 28854 11228 28870
rect 11244 28854 11260 28870
rect 11276 28854 11292 28870
rect 11308 28854 11324 28870
rect 11340 28854 11356 28870
rect 11372 28854 11388 28870
rect 11404 28854 11420 28870
rect 11436 28854 11452 28870
rect 11468 28854 11484 28870
rect 11500 28854 11516 28870
rect 11532 28854 11548 28870
rect 11564 28854 11580 28870
rect 11596 28854 11612 28870
rect 11628 28854 11644 28870
rect 11660 28854 11676 28870
rect 11692 28854 11708 28870
rect 11724 28854 11739 28870
rect 10061 28838 11739 28854
rect 10061 28822 10076 28838
rect 10092 28822 10108 28838
rect 10124 28822 10140 28838
rect 10156 28822 10172 28838
rect 10188 28822 10204 28838
rect 10220 28822 10236 28838
rect 10252 28822 10268 28838
rect 10284 28822 10300 28838
rect 10316 28822 10332 28838
rect 10348 28822 10364 28838
rect 10380 28822 10396 28838
rect 10412 28822 10428 28838
rect 10444 28822 10460 28838
rect 10476 28822 10492 28838
rect 10508 28822 10524 28838
rect 10540 28822 10556 28838
rect 10572 28822 10588 28838
rect 10604 28822 10620 28838
rect 10636 28822 10652 28838
rect 10668 28822 10684 28838
rect 10700 28822 10716 28838
rect 10732 28822 10748 28838
rect 10764 28822 10780 28838
rect 10796 28822 10812 28838
rect 10828 28822 10844 28838
rect 10860 28822 10876 28838
rect 10892 28822 10908 28838
rect 10924 28822 10940 28838
rect 10956 28822 10972 28838
rect 10988 28822 11004 28838
rect 11020 28822 11036 28838
rect 11052 28822 11068 28838
rect 11084 28822 11100 28838
rect 11116 28822 11132 28838
rect 11148 28822 11164 28838
rect 11180 28822 11196 28838
rect 11212 28822 11228 28838
rect 11244 28822 11260 28838
rect 11276 28822 11292 28838
rect 11308 28822 11324 28838
rect 11340 28822 11356 28838
rect 11372 28822 11388 28838
rect 11404 28822 11420 28838
rect 11436 28822 11452 28838
rect 11468 28822 11484 28838
rect 11500 28822 11516 28838
rect 11532 28822 11548 28838
rect 11564 28822 11580 28838
rect 11596 28822 11612 28838
rect 11628 28822 11644 28838
rect 11660 28822 11676 28838
rect 11692 28822 11708 28838
rect 11724 28822 11739 28838
rect 10061 28806 11739 28822
rect 10061 28790 10076 28806
rect 10092 28790 10108 28806
rect 10124 28790 10140 28806
rect 10156 28790 10172 28806
rect 10188 28790 10204 28806
rect 10220 28790 10236 28806
rect 10252 28790 10268 28806
rect 10284 28790 10300 28806
rect 10316 28790 10332 28806
rect 10348 28790 10364 28806
rect 10380 28790 10396 28806
rect 10412 28790 10428 28806
rect 10444 28790 10460 28806
rect 10476 28790 10492 28806
rect 10508 28790 10524 28806
rect 10540 28790 10556 28806
rect 10572 28790 10588 28806
rect 10604 28790 10620 28806
rect 10636 28790 10652 28806
rect 10668 28790 10684 28806
rect 10700 28790 10716 28806
rect 10732 28790 10748 28806
rect 10764 28790 10780 28806
rect 10796 28790 10812 28806
rect 10828 28790 10844 28806
rect 10860 28790 10876 28806
rect 10892 28790 10908 28806
rect 10924 28790 10940 28806
rect 10956 28790 10972 28806
rect 10988 28790 11004 28806
rect 11020 28790 11036 28806
rect 11052 28790 11068 28806
rect 11084 28790 11100 28806
rect 11116 28790 11132 28806
rect 11148 28790 11164 28806
rect 11180 28790 11196 28806
rect 11212 28790 11228 28806
rect 11244 28790 11260 28806
rect 11276 28790 11292 28806
rect 11308 28790 11324 28806
rect 11340 28790 11356 28806
rect 11372 28790 11388 28806
rect 11404 28790 11420 28806
rect 11436 28790 11452 28806
rect 11468 28790 11484 28806
rect 11500 28790 11516 28806
rect 11532 28790 11548 28806
rect 11564 28790 11580 28806
rect 11596 28790 11612 28806
rect 11628 28790 11644 28806
rect 11660 28790 11676 28806
rect 11692 28790 11708 28806
rect 11724 28790 11739 28806
rect 10061 28774 11739 28790
rect 10061 28758 10076 28774
rect 10092 28758 10108 28774
rect 10124 28758 10140 28774
rect 10156 28758 10172 28774
rect 10188 28758 10204 28774
rect 10220 28758 10236 28774
rect 10252 28758 10268 28774
rect 10284 28758 10300 28774
rect 10316 28758 10332 28774
rect 10348 28758 10364 28774
rect 10380 28758 10396 28774
rect 10412 28758 10428 28774
rect 10444 28758 10460 28774
rect 10476 28758 10492 28774
rect 10508 28758 10524 28774
rect 10540 28758 10556 28774
rect 10572 28758 10588 28774
rect 10604 28758 10620 28774
rect 10636 28758 10652 28774
rect 10668 28758 10684 28774
rect 10700 28758 10716 28774
rect 10732 28758 10748 28774
rect 10764 28758 10780 28774
rect 10796 28758 10812 28774
rect 10828 28758 10844 28774
rect 10860 28758 10876 28774
rect 10892 28758 10908 28774
rect 10924 28758 10940 28774
rect 10956 28758 10972 28774
rect 10988 28758 11004 28774
rect 11020 28758 11036 28774
rect 11052 28758 11068 28774
rect 11084 28758 11100 28774
rect 11116 28758 11132 28774
rect 11148 28758 11164 28774
rect 11180 28758 11196 28774
rect 11212 28758 11228 28774
rect 11244 28758 11260 28774
rect 11276 28758 11292 28774
rect 11308 28758 11324 28774
rect 11340 28758 11356 28774
rect 11372 28758 11388 28774
rect 11404 28758 11420 28774
rect 11436 28758 11452 28774
rect 11468 28758 11484 28774
rect 11500 28758 11516 28774
rect 11532 28758 11548 28774
rect 11564 28758 11580 28774
rect 11596 28758 11612 28774
rect 11628 28758 11644 28774
rect 11660 28758 11676 28774
rect 11692 28758 11708 28774
rect 11724 28758 11739 28774
rect 10061 28742 11739 28758
rect 10061 28726 10076 28742
rect 10092 28726 10108 28742
rect 10124 28726 10140 28742
rect 10156 28726 10172 28742
rect 10188 28726 10204 28742
rect 10220 28726 10236 28742
rect 10252 28726 10268 28742
rect 10284 28726 10300 28742
rect 10316 28726 10332 28742
rect 10348 28726 10364 28742
rect 10380 28726 10396 28742
rect 10412 28726 10428 28742
rect 10444 28726 10460 28742
rect 10476 28726 10492 28742
rect 10508 28726 10524 28742
rect 10540 28726 10556 28742
rect 10572 28726 10588 28742
rect 10604 28726 10620 28742
rect 10636 28726 10652 28742
rect 10668 28726 10684 28742
rect 10700 28726 10716 28742
rect 10732 28726 10748 28742
rect 10764 28726 10780 28742
rect 10796 28726 10812 28742
rect 10828 28726 10844 28742
rect 10860 28726 10876 28742
rect 10892 28726 10908 28742
rect 10924 28726 10940 28742
rect 10956 28726 10972 28742
rect 10988 28726 11004 28742
rect 11020 28726 11036 28742
rect 11052 28726 11068 28742
rect 11084 28726 11100 28742
rect 11116 28726 11132 28742
rect 11148 28726 11164 28742
rect 11180 28726 11196 28742
rect 11212 28726 11228 28742
rect 11244 28726 11260 28742
rect 11276 28726 11292 28742
rect 11308 28726 11324 28742
rect 11340 28726 11356 28742
rect 11372 28726 11388 28742
rect 11404 28726 11420 28742
rect 11436 28726 11452 28742
rect 11468 28726 11484 28742
rect 11500 28726 11516 28742
rect 11532 28726 11548 28742
rect 11564 28726 11580 28742
rect 11596 28726 11612 28742
rect 11628 28726 11644 28742
rect 11660 28726 11676 28742
rect 11692 28726 11708 28742
rect 11724 28726 11739 28742
rect 10061 28710 11739 28726
rect 10061 28694 10076 28710
rect 10092 28694 10108 28710
rect 10124 28694 10140 28710
rect 10156 28694 10172 28710
rect 10188 28694 10204 28710
rect 10220 28694 10236 28710
rect 10252 28694 10268 28710
rect 10284 28694 10300 28710
rect 10316 28694 10332 28710
rect 10348 28694 10364 28710
rect 10380 28694 10396 28710
rect 10412 28694 10428 28710
rect 10444 28694 10460 28710
rect 10476 28694 10492 28710
rect 10508 28694 10524 28710
rect 10540 28694 10556 28710
rect 10572 28694 10588 28710
rect 10604 28694 10620 28710
rect 10636 28694 10652 28710
rect 10668 28694 10684 28710
rect 10700 28694 10716 28710
rect 10732 28694 10748 28710
rect 10764 28694 10780 28710
rect 10796 28694 10812 28710
rect 10828 28694 10844 28710
rect 10860 28694 10876 28710
rect 10892 28694 10908 28710
rect 10924 28694 10940 28710
rect 10956 28694 10972 28710
rect 10988 28694 11004 28710
rect 11020 28694 11036 28710
rect 11052 28694 11068 28710
rect 11084 28694 11100 28710
rect 11116 28694 11132 28710
rect 11148 28694 11164 28710
rect 11180 28694 11196 28710
rect 11212 28694 11228 28710
rect 11244 28694 11260 28710
rect 11276 28694 11292 28710
rect 11308 28694 11324 28710
rect 11340 28694 11356 28710
rect 11372 28694 11388 28710
rect 11404 28694 11420 28710
rect 11436 28694 11452 28710
rect 11468 28694 11484 28710
rect 11500 28694 11516 28710
rect 11532 28694 11548 28710
rect 11564 28694 11580 28710
rect 11596 28694 11612 28710
rect 11628 28694 11644 28710
rect 11660 28694 11676 28710
rect 11692 28694 11708 28710
rect 11724 28694 11739 28710
rect 10061 28681 11739 28694
rect 12480 28080 12580 29180
rect 15180 28460 15280 29180
rect 17880 28500 17980 29180
rect 17881 28474 17979 28500
rect 15181 28446 15279 28460
rect 15181 28430 15206 28446
rect 15222 28430 15238 28446
rect 15254 28430 15279 28446
rect 15181 28414 15279 28430
rect 15181 28398 15206 28414
rect 15222 28398 15238 28414
rect 15254 28398 15279 28414
rect 17881 28458 17906 28474
rect 17922 28458 17938 28474
rect 17954 28458 17979 28474
rect 17881 28442 17979 28458
rect 17881 28426 17906 28442
rect 17922 28426 17938 28442
rect 17954 28426 17979 28442
rect 17881 28401 17979 28426
rect 15181 28382 15279 28398
rect 15181 28366 15206 28382
rect 15222 28366 15238 28382
rect 15254 28366 15279 28382
rect 15181 28350 15279 28366
rect 15181 28334 15206 28350
rect 15222 28334 15238 28350
rect 15254 28334 15279 28350
rect 15181 28318 15279 28334
rect 15181 28302 15206 28318
rect 15222 28302 15238 28318
rect 15254 28302 15279 28318
rect 15181 28286 15279 28302
rect 15181 28270 15206 28286
rect 15222 28270 15238 28286
rect 15254 28270 15279 28286
rect 15181 28254 15279 28270
rect 15181 28238 15206 28254
rect 15222 28238 15238 28254
rect 15254 28238 15279 28254
rect 15181 28222 15279 28238
rect 15181 28206 15206 28222
rect 15222 28206 15238 28222
rect 15254 28206 15279 28222
rect 15181 28190 15279 28206
rect 15181 28174 15206 28190
rect 15222 28174 15238 28190
rect 15254 28174 15279 28190
rect 20580 28280 20680 29180
rect 26341 28474 26439 28499
rect 26341 28458 26366 28474
rect 26382 28458 26398 28474
rect 26414 28458 26439 28474
rect 26341 28442 26439 28458
rect 26341 28426 26366 28442
rect 26382 28426 26398 28442
rect 26414 28426 26439 28442
rect 26341 28400 26439 28426
rect 20580 28180 25360 28280
rect 15181 28161 15279 28174
rect 12480 27980 23517 28080
rect 25260 28000 25360 28180
rect 26340 28000 26440 28400
rect 8800 27679 9080 27680
rect 8800 27668 9659 27679
rect 8800 27652 9106 27668
rect 9122 27652 9138 27668
rect 9154 27652 9170 27668
rect 9186 27652 9202 27668
rect 9218 27652 9234 27668
rect 9250 27652 9266 27668
rect 9282 27652 9298 27668
rect 9314 27652 9330 27668
rect 9346 27652 9362 27668
rect 9378 27652 9394 27668
rect 9410 27652 9426 27668
rect 9442 27652 9458 27668
rect 9474 27652 9490 27668
rect 9506 27652 9522 27668
rect 9538 27652 9554 27668
rect 9570 27652 9586 27668
rect 9602 27652 9618 27668
rect 9634 27652 9659 27668
rect 8800 27636 9659 27652
rect 8800 27620 9106 27636
rect 9122 27620 9138 27636
rect 9154 27620 9170 27636
rect 9186 27620 9202 27636
rect 9218 27620 9234 27636
rect 9250 27620 9266 27636
rect 9282 27620 9298 27636
rect 9314 27620 9330 27636
rect 9346 27620 9362 27636
rect 9378 27620 9394 27636
rect 9410 27620 9426 27636
rect 9442 27620 9458 27636
rect 9474 27620 9490 27636
rect 9506 27620 9522 27636
rect 9538 27620 9554 27636
rect 9570 27620 9586 27636
rect 9602 27620 9618 27636
rect 9634 27620 9659 27636
rect 8800 27604 9659 27620
rect 8800 27588 9106 27604
rect 9122 27588 9138 27604
rect 9154 27588 9170 27604
rect 9186 27588 9202 27604
rect 9218 27588 9234 27604
rect 9250 27588 9266 27604
rect 9282 27588 9298 27604
rect 9314 27588 9330 27604
rect 9346 27588 9362 27604
rect 9378 27588 9394 27604
rect 9410 27588 9426 27604
rect 9442 27588 9458 27604
rect 9474 27588 9490 27604
rect 9506 27588 9522 27604
rect 9538 27588 9554 27604
rect 9570 27588 9586 27604
rect 9602 27588 9618 27604
rect 9634 27588 9659 27604
rect 8800 27572 9659 27588
rect 8800 27556 9106 27572
rect 9122 27556 9138 27572
rect 9154 27556 9170 27572
rect 9186 27556 9202 27572
rect 9218 27556 9234 27572
rect 9250 27556 9266 27572
rect 9282 27556 9298 27572
rect 9314 27556 9330 27572
rect 9346 27556 9362 27572
rect 9378 27556 9394 27572
rect 9410 27556 9426 27572
rect 9442 27556 9458 27572
rect 9474 27556 9490 27572
rect 9506 27556 9522 27572
rect 9538 27556 9554 27572
rect 9570 27556 9586 27572
rect 9602 27556 9618 27572
rect 9634 27556 9659 27572
rect 8800 27540 9659 27556
rect 8800 27524 9106 27540
rect 9122 27524 9138 27540
rect 9154 27524 9170 27540
rect 9186 27524 9202 27540
rect 9218 27524 9234 27540
rect 9250 27524 9266 27540
rect 9282 27524 9298 27540
rect 9314 27524 9330 27540
rect 9346 27524 9362 27540
rect 9378 27524 9394 27540
rect 9410 27524 9426 27540
rect 9442 27524 9458 27540
rect 9474 27524 9490 27540
rect 9506 27524 9522 27540
rect 9538 27524 9554 27540
rect 9570 27524 9586 27540
rect 9602 27524 9618 27540
rect 9634 27524 9659 27540
rect 8800 27508 9659 27524
rect 8800 27492 9106 27508
rect 9122 27492 9138 27508
rect 9154 27492 9170 27508
rect 9186 27492 9202 27508
rect 9218 27492 9234 27508
rect 9250 27492 9266 27508
rect 9282 27492 9298 27508
rect 9314 27492 9330 27508
rect 9346 27492 9362 27508
rect 9378 27492 9394 27508
rect 9410 27492 9426 27508
rect 9442 27492 9458 27508
rect 9474 27492 9490 27508
rect 9506 27492 9522 27508
rect 9538 27492 9554 27508
rect 9570 27492 9586 27508
rect 9602 27492 9618 27508
rect 9634 27492 9659 27508
rect 8800 27476 9659 27492
rect 8800 27460 9106 27476
rect 9122 27460 9138 27476
rect 9154 27460 9170 27476
rect 9186 27460 9202 27476
rect 9218 27460 9234 27476
rect 9250 27460 9266 27476
rect 9282 27460 9298 27476
rect 9314 27460 9330 27476
rect 9346 27460 9362 27476
rect 9378 27460 9394 27476
rect 9410 27460 9426 27476
rect 9442 27460 9458 27476
rect 9474 27460 9490 27476
rect 9506 27460 9522 27476
rect 9538 27460 9554 27476
rect 9570 27460 9586 27476
rect 9602 27460 9618 27476
rect 9634 27460 9659 27476
rect 8800 27444 9659 27460
rect 8800 27428 9106 27444
rect 9122 27428 9138 27444
rect 9154 27428 9170 27444
rect 9186 27428 9202 27444
rect 9218 27428 9234 27444
rect 9250 27428 9266 27444
rect 9282 27428 9298 27444
rect 9314 27428 9330 27444
rect 9346 27428 9362 27444
rect 9378 27428 9394 27444
rect 9410 27428 9426 27444
rect 9442 27428 9458 27444
rect 9474 27428 9490 27444
rect 9506 27428 9522 27444
rect 9538 27428 9554 27444
rect 9570 27428 9586 27444
rect 9602 27428 9618 27444
rect 9634 27428 9659 27444
rect 8800 27412 9659 27428
rect 8800 27396 9106 27412
rect 9122 27396 9138 27412
rect 9154 27396 9170 27412
rect 9186 27396 9202 27412
rect 9218 27396 9234 27412
rect 9250 27396 9266 27412
rect 9282 27396 9298 27412
rect 9314 27396 9330 27412
rect 9346 27396 9362 27412
rect 9378 27396 9394 27412
rect 9410 27396 9426 27412
rect 9442 27396 9458 27412
rect 9474 27396 9490 27412
rect 9506 27396 9522 27412
rect 9538 27396 9554 27412
rect 9570 27396 9586 27412
rect 9602 27396 9618 27412
rect 9634 27396 9659 27412
rect 8800 27380 9659 27396
rect 8800 27364 9106 27380
rect 9122 27364 9138 27380
rect 9154 27364 9170 27380
rect 9186 27364 9202 27380
rect 9218 27364 9234 27380
rect 9250 27364 9266 27380
rect 9282 27364 9298 27380
rect 9314 27364 9330 27380
rect 9346 27364 9362 27380
rect 9378 27364 9394 27380
rect 9410 27364 9426 27380
rect 9442 27364 9458 27380
rect 9474 27364 9490 27380
rect 9506 27364 9522 27380
rect 9538 27364 9554 27380
rect 9570 27364 9586 27380
rect 9602 27364 9618 27380
rect 9634 27364 9659 27380
rect 8800 27348 9659 27364
rect 8800 27332 9106 27348
rect 9122 27332 9138 27348
rect 9154 27332 9170 27348
rect 9186 27332 9202 27348
rect 9218 27332 9234 27348
rect 9250 27332 9266 27348
rect 9282 27332 9298 27348
rect 9314 27332 9330 27348
rect 9346 27332 9362 27348
rect 9378 27332 9394 27348
rect 9410 27332 9426 27348
rect 9442 27332 9458 27348
rect 9474 27332 9490 27348
rect 9506 27332 9522 27348
rect 9538 27332 9554 27348
rect 9570 27332 9586 27348
rect 9602 27332 9618 27348
rect 9634 27332 9659 27348
rect 8800 27316 9659 27332
rect 8800 27300 9106 27316
rect 9122 27300 9138 27316
rect 9154 27300 9170 27316
rect 9186 27300 9202 27316
rect 9218 27300 9234 27316
rect 9250 27300 9266 27316
rect 9282 27300 9298 27316
rect 9314 27300 9330 27316
rect 9346 27300 9362 27316
rect 9378 27300 9394 27316
rect 9410 27300 9426 27316
rect 9442 27300 9458 27316
rect 9474 27300 9490 27316
rect 9506 27300 9522 27316
rect 9538 27300 9554 27316
rect 9570 27300 9586 27316
rect 9602 27300 9618 27316
rect 9634 27300 9659 27316
rect 8800 27284 9659 27300
rect 8800 27268 9106 27284
rect 9122 27268 9138 27284
rect 9154 27268 9170 27284
rect 9186 27268 9202 27284
rect 9218 27268 9234 27284
rect 9250 27268 9266 27284
rect 9282 27268 9298 27284
rect 9314 27268 9330 27284
rect 9346 27268 9362 27284
rect 9378 27268 9394 27284
rect 9410 27268 9426 27284
rect 9442 27268 9458 27284
rect 9474 27268 9490 27284
rect 9506 27268 9522 27284
rect 9538 27268 9554 27284
rect 9570 27268 9586 27284
rect 9602 27268 9618 27284
rect 9634 27268 9659 27284
rect 8800 27252 9659 27268
rect 8800 27236 9106 27252
rect 9122 27236 9138 27252
rect 9154 27236 9170 27252
rect 9186 27236 9202 27252
rect 9218 27236 9234 27252
rect 9250 27236 9266 27252
rect 9282 27236 9298 27252
rect 9314 27236 9330 27252
rect 9346 27236 9362 27252
rect 9378 27236 9394 27252
rect 9410 27236 9426 27252
rect 9442 27236 9458 27252
rect 9474 27236 9490 27252
rect 9506 27236 9522 27252
rect 9538 27236 9554 27252
rect 9570 27236 9586 27252
rect 9602 27236 9618 27252
rect 9634 27236 9659 27252
rect 8800 27220 9659 27236
rect 8800 27204 9106 27220
rect 9122 27204 9138 27220
rect 9154 27204 9170 27220
rect 9186 27204 9202 27220
rect 9218 27204 9234 27220
rect 9250 27204 9266 27220
rect 9282 27204 9298 27220
rect 9314 27204 9330 27220
rect 9346 27204 9362 27220
rect 9378 27204 9394 27220
rect 9410 27204 9426 27220
rect 9442 27204 9458 27220
rect 9474 27204 9490 27220
rect 9506 27204 9522 27220
rect 9538 27204 9554 27220
rect 9570 27204 9586 27220
rect 9602 27204 9618 27220
rect 9634 27204 9659 27220
rect 8800 27188 9659 27204
rect 8800 27172 9106 27188
rect 9122 27172 9138 27188
rect 9154 27172 9170 27188
rect 9186 27172 9202 27188
rect 9218 27172 9234 27188
rect 9250 27172 9266 27188
rect 9282 27172 9298 27188
rect 9314 27172 9330 27188
rect 9346 27172 9362 27188
rect 9378 27172 9394 27188
rect 9410 27172 9426 27188
rect 9442 27172 9458 27188
rect 9474 27172 9490 27188
rect 9506 27172 9522 27188
rect 9538 27172 9554 27188
rect 9570 27172 9586 27188
rect 9602 27172 9618 27188
rect 9634 27172 9659 27188
rect 8800 27156 9659 27172
rect 8800 27140 9106 27156
rect 9122 27140 9138 27156
rect 9154 27140 9170 27156
rect 9186 27140 9202 27156
rect 9218 27140 9234 27156
rect 9250 27140 9266 27156
rect 9282 27140 9298 27156
rect 9314 27140 9330 27156
rect 9346 27140 9362 27156
rect 9378 27140 9394 27156
rect 9410 27140 9426 27156
rect 9442 27140 9458 27156
rect 9474 27140 9490 27156
rect 9506 27140 9522 27156
rect 9538 27140 9554 27156
rect 9570 27140 9586 27156
rect 9602 27140 9618 27156
rect 9634 27140 9659 27156
rect 8800 27124 9659 27140
rect 8800 27108 9106 27124
rect 9122 27108 9138 27124
rect 9154 27108 9170 27124
rect 9186 27108 9202 27124
rect 9218 27108 9234 27124
rect 9250 27108 9266 27124
rect 9282 27108 9298 27124
rect 9314 27108 9330 27124
rect 9346 27108 9362 27124
rect 9378 27108 9394 27124
rect 9410 27108 9426 27124
rect 9442 27108 9458 27124
rect 9474 27108 9490 27124
rect 9506 27108 9522 27124
rect 9538 27108 9554 27124
rect 9570 27108 9586 27124
rect 9602 27108 9618 27124
rect 9634 27108 9659 27124
rect 8800 27092 9659 27108
rect 8800 27076 9106 27092
rect 9122 27076 9138 27092
rect 9154 27076 9170 27092
rect 9186 27076 9202 27092
rect 9218 27076 9234 27092
rect 9250 27076 9266 27092
rect 9282 27076 9298 27092
rect 9314 27076 9330 27092
rect 9346 27076 9362 27092
rect 9378 27076 9394 27092
rect 9410 27076 9426 27092
rect 9442 27076 9458 27092
rect 9474 27076 9490 27092
rect 9506 27076 9522 27092
rect 9538 27076 9554 27092
rect 9570 27076 9586 27092
rect 9602 27076 9618 27092
rect 9634 27076 9659 27092
rect 8800 27060 9659 27076
rect 8800 27044 9106 27060
rect 9122 27044 9138 27060
rect 9154 27044 9170 27060
rect 9186 27044 9202 27060
rect 9218 27044 9234 27060
rect 9250 27044 9266 27060
rect 9282 27044 9298 27060
rect 9314 27044 9330 27060
rect 9346 27044 9362 27060
rect 9378 27044 9394 27060
rect 9410 27044 9426 27060
rect 9442 27044 9458 27060
rect 9474 27044 9490 27060
rect 9506 27044 9522 27060
rect 9538 27044 9554 27060
rect 9570 27044 9586 27060
rect 9602 27044 9618 27060
rect 9634 27044 9659 27060
rect 8800 27028 9659 27044
rect 8800 27012 9106 27028
rect 9122 27012 9138 27028
rect 9154 27012 9170 27028
rect 9186 27012 9202 27028
rect 9218 27012 9234 27028
rect 9250 27012 9266 27028
rect 9282 27012 9298 27028
rect 9314 27012 9330 27028
rect 9346 27012 9362 27028
rect 9378 27012 9394 27028
rect 9410 27012 9426 27028
rect 9442 27012 9458 27028
rect 9474 27012 9490 27028
rect 9506 27012 9522 27028
rect 9538 27012 9554 27028
rect 9570 27012 9586 27028
rect 9602 27012 9618 27028
rect 9634 27012 9659 27028
rect 8800 26996 9659 27012
rect 8800 26980 9106 26996
rect 9122 26980 9138 26996
rect 9154 26980 9170 26996
rect 9186 26980 9202 26996
rect 9218 26980 9234 26996
rect 9250 26980 9266 26996
rect 9282 26980 9298 26996
rect 9314 26980 9330 26996
rect 9346 26980 9362 26996
rect 9378 26980 9394 26996
rect 9410 26980 9426 26996
rect 9442 26980 9458 26996
rect 9474 26980 9490 26996
rect 9506 26980 9522 26996
rect 9538 26980 9554 26996
rect 9570 26980 9586 26996
rect 9602 26980 9618 26996
rect 9634 26980 9659 26996
rect 8800 26964 9659 26980
rect 8800 26948 9106 26964
rect 9122 26948 9138 26964
rect 9154 26948 9170 26964
rect 9186 26948 9202 26964
rect 9218 26948 9234 26964
rect 9250 26948 9266 26964
rect 9282 26948 9298 26964
rect 9314 26948 9330 26964
rect 9346 26948 9362 26964
rect 9378 26948 9394 26964
rect 9410 26948 9426 26964
rect 9442 26948 9458 26964
rect 9474 26948 9490 26964
rect 9506 26948 9522 26964
rect 9538 26948 9554 26964
rect 9570 26948 9586 26964
rect 9602 26948 9618 26964
rect 9634 26948 9659 26964
rect 8800 26932 9659 26948
rect 8800 26916 9106 26932
rect 9122 26916 9138 26932
rect 9154 26916 9170 26932
rect 9186 26916 9202 26932
rect 9218 26916 9234 26932
rect 9250 26916 9266 26932
rect 9282 26916 9298 26932
rect 9314 26916 9330 26932
rect 9346 26916 9362 26932
rect 9378 26916 9394 26932
rect 9410 26916 9426 26932
rect 9442 26916 9458 26932
rect 9474 26916 9490 26932
rect 9506 26916 9522 26932
rect 9538 26916 9554 26932
rect 9570 26916 9586 26932
rect 9602 26916 9618 26932
rect 9634 26916 9659 26932
rect 8800 26900 9659 26916
rect 8800 26884 9106 26900
rect 9122 26884 9138 26900
rect 9154 26884 9170 26900
rect 9186 26884 9202 26900
rect 9218 26884 9234 26900
rect 9250 26884 9266 26900
rect 9282 26884 9298 26900
rect 9314 26884 9330 26900
rect 9346 26884 9362 26900
rect 9378 26884 9394 26900
rect 9410 26884 9426 26900
rect 9442 26884 9458 26900
rect 9474 26884 9490 26900
rect 9506 26884 9522 26900
rect 9538 26884 9554 26900
rect 9570 26884 9586 26900
rect 9602 26884 9618 26900
rect 9634 26884 9659 26900
rect 8800 26868 9659 26884
rect 8800 26852 9106 26868
rect 9122 26852 9138 26868
rect 9154 26852 9170 26868
rect 9186 26852 9202 26868
rect 9218 26852 9234 26868
rect 9250 26852 9266 26868
rect 9282 26852 9298 26868
rect 9314 26852 9330 26868
rect 9346 26852 9362 26868
rect 9378 26852 9394 26868
rect 9410 26852 9426 26868
rect 9442 26852 9458 26868
rect 9474 26852 9490 26868
rect 9506 26852 9522 26868
rect 9538 26852 9554 26868
rect 9570 26852 9586 26868
rect 9602 26852 9618 26868
rect 9634 26852 9659 26868
rect 8800 26836 9659 26852
rect 8800 26820 9106 26836
rect 9122 26820 9138 26836
rect 9154 26820 9170 26836
rect 9186 26820 9202 26836
rect 9218 26820 9234 26836
rect 9250 26820 9266 26836
rect 9282 26820 9298 26836
rect 9314 26820 9330 26836
rect 9346 26820 9362 26836
rect 9378 26820 9394 26836
rect 9410 26820 9426 26836
rect 9442 26820 9458 26836
rect 9474 26820 9490 26836
rect 9506 26820 9522 26836
rect 9538 26820 9554 26836
rect 9570 26820 9586 26836
rect 9602 26820 9618 26836
rect 9634 26820 9659 26836
rect 8800 26804 9659 26820
rect 8800 26788 9106 26804
rect 9122 26788 9138 26804
rect 9154 26788 9170 26804
rect 9186 26788 9202 26804
rect 9218 26788 9234 26804
rect 9250 26788 9266 26804
rect 9282 26788 9298 26804
rect 9314 26788 9330 26804
rect 9346 26788 9362 26804
rect 9378 26788 9394 26804
rect 9410 26788 9426 26804
rect 9442 26788 9458 26804
rect 9474 26788 9490 26804
rect 9506 26788 9522 26804
rect 9538 26788 9554 26804
rect 9570 26788 9586 26804
rect 9602 26788 9618 26804
rect 9634 26788 9659 26804
rect 8800 26772 9659 26788
rect 8800 26756 9106 26772
rect 9122 26756 9138 26772
rect 9154 26756 9170 26772
rect 9186 26756 9202 26772
rect 9218 26756 9234 26772
rect 9250 26756 9266 26772
rect 9282 26756 9298 26772
rect 9314 26756 9330 26772
rect 9346 26756 9362 26772
rect 9378 26756 9394 26772
rect 9410 26756 9426 26772
rect 9442 26756 9458 26772
rect 9474 26756 9490 26772
rect 9506 26756 9522 26772
rect 9538 26756 9554 26772
rect 9570 26756 9586 26772
rect 9602 26756 9618 26772
rect 9634 26756 9659 26772
rect 8800 26740 9659 26756
rect 8800 26724 9106 26740
rect 9122 26724 9138 26740
rect 9154 26724 9170 26740
rect 9186 26724 9202 26740
rect 9218 26724 9234 26740
rect 9250 26724 9266 26740
rect 9282 26724 9298 26740
rect 9314 26724 9330 26740
rect 9346 26724 9362 26740
rect 9378 26724 9394 26740
rect 9410 26724 9426 26740
rect 9442 26724 9458 26740
rect 9474 26724 9490 26740
rect 9506 26724 9522 26740
rect 9538 26724 9554 26740
rect 9570 26724 9586 26740
rect 9602 26724 9618 26740
rect 9634 26724 9659 26740
rect 8800 26708 9659 26724
rect 8800 26692 9106 26708
rect 9122 26692 9138 26708
rect 9154 26692 9170 26708
rect 9186 26692 9202 26708
rect 9218 26692 9234 26708
rect 9250 26692 9266 26708
rect 9282 26692 9298 26708
rect 9314 26692 9330 26708
rect 9346 26692 9362 26708
rect 9378 26692 9394 26708
rect 9410 26692 9426 26708
rect 9442 26692 9458 26708
rect 9474 26692 9490 26708
rect 9506 26692 9522 26708
rect 9538 26692 9554 26708
rect 9570 26692 9586 26708
rect 9602 26692 9618 26708
rect 9634 26692 9659 26708
rect 8800 26676 9659 26692
rect 8800 26660 9106 26676
rect 9122 26660 9138 26676
rect 9154 26660 9170 26676
rect 9186 26660 9202 26676
rect 9218 26660 9234 26676
rect 9250 26660 9266 26676
rect 9282 26660 9298 26676
rect 9314 26660 9330 26676
rect 9346 26660 9362 26676
rect 9378 26660 9394 26676
rect 9410 26660 9426 26676
rect 9442 26660 9458 26676
rect 9474 26660 9490 26676
rect 9506 26660 9522 26676
rect 9538 26660 9554 26676
rect 9570 26660 9586 26676
rect 9602 26660 9618 26676
rect 9634 26660 9659 26676
rect 8800 26644 9659 26660
rect 8800 26628 9106 26644
rect 9122 26628 9138 26644
rect 9154 26628 9170 26644
rect 9186 26628 9202 26644
rect 9218 26628 9234 26644
rect 9250 26628 9266 26644
rect 9282 26628 9298 26644
rect 9314 26628 9330 26644
rect 9346 26628 9362 26644
rect 9378 26628 9394 26644
rect 9410 26628 9426 26644
rect 9442 26628 9458 26644
rect 9474 26628 9490 26644
rect 9506 26628 9522 26644
rect 9538 26628 9554 26644
rect 9570 26628 9586 26644
rect 9602 26628 9618 26644
rect 9634 26628 9659 26644
rect 8800 26612 9659 26628
rect 8800 26596 9106 26612
rect 9122 26596 9138 26612
rect 9154 26596 9170 26612
rect 9186 26596 9202 26612
rect 9218 26596 9234 26612
rect 9250 26596 9266 26612
rect 9282 26596 9298 26612
rect 9314 26596 9330 26612
rect 9346 26596 9362 26612
rect 9378 26596 9394 26612
rect 9410 26596 9426 26612
rect 9442 26596 9458 26612
rect 9474 26596 9490 26612
rect 9506 26596 9522 26612
rect 9538 26596 9554 26612
rect 9570 26596 9586 26612
rect 9602 26596 9618 26612
rect 9634 26596 9659 26612
rect 8800 26580 9659 26596
rect 8800 26564 9106 26580
rect 9122 26564 9138 26580
rect 9154 26564 9170 26580
rect 9186 26564 9202 26580
rect 9218 26564 9234 26580
rect 9250 26564 9266 26580
rect 9282 26564 9298 26580
rect 9314 26564 9330 26580
rect 9346 26564 9362 26580
rect 9378 26564 9394 26580
rect 9410 26564 9426 26580
rect 9442 26564 9458 26580
rect 9474 26564 9490 26580
rect 9506 26564 9522 26580
rect 9538 26564 9554 26580
rect 9570 26564 9586 26580
rect 9602 26564 9618 26580
rect 9634 26564 9659 26580
rect 8800 26548 9659 26564
rect 8800 26532 9106 26548
rect 9122 26532 9138 26548
rect 9154 26532 9170 26548
rect 9186 26532 9202 26548
rect 9218 26532 9234 26548
rect 9250 26532 9266 26548
rect 9282 26532 9298 26548
rect 9314 26532 9330 26548
rect 9346 26532 9362 26548
rect 9378 26532 9394 26548
rect 9410 26532 9426 26548
rect 9442 26532 9458 26548
rect 9474 26532 9490 26548
rect 9506 26532 9522 26548
rect 9538 26532 9554 26548
rect 9570 26532 9586 26548
rect 9602 26532 9618 26548
rect 9634 26532 9659 26548
rect 8800 26521 9659 26532
rect 8800 26520 9080 26521
rect 28840 26079 29180 26080
rect 28541 26054 29180 26079
rect 28541 26038 28554 26054
rect 28570 26038 28586 26054
rect 28602 26038 28618 26054
rect 28634 26038 28650 26054
rect 28666 26038 28682 26054
rect 28698 26038 28714 26054
rect 28730 26038 28746 26054
rect 28762 26038 28778 26054
rect 28794 26038 28810 26054
rect 28826 26038 29180 26054
rect 28541 26022 29180 26038
rect 28541 26006 28554 26022
rect 28570 26006 28586 26022
rect 28602 26006 28618 26022
rect 28634 26006 28650 26022
rect 28666 26006 28682 26022
rect 28698 26006 28714 26022
rect 28730 26006 28746 26022
rect 28762 26006 28778 26022
rect 28794 26006 28810 26022
rect 28826 26006 29180 26022
rect 28541 25981 29180 26006
rect 28840 25980 29180 25981
rect 28640 23379 29180 23380
rect 8820 23359 9020 23360
rect 8820 23346 9119 23359
rect 8820 23330 9046 23346
rect 9062 23330 9078 23346
rect 9094 23330 9119 23346
rect 8820 23314 9119 23330
rect 8820 23298 9046 23314
rect 9062 23298 9078 23314
rect 9094 23298 9119 23314
rect 8820 23282 9119 23298
rect 8820 23266 9046 23282
rect 9062 23266 9078 23282
rect 9094 23266 9119 23282
rect 28341 23354 29180 23379
rect 28341 23338 28354 23354
rect 28370 23338 28386 23354
rect 28402 23338 28418 23354
rect 28434 23338 28450 23354
rect 28466 23338 28482 23354
rect 28498 23338 28514 23354
rect 28530 23338 28546 23354
rect 28562 23338 28578 23354
rect 28594 23338 28610 23354
rect 28626 23338 29180 23354
rect 28341 23322 29180 23338
rect 28341 23306 28354 23322
rect 28370 23306 28386 23322
rect 28402 23306 28418 23322
rect 28434 23306 28450 23322
rect 28466 23306 28482 23322
rect 28498 23306 28514 23322
rect 28530 23306 28546 23322
rect 28562 23306 28578 23322
rect 28594 23306 28610 23322
rect 28626 23306 29180 23322
rect 28341 23281 29180 23306
rect 28640 23280 29180 23281
rect 8820 23260 9119 23266
rect 9019 23250 9119 23260
rect 9019 23234 9046 23250
rect 9062 23234 9078 23250
rect 9094 23234 9119 23250
rect 9019 23218 9119 23234
rect 9019 23202 9046 23218
rect 9062 23202 9078 23218
rect 9094 23202 9119 23218
rect 9019 23186 9119 23202
rect 9019 23170 9046 23186
rect 9062 23170 9078 23186
rect 9094 23170 9119 23186
rect 9019 23154 9119 23170
rect 9019 23138 9046 23154
rect 9062 23138 9078 23154
rect 9094 23138 9119 23154
rect 9019 23122 9119 23138
rect 9019 23106 9046 23122
rect 9062 23106 9078 23122
rect 9094 23106 9119 23122
rect 9019 23090 9119 23106
rect 9019 23074 9046 23090
rect 9062 23074 9078 23090
rect 9094 23074 9119 23090
rect 9019 23061 9119 23074
rect 9421 22686 9519 22699
rect 9421 22670 9446 22686
rect 9462 22670 9478 22686
rect 9494 22670 9519 22686
rect 9421 22654 9519 22670
rect 9421 22638 9446 22654
rect 9462 22638 9478 22654
rect 9494 22638 9519 22654
rect 9421 22622 9519 22638
rect 9421 22606 9446 22622
rect 9462 22606 9478 22622
rect 9494 22606 9519 22622
rect 9421 22590 9519 22606
rect 9421 22574 9446 22590
rect 9462 22574 9478 22590
rect 9494 22574 9519 22590
rect 9421 22558 9519 22574
rect 9421 22542 9446 22558
rect 9462 22542 9478 22558
rect 9494 22542 9519 22558
rect 9421 22526 9519 22542
rect 9421 22510 9446 22526
rect 9462 22510 9478 22526
rect 9494 22510 9519 22526
rect 9421 22494 9519 22510
rect 9421 22478 9446 22494
rect 9462 22478 9478 22494
rect 9494 22478 9519 22494
rect 9421 22462 9519 22478
rect 9421 22446 9446 22462
rect 9462 22446 9478 22462
rect 9494 22446 9519 22462
rect 9421 22430 9519 22446
rect 9421 22414 9446 22430
rect 9462 22414 9478 22430
rect 9494 22414 9519 22430
rect 9421 22400 9519 22414
rect 9621 22546 9719 22559
rect 9621 22530 9646 22546
rect 9662 22530 9678 22546
rect 9694 22530 9719 22546
rect 9621 22514 9719 22530
rect 9621 22498 9646 22514
rect 9662 22498 9678 22514
rect 9694 22498 9719 22514
rect 9621 22482 9719 22498
rect 9621 22466 9646 22482
rect 9662 22466 9678 22482
rect 9694 22466 9719 22482
rect 9621 22450 9719 22466
rect 9621 22434 9646 22450
rect 9662 22434 9678 22450
rect 9694 22434 9719 22450
rect 9621 22418 9719 22434
rect 9621 22402 9646 22418
rect 9662 22402 9678 22418
rect 9694 22402 9719 22418
rect 9219 20846 9319 20859
rect 9219 20830 9246 20846
rect 9262 20830 9278 20846
rect 9294 20830 9319 20846
rect 9219 20814 9319 20830
rect 9219 20798 9246 20814
rect 9262 20798 9278 20814
rect 9294 20798 9319 20814
rect 9219 20782 9319 20798
rect 9219 20766 9246 20782
rect 9262 20766 9278 20782
rect 9294 20766 9319 20782
rect 9219 20750 9319 20766
rect 9219 20734 9246 20750
rect 9262 20734 9278 20750
rect 9294 20734 9319 20750
rect 9219 20718 9319 20734
rect 9219 20702 9246 20718
rect 9262 20702 9278 20718
rect 9294 20702 9319 20718
rect 9219 20686 9319 20702
rect 9219 20670 9246 20686
rect 9262 20670 9278 20686
rect 9294 20670 9319 20686
rect 9219 20660 9319 20670
rect 8820 20654 9319 20660
rect 8820 20638 9246 20654
rect 9262 20638 9278 20654
rect 9294 20638 9319 20654
rect 8820 20622 9319 20638
rect 8820 20606 9246 20622
rect 9262 20606 9278 20622
rect 9294 20606 9319 20622
rect 8820 20590 9319 20606
rect 8820 20574 9246 20590
rect 9262 20574 9278 20590
rect 9294 20574 9319 20590
rect 8820 20561 9319 20574
rect 8820 20560 9220 20561
rect 9420 17960 9520 22400
rect 9621 22386 9719 22402
rect 9621 22370 9646 22386
rect 9662 22370 9678 22386
rect 9694 22370 9719 22386
rect 9621 22354 9719 22370
rect 9621 22338 9646 22354
rect 9662 22338 9678 22354
rect 9694 22338 9719 22354
rect 9621 22322 9719 22338
rect 9621 22306 9646 22322
rect 9662 22306 9678 22322
rect 9694 22306 9719 22322
rect 9621 22290 9719 22306
rect 9621 22274 9646 22290
rect 9662 22274 9678 22290
rect 9694 22274 9719 22290
rect 9621 22260 9719 22274
rect 8820 17860 9520 17960
rect 9620 15260 9720 22260
rect 28660 20679 29180 20680
rect 28361 20654 29180 20679
rect 28361 20638 28374 20654
rect 28390 20638 28406 20654
rect 28422 20638 28438 20654
rect 28454 20638 28470 20654
rect 28486 20638 28502 20654
rect 28518 20638 28534 20654
rect 28550 20638 28566 20654
rect 28582 20638 28598 20654
rect 28614 20638 28630 20654
rect 28646 20638 29180 20654
rect 28361 20622 29180 20638
rect 28361 20606 28374 20622
rect 28390 20606 28406 20622
rect 28422 20606 28438 20622
rect 28454 20606 28470 20622
rect 28486 20606 28502 20622
rect 28518 20606 28534 20622
rect 28550 20606 28566 20622
rect 28582 20606 28598 20622
rect 28614 20606 28630 20622
rect 28646 20606 29180 20622
rect 28361 20581 29180 20606
rect 28660 20580 29180 20581
rect 28860 17979 29180 17980
rect 28561 17954 29180 17979
rect 28561 17938 28574 17954
rect 28590 17938 28606 17954
rect 28622 17938 28638 17954
rect 28654 17938 28670 17954
rect 28686 17938 28702 17954
rect 28718 17938 28734 17954
rect 28750 17938 28766 17954
rect 28782 17938 28798 17954
rect 28814 17938 28830 17954
rect 28846 17938 29180 17954
rect 28561 17922 29180 17938
rect 28561 17906 28574 17922
rect 28590 17906 28606 17922
rect 28622 17906 28638 17922
rect 28654 17906 28670 17922
rect 28686 17906 28702 17922
rect 28718 17906 28734 17922
rect 28750 17906 28766 17922
rect 28782 17906 28798 17922
rect 28814 17906 28830 17922
rect 28846 17906 29180 17922
rect 28561 17881 29180 17906
rect 28860 17880 29180 17881
rect 8820 15160 9720 15260
rect 8820 9879 9380 9880
rect 8820 9866 9799 9879
rect 8820 9850 9406 9866
rect 9422 9850 9438 9866
rect 9454 9850 9470 9866
rect 9486 9850 9502 9866
rect 9518 9850 9534 9866
rect 9550 9850 9566 9866
rect 9582 9850 9598 9866
rect 9614 9850 9630 9866
rect 9646 9850 9662 9866
rect 9678 9850 9694 9866
rect 9710 9850 9726 9866
rect 9742 9850 9758 9866
rect 9774 9850 9799 9866
rect 8820 9834 9799 9850
rect 8820 9818 9406 9834
rect 9422 9818 9438 9834
rect 9454 9818 9470 9834
rect 9486 9818 9502 9834
rect 9518 9818 9534 9834
rect 9550 9818 9566 9834
rect 9582 9818 9598 9834
rect 9614 9818 9630 9834
rect 9646 9818 9662 9834
rect 9678 9818 9694 9834
rect 9710 9818 9726 9834
rect 9742 9818 9758 9834
rect 9774 9818 9799 9834
rect 8820 9802 9799 9818
rect 8820 9786 9406 9802
rect 9422 9786 9438 9802
rect 9454 9786 9470 9802
rect 9486 9786 9502 9802
rect 9518 9786 9534 9802
rect 9550 9786 9566 9802
rect 9582 9786 9598 9802
rect 9614 9786 9630 9802
rect 9646 9786 9662 9802
rect 9678 9786 9694 9802
rect 9710 9786 9726 9802
rect 9742 9786 9758 9802
rect 9774 9786 9799 9802
rect 8820 9770 9799 9786
rect 8820 9754 9406 9770
rect 9422 9754 9438 9770
rect 9454 9754 9470 9770
rect 9486 9754 9502 9770
rect 9518 9754 9534 9770
rect 9550 9754 9566 9770
rect 9582 9754 9598 9770
rect 9614 9754 9630 9770
rect 9646 9754 9662 9770
rect 9678 9754 9694 9770
rect 9710 9754 9726 9770
rect 9742 9754 9758 9770
rect 9774 9754 9799 9770
rect 8820 9741 9799 9754
rect 8820 9740 9380 9741
rect 15160 9660 15240 9780
rect 15161 9644 15239 9660
rect 15161 9628 15176 9644
rect 15192 9628 15208 9644
rect 15224 9628 15239 9644
rect 15161 9612 15239 9628
rect 15161 9596 15176 9612
rect 15192 9596 15208 9612
rect 15224 9596 15239 9612
rect 15161 9581 15239 9596
rect 15320 9500 15400 9780
rect 15321 9484 15399 9500
rect 15321 9468 15336 9484
rect 15352 9468 15368 9484
rect 15384 9468 15399 9484
rect 15321 9452 15399 9468
rect 15321 9436 15336 9452
rect 15352 9436 15368 9452
rect 15384 9436 15399 9452
rect 15321 9421 15399 9436
rect 14661 9404 14739 9419
rect 14661 9388 14676 9404
rect 14692 9388 14708 9404
rect 14724 9388 14739 9404
rect 14661 9372 14739 9388
rect 14661 9356 14676 9372
rect 14692 9356 14708 9372
rect 14724 9356 14739 9372
rect 14661 9340 14739 9356
rect 15720 9340 15800 9780
rect 11961 9244 12039 9259
rect 11961 9228 11976 9244
rect 11992 9228 12008 9244
rect 12024 9228 12039 9244
rect 11961 9212 12039 9228
rect 11961 9196 11976 9212
rect 11992 9196 12008 9212
rect 12024 9196 12039 9212
rect 11961 9180 12039 9196
rect 11960 8820 12040 9180
rect 14660 8820 14740 9340
rect 15721 9324 15799 9340
rect 15721 9308 15736 9324
rect 15752 9308 15768 9324
rect 15784 9308 15799 9324
rect 15721 9292 15799 9308
rect 15721 9276 15736 9292
rect 15752 9276 15768 9292
rect 15784 9276 15799 9292
rect 15721 9261 15799 9276
rect 16060 9180 16140 9780
rect 16061 9164 16139 9180
rect 16061 9148 16076 9164
rect 16092 9148 16108 9164
rect 16124 9148 16139 9164
rect 16061 9132 16139 9148
rect 16061 9116 16076 9132
rect 16092 9116 16108 9132
rect 16124 9116 16139 9132
rect 16061 9101 16139 9116
rect 16220 8980 16300 9780
rect 23940 9420 24020 9780
rect 23941 9404 24019 9420
rect 23941 9388 23956 9404
rect 23972 9388 23988 9404
rect 24004 9388 24019 9404
rect 23941 9372 24019 9388
rect 23941 9356 23956 9372
rect 23972 9356 23988 9372
rect 24004 9356 24019 9372
rect 23941 9341 24019 9356
rect 22741 9324 22819 9339
rect 22741 9308 22756 9324
rect 22772 9308 22788 9324
rect 22804 9308 22819 9324
rect 22741 9292 22819 9308
rect 22741 9276 22756 9292
rect 22772 9276 22788 9292
rect 22804 9276 22819 9292
rect 22741 9260 22819 9276
rect 24100 9260 24180 9780
rect 28161 9644 28239 9659
rect 28161 9628 28176 9644
rect 28192 9628 28208 9644
rect 28224 9628 28239 9644
rect 28161 9612 28239 9628
rect 28161 9596 28176 9612
rect 28192 9596 28208 9612
rect 28224 9596 28239 9612
rect 28161 9580 28239 9596
rect 25461 9484 25539 9499
rect 25461 9468 25476 9484
rect 25492 9468 25508 9484
rect 25524 9468 25539 9484
rect 25461 9452 25539 9468
rect 25461 9436 25476 9452
rect 25492 9436 25508 9452
rect 25524 9436 25539 9452
rect 25461 9420 25539 9436
rect 20061 9164 20139 9179
rect 20061 9148 20076 9164
rect 20092 9148 20108 9164
rect 20124 9148 20139 9164
rect 20061 9132 20139 9148
rect 20061 9116 20076 9132
rect 20092 9116 20108 9132
rect 20124 9116 20139 9132
rect 20061 9100 20139 9116
rect 16220 8900 17440 8980
rect 17360 8820 17440 8900
rect 20060 8820 20140 9100
rect 22740 8820 22820 9260
rect 24101 9244 24179 9260
rect 24101 9228 24116 9244
rect 24132 9228 24148 9244
rect 24164 9228 24179 9244
rect 24101 9212 24179 9228
rect 24101 9196 24116 9212
rect 24132 9196 24148 9212
rect 24164 9196 24179 9212
rect 24101 9181 24179 9196
rect 25460 8820 25540 9420
rect 28160 8820 28240 9580
<< m3contact >>
rect 15206 28430 15222 28446
rect 15238 28430 15254 28446
rect 15206 28398 15222 28414
rect 15238 28398 15254 28414
rect 17906 28458 17922 28474
rect 17938 28458 17954 28474
rect 17906 28426 17922 28442
rect 17938 28426 17954 28442
rect 15206 28366 15222 28382
rect 15238 28366 15254 28382
rect 15206 28334 15222 28350
rect 15238 28334 15254 28350
rect 15206 28302 15222 28318
rect 15238 28302 15254 28318
rect 15206 28270 15222 28286
rect 15238 28270 15254 28286
rect 15206 28238 15222 28254
rect 15238 28238 15254 28254
rect 15206 28206 15222 28222
rect 15238 28206 15254 28222
rect 15206 28174 15222 28190
rect 15238 28174 15254 28190
rect 26366 28458 26382 28474
rect 26398 28458 26414 28474
rect 26366 28426 26382 28442
rect 26398 28426 26414 28442
rect 28554 26038 28570 26054
rect 28586 26038 28602 26054
rect 28618 26038 28634 26054
rect 28650 26038 28666 26054
rect 28682 26038 28698 26054
rect 28714 26038 28730 26054
rect 28746 26038 28762 26054
rect 28778 26038 28794 26054
rect 28810 26038 28826 26054
rect 28554 26006 28570 26022
rect 28586 26006 28602 26022
rect 28618 26006 28634 26022
rect 28650 26006 28666 26022
rect 28682 26006 28698 26022
rect 28714 26006 28730 26022
rect 28746 26006 28762 26022
rect 28778 26006 28794 26022
rect 28810 26006 28826 26022
rect 9046 23330 9062 23346
rect 9078 23330 9094 23346
rect 9046 23298 9062 23314
rect 9078 23298 9094 23314
rect 9046 23266 9062 23282
rect 9078 23266 9094 23282
rect 28354 23338 28370 23354
rect 28386 23338 28402 23354
rect 28418 23338 28434 23354
rect 28450 23338 28466 23354
rect 28482 23338 28498 23354
rect 28514 23338 28530 23354
rect 28546 23338 28562 23354
rect 28578 23338 28594 23354
rect 28610 23338 28626 23354
rect 28354 23306 28370 23322
rect 28386 23306 28402 23322
rect 28418 23306 28434 23322
rect 28450 23306 28466 23322
rect 28482 23306 28498 23322
rect 28514 23306 28530 23322
rect 28546 23306 28562 23322
rect 28578 23306 28594 23322
rect 28610 23306 28626 23322
rect 9046 23234 9062 23250
rect 9078 23234 9094 23250
rect 9046 23202 9062 23218
rect 9078 23202 9094 23218
rect 9046 23170 9062 23186
rect 9078 23170 9094 23186
rect 9046 23138 9062 23154
rect 9078 23138 9094 23154
rect 9046 23106 9062 23122
rect 9078 23106 9094 23122
rect 9046 23074 9062 23090
rect 9078 23074 9094 23090
rect 9446 22670 9462 22686
rect 9478 22670 9494 22686
rect 9446 22638 9462 22654
rect 9478 22638 9494 22654
rect 9446 22606 9462 22622
rect 9478 22606 9494 22622
rect 9446 22574 9462 22590
rect 9478 22574 9494 22590
rect 9446 22542 9462 22558
rect 9478 22542 9494 22558
rect 9446 22510 9462 22526
rect 9478 22510 9494 22526
rect 9446 22478 9462 22494
rect 9478 22478 9494 22494
rect 9446 22446 9462 22462
rect 9478 22446 9494 22462
rect 9446 22414 9462 22430
rect 9478 22414 9494 22430
rect 9646 22530 9662 22546
rect 9678 22530 9694 22546
rect 9646 22498 9662 22514
rect 9678 22498 9694 22514
rect 9646 22466 9662 22482
rect 9678 22466 9694 22482
rect 9646 22434 9662 22450
rect 9678 22434 9694 22450
rect 9646 22402 9662 22418
rect 9678 22402 9694 22418
rect 9246 20830 9262 20846
rect 9278 20830 9294 20846
rect 9246 20798 9262 20814
rect 9278 20798 9294 20814
rect 9246 20766 9262 20782
rect 9278 20766 9294 20782
rect 9246 20734 9262 20750
rect 9278 20734 9294 20750
rect 9246 20702 9262 20718
rect 9278 20702 9294 20718
rect 9246 20670 9262 20686
rect 9278 20670 9294 20686
rect 9246 20638 9262 20654
rect 9278 20638 9294 20654
rect 9246 20606 9262 20622
rect 9278 20606 9294 20622
rect 9246 20574 9262 20590
rect 9278 20574 9294 20590
rect 9646 22370 9662 22386
rect 9678 22370 9694 22386
rect 9646 22338 9662 22354
rect 9678 22338 9694 22354
rect 9646 22306 9662 22322
rect 9678 22306 9694 22322
rect 9646 22274 9662 22290
rect 9678 22274 9694 22290
rect 28374 20638 28390 20654
rect 28406 20638 28422 20654
rect 28438 20638 28454 20654
rect 28470 20638 28486 20654
rect 28502 20638 28518 20654
rect 28534 20638 28550 20654
rect 28566 20638 28582 20654
rect 28598 20638 28614 20654
rect 28630 20638 28646 20654
rect 28374 20606 28390 20622
rect 28406 20606 28422 20622
rect 28438 20606 28454 20622
rect 28470 20606 28486 20622
rect 28502 20606 28518 20622
rect 28534 20606 28550 20622
rect 28566 20606 28582 20622
rect 28598 20606 28614 20622
rect 28630 20606 28646 20622
rect 28574 17938 28590 17954
rect 28606 17938 28622 17954
rect 28638 17938 28654 17954
rect 28670 17938 28686 17954
rect 28702 17938 28718 17954
rect 28734 17938 28750 17954
rect 28766 17938 28782 17954
rect 28798 17938 28814 17954
rect 28830 17938 28846 17954
rect 28574 17906 28590 17922
rect 28606 17906 28622 17922
rect 28638 17906 28654 17922
rect 28670 17906 28686 17922
rect 28702 17906 28718 17922
rect 28734 17906 28750 17922
rect 28766 17906 28782 17922
rect 28798 17906 28814 17922
rect 28830 17906 28846 17922
rect 9406 9850 9422 9866
rect 9438 9850 9454 9866
rect 9470 9850 9486 9866
rect 9502 9850 9518 9866
rect 9534 9850 9550 9866
rect 9566 9850 9582 9866
rect 9598 9850 9614 9866
rect 9630 9850 9646 9866
rect 9662 9850 9678 9866
rect 9694 9850 9710 9866
rect 9726 9850 9742 9866
rect 9758 9850 9774 9866
rect 9406 9818 9422 9834
rect 9438 9818 9454 9834
rect 9470 9818 9486 9834
rect 9502 9818 9518 9834
rect 9534 9818 9550 9834
rect 9566 9818 9582 9834
rect 9598 9818 9614 9834
rect 9630 9818 9646 9834
rect 9662 9818 9678 9834
rect 9694 9818 9710 9834
rect 9726 9818 9742 9834
rect 9758 9818 9774 9834
rect 9406 9786 9422 9802
rect 9438 9786 9454 9802
rect 9470 9786 9486 9802
rect 9502 9786 9518 9802
rect 9534 9786 9550 9802
rect 9566 9786 9582 9802
rect 9598 9786 9614 9802
rect 9630 9786 9646 9802
rect 9662 9786 9678 9802
rect 9694 9786 9710 9802
rect 9726 9786 9742 9802
rect 9758 9786 9774 9802
rect 9406 9754 9422 9770
rect 9438 9754 9454 9770
rect 9470 9754 9486 9770
rect 9502 9754 9518 9770
rect 9534 9754 9550 9770
rect 9566 9754 9582 9770
rect 9598 9754 9614 9770
rect 9630 9754 9646 9770
rect 9662 9754 9678 9770
rect 9694 9754 9710 9770
rect 9726 9754 9742 9770
rect 9758 9754 9774 9770
rect 15176 9628 15192 9644
rect 15208 9628 15224 9644
rect 15176 9596 15192 9612
rect 15208 9596 15224 9612
rect 15336 9468 15352 9484
rect 15368 9468 15384 9484
rect 15336 9436 15352 9452
rect 15368 9436 15384 9452
rect 15736 9308 15752 9324
rect 15768 9308 15784 9324
rect 15736 9276 15752 9292
rect 15768 9276 15784 9292
rect 16076 9148 16092 9164
rect 16108 9148 16124 9164
rect 16076 9116 16092 9132
rect 16108 9116 16124 9132
rect 22756 9308 22772 9324
rect 22788 9308 22804 9324
rect 22756 9276 22772 9292
rect 22788 9276 22804 9292
rect 28176 9628 28192 9644
rect 28208 9628 28224 9644
rect 28176 9596 28192 9612
rect 28208 9596 28224 9612
rect 25476 9468 25492 9484
rect 25508 9468 25524 9484
rect 25476 9436 25492 9452
rect 25508 9436 25524 9452
rect 20076 9148 20092 9164
rect 20108 9148 20124 9164
rect 20076 9116 20092 9132
rect 20108 9116 20124 9132
<< metal3 >>
rect 17980 28499 26340 28500
rect 17881 28474 26439 28499
rect 15181 28446 15280 28459
rect 15181 28430 15206 28446
rect 15222 28430 15238 28446
rect 15254 28430 15280 28446
rect 15181 28414 15280 28430
rect 15181 28398 15206 28414
rect 15222 28398 15238 28414
rect 15254 28398 15280 28414
rect 17881 28458 17906 28474
rect 17922 28458 17938 28474
rect 17954 28458 26366 28474
rect 26382 28458 26398 28474
rect 26414 28458 26439 28474
rect 17881 28442 26439 28458
rect 17881 28426 17906 28442
rect 17922 28426 17938 28442
rect 17954 28426 26366 28442
rect 26382 28426 26398 28442
rect 26414 28426 26439 28442
rect 17881 28401 26439 28426
rect 17980 28400 26340 28401
rect 15181 28382 15280 28398
rect 15181 28366 15206 28382
rect 15222 28366 15238 28382
rect 15254 28366 15280 28382
rect 15181 28350 15280 28366
rect 15181 28334 15206 28350
rect 15222 28334 15238 28350
rect 15254 28334 15280 28350
rect 15181 28318 15280 28334
rect 15181 28302 15206 28318
rect 15222 28302 15238 28318
rect 15254 28302 15280 28318
rect 15181 28286 15280 28302
rect 15181 28270 15206 28286
rect 15222 28270 15238 28286
rect 15254 28270 15280 28286
rect 15181 28260 15280 28270
rect 15181 28254 17340 28260
rect 15181 28238 15206 28254
rect 15222 28238 15238 28254
rect 15254 28238 17340 28254
rect 15181 28222 17340 28238
rect 15181 28206 15206 28222
rect 15222 28206 15238 28222
rect 15254 28206 17340 28222
rect 15181 28190 17340 28206
rect 15181 28174 15206 28190
rect 15222 28174 15238 28190
rect 15254 28174 17340 28190
rect 15181 28161 17340 28174
rect 15280 28160 17340 28161
rect 17240 27900 17340 28160
rect 28060 27580 28640 27680
rect 9740 27420 10080 27520
rect 9740 26260 9820 27420
rect 28060 27400 28440 27500
rect 9220 26160 9820 26260
rect 9021 23346 9119 23359
rect 9021 23330 9046 23346
rect 9062 23330 9078 23346
rect 9094 23330 9119 23346
rect 9021 23314 9119 23330
rect 9021 23298 9046 23314
rect 9062 23298 9078 23314
rect 9094 23298 9119 23314
rect 9021 23282 9119 23298
rect 9021 23266 9046 23282
rect 9062 23266 9078 23282
rect 9094 23266 9119 23282
rect 9021 23250 9119 23266
rect 9021 23234 9046 23250
rect 9062 23234 9078 23250
rect 9094 23234 9119 23250
rect 9021 23218 9119 23234
rect 9021 23202 9046 23218
rect 9062 23202 9078 23218
rect 9094 23202 9119 23218
rect 9021 23186 9119 23202
rect 9021 23170 9046 23186
rect 9062 23170 9078 23186
rect 9094 23170 9119 23186
rect 9021 23154 9119 23170
rect 9021 23138 9046 23154
rect 9062 23138 9078 23154
rect 9094 23138 9119 23154
rect 9021 23122 9119 23138
rect 9021 23106 9046 23122
rect 9062 23106 9078 23122
rect 9094 23106 9119 23122
rect 9021 23090 9119 23106
rect 9021 23074 9046 23090
rect 9062 23074 9078 23090
rect 9094 23074 9119 23090
rect 9021 23060 9119 23074
rect 9020 19600 9120 23060
rect 9220 20860 9320 26160
rect 28340 23380 28440 27400
rect 28540 26080 28640 27580
rect 28541 26054 28839 26080
rect 28541 26038 28554 26054
rect 28570 26038 28586 26054
rect 28602 26038 28618 26054
rect 28634 26038 28650 26054
rect 28666 26038 28682 26054
rect 28698 26038 28714 26054
rect 28730 26038 28746 26054
rect 28762 26038 28778 26054
rect 28794 26038 28810 26054
rect 28826 26038 28839 26054
rect 28541 26022 28839 26038
rect 28541 26006 28554 26022
rect 28570 26006 28586 26022
rect 28602 26006 28618 26022
rect 28634 26006 28650 26022
rect 28666 26006 28682 26022
rect 28698 26006 28714 26022
rect 28730 26006 28746 26022
rect 28762 26006 28778 26022
rect 28794 26006 28810 26022
rect 28826 26006 28839 26022
rect 28541 25981 28839 26006
rect 28341 23354 28639 23380
rect 28341 23338 28354 23354
rect 28370 23338 28386 23354
rect 28402 23338 28418 23354
rect 28434 23338 28450 23354
rect 28466 23338 28482 23354
rect 28498 23338 28514 23354
rect 28530 23338 28546 23354
rect 28562 23338 28578 23354
rect 28594 23338 28610 23354
rect 28626 23338 28639 23354
rect 28341 23322 28639 23338
rect 28341 23306 28354 23322
rect 28370 23306 28386 23322
rect 28402 23306 28418 23322
rect 28434 23306 28450 23322
rect 28466 23306 28482 23322
rect 28498 23306 28514 23322
rect 28530 23306 28546 23322
rect 28562 23306 28578 23322
rect 28594 23306 28610 23322
rect 28626 23306 28639 23322
rect 28341 23281 28639 23306
rect 9520 22699 10100 22700
rect 9421 22686 10100 22699
rect 9421 22670 9446 22686
rect 9462 22670 9478 22686
rect 9494 22670 10100 22686
rect 9421 22654 10100 22670
rect 9421 22638 9446 22654
rect 9462 22638 9478 22654
rect 9494 22638 10100 22654
rect 9421 22622 10100 22638
rect 9421 22606 9446 22622
rect 9462 22606 9478 22622
rect 9494 22620 10100 22622
rect 9494 22606 9520 22620
rect 9421 22590 9520 22606
rect 9421 22574 9446 22590
rect 9462 22574 9478 22590
rect 9494 22574 9520 22590
rect 9421 22558 9520 22574
rect 9720 22559 10100 22560
rect 9421 22542 9446 22558
rect 9462 22542 9478 22558
rect 9494 22542 9520 22558
rect 9421 22526 9520 22542
rect 9421 22510 9446 22526
rect 9462 22510 9478 22526
rect 9494 22510 9520 22526
rect 9421 22494 9520 22510
rect 9421 22478 9446 22494
rect 9462 22478 9478 22494
rect 9494 22478 9520 22494
rect 9421 22462 9520 22478
rect 9421 22446 9446 22462
rect 9462 22446 9478 22462
rect 9494 22446 9520 22462
rect 9421 22430 9520 22446
rect 9421 22414 9446 22430
rect 9462 22414 9478 22430
rect 9494 22414 9520 22430
rect 9421 22401 9520 22414
rect 9621 22546 10100 22559
rect 9621 22530 9646 22546
rect 9662 22530 9678 22546
rect 9694 22530 10100 22546
rect 9621 22514 10100 22530
rect 9621 22498 9646 22514
rect 9662 22498 9678 22514
rect 9694 22498 10100 22514
rect 9621 22482 10100 22498
rect 9621 22466 9646 22482
rect 9662 22466 9678 22482
rect 9694 22480 10100 22482
rect 9694 22466 9720 22480
rect 9621 22450 9720 22466
rect 9621 22434 9646 22450
rect 9662 22434 9678 22450
rect 9694 22434 9720 22450
rect 9621 22418 9720 22434
rect 9621 22402 9646 22418
rect 9662 22402 9678 22418
rect 9694 22402 9720 22418
rect 9621 22386 9720 22402
rect 9621 22370 9646 22386
rect 9662 22370 9678 22386
rect 9694 22370 9720 22386
rect 9621 22354 9720 22370
rect 9621 22338 9646 22354
rect 9662 22338 9678 22354
rect 9694 22338 9720 22354
rect 9621 22322 9720 22338
rect 9621 22306 9646 22322
rect 9662 22306 9678 22322
rect 9694 22306 9720 22322
rect 9621 22290 9720 22306
rect 9621 22274 9646 22290
rect 9662 22274 9678 22290
rect 9694 22274 9720 22290
rect 9621 22261 9720 22274
rect 9221 20846 9319 20860
rect 9221 20830 9246 20846
rect 9262 20830 9278 20846
rect 9294 20830 9319 20846
rect 9221 20814 9319 20830
rect 9221 20798 9246 20814
rect 9262 20798 9278 20814
rect 9294 20798 9319 20814
rect 9221 20782 9319 20798
rect 9221 20766 9246 20782
rect 9262 20766 9278 20782
rect 9294 20766 9319 20782
rect 9221 20750 9319 20766
rect 9221 20734 9246 20750
rect 9262 20734 9278 20750
rect 9294 20734 9319 20750
rect 9221 20718 9319 20734
rect 9221 20702 9246 20718
rect 9262 20702 9278 20718
rect 9294 20702 9319 20718
rect 9221 20686 9319 20702
rect 9221 20670 9246 20686
rect 9262 20670 9278 20686
rect 9294 20670 9319 20686
rect 9221 20654 9319 20670
rect 9221 20638 9246 20654
rect 9262 20638 9278 20654
rect 9294 20638 9319 20654
rect 9221 20622 9319 20638
rect 9221 20606 9246 20622
rect 9262 20606 9278 20622
rect 9294 20606 9319 20622
rect 9221 20590 9319 20606
rect 9221 20574 9246 20590
rect 9262 20574 9278 20590
rect 9294 20574 9319 20590
rect 28361 20654 28659 20679
rect 28361 20638 28374 20654
rect 28390 20638 28406 20654
rect 28422 20638 28438 20654
rect 28454 20638 28470 20654
rect 28486 20638 28502 20654
rect 28518 20638 28534 20654
rect 28550 20638 28566 20654
rect 28582 20638 28598 20654
rect 28614 20638 28630 20654
rect 28646 20638 28659 20654
rect 28361 20622 28659 20638
rect 28361 20606 28374 20622
rect 28390 20606 28406 20622
rect 28422 20606 28438 20622
rect 28454 20606 28470 20622
rect 28486 20606 28502 20622
rect 28518 20606 28534 20622
rect 28550 20606 28566 20622
rect 28582 20606 28598 20622
rect 28614 20606 28630 20622
rect 28646 20606 28659 20622
rect 28361 20580 28659 20606
rect 9221 20561 9319 20574
rect 9020 19500 10080 19600
rect 28360 16720 28460 20580
rect 28561 17954 28859 17979
rect 28561 17938 28574 17954
rect 28590 17938 28606 17954
rect 28622 17938 28638 17954
rect 28654 17938 28670 17954
rect 28686 17938 28702 17954
rect 28718 17938 28734 17954
rect 28750 17938 28766 17954
rect 28782 17938 28798 17954
rect 28814 17938 28830 17954
rect 28846 17938 28859 17954
rect 28561 17922 28859 17938
rect 28561 17906 28574 17922
rect 28590 17906 28606 17922
rect 28622 17906 28638 17922
rect 28654 17906 28670 17922
rect 28686 17906 28702 17922
rect 28718 17906 28734 17922
rect 28750 17906 28766 17922
rect 28782 17906 28798 17922
rect 28814 17906 28830 17922
rect 28846 17906 28859 17922
rect 28561 17880 28859 17906
rect 28040 16620 28460 16720
rect 28560 16040 28660 17880
rect 28040 15940 28660 16040
rect 9660 13780 10080 13920
rect 9660 9880 9800 13780
rect 9381 9866 9799 9880
rect 9381 9850 9406 9866
rect 9422 9850 9438 9866
rect 9454 9850 9470 9866
rect 9486 9850 9502 9866
rect 9518 9850 9534 9866
rect 9550 9850 9566 9866
rect 9582 9850 9598 9866
rect 9614 9850 9630 9866
rect 9646 9850 9662 9866
rect 9678 9850 9694 9866
rect 9710 9850 9726 9866
rect 9742 9850 9758 9866
rect 9774 9850 9799 9866
rect 9381 9834 9799 9850
rect 9381 9818 9406 9834
rect 9422 9818 9438 9834
rect 9454 9818 9470 9834
rect 9486 9818 9502 9834
rect 9518 9818 9534 9834
rect 9550 9818 9566 9834
rect 9582 9818 9598 9834
rect 9614 9818 9630 9834
rect 9646 9818 9662 9834
rect 9678 9818 9694 9834
rect 9710 9818 9726 9834
rect 9742 9818 9758 9834
rect 9774 9818 9799 9834
rect 9381 9802 9799 9818
rect 9381 9786 9406 9802
rect 9422 9786 9438 9802
rect 9454 9786 9470 9802
rect 9486 9786 9502 9802
rect 9518 9786 9534 9802
rect 9550 9786 9566 9802
rect 9582 9786 9598 9802
rect 9614 9786 9630 9802
rect 9646 9786 9662 9802
rect 9678 9786 9694 9802
rect 9710 9786 9726 9802
rect 9742 9786 9758 9802
rect 9774 9786 9799 9802
rect 9381 9770 9799 9786
rect 9381 9754 9406 9770
rect 9422 9754 9438 9770
rect 9454 9754 9470 9770
rect 9486 9754 9502 9770
rect 9518 9754 9534 9770
rect 9550 9754 9566 9770
rect 9582 9754 9598 9770
rect 9614 9754 9630 9770
rect 9646 9754 9662 9770
rect 9678 9754 9694 9770
rect 9710 9754 9726 9770
rect 9742 9754 9758 9770
rect 9774 9754 9799 9770
rect 9381 9741 9799 9754
rect 15240 9659 28160 9660
rect 15161 9644 28239 9659
rect 15161 9628 15176 9644
rect 15192 9628 15208 9644
rect 15224 9628 28176 9644
rect 28192 9628 28208 9644
rect 28224 9628 28239 9644
rect 15161 9612 28239 9628
rect 15161 9596 15176 9612
rect 15192 9596 15208 9612
rect 15224 9596 28176 9612
rect 28192 9596 28208 9612
rect 28224 9596 28239 9612
rect 15161 9581 28239 9596
rect 15240 9580 28160 9581
rect 15400 9499 25460 9500
rect 15321 9484 25539 9499
rect 15321 9468 15336 9484
rect 15352 9468 15368 9484
rect 15384 9468 25476 9484
rect 25492 9468 25508 9484
rect 25524 9468 25539 9484
rect 15321 9452 25539 9468
rect 15321 9436 15336 9452
rect 15352 9436 15368 9452
rect 15384 9436 25476 9452
rect 25492 9436 25508 9452
rect 25524 9436 25539 9452
rect 15321 9421 25539 9436
rect 15400 9420 25460 9421
rect 15800 9339 22740 9340
rect 15721 9324 22819 9339
rect 15721 9308 15736 9324
rect 15752 9308 15768 9324
rect 15784 9308 22756 9324
rect 22772 9308 22788 9324
rect 22804 9308 22819 9324
rect 15721 9292 22819 9308
rect 15721 9276 15736 9292
rect 15752 9276 15768 9292
rect 15784 9276 22756 9292
rect 22772 9276 22788 9292
rect 22804 9276 22819 9292
rect 15721 9261 22819 9276
rect 15800 9260 22740 9261
rect 16140 9179 20060 9180
rect 16061 9164 20139 9179
rect 16061 9148 16076 9164
rect 16092 9148 16108 9164
rect 16124 9148 20076 9164
rect 20092 9148 20108 9164
rect 20124 9148 20139 9164
rect 16061 9132 20139 9148
rect 16061 9116 16076 9132
rect 16092 9116 16108 9132
rect 16124 9116 20076 9132
rect 20092 9116 20108 9132
rect 20124 9116 20139 9132
rect 16061 9101 20139 9116
rect 16140 9100 20060 9101
<< end >>
