/* Verilog module written by DEF2Verilog (qflow) */
module cordic_element (
    input [1:0] Ain,
    output [1:0] Aout,
    input ISin,
    output ISout,
    input Rdy,
    input [2:0] Stg,
    output Vld,
    input [1:0] Xin,
    output [1:0] Xout,
    input [1:0] Yin,
    output [1:0] Yout,
    input clk
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [6:0] LoadCtl ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire ISin ;
wire _506_ ;
wire [11:0] Acalc ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire ISout ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire [1:0] _861_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire _285_ ;
wire _1_ ;
wire [2:0] Stg ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire Stg_0_bF$buf0 ;
wire Stg_0_bF$buf1 ;
wire Stg_0_bF$buf2 ;
wire Stg_0_bF$buf3 ;
wire Stg_0_bF$buf4 ;
wire Stg_0_bF$buf5 ;
wire Stg_0_bF$buf6 ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire [11:0] Ycalc ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _188__bF$buf0 ;
wire _188__bF$buf1 ;
wire _188__bF$buf2 ;
wire _188__bF$buf3 ;
wire _188__bF$buf4 ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire [1:0] Ain0 ;
wire [1:0] Ain1 ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire Stg_2_bF$buf0 ;
wire Stg_2_bF$buf1 ;
wire Stg_2_bF$buf2 ;
wire Stg_2_bF$buf3 ;
wire Stg_2_bF$buf4 ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [11:4] Xin12b ;
wire [1:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire [11:0] Xcalc ;
wire [1:0] Yin0 ;
wire [1:0] Yin1 ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire [1:0] Aout ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _201__bF$buf0 ;
wire _201__bF$buf1 ;
wire _201__bF$buf2 ;
wire _201__bF$buf3 ;
wire _201__bF$buf4 ;
wire _201__bF$buf5 ;
wire _201__bF$buf6 ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire [1:0] Xin0 ;
wire [1:0] Xin1 ;
wire _534_ ;
wire _114_ ;
wire Ain12b_11_bF$buf0 ;
wire Ain12b_11_bF$buf1 ;
wire Ain12b_11_bF$buf2 ;
wire Ain12b_11_bF$buf3 ;
wire Ain12b_11_bF$buf4 ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire [1:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire [1:0] Ain ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [1:0] Xout ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire [11:4] Ain12b ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _164__bF$buf0 ;
wire _164__bF$buf1 ;
wire _164__bF$buf2 ;
wire _164__bF$buf3 ;
wire _164__bF$buf4 ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _183__bF$buf0 ;
wire _183__bF$buf1 ;
wire _183__bF$buf2 ;
wire _183__bF$buf3 ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire LoadCtl_6_bF$buf0 ;
wire LoadCtl_6_bF$buf1 ;
wire LoadCtl_6_bF$buf2 ;
wire LoadCtl_6_bF$buf3 ;
wire LoadCtl_6_bF$buf4 ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire [11:4] Yin12b ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire [1:0] _862_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire gnd = 1'b0 ;
wire [1:0] _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire Stg_1_bF$buf0 ;
wire Stg_1_bF$buf1 ;
wire Stg_1_bF$buf2 ;
wire Stg_1_bF$buf3 ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire [1:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire vdd = 1'b1 ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_0__1661_ (
);

FILL FILL_0__1241_ (
);

FILL FILL_1__1402_ (
);

INVX1 _1677_ (
    .A(_843_),
    .Y(_844_)
);

NAND3X1 _1257_ (
    .A(_457_),
    .B(_479_),
    .C(_466_),
    .Y(_481_)
);

FILL FILL_0__1717_ (
);

FILL FILL_0__1470_ (
);

FILL FILL_0__1050_ (
);

FILL FILL_2__1068_ (
);

FILL FILL_1__1631_ (
);

FILL FILL_1__1211_ (
);

INVX1 _1486_ (
    .A(_119_),
    .Y(_665_)
);

OAI21X1 _1066_ (
    .A(Ain12b_11_bF$buf0),
    .B(_298_),
    .C(_295_),
    .Y(_299_)
);

FILL FILL_2__1700_ (
);

FILL FILL_0__1526_ (
);

FILL FILL_0__1106_ (
);

FILL FILL_2__1297_ (
);

FILL FILL_1__1440_ (
);

FILL FILL_1__1020_ (
);

OAI21X1 _1295_ (
    .A(_513_),
    .B(_515_),
    .C(_503_),
    .Y(_16_)
);

FILL FILL_0__1335_ (
);

FILL FILL_1__886_ (
);

FILL FILL_0__1564_ (
);

FILL FILL_0__1144_ (
);

FILL FILL_1__1725_ (
);

FILL FILL_1__1305_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_0_BUFX2_insert21 (
);

FILL FILL_0_BUFX2_insert22 (
);

FILL FILL_0_BUFX2_insert23 (
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_0_BUFX2_insert26 (
);

FILL FILL_0_BUFX2_insert27 (
);

FILL FILL_0_BUFX2_insert28 (
);

FILL FILL_0_BUFX2_insert29 (
);

FILL FILL_0__1373_ (
);

FILL FILL_1__1534_ (
);

FILL FILL_1__1114_ (
);

NAND2X1 _1389_ (
    .A(Acalc[9]),
    .B(_188__bF$buf4),
    .Y(_603_)
);

FILL FILL88350x75750 (
);

FILL FILL_2__1603_ (
);

FILL FILL_0__1429_ (
);

FILL FILL_0__1009_ (
);

FILL FILL_2__958_ (
);

FILL FILL_0__1182_ (
);

OAI21X1 _1601_ (
    .A(Stg_2_bF$buf0),
    .B(_484_),
    .C(_771_),
    .Y(_772_)
);

NAND2X1 _932_ (
    .A(Xin0[1]),
    .B(Stg_0_bF$buf6),
    .Y(_169_)
);

FILL FILL_1__1343_ (
);

NAND3X1 _1198_ (
    .A(_422_),
    .B(_423_),
    .C(_424_),
    .Y(_425_)
);

FILL FILL_0__1658_ (
);

FILL FILL_0__1238_ (
);

NAND2X1 _1410_ (
    .A(Acalc[11]),
    .B(_188__bF$buf4),
    .Y(_622_)
);

FILL FILL_1__1572_ (
);

FILL FILL_1__1152_ (
);

BUFX2 BUFX2_insert30 (
    .A(Stg[2]),
    .Y(Stg_2_bF$buf4)
);

BUFX2 BUFX2_insert31 (
    .A(Stg[2]),
    .Y(Stg_2_bF$buf3)
);

BUFX2 BUFX2_insert32 (
    .A(Stg[2]),
    .Y(Stg_2_bF$buf2)
);

BUFX2 BUFX2_insert33 (
    .A(Stg[2]),
    .Y(Stg_2_bF$buf1)
);

BUFX2 BUFX2_insert34 (
    .A(Stg[2]),
    .Y(Stg_2_bF$buf0)
);

BUFX2 BUFX2_insert35 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert36 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert37 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

BUFX2 BUFX2_insert38 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

BUFX2 BUFX2_insert39 (
    .A(Stg[1]),
    .Y(Stg_1_bF$buf3)
);

FILL FILL_2__1221_ (
);

FILL FILL_0__1467_ (
);

FILL FILL_0__1047_ (
);

FILL FILL_1__1628_ (
);

FILL FILL_1__1208_ (
);

NAND2X1 _970_ (
    .A(Stg_0_bF$buf6),
    .B(Xin1[0]),
    .Y(_206_)
);

FILL FILL_1__1381_ (
);

FILL FILL_2__1450_ (
);

FILL FILL_2__1030_ (
);

FILL FILL_0__1696_ (
);

FILL FILL_0__1276_ (
);

FILL FILL_1__1437_ (
);

FILL FILL_1__1017_ (
);

FILL FILL_1__1190_ (
);

FILL FILL_0__1085_ (
);

AOI21X1 _1504_ (
    .A(Stg_2_bF$buf1),
    .B(_676_),
    .C(_677_),
    .Y(_678_)
);

FILL FILL_1__1666_ (
);

FILL FILL_1__1246_ (
);

DFFPOSX1 _1733_ (
    .D(_5_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[3])
);

NOR2X1 _1313_ (
    .A(Ain12b_11_bF$buf0),
    .B(_494_),
    .Y(_532_)
);

FILL FILL_1__1475_ (
);

FILL FILL_1__1055_ (
);

FILL FILL_2__1544_ (
);

FILL FILL_2__1124_ (
);

FILL FILL_2__899_ (
);

NAND2X1 _1542_ (
    .A(_164__bF$buf4),
    .B(_221_),
    .Y(_715_)
);

OAI21X1 _1122_ (
    .A(_348_),
    .B(_331_),
    .C(_343_),
    .Y(_352_)
);

FILL FILL_0__870_ (
);

FILL FILL_1__904_ (
);

NOR2X1 _873_ (
    .A(LoadCtl_0_bF$buf2),
    .B(LoadCtl[1]),
    .Y(_116_)
);

FILL FILL_1__1284_ (
);

FILL FILL_0__1599_ (
);

FILL FILL_0__1179_ (
);

FILL FILL_0__926_ (
);

NAND2X1 _929_ (
    .A(Stg_0_bF$buf1),
    .B(Xin1[1]),
    .Y(_166_)
);

DFFPOSX1 _1771_ (
    .D(_43_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[7])
);

INVX1 _1351_ (
    .A(Ain12b[6]),
    .Y(_568_)
);

FILL FILL_1__1093_ (
);

FILL FILL_0__1811_ (
);

AND2X2 _1407_ (
    .A(_615_),
    .B(_619_),
    .Y(_620_)
);

FILL FILL_1__1569_ (
);

FILL FILL_1__1149_ (
);

AND2X2 _1580_ (
    .A(_751_),
    .B(_729_),
    .Y(_752_)
);

NOR2X1 _1160_ (
    .A(_382_),
    .B(_387_),
    .Y(_389_)
);

FILL FILL_1__942_ (
);

FILL FILL_0__1620_ (
);

FILL FILL_0__1200_ (
);

FILL FILL_2__1391_ (
);

NAND2X1 _1636_ (
    .A(_803_),
    .B(_804_),
    .Y(_805_)
);

AND2X2 _1216_ (
    .A(_437_),
    .B(_436_),
    .Y(_442_)
);

FILL FILL_0__964_ (
);

NAND2X1 _967_ (
    .A(Stg_0_bF$buf4),
    .B(Xin12b[4]),
    .Y(_203_)
);

FILL FILL_1__1378_ (
);

FILL FILL_2__1447_ (
);

FILL FILL_2__1027_ (
);

NAND2X1 _1445_ (
    .A(Yin[1]),
    .B(_625_),
    .Y(_643_)
);

NAND2X1 _1025_ (
    .A(Stg_0_bF$buf2),
    .B(Yin1[0]),
    .Y(_259_)
);

FILL FILL_1__1187_ (
);

FILL FILL_1__980_ (
);

NOR2X1 _1674_ (
    .A(_840_),
    .B(_837_),
    .Y(_841_)
);

OAI21X1 _1254_ (
    .A(_477_),
    .B(_455_),
    .C(_474_),
    .Y(_478_)
);

FILL FILL_0__1714_ (
);

NAND2X1 _1483_ (
    .A(Ain[1]),
    .B(_635_),
    .Y(_663_)
);

OAI21X1 _1063_ (
    .A(_269_),
    .B(_249_),
    .C(_201__bF$buf3),
    .Y(_296_)
);

FILL FILL_0__1523_ (
);

FILL FILL_0__1103_ (
);

FILL FILL_2__1294_ (
);

NAND3X1 _1539_ (
    .A(_678_),
    .B(_199_),
    .C(_224_),
    .Y(_712_)
);

NAND2X1 _1119_ (
    .A(_348_),
    .B(_331_),
    .Y(_350_)
);

FILL FILL_0__867_ (
);

NOR2X1 _1292_ (
    .A(_512_),
    .B(_505_),
    .Y(_513_)
);

FILL FILL_0__1332_ (
);

DFFPOSX1 _1768_ (
    .D(_40_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[8])
);

AND2X2 _1348_ (
    .A(_563_),
    .B(_201__bF$buf0),
    .Y(_565_)
);

FILL FILL_0__1808_ (
);

FILL FILL_1__883_ (
);

FILL FILL_0__1561_ (
);

FILL FILL_0__1141_ (
);

FILL FILL_1__1722_ (
);

FILL FILL_1__1302_ (
);

OAI21X1 _1577_ (
    .A(_748_),
    .B(_747_),
    .C(Yin12b[4]),
    .Y(_749_)
);

AOI21X1 _1157_ (
    .A(_384_),
    .B(_366_),
    .C(_385_),
    .Y(_386_)
);

FILL FILL_1__939_ (
);

FILL FILL_0__1617_ (
);

FILL FILL_0__1370_ (
);

FILL FILL_2__1388_ (
);

FILL FILL_1__1531_ (
);

FILL FILL_1__1111_ (
);

INVX1 _1386_ (
    .A(_599_),
    .Y(_601_)
);

FILL FILL_2__1600_ (
);

FILL FILL_0__1426_ (
);

FILL FILL_0__1006_ (
);

FILL FILL_2__955_ (
);

FILL FILL_1__1340_ (
);

INVX1 _1195_ (
    .A(Xin12b[8]),
    .Y(_422_)
);

FILL FILL_1__977_ (
);

FILL FILL_0__1655_ (
);

FILL FILL_0__1235_ (
);

FILL FILL_0__999_ (
);

FILL FILL_0__1464_ (
);

FILL FILL_0__1044_ (
);

FILL FILL_1__1625_ (
);

FILL FILL_1__1205_ (
);

FILL FILL_0__1693_ (
);

FILL FILL_0__1273_ (
);

FILL FILL_1__1434_ (
);

FILL FILL_1__1014_ (
);

OR2X2 _1289_ (
    .A(_508_),
    .B(Ain1[0]),
    .Y(_510_)
);

FILL FILL_0__1329_ (
);

FILL FILL_0__1082_ (
);

MUX2X1 _1501_ (
    .A(Xin12b[9]),
    .B(Xin12b[8]),
    .S(Stg_0_bF$buf3),
    .Y(_675_)
);

FILL FILL_1__1663_ (
);

FILL FILL_1__1243_ (
);

AOI21X1 _1098_ (
    .A(_328_),
    .B(_329_),
    .C(_192_),
    .Y(_330_)
);

FILL FILL_0__1558_ (
);

FILL FILL_0__1138_ (
);

FILL FILL_1__1719_ (
);

FILL FILL88350x61350 (
);

DFFPOSX1 _1730_ (
    .D(_2_),
    .CLK(clk_bF$buf7),
    .Q(Xcalc[0])
);

NAND2X1 _1310_ (
    .A(Acalc[3]),
    .B(_188__bF$buf0),
    .Y(_530_)
);

FILL FILL_1__1472_ (
);

FILL FILL_1__1052_ (
);

FILL FILL_2__1541_ (
);

FILL FILL_2__1121_ (
);

FILL FILL_0__1367_ (
);

FILL FILL_1__1528_ (
);

FILL FILL_1__1108_ (
);

FILL FILL_1__901_ (
);

NAND2X1 _870_ (
    .A(LoadCtl[3]),
    .B(_112_),
    .Y(_113_)
);

FILL FILL_1__1281_ (
);

FILL FILL_0__1596_ (
);

FILL FILL_0__1176_ (
);

FILL FILL_0__923_ (
);

INVX1 _926_ (
    .A(Yin0[0]),
    .Y(_163_)
);

FILL FILL_1__1337_ (
);

FILL FILL_1__1090_ (
);

NAND2X1 _1404_ (
    .A(Ain12b_11_bF$buf2),
    .B(_616_),
    .Y(_617_)
);

FILL FILL_1__1566_ (
);

FILL FILL_1__1146_ (
);

FILL FILL87450x86550 (
);

NAND3X1 _1633_ (
    .A(_201__bF$buf5),
    .B(_801_),
    .C(_799_),
    .Y(_802_)
);

OR2X2 _1213_ (
    .A(_437_),
    .B(_436_),
    .Y(_439_)
);

FILL FILL_0__961_ (
);

INVX1 _964_ (
    .A(Yin0[1]),
    .Y(_200_)
);

FILL FILL_1__1375_ (
);

FILL FILL_2__1444_ (
);

FILL FILL_2__1024_ (
);

OAI21X1 _1442_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_205_),
    .C(_641_),
    .Y(_37_)
);

INVX1 _1022_ (
    .A(Yin1[1]),
    .Y(_256_)
);

FILL FILL_1__1184_ (
);

FILL FILL_0__1499_ (
);

FILL FILL_0__1079_ (
);

OR2X2 _1671_ (
    .A(_837_),
    .B(_838_),
    .Y(_839_)
);

INVX1 _1251_ (
    .A(_474_),
    .Y(_475_)
);

FILL FILL_0__1711_ (
);

NAND2X1 _1727_ (
    .A(_95_),
    .B(_105_),
    .Y(_72_)
);

INVX1 _1307_ (
    .A(_523_),
    .Y(_527_)
);

FILL FILL_1__1469_ (
);

FILL FILL_1__1049_ (
);

AOI21X1 _1480_ (
    .A(_660_),
    .B(_632_),
    .C(_661_),
    .Y(_55_)
);

NAND2X1 _1060_ (
    .A(_236_),
    .B(_292_),
    .Y(_293_)
);

FILL FILL_0__1520_ (
);

FILL FILL_0__1100_ (
);

FILL FILL_2__1291_ (
);

INVX2 _1536_ (
    .A(_707_),
    .Y(_709_)
);

AND2X2 _1116_ (
    .A(_343_),
    .B(_346_),
    .Y(_347_)
);

FILL FILL_0__864_ (
);

INVX1 _867_ (
    .A(Acalc[6]),
    .Y(_110_)
);

FILL FILL88650x36150 (
);

FILL FILL_1__1698_ (
);

FILL FILL_1__1278_ (
);

FILL FILL_2__1347_ (
);

DFFPOSX1 _1765_ (
    .D(_37_),
    .CLK(clk_bF$buf5),
    .Q(Xin0[1])
);

AOI21X1 _1345_ (
    .A(_539_),
    .B(_560_),
    .C(_561_),
    .Y(_562_)
);

FILL FILL_1__1087_ (
);

FILL FILL_1__880_ (
);

NAND3X1 _1574_ (
    .A(_244_),
    .B(_742_),
    .C(_745_),
    .Y(_746_)
);

NAND3X1 _1154_ (
    .A(_363_),
    .B(_366_),
    .C(_347_),
    .Y(_383_)
);

FILL FILL_1__936_ (
);

FILL FILL_0__1614_ (
);

FILL FILL_0__958_ (
);

NAND2X1 _1383_ (
    .A(_596_),
    .B(_560_),
    .Y(_598_)
);

FILL FILL_0__1423_ (
);

FILL FILL_0__1003_ (
);

FILL FILL_2__952_ (
);

FILL FILL_2__1194_ (
);

NAND2X1 _1439_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[0]),
    .Y(_640_)
);

OAI21X1 _1019_ (
    .A(_253_),
    .B(_250_),
    .C(_233_),
    .Y(_2_)
);

OAI21X1 _1192_ (
    .A(_401_),
    .B(_394_),
    .C(_201__bF$buf4),
    .Y(_419_)
);

FILL FILL_1__974_ (
);

FILL FILL_0__1652_ (
);

FILL FILL_0__1232_ (
);

FILL FILL_1__1813_ (
);

AND2X2 _1668_ (
    .A(_832_),
    .B(_835_),
    .Y(_836_)
);

NAND2X1 _1248_ (
    .A(Yin12b[11]),
    .B(_471_),
    .Y(_472_)
);

FILL FILL_0__996_ (
);

INVX1 _999_ (
    .A(Yin1[0]),
    .Y(_234_)
);

FILL FILL_0__1708_ (
);

FILL FILL_0__1461_ (
);

FILL FILL_0__1041_ (
);

FILL FILL_1__1622_ (
);

FILL FILL_1__1202_ (
);

OAI21X1 _1477_ (
    .A(_568_),
    .B(_632_),
    .C(_659_),
    .Y(_54_)
);

INVX1 _1057_ (
    .A(_289_),
    .Y(_290_)
);

FILL FILL_0__1517_ (
);

FILL FILL_0__1690_ (
);

FILL FILL_2__1288_ (
);

FILL FILL_0__1270_ (
);

FILL FILL_1__1431_ (
);

FILL FILL_1__1011_ (
);

NAND3X1 _1286_ (
    .A(Stg_2_bF$buf0),
    .B(_484_),
    .C(_506_),
    .Y(_507_)
);

FILL FILL_2__1500_ (
);

FILL FILL_0__1326_ (
);

FILL FILL_1_BUFX2_insert30 (
);

FILL FILL_1_BUFX2_insert31 (
);

FILL FILL_1_BUFX2_insert32 (
);

FILL FILL_1_BUFX2_insert33 (
);

FILL FILL_1_BUFX2_insert34 (
);

FILL FILL_1_BUFX2_insert35 (
);

FILL FILL_1_BUFX2_insert36 (
);

FILL FILL_1_BUFX2_insert37 (
);

FILL FILL_1_BUFX2_insert38 (
);

FILL FILL_1_BUFX2_insert39 (
);

FILL FILL_0_CLKBUF1_insert12 (
);

FILL FILL_0_CLKBUF1_insert13 (
);

FILL FILL_0_CLKBUF1_insert14 (
);

FILL FILL_0_CLKBUF1_insert15 (
);

FILL FILL_0_CLKBUF1_insert16 (
);

FILL FILL_0_CLKBUF1_insert17 (
);

FILL FILL_0_CLKBUF1_insert18 (
);

FILL FILL_0_CLKBUF1_insert19 (
);

FILL FILL_1__1660_ (
);

FILL FILL_1__1240_ (
);

NAND2X1 _1095_ (
    .A(_326_),
    .B(_325_),
    .Y(_327_)
);

FILL FILL_1__877_ (
);

FILL FILL_0__1555_ (
);

FILL FILL_0__1135_ (
);

FILL FILL_1__1716_ (
);

FILL FILL_0__899_ (
);

FILL FILL88350x82950 (
);

FILL FILL_0__1364_ (
);

FILL FILL_1__1525_ (
);

FILL FILL_1__1105_ (
);

FILL FILL87150x64950 (
);

FILL FILL_2__949_ (
);

FILL FILL_0__1593_ (
);

FILL FILL_0__1173_ (
);

FILL FILL_0__920_ (
);

AOI22X1 _923_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Xcalc[1]),
    .C(_119_),
    .D(Xcalc[3]),
    .Y(_161_)
);

FILL FILL_1__1334_ (
);

OAI21X1 _1189_ (
    .A(Stg_2_bF$buf4),
    .B(_414_),
    .C(_415_),
    .Y(_416_)
);

FILL FILL_0__1649_ (
);

FILL FILL_0__1229_ (
);

INVX1 _1401_ (
    .A(_613_),
    .Y(_614_)
);

FILL FILL_1__1563_ (
);

FILL FILL_1__1143_ (
);

FILL FILL_0__1458_ (
);

FILL FILL_0__1038_ (
);

FILL FILL_1__1619_ (
);

NAND2X1 _1630_ (
    .A(_780_),
    .B(_779_),
    .Y(_799_)
);

AOI21X1 _1210_ (
    .A(_435_),
    .B(_183__bF$buf2),
    .C(_395_),
    .Y(_436_)
);

MUX2X1 _961_ (
    .A(Xin12b[5]),
    .B(Xin12b[4]),
    .S(Stg_0_bF$buf4),
    .Y(_197_)
);

FILL FILL_1__1372_ (
);

FILL FILL_2__1441_ (
);

FILL FILL_2__1021_ (
);

FILL FILL_0__1687_ (
);

FILL FILL_0__1267_ (
);

FILL FILL_1__1428_ (
);

FILL FILL_1__1008_ (
);

FILL FILL_1__1181_ (
);

FILL FILL_0__1496_ (
);

FILL FILL_0__1076_ (
);

FILL FILL_1_BUFX2_insert0 (
);

FILL FILL_1_BUFX2_insert1 (
);

FILL FILL_1_BUFX2_insert2 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert4 (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

FILL FILL_1__1657_ (
);

FILL FILL_1__1237_ (
);

AOI21X1 _1724_ (
    .A(_92_),
    .B(_87_),
    .C(_96_),
    .Y(_103_)
);

NAND2X1 _1304_ (
    .A(_518_),
    .B(_522_),
    .Y(_524_)
);

FILL FILL_1__1466_ (
);

FILL FILL_1__1046_ (
);

OAI21X1 _1533_ (
    .A(Stg_1_bF$buf1),
    .B(_574_),
    .C(LoadCtl_6_bF$buf3),
    .Y(_707_)
);

OAI21X1 _1113_ (
    .A(_322_),
    .B(_310_),
    .C(_201__bF$buf0),
    .Y(_344_)
);

NAND2X1 _864_ (
    .A(LoadCtl[4]),
    .B(Acalc[8]),
    .Y(_107_)
);

FILL FILL_1__1695_ (
);

FILL FILL_1__1275_ (
);

FILL FILL_2__1344_ (
);

FILL FILL_0__917_ (
);

FILL FILL88650x57750 (
);

DFFPOSX1 _1762_ (
    .D(_34_),
    .CLK(clk_bF$buf2),
    .Q(Xin1[0])
);

OAI21X1 _1342_ (
    .A(_557_),
    .B(_559_),
    .C(_544_),
    .Y(_19_)
);

FILL FILL_1__1084_ (
);

FILL FILL87450x39750 (
);

FILL FILL_0__1399_ (
);

NOR2X1 _1571_ (
    .A(_719_),
    .B(_712_),
    .Y(_743_)
);

NAND2X1 _1151_ (
    .A(Xin12b[6]),
    .B(_379_),
    .Y(_380_)
);

FILL FILL_1__933_ (
);

FILL FILL_0__1611_ (
);

AOI21X1 _1627_ (
    .A(_794_),
    .B(_766_),
    .C(_795_),
    .Y(_796_)
);

INVX1 _1207_ (
    .A(Xcalc[9]),
    .Y(_433_)
);

FILL FILL_0__955_ (
);

MUX2X1 _958_ (
    .A(Xin0[1]),
    .B(Xin0[0]),
    .S(Stg_0_bF$buf6),
    .Y(_194_)
);

FILL FILL_1__1369_ (
);

OR2X2 _1380_ (
    .A(_570_),
    .B(_582_),
    .Y(_595_)
);

FILL FILL_2__1438_ (
);

FILL FILL_0__1420_ (
);

FILL FILL_2__1018_ (
);

FILL FILL_0__1000_ (
);

FILL FILL_2__1191_ (
);

OAI21X1 _1436_ (
    .A(_165_),
    .B(_119_),
    .C(_638_),
    .Y(_34_)
);

INVX1 _1016_ (
    .A(_247_),
    .Y(_251_)
);

FILL FILL_1__1598_ (
);

FILL FILL_1__1178_ (
);

FILL FILL_1__971_ (
);

FILL FILL_2__1667_ (
);

FILL FILL_2__1247_ (
);

FILL FILL_1__1810_ (
);

OAI21X1 _1665_ (
    .A(_803_),
    .B(_799_),
    .C(_201__bF$buf5),
    .Y(_833_)
);

NAND2X1 _1245_ (
    .A(_466_),
    .B(_469_),
    .Y(_470_)
);

FILL FILL_0__993_ (
);

AOI21X1 _996_ (
    .A(_231_),
    .B(_230_),
    .C(_192_),
    .Y(_232_)
);

FILL FILL_0__1705_ (
);

NAND2X1 _1474_ (
    .A(Ain[1]),
    .B(_629_),
    .Y(_658_)
);

NAND2X1 _1054_ (
    .A(_164__bF$buf4),
    .B(_243_),
    .Y(_287_)
);

FILL FILL_0__1514_ (
);

FILL FILL_2__1285_ (
);

INVX1 _1283_ (
    .A(Ain0[1]),
    .Y(_504_)
);

FILL FILL_0__1323_ (
);

FILL FILL_2__1094_ (
);

DFFPOSX1 _1759_ (
    .D(_31_),
    .CLK(clk_bF$buf6),
    .Q(Xin12b[7])
);

NOR2X1 _1339_ (
    .A(_556_),
    .B(_545_),
    .Y(_557_)
);

AOI21X1 _1092_ (
    .A(_323_),
    .B(_320_),
    .C(_202_),
    .Y(_324_)
);

FILL FILL_1__874_ (
);

FILL FILL_2__908_ (
);

FILL FILL_0__1552_ (
);

FILL FILL_0__1132_ (
);

FILL FILL_1__1713_ (
);

NAND2X1 _1568_ (
    .A(Stg_2_bF$buf3),
    .B(_739_),
    .Y(_740_)
);

NAND3X1 _1148_ (
    .A(_201__bF$buf1),
    .B(_376_),
    .C(_372_),
    .Y(_377_)
);

FILL FILL_0__896_ (
);

NAND2X1 _899_ (
    .A(Ycalc[11]),
    .B(_137_),
    .Y(_139_)
);

FILL FILL_0__1608_ (
);

FILL FILL_0__1361_ (
);

FILL FILL_1__1522_ (
);

FILL FILL_1__1102_ (
);

FILL FILL_2_BUFX2_insert50 (
);

FILL FILL_2_BUFX2_insert53 (
);

FILL FILL_2_BUFX2_insert56 (
);

FILL FILL_2_BUFX2_insert58 (
);

DFFPOSX1 _1797_ (
    .D(_62_),
    .CLK(clk_bF$buf3),
    .Q(_860_)
);

NAND2X1 _1377_ (
    .A(_591_),
    .B(_589_),
    .Y(_592_)
);

FILL FILL_0__1417_ (
);

FILL FILL_0__1590_ (
);

FILL FILL_0__1170_ (
);

FILL FILL_2__1188_ (
);

INVX1 _920_ (
    .A(Xcalc[5]),
    .Y(_158_)
);

FILL FILL_1__1331_ (
);

NAND3X1 _1186_ (
    .A(_376_),
    .B(_396_),
    .C(_371_),
    .Y(_413_)
);

FILL FILL_1__968_ (
);

FILL FILL_2__1400_ (
);

FILL FILL_0__1646_ (
);

FILL FILL_0__1226_ (
);

FILL FILL_1__1560_ (
);

FILL FILL_1__1140_ (
);

FILL FILL_0__1455_ (
);

FILL FILL_0__1035_ (
);

FILL FILL_1__1616_ (
);

FILL FILL_0__1684_ (
);

FILL FILL_0__1264_ (
);

FILL FILL_1__1425_ (
);

FILL FILL_1__1005_ (
);

FILL FILL_0__1493_ (
);

FILL FILL_0__1073_ (
);

FILL FILL_1__1654_ (
);

FILL FILL_1__1234_ (
);

INVX1 _1089_ (
    .A(_310_),
    .Y(_321_)
);

FILL FILL_0__1549_ (
);

FILL FILL_0__1129_ (
);

NAND2X1 _1721_ (
    .A(_98_),
    .B(_99_),
    .Y(_100_)
);

OAI21X1 _1301_ (
    .A(Stg_2_bF$buf0),
    .B(Stg_1_bF$buf1),
    .C(Ain12b_11_bF$buf4),
    .Y(_521_)
);

FILL FILL_1__1463_ (
);

FILL FILL_1__1043_ (
);

FILL FILL_0__1358_ (
);

FILL FILL_1__1519_ (
);

INVX1 _1530_ (
    .A(_703_),
    .Y(_704_)
);

INVX1 _1110_ (
    .A(_340_),
    .Y(_341_)
);

FILL FILL_1__1692_ (
);

FILL FILL_1__1272_ (
);

FILL FILL_2__1341_ (
);

FILL FILL_0__1587_ (
);

FILL FILL_0__1167_ (
);

FILL FILL_0__914_ (
);

NAND2X1 _917_ (
    .A(LoadCtl[4]),
    .B(Xcalc[9]),
    .Y(_155_)
);

FILL FILL_1__1328_ (
);

FILL FILL_1__1081_ (
);

FILL FILL_0__1396_ (
);

BUFX2 _1815_ (
    .A(_862_[1]),
    .Y(Yout[1])
);

FILL FILL_1__1557_ (
);

FILL FILL_1__1137_ (
);

FILL FILL_1__930_ (
);

NAND3X1 _1624_ (
    .A(_768_),
    .B(_766_),
    .C(_792_),
    .Y(_793_)
);

INVX1 _1204_ (
    .A(_430_),
    .Y(_431_)
);

FILL FILL_0__952_ (
);

NAND2X1 _955_ (
    .A(_183__bF$buf3),
    .B(_190_),
    .Y(_191_)
);

FILL FILL_1__1366_ (
);

NAND2X1 _1433_ (
    .A(Xin[1]),
    .B(_635_),
    .Y(_637_)
);

NAND2X1 _1013_ (
    .A(Stg_2_bF$buf2),
    .B(_247_),
    .Y(_248_)
);

FILL FILL_1__1595_ (
);

FILL FILL_1__1175_ (
);

FILL FILL_2__1664_ (
);

FILL FILL_2__1244_ (
);

INVX1 _1662_ (
    .A(_829_),
    .Y(_830_)
);

INVX1 _1242_ (
    .A(_462_),
    .Y(_467_)
);

FILL FILL_0__990_ (
);

AND2X2 _993_ (
    .A(_227_),
    .B(_228_),
    .Y(_229_)
);

FILL FILL_0__1702_ (
);

FILL FILL_0__1299_ (
);

OAI21X1 _1718_ (
    .A(_858_),
    .B(_76_),
    .C(_201__bF$buf2),
    .Y(_97_)
);

OAI21X1 _1471_ (
    .A(_201__bF$buf1),
    .B(_625_),
    .C(_656_),
    .Y(_51_)
);

INVX1 _1051_ (
    .A(Yin12b[9]),
    .Y(_284_)
);

FILL FILL_0__1511_ (
);

FILL FILL88650x43350 (
);

INVX1 _1527_ (
    .A(_700_),
    .Y(_701_)
);

OAI21X1 _1107_ (
    .A(Stg_2_bF$buf4),
    .B(_247_),
    .C(_337_),
    .Y(_338_)
);

FILL FILL_1__1689_ (
);

FILL FILL_1__1269_ (
);

NAND2X1 _1280_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_501_),
    .Y(_502_)
);

FILL FILL_2__1338_ (
);

FILL FILL_0__1320_ (
);

FILL FILL_2__1091_ (
);

DFFPOSX1 _1756_ (
    .D(_28_),
    .CLK(clk_bF$buf4),
    .Q(Xin12b[8])
);

OAI21X1 _1336_ (
    .A(_549_),
    .B(_547_),
    .C(_553_),
    .Y(_554_)
);

FILL FILL_1__1498_ (
);

FILL FILL_1__1078_ (
);

FILL FILL_1__871_ (
);

FILL FILL_2__905_ (
);

FILL FILL_1__1710_ (
);

OAI21X1 _1565_ (
    .A(Stg_0_bF$buf5),
    .B(_458_),
    .C(_736_),
    .Y(_737_)
);

NAND2X1 _1145_ (
    .A(_183__bF$buf1),
    .B(_288_),
    .Y(_374_)
);

FILL FILL_0__893_ (
);

FILL FILL_1__927_ (
);

OAI21X1 _896_ (
    .A(_117_),
    .B(_135_),
    .C(_136_),
    .Y(_862_[0])
);

FILL FILL_0__1605_ (
);

FILL FILL_0__949_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_2_BUFX2_insert22 (
);

FILL FILL_2_BUFX2_insert25 (
);

FILL FILL_2_BUFX2_insert28 (
);

DFFPOSX1 _1794_ (
    .D(LoadCtl[3]),
    .CLK(clk_bF$buf7),
    .Q(LoadCtl[4])
);

NAND2X1 _1374_ (
    .A(Ain12b[8]),
    .B(_588_),
    .Y(_589_)
);

FILL FILL_0__1414_ (
);

FILL FILL_2__1185_ (
);

AND2X2 _1183_ (
    .A(_409_),
    .B(_400_),
    .Y(_410_)
);

FILL FILL_1__965_ (
);

FILL FILL_0__1643_ (
);

FILL FILL_0__1223_ (
);

OAI21X1 _1659_ (
    .A(Stg_2_bF$buf3),
    .B(_825_),
    .C(_826_),
    .Y(_827_)
);

NAND3X1 _1239_ (
    .A(_440_),
    .B(_444_),
    .C(_426_),
    .Y(_464_)
);

FILL FILL_0__987_ (
);

FILL FILL_0__1452_ (
);

FILL FILL_0__1032_ (
);

FILL FILL_1__1613_ (
);

NAND2X1 _1468_ (
    .A(Ain[0]),
    .B(_625_),
    .Y(_655_)
);

NAND2X1 _1048_ (
    .A(Xcalc[2]),
    .B(_188__bF$buf4),
    .Y(_281_)
);

FILL FILL_0__1508_ (
);

FILL FILL_0__1681_ (
);

FILL FILL_0__1261_ (
);

FILL FILL_1__1422_ (
);

FILL FILL_1__1002_ (
);

AOI21X1 _1697_ (
    .A(_76_),
    .B(_201__bF$buf2),
    .C(_858_),
    .Y(_77_)
);

NAND2X1 _1277_ (
    .A(_498_),
    .B(_497_),
    .Y(_499_)
);

FILL FILL_0__1317_ (
);

FILL FILL_0__1490_ (
);

FILL FILL_0__1070_ (
);

FILL FILL_2__1088_ (
);

FILL FILL_1__1651_ (
);

FILL FILL_1__1231_ (
);

NAND2X1 _1086_ (
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

FILL FILL_1__868_ (
);

FILL FILL_0__1546_ (
);

FILL FILL_0__1126_ (
);

FILL FILL_1__1707_ (
);

FILL FILL_1__1460_ (
);

FILL FILL_1__1040_ (
);

FILL FILL_0__1355_ (
);

FILL FILL_1__1516_ (
);

FILL FILL_0__1584_ (
);

FILL FILL_0__1164_ (
);

FILL FILL_0__911_ (
);

AOI22X1 _914_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Xcalc[0]),
    .C(_119_),
    .D(Xcalc[2]),
    .Y(_153_)
);

FILL FILL_1__1325_ (
);

FILL FILL_0__1393_ (
);

BUFX2 _1812_ (
    .A(_861_[0]),
    .Y(Xout[0])
);

FILL FILL_1__1554_ (
);

FILL FILL_1__1134_ (
);

FILL FILL_0__1449_ (
);

FILL FILL_0__1029_ (
);

AOI22X1 _1621_ (
    .A(_132_),
    .B(_188__bF$buf2),
    .C(_790_),
    .D(_709_),
    .Y(_67_)
);

INVX1 _1201_ (
    .A(_427_),
    .Y(_428_)
);

INVX8 _952_ (
    .A(LoadCtl_6_bF$buf4),
    .Y(_188_)
);

FILL FILL_1__1363_ (
);

FILL FILL_0__1678_ (
);

FILL FILL_0__1258_ (
);

FILL FILL_1__1419_ (
);

NOR2X1 _1430_ (
    .A(_112_),
    .B(_117_),
    .Y(_635_)
);

NAND2X1 _1010_ (
    .A(Stg_0_bF$buf2),
    .B(Yin12b[5]),
    .Y(_245_)
);

FILL FILL88350x21750 (
);

FILL FILL_1__1592_ (
);

FILL FILL_1__1172_ (
);

FILL FILL_2__1661_ (
);

FILL FILL_2__1241_ (
);

FILL FILL_0__1487_ (
);

FILL FILL_0__1067_ (
);

FILL FILL_1__1648_ (
);

FILL FILL_1__1228_ (
);

AOI21X1 _990_ (
    .A(_225_),
    .B(_217_),
    .C(_200_),
    .Y(_226_)
);

FILL FILL_2__1717_ (
);

FILL FILL_0__1296_ (
);

AOI22X1 _1715_ (
    .A(_129_),
    .B(_188__bF$buf2),
    .C(_94_),
    .D(_709_),
    .Y(_71_)
);

FILL FILL_1__1457_ (
);

FILL FILL_1__1037_ (
);

OAI21X1 _1524_ (
    .A(Ain12b_11_bF$buf4),
    .B(_696_),
    .C(_697_),
    .Y(_698_)
);

NAND2X1 _1104_ (
    .A(Stg_1_bF$buf3),
    .B(_334_),
    .Y(_335_)
);

FILL FILL_1__1686_ (
);

FILL FILL_1__1266_ (
);

FILL FILL88650x64950 (
);

FILL FILL_0__908_ (
);

FILL FILL87450x46950 (
);

DFFPOSX1 _1753_ (
    .D(_25_),
    .CLK(clk_bF$buf7),
    .Q(Acalc[11])
);

AND2X2 _1333_ (
    .A(_550_),
    .B(Ain12b[5]),
    .Y(_551_)
);

FILL FILL_1__1495_ (
);

FILL FILL_1__1075_ (
);

FILL FILL_2__902_ (
);

FILL FILL_2__1564_ (
);

FILL FILL_2__1144_ (
);

BUFX2 _1809_ (
    .A(_859_[1]),
    .Y(Aout[1])
);

AOI22X1 _1562_ (
    .A(_708_),
    .B(_188__bF$buf2),
    .C(_734_),
    .D(_709_),
    .Y(_64_)
);

NOR3X1 _1142_ (
    .A(_338_),
    .B(_359_),
    .C(_332_),
    .Y(_371_)
);

FILL FILL_0__890_ (
);

FILL FILL_1__924_ (
);

OAI22X1 _893_ (
    .A(_112_),
    .B(_133_),
    .C(_132_),
    .D(_113_),
    .Y(_134_)
);

FILL FILL_0__1602_ (
);

FILL FILL_0__1199_ (
);

OAI21X1 _1618_ (
    .A(_787_),
    .B(_755_),
    .C(_766_),
    .Y(_788_)
);

FILL FILL_0__946_ (
);

INVX2 _949_ (
    .A(_185_),
    .Y(_186_)
);

DFFPOSX1 _1791_ (
    .D(LoadCtl_0_bF$buf0),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[1])
);

NAND2X1 _1371_ (
    .A(_201__bF$buf3),
    .B(_292_),
    .Y(_586_)
);

FILL FILL_0__1411_ (
);

OAI21X1 _1427_ (
    .A(_172_),
    .B(_632_),
    .C(_633_),
    .Y(_30_)
);

NAND2X1 _1007_ (
    .A(Stg_0_bF$buf0),
    .B(Yin12b[7]),
    .Y(_242_)
);

FILL FILL_1__1589_ (
);

FILL FILL_1__1169_ (
);

AOI22X1 _1180_ (
    .A(_157_),
    .B(_188__bF$buf3),
    .C(_406_),
    .D(_407_),
    .Y(_9_)
);

FILL FILL_1__962_ (
);

FILL FILL_2__1658_ (
);

FILL FILL_0__1640_ (
);

FILL FILL_0__1220_ (
);

FILL FILL_2__1238_ (
);

NAND3X1 _1656_ (
    .A(_780_),
    .B(_801_),
    .C(_779_),
    .Y(_824_)
);

OAI21X1 _1236_ (
    .A(_459_),
    .B(_460_),
    .C(_458_),
    .Y(_461_)
);

FILL FILL_0__984_ (
);

MUX2X1 _987_ (
    .A(_222_),
    .B(_221_),
    .S(_164__bF$buf4),
    .Y(_223_)
);

FILL FILL_1__1398_ (
);

FILL FILL_1__1610_ (
);

OAI21X1 _1465_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_163_),
    .C(_653_),
    .Y(_48_)
);

OAI21X1 _1045_ (
    .A(_273_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

FILL FILL_0__1505_ (
);

OAI21X1 _1694_ (
    .A(_843_),
    .B(_847_),
    .C(_201__bF$buf2),
    .Y(_74_)
);

OAI21X1 _1274_ (
    .A(Ain12b_11_bF$buf2),
    .B(_494_),
    .C(_495_),
    .Y(_496_)
);

FILL FILL_0__1314_ (
);

FILL FILL_2__1085_ (
);

OAI21X1 _1083_ (
    .A(_164__bF$buf3),
    .B(_313_),
    .C(_314_),
    .Y(_315_)
);

FILL FILL_1__865_ (
);

FILL FILL_0__1543_ (
);

FILL FILL_0__1123_ (
);

FILL FILL_1__1704_ (
);

FILL FILL87750x54150 (
);

NAND2X1 _1559_ (
    .A(_729_),
    .B(_731_),
    .Y(_732_)
);

AND2X2 _1139_ (
    .A(_352_),
    .B(_368_),
    .Y(_369_)
);

FILL FILL_0__887_ (
);

FILL FILL_0__1352_ (
);

FILL FILL_1__1513_ (
);

DFFPOSX1 _1788_ (
    .D(_60_),
    .CLK(clk_bF$buf0),
    .Q(Ain0[0])
);

AOI21X1 _1368_ (
    .A(_573_),
    .B(_582_),
    .C(_188__bF$buf3),
    .Y(_584_)
);

FILL FILL_0__1408_ (
);

FILL FILL_0__1581_ (
);

FILL FILL_0__1161_ (
);

INVX1 _911_ (
    .A(Xcalc[4]),
    .Y(_150_)
);

FILL FILL_1__1322_ (
);

OAI21X1 _1597_ (
    .A(_763_),
    .B(_767_),
    .C(Yin12b[5]),
    .Y(_768_)
);

AND2X2 _1177_ (
    .A(_400_),
    .B(_404_),
    .Y(_405_)
);

FILL FILL_1__959_ (
);

FILL FILL_2__1811_ (
);

FILL FILL_0__1637_ (
);

FILL FILL_0__1217_ (
);

FILL FILL_0__1390_ (
);

FILL FILL_1__1551_ (
);

FILL FILL_1__1131_ (
);

FILL FILL_0__1446_ (
);

FILL FILL_0__1026_ (
);

FILL FILL_1__1607_ (
);

FILL FILL_1__1360_ (
);

FILL FILL_1__997_ (
);

FILL FILL_0__1675_ (
);

FILL FILL_0__1255_ (
);

FILL FILL_1__1416_ (
);

FILL FILL_0__1484_ (
);

FILL FILL_0__1064_ (
);

FILL FILL_1__1645_ (
);

FILL FILL_1__1225_ (
);

FILL FILL_2__1714_ (
);

FILL FILL_0__1293_ (
);

OAI21X1 _1712_ (
    .A(_91_),
    .B(_90_),
    .C(_84_),
    .Y(_92_)
);

FILL FILL_1__1454_ (
);

FILL FILL_1__1034_ (
);

FILL FILL88050x54150 (
);

FILL FILL_0__1349_ (
);

NAND3X1 _1521_ (
    .A(Stg_2_bF$buf1),
    .B(_693_),
    .C(_694_),
    .Y(_695_)
);

NAND3X1 _1101_ (
    .A(_295_),
    .B(_319_),
    .C(_298_),
    .Y(_332_)
);

FILL FILL_1__1683_ (
);

FILL FILL_1__1263_ (
);

FILL FILL_0__1578_ (
);

FILL FILL_0__1158_ (
);

FILL FILL_0__905_ (
);

NAND2X1 _908_ (
    .A(LoadCtl[4]),
    .B(Xcalc[8]),
    .Y(_147_)
);

FILL FILL_1__1319_ (
);

DFFPOSX1 _1750_ (
    .D(_22_),
    .CLK(clk_bF$buf7),
    .Q(Acalc[8])
);

OAI21X1 _1330_ (
    .A(Stg_0_bF$buf1),
    .B(Stg_1_bF$buf2),
    .C(_184_),
    .Y(_548_)
);

FILL FILL_1__1492_ (
);

FILL FILL_1__1072_ (
);

FILL FILL_2__1808_ (
);

FILL FILL_2__1561_ (
);

FILL FILL_2__1141_ (
);

FILL FILL_0__1387_ (
);

DFFPOSX1 _1806_ (
    .D(_71_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[10])
);

FILL FILL_1__1548_ (
);

FILL FILL_1__1128_ (
);

FILL FILL_1__921_ (
);

OAI21X1 _890_ (
    .A(LoadCtl[4]),
    .B(_129_),
    .C(_130_),
    .Y(_131_)
);

FILL FILL_2__1617_ (
);

FILL FILL_0__1196_ (
);

NAND3X1 _1615_ (
    .A(Yin12b[6]),
    .B(_783_),
    .C(_784_),
    .Y(_785_)
);

FILL FILL_0__943_ (
);

INVX4 _946_ (
    .A(Stg_2_bF$buf3),
    .Y(_183_)
);

FILL FILL_1__1357_ (
);

OAI21X1 _1424_ (
    .A(_441_),
    .B(_629_),
    .C(_631_),
    .Y(_29_)
);

MUX2X1 _1004_ (
    .A(_238_),
    .B(_236_),
    .S(_164__bF$buf1),
    .Y(_239_)
);

FILL FILL_1__1586_ (
);

FILL FILL_1__1166_ (
);

FILL FILL_2__1655_ (
);

FILL FILL_2__1235_ (
);

NAND3X1 _1653_ (
    .A(Yin12b[7]),
    .B(_802_),
    .C(_805_),
    .Y(_821_)
);

INVX1 _1233_ (
    .A(Xin12b[10]),
    .Y(_458_)
);

FILL FILL_0__981_ (
);

MUX2X1 _984_ (
    .A(_219_),
    .B(_218_),
    .S(_164__bF$buf2),
    .Y(_220_)
);

FILL FILL_1__1395_ (
);

FILL FILL_2__1464_ (
);

NOR3X1 _1709_ (
    .A(_786_),
    .B(_806_),
    .C(_809_),
    .Y(_89_)
);

FILL FILL88650x50550 (
);

NAND2X1 _1462_ (
    .A(Yin[1]),
    .B(_119_),
    .Y(_652_)
);

NAND3X1 _1042_ (
    .A(_255_),
    .B(_275_),
    .C(_274_),
    .Y(_276_)
);

FILL FILL_0__1502_ (
);

FILL FILL_0__1099_ (
);

NAND3X1 _1518_ (
    .A(_183__bF$buf1),
    .B(_690_),
    .C(_691_),
    .Y(_692_)
);

OAI21X1 _1691_ (
    .A(_138_),
    .B(LoadCtl_6_bF$buf3),
    .C(_857_),
    .Y(_70_)
);

OAI21X1 _1271_ (
    .A(Stg_1_bF$buf1),
    .B(_492_),
    .C(Stg_2_bF$buf2),
    .Y(_493_)
);

FILL FILL_0__1311_ (
);

FILL FILL_2__1082_ (
);

DFFPOSX1 _1747_ (
    .D(_19_),
    .CLK(clk_bF$buf3),
    .Q(Acalc[5])
);

OAI21X1 _1327_ (
    .A(_541_),
    .B(_542_),
    .C(_536_),
    .Y(_545_)
);

FILL FILL_1__1489_ (
);

FILL FILL_1__1069_ (
);

NAND2X1 _1080_ (
    .A(Stg_0_bF$buf5),
    .B(_311_),
    .Y(_312_)
);

FILL FILL_0__1540_ (
);

FILL FILL_2__1558_ (
);

FILL FILL_2__1138_ (
);

FILL FILL_0__1120_ (
);

FILL FILL_1__1701_ (
);

NAND2X1 _1556_ (
    .A(Yin1[1]),
    .B(_728_),
    .Y(_729_)
);

NAND3X1 _1136_ (
    .A(_212_),
    .B(_365_),
    .C(_364_),
    .Y(_366_)
);

FILL FILL_0__884_ (
);

FILL FILL_1__918_ (
);

OAI21X1 _887_ (
    .A(_117_),
    .B(_127_),
    .C(_128_),
    .Y(_859_[1])
);

FILL FILL_1__1298_ (
);

FILL FILL_1__1510_ (
);

DFFPOSX1 _1785_ (
    .D(_57_),
    .CLK(clk_bF$buf6),
    .Q(Ain12b[5])
);

NOR2X1 _1365_ (
    .A(_580_),
    .B(_579_),
    .Y(_581_)
);

FILL FILL_0__1405_ (
);

NAND2X1 _1594_ (
    .A(_761_),
    .B(_762_),
    .Y(_765_)
);

NAND2X1 _1174_ (
    .A(_201__bF$buf4),
    .B(_394_),
    .Y(_402_)
);

FILL FILL_1__956_ (
);

FILL FILL_0__1634_ (
);

FILL FILL_0__1214_ (
);

FILL FILL_0__978_ (
);

FILL FILL_0__1443_ (
);

FILL FILL_0__1023_ (
);

FILL FILL_2__972_ (
);

FILL FILL_1__1604_ (
);

OAI21X1 _1459_ (
    .A(_265_),
    .B(_635_),
    .C(_650_),
    .Y(_45_)
);

AOI21X1 _1039_ (
    .A(_270_),
    .B(_272_),
    .C(_205_),
    .Y(_273_)
);

FILL FILL_1__994_ (
);

FILL FILL_0__1672_ (
);

FILL FILL_0__1252_ (
);

FILL FILL_1__1413_ (
);

AND2X2 _1688_ (
    .A(_841_),
    .B(_854_),
    .Y(_855_)
);

OAI21X1 _1268_ (
    .A(_188__bF$buf0),
    .B(_489_),
    .C(_490_),
    .Y(_14_)
);

FILL FILL_0__1308_ (
);

FILL FILL_0__1481_ (
);

FILL FILL_0__1061_ (
);

FILL FILL_1__1642_ (
);

FILL FILL_1__1222_ (
);

OAI21X1 _1497_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_670_),
    .C(_671_),
    .Y(_62_)
);

INVX1 _1077_ (
    .A(_308_),
    .Y(_309_)
);

FILL FILL_2__1711_ (
);

FILL FILL_0__1537_ (
);

FILL FILL_0__1117_ (
);

FILL FILL_0__1290_ (
);

FILL FILL_1__1451_ (
);

FILL FILL_1__1031_ (
);

FILL FILL_0__1346_ (
);

FILL FILL_1__1507_ (
);

FILL FILL88050x75750 (
);

FILL FILL_1__1680_ (
);

FILL FILL_1__1260_ (
);

FILL FILL_1__897_ (
);

FILL FILL_0__1575_ (
);

FILL FILL_0__1155_ (
);

FILL FILL_0__902_ (
);

AOI22X1 _905_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Ycalc[1]),
    .C(_119_),
    .D(Ycalc[3]),
    .Y(_145_)
);

FILL FILL_1__1316_ (
);

FILL FILL_0__1384_ (
);

DFFPOSX1 _1803_ (
    .D(_68_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[7])
);

FILL FILL_1__1545_ (
);

FILL FILL_1__1125_ (
);

FILL FILL_2__1614_ (
);

FILL FILL_2__969_ (
);

FILL FILL_0__1193_ (
);

NAND3X1 _1612_ (
    .A(_241_),
    .B(_778_),
    .C(_781_),
    .Y(_782_)
);

FILL FILL_0__940_ (
);

NOR2X1 _943_ (
    .A(_163_),
    .B(_179_),
    .Y(_180_)
);

FILL FILL_1__1354_ (
);

FILL FILL_0__1669_ (
);

FILL FILL_0__1249_ (
);

NAND2X1 _1421_ (
    .A(Xin[0]),
    .B(_629_),
    .Y(_630_)
);

OAI21X1 _1001_ (
    .A(Stg_0_bF$buf2),
    .B(_234_),
    .C(_235_),
    .Y(_236_)
);

FILL FILL_1__1583_ (
);

FILL FILL_1__1163_ (
);

FILL FILL_0__1478_ (
);

FILL FILL_0__1058_ (
);

FILL FILL_1__1639_ (
);

FILL FILL_1__1219_ (
);

NAND3X1 _1650_ (
    .A(_262_),
    .B(_807_),
    .C(_808_),
    .Y(_818_)
);

OAI21X1 _1230_ (
    .A(Ain12b_11_bF$buf3),
    .B(_436_),
    .C(_437_),
    .Y(_455_)
);

NAND3X1 _981_ (
    .A(_201__bF$buf6),
    .B(_179_),
    .C(_216_),
    .Y(_217_)
);

FILL FILL_1__1392_ (
);

FILL FILL_2__1708_ (
);

FILL FILL_2__1461_ (
);

FILL FILL_2__1041_ (
);

FILL FILL_0__1287_ (
);

AOI21X1 _1706_ (
    .A(_85_),
    .B(_84_),
    .C(_82_),
    .Y(_86_)
);

FILL FILL_1__1448_ (
);

FILL FILL_1__1028_ (
);

FILL FILL_0__1096_ (
);

NAND3X1 _1515_ (
    .A(Stg_2_bF$buf4),
    .B(_687_),
    .C(_688_),
    .Y(_689_)
);

FILL FILL_1__1677_ (
);

FILL FILL_1__1257_ (
);

DFFPOSX1 _1744_ (
    .D(_16_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[2])
);

OAI21X1 _1324_ (
    .A(_541_),
    .B(_542_),
    .C(LoadCtl_6_bF$buf2),
    .Y(_543_)
);

FILL FILL_1__1486_ (
);

FILL FILL_1__1066_ (
);

FILL FILL_2__1555_ (
);

FILL FILL_2__1135_ (
);

AOI21X1 _1553_ (
    .A(_725_),
    .B(Stg_2_bF$buf3),
    .C(_717_),
    .Y(_726_)
);

NAND3X1 _1133_ (
    .A(Xin12b[5]),
    .B(_362_),
    .C(_360_),
    .Y(_363_)
);

FILL FILL_0__881_ (
);

FILL FILL_1__915_ (
);

OAI21X1 _884_ (
    .A(_124_),
    .B(_113_),
    .C(_125_),
    .Y(_126_)
);

FILL FILL_1__1295_ (
);

NOR3X1 _1609_ (
    .A(_741_),
    .B(_760_),
    .C(_735_),
    .Y(_779_)
);

FILL FILL_0__937_ (
);

DFFPOSX1 _1782_ (
    .D(_54_),
    .CLK(clk_bF$buf2),
    .Q(Ain12b[6])
);

NAND2X1 _1362_ (
    .A(Ain12b[7]),
    .B(_577_),
    .Y(_578_)
);

FILL FILL_0__1402_ (
);

OAI21X1 _1418_ (
    .A(_471_),
    .B(_625_),
    .C(_627_),
    .Y(_27_)
);

OAI21X1 _1591_ (
    .A(_741_),
    .B(_735_),
    .C(_201__bF$buf6),
    .Y(_762_)
);

AOI21X1 _1171_ (
    .A(_394_),
    .B(_201__bF$buf1),
    .C(_396_),
    .Y(_399_)
);

FILL FILL_1__953_ (
);

FILL FILL_0__1631_ (
);

FILL FILL_0__1211_ (
);

FILL FILL88350x3750 (
);

OAI21X1 _1647_ (
    .A(_811_),
    .B(_813_),
    .C(_815_),
    .Y(_816_)
);

OAI21X1 _1227_ (
    .A(_451_),
    .B(_450_),
    .C(_201__bF$buf4),
    .Y(_452_)
);

FILL FILL_0__975_ (
);

OAI21X1 _978_ (
    .A(Stg_0_bF$buf4),
    .B(_212_),
    .C(_213_),
    .Y(_214_)
);

FILL FILL_1__1389_ (
);

FILL FILL_0__1440_ (
);

FILL FILL_2__1458_ (
);

FILL FILL_0__1020_ (
);

FILL FILL_2__1038_ (
);

FILL FILL_1__1601_ (
);

NAND2X1 _1456_ (
    .A(Yin[0]),
    .B(_635_),
    .Y(_649_)
);

OAI21X1 _1036_ (
    .A(Ain12b_11_bF$buf2),
    .B(_252_),
    .C(_269_),
    .Y(_270_)
);

FILL FILL_1__1198_ (
);

FILL FILL_1__991_ (
);

FILL FILL_1__1410_ (
);

NOR2X1 _1685_ (
    .A(_844_),
    .B(_851_),
    .Y(_852_)
);

AND2X2 _1265_ (
    .A(_486_),
    .B(_483_),
    .Y(_488_)
);

FILL FILL_0__1725_ (
);

FILL FILL_0__1305_ (
);

OAI21X1 _1494_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_504_),
    .C(_669_),
    .Y(_61_)
);

OAI21X1 _1074_ (
    .A(_304_),
    .B(_306_),
    .C(_281_),
    .Y(_4_)
);

FILL FILL87750x61350 (
);

FILL FILL_0__1534_ (
);

FILL FILL_0__1114_ (
);

FILL FILL_0__878_ (
);

BUFX2 BUFX2_insert0 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf6)
);

BUFX2 BUFX2_insert1 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf5)
);

BUFX2 BUFX2_insert2 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf4)
);

BUFX2 BUFX2_insert3 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf3)
);

BUFX2 BUFX2_insert4 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf2)
);

BUFX2 BUFX2_insert5 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf1)
);

BUFX2 BUFX2_insert6 (
    .A(Stg[0]),
    .Y(Stg_0_bF$buf0)
);

BUFX2 BUFX2_insert7 (
    .A(_188_),
    .Y(_188__bF$buf4)
);

BUFX2 BUFX2_insert8 (
    .A(_188_),
    .Y(_188__bF$buf3)
);

BUFX2 BUFX2_insert9 (
    .A(_188_),
    .Y(_188__bF$buf2)
);

FILL FILL_0__1343_ (
);

FILL FILL_2__872_ (
);

FILL FILL_1__1504_ (
);

DFFPOSX1 _1779_ (
    .D(_51_),
    .CLK(clk_bF$buf6),
    .Q(Ain12b[11])
);

OAI21X1 _1359_ (
    .A(Stg_2_bF$buf0),
    .B(Stg_0_bF$buf6),
    .C(Ain12b_11_bF$buf4),
    .Y(_575_)
);

FILL FILL_1__894_ (
);

FILL FILL_0__1572_ (
);

FILL FILL_0__1152_ (
);

INVX1 _902_ (
    .A(Ycalc[5]),
    .Y(_142_)
);

FILL FILL_1__1313_ (
);

NAND2X1 _1588_ (
    .A(_183__bF$buf0),
    .B(_223_),
    .Y(_759_)
);

AOI21X1 _1168_ (
    .A(_315_),
    .B(_183__bF$buf2),
    .C(_395_),
    .Y(_396_)
);

FILL FILL_0__1628_ (
);

FILL FILL_0__1208_ (
);

FILL FILL_0__1381_ (
);

DFFPOSX1 _1800_ (
    .D(_65_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[4])
);

FILL FILL_1__1542_ (
);

FILL FILL_1__1122_ (
);

OAI21X1 _1397_ (
    .A(_609_),
    .B(_605_),
    .C(LoadCtl_6_bF$buf0),
    .Y(_611_)
);

FILL FILL_2__1611_ (
);

FILL FILL_0__1437_ (
);

FILL FILL_0__1017_ (
);

FILL FILL_2__966_ (
);

FILL FILL_0__1190_ (
);

OAI21X1 _940_ (
    .A(Stg_0_bF$buf4),
    .B(_175_),
    .C(_176_),
    .Y(_177_)
);

FILL FILL_1__1351_ (
);

FILL FILL_1__988_ (
);

FILL FILL_0__1666_ (
);

FILL FILL_0__1246_ (
);

FILL FILL_1__1407_ (
);

FILL FILL_1__1580_ (
);

FILL FILL_1__1160_ (
);

FILL FILL_0__1475_ (
);

FILL FILL_0__1055_ (
);

FILL FILL_1__1636_ (
);

FILL FILL_1__1216_ (
);

FILL FILL_0__1284_ (
);

AOI21X1 _1703_ (
    .A(_845_),
    .B(_848_),
    .C(_284_),
    .Y(_83_)
);

FILL FILL88050x61350 (
);

FILL FILL_1__1445_ (
);

FILL FILL_1__1025_ (
);

FILL FILL_2__1514_ (
);

FILL FILL_2__869_ (
);

FILL FILL_0__1093_ (
);

NAND2X1 _1512_ (
    .A(Stg_0_bF$buf4),
    .B(_212_),
    .Y(_686_)
);

FILL FILL_1__1674_ (
);

FILL FILL_1__1254_ (
);

FILL FILL_0__1569_ (
);

FILL FILL_0__1149_ (
);

DFFPOSX1 _1741_ (
    .D(_13_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[11])
);

AOI21X1 _1321_ (
    .A(_536_),
    .B(_538_),
    .C(_539_),
    .Y(_540_)
);

FILL FILL_1__1483_ (
);

FILL FILL_1__1063_ (
);

FILL FILL_2__1132_ (
);

FILL FILL_0__1378_ (
);

FILL FILL_1__1539_ (
);

FILL FILL_1__1119_ (
);

OAI21X1 _1550_ (
    .A(Stg_0_bF$buf3),
    .B(Xin12b[9]),
    .C(_722_),
    .Y(_723_)
);

NAND3X1 _1130_ (
    .A(_201__bF$buf1),
    .B(_359_),
    .C(_354_),
    .Y(_360_)
);

FILL FILL_1__912_ (
);

OAI21X1 _881_ (
    .A(LoadCtl[4]),
    .B(_121_),
    .C(_122_),
    .Y(_123_)
);

FILL FILL_1__1292_ (
);

FILL FILL_2__1608_ (
);

FILL FILL_2__1361_ (
);

FILL FILL_0__1187_ (
);

NAND2X1 _1606_ (
    .A(_183__bF$buf0),
    .B(_676_),
    .Y(_776_)
);

FILL FILL_0__934_ (
);

OAI21X1 _937_ (
    .A(Stg_0_bF$buf3),
    .B(_172_),
    .C(_173_),
    .Y(_174_)
);

FILL FILL_1__1348_ (
);

NAND2X1 _1415_ (
    .A(Xin[0]),
    .B(_625_),
    .Y(_626_)
);

FILL FILL_1__1577_ (
);

FILL FILL_1__1157_ (
);

FILL FILL_1__950_ (
);

OAI21X1 _1644_ (
    .A(Stg_2_bF$buf0),
    .B(_484_),
    .C(_812_),
    .Y(_813_)
);

OAI21X1 _1224_ (
    .A(Stg_2_bF$buf4),
    .B(_373_),
    .C(_415_),
    .Y(_449_)
);

FILL FILL_0__972_ (
);

OAI21X1 _975_ (
    .A(Stg_0_bF$buf3),
    .B(_209_),
    .C(_210_),
    .Y(_211_)
);

FILL FILL_1__1386_ (
);

FILL FILL_2__1455_ (
);

FILL FILL_2__1035_ (
);

OAI21X1 _1453_ (
    .A(_241_),
    .B(_632_),
    .C(_647_),
    .Y(_42_)
);

OAI21X1 _1033_ (
    .A(Stg_0_bF$buf0),
    .B(_265_),
    .C(_266_),
    .Y(_267_)
);

FILL FILL_1__1195_ (
);

NAND2X1 _1509_ (
    .A(_164__bF$buf2),
    .B(_170_),
    .Y(_683_)
);

FILL FILL88350x36150 (
);

NAND3X1 _1682_ (
    .A(_284_),
    .B(_848_),
    .C(_845_),
    .Y(_849_)
);

NAND2X1 _1262_ (
    .A(Stg_0_bF$buf1),
    .B(Stg_1_bF$buf2),
    .Y(_485_)
);

FILL FILL_0__1722_ (
);

FILL FILL_0__1302_ (
);

DFFPOSX1 _1738_ (
    .D(_10_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[8])
);

INVX1 _1318_ (
    .A(Ain12b[4]),
    .Y(_537_)
);

NAND2X1 _1491_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Ain[0]),
    .Y(_668_)
);

NOR2X1 _1071_ (
    .A(_283_),
    .B(_303_),
    .Y(_304_)
);

FILL FILL_0__1531_ (
);

FILL FILL_0__1111_ (
);

NAND3X1 _1547_ (
    .A(_201__bF$buf6),
    .B(_719_),
    .C(_712_),
    .Y(_720_)
);

NOR2X1 _1127_ (
    .A(_164__bF$buf3),
    .B(_356_),
    .Y(_357_)
);

FILL FILL_0__875_ (
);

FILL FILL_1__909_ (
);

OAI21X1 _878_ (
    .A(_117_),
    .B(_115_),
    .C(_120_),
    .Y(_859_[0])
);

FILL FILL_1__1289_ (
);

FILL FILL_0__1340_ (
);

FILL FILL_2__1358_ (
);

FILL FILL_1__1501_ (
);

FILL FILL88650x79350 (
);

DFFPOSX1 _1776_ (
    .D(_48_),
    .CLK(clk_bF$buf5),
    .Q(Yin0[0])
);

OAI22X1 _1356_ (
    .A(_110_),
    .B(LoadCtl_6_bF$buf4),
    .C(_572_),
    .D(_571_),
    .Y(_20_)
);

FILL FILL_1__1098_ (
);

FILL FILL_1__891_ (
);

FILL FILL_1__1310_ (
);

INVX1 _1585_ (
    .A(_755_),
    .Y(_756_)
);

NOR2X1 _1165_ (
    .A(_392_),
    .B(_388_),
    .Y(_393_)
);

FILL FILL_1__947_ (
);

FILL FILL_0__1625_ (
);

FILL FILL_0__1205_ (
);

FILL FILL_0__969_ (
);

NAND2X1 _1394_ (
    .A(Ain12b[9]),
    .B(_201__bF$buf0),
    .Y(_608_)
);

FILL FILL_0__1434_ (
);

FILL FILL_0__1014_ (
);

FILL FILL_2__963_ (
);

FILL FILL_1__985_ (
);

FILL FILL_0__1663_ (
);

FILL FILL_0__1243_ (
);

FILL FILL_1__1404_ (
);

NOR2X1 _1679_ (
    .A(_777_),
    .B(_774_),
    .Y(_846_)
);

OAI22X1 _1259_ (
    .A(_154_),
    .B(LoadCtl_6_bF$buf1),
    .C(_480_),
    .D(_482_),
    .Y(_13_)
);

FILL FILL_0__1719_ (
);

FILL FILL_0__1472_ (
);

FILL FILL_0__1052_ (
);

FILL FILL_1__1633_ (
);

FILL FILL_1__1213_ (
);

OAI21X1 _1488_ (
    .A(_664_),
    .B(_665_),
    .C(_666_),
    .Y(_58_)
);

INVX1 _1068_ (
    .A(_300_),
    .Y(_301_)
);

FILL FILL_0__1528_ (
);

FILL FILL_0__1108_ (
);

FILL FILL_0__1281_ (
);

FILL FILL_2__1299_ (
);

NOR2X1 _1700_ (
    .A(_73_),
    .B(_74_),
    .Y(_80_)
);

FILL FILL_1__1442_ (
);

FILL FILL_1__1022_ (
);

INVX1 _1297_ (
    .A(_516_),
    .Y(_517_)
);

FILL FILL_2__1511_ (
);

FILL FILL_0__1337_ (
);

FILL FILL_2__866_ (
);

FILL FILL_0__1090_ (
);

FILL FILL_1__1671_ (
);

FILL FILL_1__1251_ (
);

FILL FILL_1__888_ (
);

FILL FILL_0__1566_ (
);

FILL FILL_0__1146_ (
);

FILL FILL_1__1727_ (
);

FILL FILL_1__1307_ (
);

FILL FILL_0_BUFX2_insert40 (
);

FILL FILL_0_BUFX2_insert41 (
);

FILL FILL_0_BUFX2_insert42 (
);

FILL FILL_0_BUFX2_insert43 (
);

FILL FILL_0_BUFX2_insert44 (
);

FILL FILL_0_BUFX2_insert45 (
);

FILL FILL_0_BUFX2_insert46 (
);

FILL FILL_0_BUFX2_insert47 (
);

FILL FILL_0_BUFX2_insert48 (
);

FILL FILL_0_BUFX2_insert49 (
);

FILL FILL_1__1480_ (
);

FILL FILL_1__1060_ (
);

FILL FILL_0__1375_ (
);

FILL FILL_1__1536_ (
);

FILL FILL_1__1116_ (
);

FILL FILL_2__1605_ (
);

FILL FILL_0__1184_ (
);

OAI21X1 _1603_ (
    .A(_142_),
    .B(LoadCtl_6_bF$buf3),
    .C(_773_),
    .Y(_66_)
);

FILL FILL_0__931_ (
);

MUX2X1 _934_ (
    .A(_170_),
    .B(_167_),
    .S(_164__bF$buf1),
    .Y(_171_)
);

FILL FILL_1__1345_ (
);

OAI21X1 _1412_ (
    .A(_188__bF$buf4),
    .B(_623_),
    .C(_622_),
    .Y(_25_)
);

FILL FILL_1__1574_ (
);

FILL FILL_1__1154_ (
);

BUFX2 BUFX2_insert50 (
    .A(Ain12b[11]),
    .Y(Ain12b_11_bF$buf1)
);

BUFX2 BUFX2_insert51 (
    .A(Ain12b[11]),
    .Y(Ain12b_11_bF$buf0)
);

BUFX2 BUFX2_insert52 (
    .A(_201_),
    .Y(_201__bF$buf6)
);

BUFX2 BUFX2_insert53 (
    .A(_201_),
    .Y(_201__bF$buf5)
);

BUFX2 BUFX2_insert54 (
    .A(_201_),
    .Y(_201__bF$buf4)
);

BUFX2 BUFX2_insert55 (
    .A(_201_),
    .Y(_201__bF$buf3)
);

BUFX2 BUFX2_insert56 (
    .A(_201_),
    .Y(_201__bF$buf2)
);

BUFX2 BUFX2_insert57 (
    .A(_201_),
    .Y(_201__bF$buf1)
);

BUFX2 BUFX2_insert58 (
    .A(_201_),
    .Y(_201__bF$buf0)
);

FILL FILL_0__1469_ (
);

FILL FILL_0__1049_ (
);

NOR2X1 _1641_ (
    .A(_806_),
    .B(_809_),
    .Y(_810_)
);

AOI22X1 _1221_ (
    .A(_440_),
    .B(_444_),
    .C(_431_),
    .D(_421_),
    .Y(_447_)
);

MUX2X1 _972_ (
    .A(_207_),
    .B(_204_),
    .S(_164__bF$buf2),
    .Y(_208_)
);

FILL FILL_1__1383_ (
);

FILL FILL_2__1452_ (
);

FILL FILL_2__1032_ (
);

FILL FILL_0__1698_ (
);

FILL FILL_0__1278_ (
);

FILL FILL_1__1439_ (
);

FILL FILL_1__1019_ (
);

NAND2X1 _1450_ (
    .A(Yin[1]),
    .B(_629_),
    .Y(_646_)
);

OAI21X1 _1030_ (
    .A(Stg_0_bF$buf0),
    .B(_262_),
    .C(_263_),
    .Y(_264_)
);

FILL FILL_1__1192_ (
);

FILL FILL_2__1508_ (
);

FILL FILL_2__1681_ (
);

FILL FILL_0__1087_ (
);

NAND2X1 _1506_ (
    .A(_492_),
    .B(_165_),
    .Y(_680_)
);

FILL FILL_1__1668_ (
);

FILL FILL_1__1248_ (
);

FILL FILL88350x57750 (
);

DFFPOSX1 _1735_ (
    .D(_7_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[5])
);

AOI21X1 _1315_ (
    .A(_493_),
    .B(_533_),
    .C(_201__bF$buf3),
    .Y(_534_)
);

FILL FILL_1__1477_ (
);

FILL FILL_1__1057_ (
);

OAI22X1 _1544_ (
    .A(_184_),
    .B(_218_),
    .C(_222_),
    .D(_289_),
    .Y(_717_)
);

INVX1 _1124_ (
    .A(_353_),
    .Y(_354_)
);

FILL FILL_0__872_ (
);

FILL FILL_1__906_ (
);

INVX1 _875_ (
    .A(LoadCtl[1]),
    .Y(_118_)
);

FILL FILL_1__1286_ (
);

FILL FILL_2__1355_ (
);

FILL FILL_0__928_ (
);

DFFPOSX1 _1773_ (
    .D(_45_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[5])
);

NAND2X1 _1353_ (
    .A(_569_),
    .B(_567_),
    .Y(_570_)
);

FILL FILL_1__1095_ (
);

FILL FILL_0__1813_ (
);

FILL FILL_2__922_ (
);

OAI22X1 _1409_ (
    .A(_106_),
    .B(LoadCtl_6_bF$buf0),
    .C(_621_),
    .D(_620_),
    .Y(_24_)
);

FILL FILL88650x10950 (
);

OAI21X1 _1582_ (
    .A(_750_),
    .B(_752_),
    .C(_753_),
    .Y(_754_)
);

NAND2X1 _1162_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_390_),
    .Y(_391_)
);

FILL FILL_1__944_ (
);

FILL FILL_0__1622_ (
);

FILL FILL_0__1202_ (
);

NAND3X1 _1638_ (
    .A(_201__bF$buf5),
    .B(_803_),
    .C(_799_),
    .Y(_807_)
);

OAI21X1 _1218_ (
    .A(_443_),
    .B(_442_),
    .C(_441_),
    .Y(_444_)
);

FILL FILL_0__966_ (
);

INVX1 _969_ (
    .A(Xin0[1]),
    .Y(_205_)
);

AOI21X1 _1391_ (
    .A(_599_),
    .B(_593_),
    .C(_604_),
    .Y(_605_)
);

FILL FILL_0__1431_ (
);

FILL FILL_0__1011_ (
);

INVX1 _1447_ (
    .A(Yin12b[8]),
    .Y(_644_)
);

MUX2X1 _1027_ (
    .A(_260_),
    .B(_258_),
    .S(_164__bF$buf1),
    .Y(_261_)
);

FILL FILL_1__1189_ (
);

FILL FILL_1__982_ (
);

FILL FILL_0__1660_ (
);

FILL FILL_2__1678_ (
);

FILL FILL_2__1258_ (
);

FILL FILL_0__1240_ (
);

FILL FILL_1__1401_ (
);

OAI21X1 _1676_ (
    .A(Stg_2_bF$buf3),
    .B(_758_),
    .C(_826_),
    .Y(_843_)
);

AOI21X1 _1256_ (
    .A(_466_),
    .B(_457_),
    .C(_479_),
    .Y(_480_)
);

FILL FILL_0__1716_ (
);

FILL FILL_1__1630_ (
);

FILL FILL_1__1210_ (
);

INVX1 _1485_ (
    .A(Ain[0]),
    .Y(_664_)
);

AOI21X1 _1065_ (
    .A(_240_),
    .B(_248_),
    .C(_269_),
    .Y(_298_)
);

FILL FILL_0__1525_ (
);

FILL FILL_0__1105_ (
);

FILL FILL_0__869_ (
);

NAND2X1 _1294_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_514_),
    .Y(_515_)
);

FILL FILL_0__1334_ (
);

FILL FILL_2__863_ (
);

FILL FILL_1__885_ (
);

FILL FILL_2__919_ (
);

FILL FILL_0__1563_ (
);

FILL FILL_0__1143_ (
);

FILL FILL_1__1724_ (
);

FILL FILL_1__1304_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

OAI21X1 _1579_ (
    .A(Yin1[1]),
    .B(_728_),
    .C(_710_),
    .Y(_751_)
);

AND2X2 _1159_ (
    .A(_387_),
    .B(_382_),
    .Y(_388_)
);

FILL FILL_0__1619_ (
);

FILL FILL_0__1372_ (
);

FILL FILL_1__1533_ (
);

FILL FILL_1__1113_ (
);

OAI21X1 _1388_ (
    .A(_600_),
    .B(_602_),
    .C(_585_),
    .Y(_22_)
);

FILL FILL_0__1428_ (
);

FILL FILL_0__1008_ (
);

FILL FILL_0__1181_ (
);

FILL FILL_2__1199_ (
);

NAND3X1 _1600_ (
    .A(_749_),
    .B(_769_),
    .C(_756_),
    .Y(_771_)
);

INVX1 _931_ (
    .A(Xin0[0]),
    .Y(_168_)
);

FILL FILL_1__1342_ (
);

NAND2X1 _1197_ (
    .A(_416_),
    .B(_419_),
    .Y(_424_)
);

FILL FILL_1__979_ (
);

FILL FILL_2__1411_ (
);

FILL FILL_0__1657_ (
);

FILL FILL_0__1237_ (
);

FILL FILL_1__1571_ (
);

FILL FILL_1__1151_ (
);

BUFX2 BUFX2_insert20 (
    .A(_164_),
    .Y(_164__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(_164_),
    .Y(_164__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(_164_),
    .Y(_164__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(_164_),
    .Y(_164__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(_164_),
    .Y(_164__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf0)
);

FILL FILL_0__1466_ (
);

FILL FILL_0__1046_ (
);

FILL FILL_1__1627_ (
);

FILL FILL_1__1207_ (
);

FILL FILL_1__1380_ (
);

FILL FILL_0__1695_ (
);

FILL FILL_0__1275_ (
);

FILL FILL_1__1436_ (
);

FILL FILL_1__1016_ (
);

FILL FILL_2__1505_ (
);

FILL FILL_0__1084_ (
);

OAI22X1 _1503_ (
    .A(_184_),
    .B(_193_),
    .C(_197_),
    .D(_289_),
    .Y(_677_)
);

FILL FILL_1__1665_ (
);

FILL FILL_1__1245_ (
);

DFFPOSX1 _1732_ (
    .D(_4_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[2])
);

NAND2X1 _1312_ (
    .A(Acalc[4]),
    .B(_188__bF$buf4),
    .Y(_531_)
);

FILL FILL_1__1474_ (
);

FILL FILL_1__1054_ (
);

FILL FILL_0__1369_ (
);

OAI21X1 _1541_ (
    .A(Stg_0_bF$buf5),
    .B(_441_),
    .C(_713_),
    .Y(_714_)
);

AOI22X1 _1121_ (
    .A(_150_),
    .B(_188__bF$buf3),
    .C(_351_),
    .D(_186_),
    .Y(_6_)
);

FILL FILL_1__903_ (
);

AOI21X1 _872_ (
    .A(_108_),
    .B(_109_),
    .C(_114_),
    .Y(_115_)
);

FILL FILL_1__1283_ (
);

FILL FILL_2__1352_ (
);

FILL FILL_0__1598_ (
);

FILL FILL_0__1178_ (
);

FILL FILL_0__925_ (
);

INVX1 _928_ (
    .A(Xin1[0]),
    .Y(_165_)
);

FILL FILL_1__1339_ (
);

DFFPOSX1 _1770_ (
    .D(_42_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[6])
);

NAND2X1 _1350_ (
    .A(Ain12b[6]),
    .B(_566_),
    .Y(_567_)
);

FILL FILL_1__1092_ (
);

FILL FILL_0__1810_ (
);

FILL FILL_2__1408_ (
);

NAND2X1 _1406_ (
    .A(_617_),
    .B(_618_),
    .Y(_619_)
);

FILL FILL_1__1568_ (
);

FILL FILL_1__1148_ (
);

FILL FILL_1__941_ (
);

OAI21X1 _1635_ (
    .A(_777_),
    .B(_774_),
    .C(_201__bF$buf5),
    .Y(_804_)
);

INVX1 _1215_ (
    .A(Xin12b[9]),
    .Y(_441_)
);

FILL FILL_0__963_ (
);

INVX1 _966_ (
    .A(Xin1[1]),
    .Y(_202_)
);

FILL FILL_2_CLKBUF1_insert14 (
);

FILL FILL_2_CLKBUF1_insert17 (
);

FILL FILL_1__1377_ (
);

OAI21X1 _1444_ (
    .A(_311_),
    .B(_625_),
    .C(_642_),
    .Y(_38_)
);

OAI21X1 _1024_ (
    .A(Stg_0_bF$buf2),
    .B(_256_),
    .C(_257_),
    .Y(_258_)
);

FILL FILL_1__1186_ (
);

FILL FILL88350x43350 (
);

FILL FILL_2__1675_ (
);

FILL FILL_2__1255_ (
);

INVX1 _1673_ (
    .A(_835_),
    .Y(_840_)
);

NOR2X1 _1253_ (
    .A(Ain12b_11_bF$buf3),
    .B(_454_),
    .Y(_477_)
);

FILL FILL_0__1713_ (
);

DFFPOSX1 _1729_ (
    .D(_1_),
    .CLK(clk_bF$buf5),
    .Q(Ycalc[1])
);

NAND2X1 _1309_ (
    .A(_528_),
    .B(_526_),
    .Y(_529_)
);

OAI21X1 _1482_ (
    .A(_537_),
    .B(_635_),
    .C(_662_),
    .Y(_56_)
);

AOI21X1 _1062_ (
    .A(_288_),
    .B(Stg_2_bF$buf1),
    .C(_294_),
    .Y(_295_)
);

FILL FILL_0__1522_ (
);

FILL FILL_0__1102_ (
);

INVX1 _1538_ (
    .A(_710_),
    .Y(_711_)
);

OR2X2 _1118_ (
    .A(_331_),
    .B(_348_),
    .Y(_349_)
);

FILL FILL_0__866_ (
);

INVX2 _869_ (
    .A(LoadCtl[2]),
    .Y(_112_)
);

INVX1 _1291_ (
    .A(_511_),
    .Y(_512_)
);

FILL FILL88650x86550 (
);

FILL FILL_0__1331_ (
);

FILL FILL_2__1349_ (
);

DFFPOSX1 _1767_ (
    .D(_39_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[11])
);

NOR2X1 _1347_ (
    .A(_201__bF$buf0),
    .B(_563_),
    .Y(_564_)
);

FILL FILL_1__1089_ (
);

FILL FILL_1__882_ (
);

FILL FILL_2__916_ (
);

FILL FILL_0__1560_ (
);

FILL FILL_2__1578_ (
);

FILL FILL_0__1140_ (
);

FILL FILL_2__1158_ (
);

FILL FILL_1__1721_ (
);

FILL FILL_1__1301_ (
);

AOI21X1 _1576_ (
    .A(_735_),
    .B(_201__bF$buf6),
    .C(_741_),
    .Y(_748_)
);

AOI21X1 _1156_ (
    .A(_364_),
    .B(_365_),
    .C(_212_),
    .Y(_385_)
);

FILL FILL_1__938_ (
);

FILL FILL_0__1616_ (
);

FILL FILL_1__1530_ (
);

FILL FILL_1__1110_ (
);

NOR2X1 _1385_ (
    .A(_593_),
    .B(_599_),
    .Y(_600_)
);

FILL FILL_0__1425_ (
);

FILL FILL_0__1005_ (
);

FILL FILL_2__1196_ (
);

NAND3X1 _1194_ (
    .A(Xin12b[8]),
    .B(_417_),
    .C(_420_),
    .Y(_421_)
);

FILL FILL_1__976_ (
);

FILL FILL_0__1654_ (
);

FILL FILL_0__1234_ (
);

FILL FILL87750x21750 (
);

FILL FILL_1__1815_ (
);

FILL FILL_0__998_ (
);

FILL FILL_0__1463_ (
);

FILL FILL_0__1043_ (
);

FILL FILL88650x18150 (
);

FILL FILL_1__1624_ (
);

FILL FILL_1__1204_ (
);

NOR2X1 _1479_ (
    .A(Ain12b[7]),
    .B(_632_),
    .Y(_661_)
);

INVX1 _1059_ (
    .A(_184_),
    .Y(_292_)
);

FILL FILL_0__1519_ (
);

FILL FILL_0__1692_ (
);

FILL FILL_0__1272_ (
);

FILL FILL_1__1433_ (
);

FILL FILL_1__1013_ (
);

NAND2X1 _1288_ (
    .A(Ain1[0]),
    .B(_508_),
    .Y(_509_)
);

FILL FILL_2__1502_ (
);

FILL FILL_0__1328_ (
);

FILL FILL_1_BUFX2_insert50 (
);

FILL FILL_1_BUFX2_insert51 (
);

FILL FILL_1_BUFX2_insert52 (
);

FILL FILL_1_BUFX2_insert53 (
);

FILL FILL_1_BUFX2_insert54 (
);

FILL FILL_1_BUFX2_insert55 (
);

FILL FILL_1_BUFX2_insert56 (
);

FILL FILL_1_BUFX2_insert57 (
);

FILL FILL_1_BUFX2_insert58 (
);

FILL FILL88650x7350 (
);

FILL FILL_2__1099_ (
);

FILL FILL_0__1081_ (
);

NAND2X1 _1500_ (
    .A(_199_),
    .B(_224_),
    .Y(_674_)
);

FILL FILL_1__1662_ (
);

FILL FILL_1__1242_ (
);

NAND2X1 _1097_ (
    .A(_309_),
    .B(_327_),
    .Y(_329_)
);

FILL FILL_1__879_ (
);

FILL FILL_2__1311_ (
);

FILL FILL_0__1557_ (
);

FILL FILL_0__1137_ (
);

FILL FILL_1__1718_ (
);

FILL FILL_1__1471_ (
);

FILL FILL_1__1051_ (
);

FILL FILL_0__1366_ (
);

FILL FILL_1__1527_ (
);

FILL FILL_1__1107_ (
);

FILL FILL_1__900_ (
);

FILL FILL_1__1280_ (
);

FILL FILL_0__1595_ (
);

FILL FILL_0__1175_ (
);

FILL FILL_0__922_ (
);

INVX1 _925_ (
    .A(Ycalc[0]),
    .Y(_162_)
);

FILL FILL_1__1336_ (
);

FILL FILL_2__1405_ (
);

INVX1 _1403_ (
    .A(Ain12b[10]),
    .Y(_616_)
);

FILL FILL_1__1565_ (
);

FILL FILL_1__1145_ (
);

FILL FILL88050x21750 (
);

AOI21X1 _1632_ (
    .A(_725_),
    .B(_183__bF$buf2),
    .C(_800_),
    .Y(_801_)
);

NAND2X1 _1212_ (
    .A(_436_),
    .B(_437_),
    .Y(_438_)
);

FILL FILL_0__960_ (
);

MUX2X1 _963_ (
    .A(_198_),
    .B(_195_),
    .S(Stg_2_bF$buf1),
    .Y(_199_)
);

FILL FILL_1__1374_ (
);

FILL FILL_0__1689_ (
);

FILL FILL_0__1269_ (
);

NAND2X1 _1441_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[1]),
    .Y(_641_)
);

NOR2X1 _1021_ (
    .A(_168_),
    .B(_252_),
    .Y(_255_)
);

FILL FILL_1__1183_ (
);

FILL FILL_2__1672_ (
);

FILL FILL_2__1252_ (
);

FILL FILL_0__1498_ (
);

FILL FILL_0__1078_ (
);

FILL FILL_1__1659_ (
);

FILL FILL_1__1239_ (
);

FILL FILL88350x64950 (
);

OAI21X1 _1670_ (
    .A(_836_),
    .B(_823_),
    .C(_191_),
    .Y(_838_)
);

NAND2X1 _1250_ (
    .A(_472_),
    .B(_473_),
    .Y(_474_)
);

FILL FILL_0__1710_ (
);

FILL FILL_2__1308_ (
);

OAI21X1 _1726_ (
    .A(_102_),
    .B(_104_),
    .C(_709_),
    .Y(_105_)
);

OAI21X1 _1306_ (
    .A(_523_),
    .B(_525_),
    .C(_517_),
    .Y(_526_)
);

FILL FILL_1__1468_ (
);

FILL FILL_1__1048_ (
);

INVX1 _1535_ (
    .A(Ycalc[3]),
    .Y(_708_)
);

NAND3X1 _1115_ (
    .A(_175_),
    .B(_340_),
    .C(_345_),
    .Y(_346_)
);

FILL FILL_0__863_ (
);

NOR2X1 _866_ (
    .A(LoadCtl[3]),
    .B(LoadCtl[2]),
    .Y(_109_)
);

FILL FILL_1__1697_ (
);

FILL FILL_1__1277_ (
);

FILL FILL_0__919_ (
);

DFFPOSX1 _1764_ (
    .D(_36_),
    .CLK(clk_bF$buf5),
    .Q(Xin0[0])
);

OAI21X1 _1344_ (
    .A(_536_),
    .B(_555_),
    .C(_552_),
    .Y(_561_)
);

FILL FILL_1__1086_ (
);

FILL FILL_2__913_ (
);

FILL FILL_2__1575_ (
);

FILL FILL_2__1155_ (
);

OAI21X1 _1573_ (
    .A(Ain12b_11_bF$buf1),
    .B(_743_),
    .C(_744_),
    .Y(_745_)
);

AND2X2 _1153_ (
    .A(_380_),
    .B(_381_),
    .Y(_382_)
);

FILL FILL_1__935_ (
);

FILL FILL_0__1613_ (
);

AOI21X1 _1629_ (
    .A(_797_),
    .B(_782_),
    .C(_791_),
    .Y(_798_)
);

OR2X2 _1209_ (
    .A(_355_),
    .B(_357_),
    .Y(_435_)
);

FILL FILL_0__957_ (
);

AOI21X1 _1382_ (
    .A(_561_),
    .B(_596_),
    .C(_594_),
    .Y(_597_)
);

FILL FILL_0__1422_ (
);

FILL FILL_0__1002_ (
);

OAI21X1 _1438_ (
    .A(_202_),
    .B(_119_),
    .C(_639_),
    .Y(_35_)
);

OAI21X1 _1018_ (
    .A(_168_),
    .B(_252_),
    .C(_186_),
    .Y(_253_)
);

INVX1 _1191_ (
    .A(_416_),
    .Y(_418_)
);

FILL FILL_1__973_ (
);

FILL FILL_0__1651_ (
);

FILL FILL_2__1669_ (
);

FILL FILL_0__1231_ (
);

FILL FILL_2__1249_ (
);

FILL FILL_1__1812_ (
);

NAND3X1 _1667_ (
    .A(Yin12b[8]),
    .B(_829_),
    .C(_834_),
    .Y(_835_)
);

INVX1 _1247_ (
    .A(Xin12b[11]),
    .Y(_471_)
);

FILL FILL_0__995_ (
);

NAND2X1 _998_ (
    .A(Xcalc[0]),
    .B(_188__bF$buf1),
    .Y(_233_)
);

FILL FILL_0__1707_ (
);

FILL FILL_0__1460_ (
);

FILL FILL_0__1040_ (
);

FILL FILL_1__1621_ (
);

FILL FILL_1__1201_ (
);

FILL FILL88650x72150 (
);

NAND2X1 _1476_ (
    .A(Ain[0]),
    .B(_632_),
    .Y(_659_)
);

NAND2X1 _1056_ (
    .A(Stg_1_bF$buf2),
    .B(_183__bF$buf1),
    .Y(_289_)
);

FILL FILL88650x39750 (
);

FILL FILL_0__1516_ (
);

FILL FILL_1__1430_ (
);

FILL FILL_1__1010_ (
);

OAI21X1 _1285_ (
    .A(_492_),
    .B(_164__bF$buf1),
    .C(Ain12b_11_bF$buf4),
    .Y(_506_)
);

FILL FILL_0__1325_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_1_BUFX2_insert21 (
);

FILL FILL_1_BUFX2_insert22 (
);

FILL FILL_1_BUFX2_insert23 (
);

FILL FILL_1_BUFX2_insert24 (
);

FILL FILL_1_BUFX2_insert25 (
);

FILL FILL_1_BUFX2_insert26 (
);

FILL FILL_1_BUFX2_insert27 (
);

FILL FILL_1_BUFX2_insert28 (
);

FILL FILL_1_BUFX2_insert29 (
);

FILL FILL_2__1096_ (
);

NAND3X1 _1094_ (
    .A(_202_),
    .B(_320_),
    .C(_323_),
    .Y(_326_)
);

FILL FILL_1__876_ (
);

FILL FILL_0__1554_ (
);

FILL FILL_0__1134_ (
);

FILL FILL_1__1715_ (
);

FILL FILL_0__898_ (
);

FILL FILL_0__1363_ (
);

FILL FILL_1__1524_ (
);

FILL FILL_1__1104_ (
);

DFFPOSX1 _1799_ (
    .D(_64_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[3])
);

OAI21X1 _1379_ (
    .A(_580_),
    .B(_567_),
    .C(_578_),
    .Y(_594_)
);

FILL FILL_0__1419_ (
);

FILL FILL_0__1592_ (
);

FILL FILL_0__1172_ (
);

AOI21X1 _922_ (
    .A(_109_),
    .B(_156_),
    .C(_159_),
    .Y(_160_)
);

FILL FILL_1__1333_ (
);

INVX1 _1188_ (
    .A(_395_),
    .Y(_415_)
);

FILL FILL_2__1402_ (
);

FILL FILL_0__1648_ (
);

FILL FILL_0__1228_ (
);

FILL FILL_1__1809_ (
);

OR2X2 _1400_ (
    .A(_592_),
    .B(_609_),
    .Y(_613_)
);

FILL FILL_1__1562_ (
);

FILL FILL_1__1142_ (
);

FILL FILL_0__1457_ (
);

FILL FILL_0__1037_ (
);

FILL FILL_2__986_ (
);

FILL FILL_1__1618_ (
);

MUX2X1 _960_ (
    .A(Xin12b[7]),
    .B(Xin12b[6]),
    .S(Stg_0_bF$buf3),
    .Y(_196_)
);

FILL FILL_1__1371_ (
);

FILL FILL_0__1686_ (
);

FILL FILL_0__1266_ (
);

FILL FILL_1__1427_ (
);

FILL FILL_1__1007_ (
);

FILL FILL_1__1180_ (
);

FILL FILL_0__1495_ (
);

FILL FILL_0__1075_ (
);

FILL FILL_1__1656_ (
);

FILL FILL_1__1236_ (
);

FILL FILL_2__1725_ (
);

FILL FILL_2__1305_ (
);

NOR3X1 _1723_ (
    .A(_96_),
    .B(_101_),
    .C(_86_),
    .Y(_102_)
);

NOR2X1 _1303_ (
    .A(_518_),
    .B(_522_),
    .Y(_523_)
);

FILL FILL_1__1465_ (
);

FILL FILL_1__1045_ (
);

AOI21X1 _1532_ (
    .A(_704_),
    .B(_705_),
    .C(_192_),
    .Y(_706_)
);

OAI21X1 _1112_ (
    .A(_342_),
    .B(_341_),
    .C(Xin12b[4]),
    .Y(_343_)
);

INVX1 _863_ (
    .A(Acalc[10]),
    .Y(_106_)
);

FILL FILL_1__1694_ (
);

FILL FILL_1__1274_ (
);

FILL FILL_0__1589_ (
);

FILL FILL_0__1169_ (
);

FILL FILL_0__916_ (
);

INVX1 _919_ (
    .A(Xcalc[7]),
    .Y(_157_)
);

DFFPOSX1 _1761_ (
    .D(_33_),
    .CLK(clk_bF$buf6),
    .Q(Xin12b[5])
);

NAND2X1 _1341_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_558_),
    .Y(_559_)
);

FILL FILL_1__1083_ (
);

FILL FILL_2__910_ (
);

FILL FILL_2__1572_ (
);

FILL FILL_2__1152_ (
);

FILL FILL_0__1398_ (
);

FILL FILL_1__1559_ (
);

FILL FILL_1__1139_ (
);

NAND3X1 _1570_ (
    .A(_201__bF$buf6),
    .B(_741_),
    .C(_735_),
    .Y(_742_)
);

NAND2X1 _1150_ (
    .A(_378_),
    .B(_377_),
    .Y(_379_)
);

FILL FILL_1__932_ (
);

FILL FILL_0__1610_ (
);

FILL FILL_2__1628_ (
);

FILL FILL_2__1208_ (
);

AOI21X1 _1626_ (
    .A(_764_),
    .B(_765_),
    .C(_265_),
    .Y(_795_)
);

OAI21X1 _1206_ (
    .A(_432_),
    .B(_428_),
    .C(_408_),
    .Y(_10_)
);

FILL FILL_0__954_ (
);

MUX2X1 _957_ (
    .A(Xin1[1]),
    .B(Xin1[0]),
    .S(Stg_0_bF$buf1),
    .Y(_193_)
);

FILL FILL_1__1368_ (
);

NAND2X1 _1435_ (
    .A(Xin[0]),
    .B(_119_),
    .Y(_638_)
);

NOR2X1 _1015_ (
    .A(Xin0[0]),
    .B(_249_),
    .Y(_250_)
);

FILL FILL_1__1597_ (
);

FILL FILL_1__1177_ (
);

FILL FILL_1__970_ (
);

OAI21X1 _1664_ (
    .A(_831_),
    .B(_830_),
    .C(_644_),
    .Y(_832_)
);

NAND2X1 _1244_ (
    .A(_467_),
    .B(_468_),
    .Y(_469_)
);

FILL FILL_0__992_ (
);

OR2X2 _995_ (
    .A(_229_),
    .B(_181_),
    .Y(_231_)
);

FILL FILL_0__1704_ (
);

FILL FILL_2__1475_ (
);

FILL FILL_2__1055_ (
);

OAI21X1 _1473_ (
    .A(_590_),
    .B(_629_),
    .C(_657_),
    .Y(_52_)
);

OAI21X1 _1053_ (
    .A(Stg_0_bF$buf0),
    .B(Yin12b[8]),
    .C(_285_),
    .Y(_286_)
);

FILL FILL_0__1513_ (
);

NOR2X1 _1529_ (
    .A(_673_),
    .B(_702_),
    .Y(_703_)
);

NAND3X1 _1109_ (
    .A(_201__bF$buf1),
    .B(_339_),
    .C(_332_),
    .Y(_340_)
);

NAND2X1 _1282_ (
    .A(Acalc[2]),
    .B(_188__bF$buf1),
    .Y(_503_)
);

FILL FILL_0__1322_ (
);

DFFPOSX1 _1758_ (
    .D(_30_),
    .CLK(clk_bF$buf4),
    .Q(Xin12b[6])
);

INVX1 _1338_ (
    .A(_555_),
    .Y(_556_)
);

OAI21X1 _1091_ (
    .A(Ain12b_11_bF$buf0),
    .B(_321_),
    .C(_322_),
    .Y(_323_)
);

FILL FILL_1__873_ (
);

FILL FILL_0__1551_ (
);

FILL FILL_2__1569_ (
);

FILL FILL_0__1131_ (
);

FILL FILL_2__1149_ (
);

FILL FILL_1__1712_ (
);

OAI21X1 _1567_ (
    .A(Stg_1_bF$buf3),
    .B(_675_),
    .C(_738_),
    .Y(_739_)
);

INVX1 _1147_ (
    .A(_375_),
    .Y(_376_)
);

FILL FILL_0__895_ (
);

FILL FILL_1__929_ (
);

INVX1 _898_ (
    .A(Ycalc[9]),
    .Y(_138_)
);

FILL FILL_0__1607_ (
);

FILL FILL_0__1360_ (
);

FILL FILL_1__1521_ (
);

FILL FILL_1__1101_ (
);

FILL FILL_2_BUFX2_insert42 (
);

FILL FILL_2_BUFX2_insert45 (
);

FILL FILL_2_BUFX2_insert47 (
);

DFFPOSX1 _1796_ (
    .D(LoadCtl[5]),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[6])
);

NAND2X1 _1376_ (
    .A(_590_),
    .B(_587_),
    .Y(_591_)
);

FILL FILL_0__1416_ (
);

FILL FILL_1__1330_ (
);

NAND2X1 _1185_ (
    .A(_410_),
    .B(_411_),
    .Y(_412_)
);

FILL FILL_1__967_ (
);

FILL FILL_0__1645_ (
);

FILL FILL_0__1225_ (
);

FILL FILL88650x25350 (
);

FILL FILL_0__989_ (
);

FILL FILL_0__1454_ (
);

FILL FILL_0__1034_ (
);

FILL FILL_2__983_ (
);

FILL FILL_1__1615_ (
);

FILL FILL_0__1683_ (
);

FILL FILL_0__1263_ (
);

FILL FILL_1__1424_ (
);

FILL FILL_1__1004_ (
);

NAND3X1 _1699_ (
    .A(_311_),
    .B(_75_),
    .C(_78_),
    .Y(_79_)
);

NAND2X1 _1279_ (
    .A(_487_),
    .B(_499_),
    .Y(_501_)
);

FILL FILL_0__1319_ (
);

FILL FILL_0__1492_ (
);

FILL FILL_0__1072_ (
);

FILL FILL_1__1653_ (
);

FILL FILL_1__1233_ (
);

NAND3X1 _1088_ (
    .A(_201__bF$buf0),
    .B(_319_),
    .C(_310_),
    .Y(_320_)
);

FILL FILL_2__1722_ (
);

FILL FILL_2__1302_ (
);

FILL FILL_0__1548_ (
);

FILL FILL_0__1128_ (
);

FILL FILL_1__1709_ (
);

OR2X2 _1720_ (
    .A(_97_),
    .B(_475_),
    .Y(_99_)
);

NAND2X1 _1300_ (
    .A(_201__bF$buf3),
    .B(_519_),
    .Y(_520_)
);

FILL FILL_1__1462_ (
);

FILL FILL_1__1042_ (
);

FILL FILL_0__1357_ (
);

FILL FILL_1__1518_ (
);

FILL FILL_1__1691_ (
);

FILL FILL_1__1271_ (
);

FILL FILL_0__1586_ (
);

FILL FILL_0__1166_ (
);

FILL FILL_0__913_ (
);

INVX1 _916_ (
    .A(Xcalc[11]),
    .Y(_154_)
);

FILL FILL_1__1327_ (
);

FILL FILL_1__1080_ (
);

FILL FILL_0__1395_ (
);

BUFX2 _1814_ (
    .A(_862_[0]),
    .Y(Yout[0])
);

FILL FILL_1__1556_ (
);

FILL FILL_1__1136_ (
);

FILL FILL_2__1625_ (
);

FILL FILL_2__1205_ (
);

AND2X2 _1623_ (
    .A(_749_),
    .B(_746_),
    .Y(_792_)
);

AOI21X1 _1203_ (
    .A(_411_),
    .B(_410_),
    .C(_429_),
    .Y(_430_)
);

FILL FILL_0__951_ (
);

NOR2X1 _954_ (
    .A(Stg_0_bF$buf6),
    .B(Stg_1_bF$buf1),
    .Y(_190_)
);

FILL FILL_1__1365_ (
);

OAI21X1 _1432_ (
    .A(_175_),
    .B(_635_),
    .C(_636_),
    .Y(_32_)
);

MUX2X1 _1012_ (
    .A(_246_),
    .B(_243_),
    .S(_164__bF$buf4),
    .Y(_247_)
);

FILL FILL_1__1594_ (
);

FILL FILL_1__1174_ (
);

FILL FILL_0__1489_ (
);

FILL FILL_0__1069_ (
);

NAND3X1 _1661_ (
    .A(_201__bF$buf5),
    .B(_828_),
    .C(_824_),
    .Y(_829_)
);

OAI21X1 _1241_ (
    .A(_463_),
    .B(_465_),
    .C(_462_),
    .Y(_466_)
);

NAND3X1 _992_ (
    .A(_200_),
    .B(_217_),
    .C(_225_),
    .Y(_228_)
);

FILL FILL_2__1719_ (
);

FILL FILL_0__1701_ (
);

FILL FILL_2__1472_ (
);

FILL FILL_2__1052_ (
);

FILL FILL_0__1298_ (
);

INVX1 _1717_ (
    .A(_81_),
    .Y(_96_)
);

FILL FILL_1__1459_ (
);

FILL FILL_1__1039_ (
);

NAND2X1 _1470_ (
    .A(Ain[1]),
    .B(_625_),
    .Y(_656_)
);

INVX1 _1050_ (
    .A(_282_),
    .Y(_283_)
);

FILL FILL_0__1510_ (
);

FILL FILL_2__1528_ (
);

FILL FILL88050x7350 (
);

NAND3X1 _1526_ (
    .A(Yin1[0]),
    .B(_679_),
    .C(_698_),
    .Y(_700_)
);

NAND2X1 _1106_ (
    .A(Stg_2_bF$buf4),
    .B(_336_),
    .Y(_337_)
);

FILL FILL_1__1688_ (
);

FILL FILL_1__1268_ (
);

DFFPOSX1 _1755_ (
    .D(_27_),
    .CLK(clk_bF$buf4),
    .Q(Xin12b[11])
);

INVX1 _1335_ (
    .A(Ain12b[5]),
    .Y(_553_)
);

FILL FILL_1__1497_ (
);

FILL FILL_1__1077_ (
);

FILL FILL_1__870_ (
);

FILL FILL_2__1566_ (
);

FILL FILL_2__1146_ (
);

NAND2X1 _1564_ (
    .A(Stg_0_bF$buf5),
    .B(Xin12b[11]),
    .Y(_736_)
);

AOI21X1 _1144_ (
    .A(_164__bF$buf3),
    .B(_334_),
    .C(_357_),
    .Y(_373_)
);

FILL FILL_0__892_ (
);

FILL FILL_1__926_ (
);

AOI22X1 _895_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Ycalc[0]),
    .C(_119_),
    .D(Ycalc[2]),
    .Y(_136_)
);

FILL FILL_0__1604_ (
);

FILL FILL_2__1375_ (
);

FILL FILL_0__948_ (
);

FILL FILL_2_BUFX2_insert11 (
);

DFFPOSX1 _1793_ (
    .D(LoadCtl[2]),
    .CLK(clk_bF$buf7),
    .Q(LoadCtl[3])
);

INVX1 _1373_ (
    .A(_587_),
    .Y(_588_)
);

FILL FILL_0__1413_ (
);

OAI21X1 _1429_ (
    .A(_209_),
    .B(_632_),
    .C(_634_),
    .Y(_31_)
);

INVX1 _1009_ (
    .A(Yin12b[4]),
    .Y(_244_)
);

NAND2X1 _1182_ (
    .A(_392_),
    .B(_404_),
    .Y(_409_)
);

FILL FILL_1__964_ (
);

FILL FILL_0__1642_ (
);

FILL FILL_0__1222_ (
);

INVX1 _1658_ (
    .A(_800_),
    .Y(_826_)
);

OAI21X1 _1238_ (
    .A(_421_),
    .B(_445_),
    .C(_440_),
    .Y(_463_)
);

FILL FILL_0__986_ (
);

OAI21X1 _989_ (
    .A(Ain12b_11_bF$buf4),
    .B(_199_),
    .C(_224_),
    .Y(_225_)
);

FILL FILL_2__1469_ (
);

FILL FILL_0__1451_ (
);

FILL FILL_2__1049_ (
);

FILL FILL_0__1031_ (
);

FILL FILL88650x46950 (
);

FILL FILL_2__980_ (
);

FILL FILL_1__1612_ (
);

OAI21X1 _1467_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_200_),
    .C(_654_),
    .Y(_49_)
);

OAI21X1 _1047_ (
    .A(_188__bF$buf1),
    .B(_280_),
    .C(_254_),
    .Y(_3_)
);

FILL FILL87450x61350 (
);

FILL FILL_0__1507_ (
);

FILL FILL_0__1680_ (
);

FILL FILL_0__1260_ (
);

FILL FILL_1__1421_ (
);

FILL FILL_1__1001_ (
);

NAND2X1 _1696_ (
    .A(_844_),
    .B(_842_),
    .Y(_76_)
);

NAND2X1 _1276_ (
    .A(Ain0[1]),
    .B(_496_),
    .Y(_498_)
);

FILL FILL_0__1316_ (
);

FILL FILL_1__1650_ (
);

FILL FILL_1__1230_ (
);

NAND2X1 _1085_ (
    .A(_258_),
    .B(_292_),
    .Y(_317_)
);

FILL FILL_1__867_ (
);

FILL FILL_0__1545_ (
);

FILL FILL_0__1125_ (
);

FILL FILL_1__1706_ (
);

FILL FILL_0__889_ (
);

FILL FILL_0__1354_ (
);

FILL FILL_2__883_ (
);

FILL FILL_1__1515_ (
);

FILL FILL_0__1583_ (
);

FILL FILL_0__1163_ (
);

FILL FILL_0__910_ (
);

AOI21X1 _913_ (
    .A(_109_),
    .B(_148_),
    .C(_151_),
    .Y(_152_)
);

FILL FILL_1__1324_ (
);

AOI21X1 _1599_ (
    .A(_756_),
    .B(_749_),
    .C(_769_),
    .Y(_770_)
);

AOI21X1 _1179_ (
    .A(_393_),
    .B(_405_),
    .C(_185_),
    .Y(_407_)
);

FILL FILL_2__1813_ (
);

FILL FILL_0__1639_ (
);

FILL FILL_0__1219_ (
);

FILL FILL_0__1392_ (
);

BUFX2 _1811_ (
    .A(LoadCtl_6_bF$buf0),
    .Y(Vld)
);

FILL FILL_1__1553_ (
);

FILL FILL_1__1133_ (
);

FILL FILL_2__1622_ (
);

FILL FILL_2__1202_ (
);

FILL FILL_0__1448_ (
);

FILL FILL_0__1028_ (
);

FILL FILL_2__977_ (
);

FILL FILL_1__1609_ (
);

OAI21X1 _1620_ (
    .A(_786_),
    .B(_788_),
    .C(_789_),
    .Y(_790_)
);

OR2X2 _1200_ (
    .A(_412_),
    .B(_426_),
    .Y(_427_)
);

OAI21X1 _951_ (
    .A(_162_),
    .B(LoadCtl_6_bF$buf4),
    .C(_187_),
    .Y(_0_)
);

FILL FILL_1__1362_ (
);

FILL FILL_1__999_ (
);

FILL FILL_0__1677_ (
);

FILL FILL_0__1257_ (
);

FILL FILL_1__1418_ (
);

FILL FILL_1__1591_ (
);

FILL FILL_1__1171_ (
);

FILL FILL_0__1486_ (
);

FILL FILL_0__1066_ (
);

FILL FILL_1__1647_ (
);

FILL FILL_1__1227_ (
);

FILL FILL_0__1295_ (
);

OR2X2 _1714_ (
    .A(_93_),
    .B(_86_),
    .Y(_94_)
);

FILL FILL_1__1456_ (
);

FILL FILL_1__1036_ (
);

FILL FILL_2__1525_ (
);

FILL FILL_2__1105_ (
);

INVX1 _1523_ (
    .A(_678_),
    .Y(_697_)
);

OAI21X1 _1103_ (
    .A(Stg_0_bF$buf5),
    .B(_311_),
    .C(_333_),
    .Y(_334_)
);

FILL FILL_1__1685_ (
);

FILL FILL_1__1265_ (
);

FILL FILL_0__907_ (
);

DFFPOSX1 _1752_ (
    .D(_24_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[10])
);

NOR2X1 _1332_ (
    .A(_549_),
    .B(_547_),
    .Y(_550_)
);

FILL FILL_1__1494_ (
);

FILL FILL_1__1074_ (
);

FILL FILL_0__1389_ (
);

BUFX2 _1808_ (
    .A(_859_[0]),
    .Y(Aout[0])
);

OAI21X1 _1561_ (
    .A(_711_),
    .B(_732_),
    .C(_733_),
    .Y(_734_)
);

OAI22X1 _1141_ (
    .A(_158_),
    .B(LoadCtl_6_bF$buf2),
    .C(_370_),
    .D(_369_),
    .Y(_7_)
);

FILL FILL_1__923_ (
);

INVX1 _892_ (
    .A(Ycalc[4]),
    .Y(_133_)
);

FILL FILL_0__1601_ (
);

FILL FILL_2__1619_ (
);

FILL FILL_2__1372_ (
);

FILL FILL_0__1198_ (
);

NAND2X1 _1617_ (
    .A(_749_),
    .B(_768_),
    .Y(_787_)
);

FILL FILL_0__945_ (
);

OAI21X1 _948_ (
    .A(Stg_0_bF$buf4),
    .B(_184_),
    .C(LoadCtl_6_bF$buf2),
    .Y(_185_)
);

FILL FILL_1__1359_ (
);

DFFPOSX1 _1790_ (
    .D(Rdy),
    .CLK(clk_bF$buf4),
    .Q(LoadCtl[0])
);

NAND2X1 _1370_ (
    .A(Acalc[8]),
    .B(_188__bF$buf4),
    .Y(_585_)
);

FILL FILL_0__1410_ (
);

NAND2X1 _1426_ (
    .A(Xin[0]),
    .B(_632_),
    .Y(_633_)
);

INVX1 _1006_ (
    .A(Yin12b[6]),
    .Y(_241_)
);

FILL FILL_1__1588_ (
);

FILL FILL_1__1168_ (
);

FILL FILL_1__961_ (
);

OAI21X1 _1655_ (
    .A(_822_),
    .B(_788_),
    .C(_819_),
    .Y(_823_)
);

NOR2X1 _1235_ (
    .A(_454_),
    .B(_452_),
    .Y(_460_)
);

FILL FILL_0__983_ (
);

MUX2X1 _986_ (
    .A(Xin12b[6]),
    .B(Xin12b[5]),
    .S(Stg_0_bF$buf4),
    .Y(_222_)
);

FILL FILL_1__1397_ (
);

FILL FILL_2__1466_ (
);

FILL FILL_2__1046_ (
);

NAND2X1 _1464_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Yin[0]),
    .Y(_653_)
);

INVX1 _1044_ (
    .A(_275_),
    .Y(_278_)
);

FILL FILL_0__1504_ (
);

INVX1 _1693_ (
    .A(_858_),
    .Y(_73_)
);

OAI21X1 _1273_ (
    .A(Ain12b_11_bF$buf2),
    .B(_486_),
    .C(_494_),
    .Y(_495_)
);

FILL FILL_0__1313_ (
);

DFFPOSX1 _1749_ (
    .D(_21_),
    .CLK(clk_bF$buf3),
    .Q(Acalc[7])
);

INVX1 _1329_ (
    .A(_546_),
    .Y(_547_)
);

FILL FILL88350x79350 (
);

NAND2X1 _1082_ (
    .A(_164__bF$buf3),
    .B(_264_),
    .Y(_314_)
);

FILL FILL_1__864_ (
);

FILL FILL_0__1542_ (
);

FILL FILL_0__1122_ (
);

FILL FILL_1__1703_ (
);

INVX1 _1558_ (
    .A(_730_),
    .Y(_731_)
);

INVX1 _1138_ (
    .A(_367_),
    .Y(_368_)
);

FILL FILL_0__886_ (
);

NAND2X1 _889_ (
    .A(LoadCtl[4]),
    .B(Ycalc[8]),
    .Y(_130_)
);

FILL FILL_2__1369_ (
);

FILL FILL_0__1351_ (
);

FILL FILL_2__880_ (
);

FILL FILL_1__1512_ (
);

DFFPOSX1 _1787_ (
    .D(_59_),
    .CLK(clk_bF$buf7),
    .Q(Ain1[1])
);

OR2X2 _1367_ (
    .A(_573_),
    .B(_582_),
    .Y(_583_)
);

FILL FILL_0__1407_ (
);

FILL FILL_2__936_ (
);

FILL FILL_0__1580_ (
);

FILL FILL_0__1160_ (
);

INVX1 _910_ (
    .A(Xcalc[6]),
    .Y(_149_)
);

FILL FILL_1__1321_ (
);

INVX1 _1596_ (
    .A(_765_),
    .Y(_767_)
);

NAND3X1 _1176_ (
    .A(_209_),
    .B(_397_),
    .C(_403_),
    .Y(_404_)
);

FILL FILL_1__958_ (
);

FILL FILL88650x32550 (
);

FILL FILL_0__1636_ (
);

FILL FILL_0__1216_ (
);

FILL FILL_1__1550_ (
);

FILL FILL_1__1130_ (
);

FILL FILL_0__1445_ (
);

FILL FILL_0__1025_ (
);

FILL FILL_2__974_ (
);

FILL FILL_1__1606_ (
);

FILL FILL_1__996_ (
);

FILL FILL_0__1674_ (
);

FILL FILL_0__1254_ (
);

FILL FILL_1__1415_ (
);

FILL FILL_0__1483_ (
);

FILL FILL_0__1063_ (
);

FILL FILL_1__1644_ (
);

FILL FILL_1__1224_ (
);

AOI21X1 _1499_ (
    .A(_181_),
    .B(_228_),
    .C(_226_),
    .Y(_673_)
);

INVX1 _1079_ (
    .A(Yin12b[10]),
    .Y(_311_)
);

FILL FILL_0__1539_ (
);

FILL FILL_0__1119_ (
);

FILL FILL_0__1292_ (
);

NAND3X1 _1711_ (
    .A(_849_),
    .B(_853_),
    .C(_836_),
    .Y(_91_)
);

FILL FILL_1__1453_ (
);

FILL FILL_1__1033_ (
);

FILL FILL_2__1522_ (
);

FILL FILL_2__1102_ (
);

FILL FILL_0__1348_ (
);

FILL FILL_2__877_ (
);

FILL FILL_1__1509_ (
);

NAND2X1 _1520_ (
    .A(Stg_1_bF$buf0),
    .B(_211_),
    .Y(_694_)
);

AOI21X1 _1100_ (
    .A(_308_),
    .B(_326_),
    .C(_324_),
    .Y(_331_)
);

FILL FILL_1__1682_ (
);

FILL FILL_1__1262_ (
);

FILL FILL_1__899_ (
);

FILL FILL_0__1577_ (
);

FILL FILL_0__1157_ (
);

FILL FILL_0__904_ (
);

INVX1 _907_ (
    .A(Xcalc[10]),
    .Y(_146_)
);

FILL FILL_1__1318_ (
);

FILL FILL_1__1491_ (
);

FILL FILL_1__1071_ (
);

FILL FILL_0__1386_ (
);

DFFPOSX1 _1805_ (
    .D(_70_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[9])
);

FILL FILL_1__1547_ (
);

FILL FILL_1__1127_ (
);

FILL FILL_1__920_ (
);

FILL FILL_0__1195_ (
);

OAI21X1 _1614_ (
    .A(Ain12b_11_bF$buf1),
    .B(_779_),
    .C(_777_),
    .Y(_784_)
);

FILL FILL_0__942_ (
);

INVX1 _945_ (
    .A(_181_),
    .Y(_182_)
);

FILL FILL_1__1356_ (
);

FILL FILL_2__1425_ (
);

NAND2X1 _1423_ (
    .A(Xin[1]),
    .B(_629_),
    .Y(_631_)
);

OAI21X1 _1003_ (
    .A(Stg_0_bF$buf2),
    .B(_163_),
    .C(_237_),
    .Y(_238_)
);

FILL FILL_1__1585_ (
);

FILL FILL_1__1165_ (
);

AND2X2 _1652_ (
    .A(_782_),
    .B(_785_),
    .Y(_820_)
);

OAI21X1 _1232_ (
    .A(_456_),
    .B(_453_),
    .C(Xin12b[10]),
    .Y(_457_)
);

FILL FILL_0__980_ (
);

MUX2X1 _983_ (
    .A(Xin1[0]),
    .B(Xin0[1]),
    .S(Stg_0_bF$buf6),
    .Y(_219_)
);

FILL FILL_1__1394_ (
);

FILL FILL_2__1043_ (
);

FILL FILL88050x57750 (
);

FILL FILL_0__1289_ (
);

OAI21X1 _1708_ (
    .A(_785_),
    .B(_806_),
    .C(_821_),
    .Y(_88_)
);

OAI21X1 _1461_ (
    .A(_234_),
    .B(_119_),
    .C(_651_),
    .Y(_46_)
);

NAND3X1 _1041_ (
    .A(_205_),
    .B(_272_),
    .C(_270_),
    .Y(_275_)
);

FILL FILL_2__1519_ (
);

FILL FILL_0__1501_ (
);

FILL FILL_2__1692_ (
);

FILL FILL_2__1272_ (
);

FILL FILL_0__1098_ (
);

NAND2X1 _1517_ (
    .A(_164__bF$buf2),
    .B(_207_),
    .Y(_691_)
);

FILL FILL_1__1679_ (
);

FILL FILL_1__1259_ (
);

OAI21X1 _1690_ (
    .A(_856_),
    .B(_855_),
    .C(_709_),
    .Y(_857_)
);

INVX2 _1270_ (
    .A(Stg_0_bF$buf4),
    .Y(_492_)
);

FILL FILL_0__1310_ (
);

DFFPOSX1 _1746_ (
    .D(_18_),
    .CLK(clk_bF$buf3),
    .Q(Acalc[4])
);

NAND2X1 _1326_ (
    .A(Acalc[5]),
    .B(_188__bF$buf3),
    .Y(_544_)
);

FILL FILL_1__1488_ (
);

FILL FILL_1__1068_ (
);

FILL FILL_1__1700_ (
);

NAND2X1 _1555_ (
    .A(_720_),
    .B(_727_),
    .Y(_728_)
);

OAI21X1 _1135_ (
    .A(Ain12b_11_bF$buf3),
    .B(_353_),
    .C(_359_),
    .Y(_365_)
);

FILL FILL_0__883_ (
);

FILL FILL_1__917_ (
);

AOI22X1 _886_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Acalc[1]),
    .C(_119_),
    .D(Acalc[3]),
    .Y(_128_)
);

FILL FILL_1__1297_ (
);

FILL FILL_2__1366_ (
);

FILL FILL_0__939_ (
);

DFFPOSX1 _1784_ (
    .D(_56_),
    .CLK(clk_bF$buf6),
    .Q(Ain12b[4])
);

NOR2X1 _1364_ (
    .A(Ain12b[7]),
    .B(_577_),
    .Y(_580_)
);

FILL FILL_0__1404_ (
);

FILL FILL_2__933_ (
);

INVX1 _1593_ (
    .A(_763_),
    .Y(_764_)
);

INVX1 _1173_ (
    .A(_396_),
    .Y(_401_)
);

FILL FILL_1__955_ (
);

FILL FILL_0__1633_ (
);

FILL FILL_0__1213_ (
);

INVX1 _1649_ (
    .A(Ycalc[8]),
    .Y(_817_)
);

INVX1 _1229_ (
    .A(_449_),
    .Y(_454_)
);

FILL FILL_0__977_ (
);

FILL FILL_0__1442_ (
);

FILL FILL_0__1022_ (
);

FILL FILL_1__1603_ (
);

NAND2X1 _1458_ (
    .A(Yin[1]),
    .B(_635_),
    .Y(_650_)
);

NAND3X1 _1038_ (
    .A(_201__bF$buf3),
    .B(_271_),
    .C(_249_),
    .Y(_272_)
);

FILL FILL_1__993_ (
);

FILL FILL_2__1689_ (
);

FILL FILL_0__1671_ (
);

FILL FILL_2__1269_ (
);

FILL FILL_0__1251_ (
);

FILL FILL_1__1412_ (
);

AND2X2 _1687_ (
    .A(_853_),
    .B(_849_),
    .Y(_854_)
);

NAND2X1 _1267_ (
    .A(Acalc[0]),
    .B(_188__bF$buf0),
    .Y(_490_)
);

FILL FILL_0__1727_ (
);

FILL FILL_0__1307_ (
);

FILL FILL_0__1480_ (
);

FILL FILL_0__1060_ (
);

FILL FILL_1__1641_ (
);

FILL FILL_1__1221_ (
);

NAND2X1 _1496_ (
    .A(LoadCtl_6_bF$buf1),
    .B(ISin),
    .Y(_671_)
);

OAI21X1 _1076_ (
    .A(_282_),
    .B(_302_),
    .C(_300_),
    .Y(_308_)
);

FILL FILL_0__1536_ (
);

FILL FILL_0__1116_ (
);

FILL FILL_1__1450_ (
);

FILL FILL_1__1030_ (
);

FILL FILL_0__1345_ (
);

FILL FILL_2__874_ (
);

FILL FILL_1__1506_ (
);

FILL FILL_1__896_ (
);

FILL FILL_0__1574_ (
);

FILL FILL_0__1154_ (
);

FILL FILL_0__901_ (
);

AOI21X1 _904_ (
    .A(_109_),
    .B(_140_),
    .C(_143_),
    .Y(_144_)
);

FILL FILL_1__1315_ (
);

FILL FILL_0__1383_ (
);

DFFPOSX1 _1802_ (
    .D(_67_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[6])
);

FILL FILL_1__1544_ (
);

FILL FILL_1__1124_ (
);

OAI21X1 _1399_ (
    .A(_609_),
    .B(_589_),
    .C(_608_),
    .Y(_612_)
);

FILL FILL_0__1439_ (
);

FILL FILL_0__1019_ (
);

FILL FILL_0__1192_ (
);

OAI21X1 _1611_ (
    .A(Ain12b_11_bF$buf1),
    .B(_779_),
    .C(_780_),
    .Y(_781_)
);

MUX2X1 _942_ (
    .A(_178_),
    .B(_171_),
    .S(Stg_2_bF$buf2),
    .Y(_179_)
);

FILL FILL_1__1353_ (
);

FILL FILL_2__1422_ (
);

FILL FILL_2__1002_ (
);

FILL FILL_0__1668_ (
);

FILL FILL_0__1248_ (
);

FILL FILL_1__1409_ (
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert16 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert17 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert18 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert19 (
    .A(clk),
    .Y(clk_bF$buf0)
);

AND2X2 _1420_ (
    .A(_628_),
    .B(_109_),
    .Y(_629_)
);

NAND2X1 _1000_ (
    .A(Stg_0_bF$buf2),
    .B(Yin1[1]),
    .Y(_235_)
);

FILL FILL_1__1582_ (
);

FILL FILL_1__1162_ (
);

FILL FILL_0__1477_ (
);

FILL FILL_0__1057_ (
);

FILL FILL_1__1638_ (
);

FILL FILL_1__1218_ (
);

MUX2X1 _980_ (
    .A(_215_),
    .B(_208_),
    .S(Stg_2_bF$buf1),
    .Y(_216_)
);

FILL FILL_1__1391_ (
);

FILL FILL_0__1286_ (
);

NAND3X1 _1705_ (
    .A(_836_),
    .B(_854_),
    .C(_823_),
    .Y(_85_)
);

FILL FILL_1__1447_ (
);

FILL FILL_1__1027_ (
);

FILL FILL_2__1516_ (
);

FILL FILL_0__1095_ (
);

NAND2X1 _1514_ (
    .A(Stg_1_bF$buf0),
    .B(_174_),
    .Y(_688_)
);

FILL FILL_1__1676_ (
);

FILL FILL_1__1256_ (
);

DFFPOSX1 _1743_ (
    .D(_15_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[1])
);

INVX1 _1323_ (
    .A(_539_),
    .Y(_542_)
);

FILL FILL_1__1485_ (
);

FILL FILL_1__1065_ (
);

OAI21X1 _1552_ (
    .A(_164__bF$buf0),
    .B(_723_),
    .C(_724_),
    .Y(_725_)
);

OAI21X1 _1132_ (
    .A(Ain12b_11_bF$buf0),
    .B(_353_),
    .C(_361_),
    .Y(_362_)
);

FILL FILL_0__880_ (
);

FILL FILL_1__914_ (
);

NAND2X1 _883_ (
    .A(LoadCtl[2]),
    .B(Acalc[5]),
    .Y(_125_)
);

FILL FILL_1__1294_ (
);

FILL FILL_2__1363_ (
);

FILL FILL_0__1189_ (
);

NAND3X1 _1608_ (
    .A(_201__bF$buf5),
    .B(_777_),
    .C(_774_),
    .Y(_778_)
);

FILL FILL_0__936_ (
);

NAND2X1 _939_ (
    .A(Stg_0_bF$buf4),
    .B(Xin12b[5]),
    .Y(_176_)
);

DFFPOSX1 _1781_ (
    .D(_53_),
    .CLK(clk_bF$buf3),
    .Q(Ain12b[9])
);

INVX1 _1361_ (
    .A(_576_),
    .Y(_577_)
);

FILL FILL_0__1401_ (
);

FILL FILL_2__1419_ (
);

FILL FILL_2__930_ (
);

FILL FILL_2__1592_ (
);

NAND2X1 _1417_ (
    .A(Xin[1]),
    .B(_625_),
    .Y(_627_)
);

FILL FILL_1__1579_ (
);

FILL FILL_1__1159_ (
);

INVX1 _1590_ (
    .A(_760_),
    .Y(_761_)
);

INVX1 _1170_ (
    .A(_397_),
    .Y(_398_)
);

FILL FILL_1__952_ (
);

FILL FILL_0__1630_ (
);

FILL FILL_0__1210_ (
);

INVX1 _1646_ (
    .A(_814_),
    .Y(_815_)
);

INVX1 _1226_ (
    .A(_436_),
    .Y(_451_)
);

FILL FILL_0__974_ (
);

NAND2X1 _977_ (
    .A(Stg_0_bF$buf3),
    .B(Xin12b[6]),
    .Y(_213_)
);

FILL FILL_1__1388_ (
);

FILL FILL_1__1600_ (
);

OAI21X1 _1455_ (
    .A(_262_),
    .B(_632_),
    .C(_648_),
    .Y(_43_)
);

MUX2X1 _1035_ (
    .A(_268_),
    .B(_261_),
    .S(Stg_2_bF$buf2),
    .Y(_269_)
);

FILL FILL_1__1197_ (
);

FILL FILL_1__990_ (
);

FILL FILL_2__1686_ (
);

FILL FILL_2__1266_ (
);

OAI21X1 _1684_ (
    .A(_827_),
    .B(_824_),
    .C(_201__bF$buf2),
    .Y(_851_)
);

NOR2X1 _1264_ (
    .A(_483_),
    .B(_486_),
    .Y(_487_)
);

FILL FILL88350x86550 (
);

FILL FILL_0__1724_ (
);

FILL FILL_0__1304_ (
);

NAND2X1 _1493_ (
    .A(LoadCtl_0_bF$buf2),
    .B(Ain[1]),
    .Y(_669_)
);

OAI21X1 _1073_ (
    .A(_282_),
    .B(_305_),
    .C(_186_),
    .Y(_306_)
);

FILL FILL_0__1533_ (
);

FILL FILL_0__1113_ (
);

NAND2X1 _1549_ (
    .A(Stg_0_bF$buf5),
    .B(_458_),
    .Y(_722_)
);

OAI21X1 _1129_ (
    .A(Stg_2_bF$buf4),
    .B(_268_),
    .C(_358_),
    .Y(_359_)
);

FILL FILL_0__877_ (
);

FILL FILL_0__1342_ (
);

FILL FILL_1__1503_ (
);

DFFPOSX1 _1778_ (
    .D(_50_),
    .CLK(clk_bF$buf3),
    .Q(Ain12b[10])
);

NAND3X1 _1358_ (
    .A(_183__bF$buf3),
    .B(_492_),
    .C(_201__bF$buf3),
    .Y(_574_)
);

FILL FILL_1__893_ (
);

FILL FILL_2__927_ (
);

FILL FILL_0__1571_ (
);

FILL FILL_2__1589_ (
);

FILL FILL_0__1151_ (
);

FILL FILL_2__1169_ (
);

INVX1 _901_ (
    .A(Ycalc[7]),
    .Y(_141_)
);

FILL FILL_1__1312_ (
);

AOI21X1 _1587_ (
    .A(_164__bF$buf3),
    .B(_714_),
    .C(_757_),
    .Y(_758_)
);

NOR2X1 _1167_ (
    .A(_183__bF$buf2),
    .B(_356_),
    .Y(_395_)
);

FILL FILL_1__949_ (
);

FILL FILL_0__1627_ (
);

FILL FILL_0__1207_ (
);

FILL FILL87450x21750 (
);

FILL FILL_0__1380_ (
);

FILL FILL_1__1541_ (
);

FILL FILL_1__1121_ (
);

AND2X2 _1396_ (
    .A(_605_),
    .B(_609_),
    .Y(_610_)
);

FILL FILL_0__1436_ (
);

FILL FILL_0__1016_ (
);

FILL FILL88350x18150 (
);

FILL FILL_1__1350_ (
);

FILL FILL_1__987_ (
);

FILL FILL_0__1665_ (
);

FILL FILL_0__1245_ (
);

FILL FILL_1__1406_ (
);

FILL FILL87750x64950 (
);

FILL FILL_0__1474_ (
);

FILL FILL_0__1054_ (
);

FILL FILL_1__1635_ (
);

FILL FILL_1__1215_ (
);

FILL FILL_0__1283_ (
);

NAND2X1 _1702_ (
    .A(_81_),
    .B(_79_),
    .Y(_82_)
);

FILL FILL_1__1444_ (
);

FILL FILL_1__1024_ (
);

OAI21X1 _1299_ (
    .A(Stg_0_bF$buf6),
    .B(_164__bF$buf1),
    .C(Stg_2_bF$buf2),
    .Y(_519_)
);

FILL FILL_0__1339_ (
);

FILL FILL_0__1092_ (
);

NAND2X1 _1511_ (
    .A(_492_),
    .B(_175_),
    .Y(_685_)
);

FILL FILL_1__1673_ (
);

FILL FILL_1__1253_ (
);

FILL FILL_2__1322_ (
);

FILL FILL_0__1568_ (
);

FILL FILL_0__1148_ (
);

FILL FILL_1__1309_ (
);

DFFPOSX1 _1740_ (
    .D(_12_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[10])
);

OAI21X1 _1320_ (
    .A(_525_),
    .B(_517_),
    .C(_527_),
    .Y(_539_)
);

FILL FILL_1__1482_ (
);

FILL FILL_1__1062_ (
);

FILL FILL_0__1377_ (
);

FILL FILL_1__1538_ (
);

FILL FILL_1__1118_ (
);

FILL FILL_1__911_ (
);

NAND2X1 _880_ (
    .A(LoadCtl[4]),
    .B(Acalc[9]),
    .Y(_122_)
);

FILL FILL_1__1291_ (
);

FILL FILL_0__1186_ (
);

AOI21X1 _1605_ (
    .A(_164__bF$buf3),
    .B(_737_),
    .C(_757_),
    .Y(_775_)
);

FILL FILL_0__933_ (
);

NAND2X1 _936_ (
    .A(Stg_0_bF$buf3),
    .B(Xin12b[7]),
    .Y(_173_)
);

FILL FILL_1__1347_ (
);

FILL FILL_2__1416_ (
);

NOR2X1 _1414_ (
    .A(_117_),
    .B(_624_),
    .Y(_625_)
);

FILL FILL_1__1576_ (
);

FILL FILL_1__1156_ (
);

FILL FILL88050x64950 (
);

NAND2X1 _1643_ (
    .A(_810_),
    .B(_798_),
    .Y(_812_)
);

OAI21X1 _1223_ (
    .A(_433_),
    .B(LoadCtl_6_bF$buf1),
    .C(_448_),
    .Y(_11_)
);

FILL FILL_0__971_ (
);

NAND2X1 _974_ (
    .A(Stg_0_bF$buf3),
    .B(Xin12b[8]),
    .Y(_210_)
);

FILL FILL_1__1385_ (
);

NAND2X1 _1452_ (
    .A(Yin[0]),
    .B(_632_),
    .Y(_647_)
);

NAND2X1 _1032_ (
    .A(Stg_0_bF$buf0),
    .B(Yin12b[6]),
    .Y(_266_)
);

FILL FILL_1__1194_ (
);

FILL FILL_2__1683_ (
);

FILL FILL_2__1263_ (
);

FILL FILL_0__1089_ (
);

NAND3X1 _1508_ (
    .A(Stg_1_bF$buf2),
    .B(_681_),
    .C(_680_),
    .Y(_682_)
);

NAND3X1 _1681_ (
    .A(_201__bF$buf2),
    .B(_843_),
    .C(_847_),
    .Y(_848_)
);

INVX1 _1261_ (
    .A(_190_),
    .Y(_484_)
);

FILL FILL_0__1721_ (
);

FILL FILL_2__1319_ (
);

FILL FILL_0__1301_ (
);

DFFPOSX1 _1737_ (
    .D(_9_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[7])
);

NAND2X1 _1317_ (
    .A(Ain12b[4]),
    .B(_535_),
    .Y(_536_)
);

FILL FILL_1__1479_ (
);

FILL FILL_1__1059_ (
);

OAI21X1 _1490_ (
    .A(_660_),
    .B(_665_),
    .C(_667_),
    .Y(_59_)
);

NOR2X1 _1070_ (
    .A(_302_),
    .B(_301_),
    .Y(_303_)
);

FILL FILL_0__1530_ (
);

FILL FILL_0__1110_ (
);

OAI21X1 _1546_ (
    .A(_183__bF$buf0),
    .B(_716_),
    .C(_718_),
    .Y(_719_)
);

INVX1 _1126_ (
    .A(Yin12b[11]),
    .Y(_356_)
);

FILL FILL_0__874_ (
);

FILL FILL_1__908_ (
);

AOI22X1 _877_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Acalc[0]),
    .C(_119_),
    .D(Acalc[2]),
    .Y(_120_)
);

FILL FILL_1__1288_ (
);

FILL FILL_1__1500_ (
);

DFFPOSX1 _1775_ (
    .D(_47_),
    .CLK(clk_bF$buf1),
    .Q(Yin1[1])
);

OAI21X1 _1355_ (
    .A(_570_),
    .B(_562_),
    .C(LoadCtl_6_bF$buf4),
    .Y(_572_)
);

FILL FILL_1__1097_ (
);

FILL FILL_0__1815_ (
);

FILL FILL_1__890_ (
);

FILL FILL_2__924_ (
);

FILL FILL_2__1586_ (
);

FILL FILL_2__1166_ (
);

AOI21X1 _1584_ (
    .A(_751_),
    .B(_729_),
    .C(_750_),
    .Y(_755_)
);

AOI21X1 _1164_ (
    .A(_377_),
    .B(_378_),
    .C(_172_),
    .Y(_392_)
);

FILL FILL_1__946_ (
);

FILL FILL_0__1624_ (
);

FILL FILL_0__1204_ (
);

FILL FILL_0__968_ (
);

NAND2X1 _1393_ (
    .A(Ain12b_11_bF$buf2),
    .B(_606_),
    .Y(_607_)
);

FILL FILL_0__1433_ (
);

FILL FILL_0__1013_ (
);

OAI21X1 _1449_ (
    .A(_644_),
    .B(_629_),
    .C(_645_),
    .Y(_40_)
);

NAND2X1 _1029_ (
    .A(Stg_0_bF$buf0),
    .B(Yin12b[8]),
    .Y(_263_)
);

FILL FILL88350x72150 (
);

FILL FILL88350x39750 (
);

FILL FILL_1__984_ (
);

FILL FILL_0__1662_ (
);

FILL FILL_0__1242_ (
);

FILL FILL_1__1403_ (
);

OAI21X1 _1678_ (
    .A(Ain12b_11_bF$buf1),
    .B(_842_),
    .C(_844_),
    .Y(_845_)
);

NAND2X1 _1258_ (
    .A(_186_),
    .B(_481_),
    .Y(_482_)
);

FILL FILL_0__1718_ (
);

FILL FILL_0__1471_ (
);

FILL FILL_2__1489_ (
);

FILL FILL_0__1051_ (
);

FILL FILL_1__1632_ (
);

FILL FILL_1__1212_ (
);

OAI21X1 _1487_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_118_),
    .C(Ain1[0]),
    .Y(_666_)
);

NAND3X1 _1067_ (
    .A(Xin1[0]),
    .B(_299_),
    .C(_297_),
    .Y(_300_)
);

FILL FILL_0__1527_ (
);

FILL FILL_0__1107_ (
);

FILL FILL_0__1280_ (
);

FILL FILL_1__1441_ (
);

FILL FILL_1__1021_ (
);

NAND2X1 _1296_ (
    .A(_509_),
    .B(_514_),
    .Y(_516_)
);

FILL FILL_0__1336_ (
);

FILL FILL_1__1670_ (
);

FILL FILL_1__1250_ (
);

FILL FILL_1__887_ (
);

FILL FILL_0__1565_ (
);

FILL FILL_0__1145_ (
);

FILL FILL_1__1726_ (
);

FILL FILL_1__1306_ (
);

FILL FILL_0_BUFX2_insert30 (
);

FILL FILL_0_BUFX2_insert31 (
);

FILL FILL_0_BUFX2_insert32 (
);

FILL FILL_0_BUFX2_insert33 (
);

FILL FILL_0_BUFX2_insert34 (
);

FILL FILL_0_BUFX2_insert35 (
);

FILL FILL_0_BUFX2_insert36 (
);

FILL FILL_0_BUFX2_insert37 (
);

FILL FILL_0_BUFX2_insert38 (
);

FILL FILL_0_BUFX2_insert39 (
);

FILL FILL_0__1374_ (
);

FILL FILL_1__1535_ (
);

FILL FILL_1__1115_ (
);

FILL FILL_0__1183_ (
);

OAI21X1 _1602_ (
    .A(_770_),
    .B(_772_),
    .C(_709_),
    .Y(_773_)
);

FILL FILL_0__930_ (
);

OAI21X1 _933_ (
    .A(Stg_0_bF$buf6),
    .B(_168_),
    .C(_169_),
    .Y(_170_)
);

FILL FILL_1__1344_ (
);

AND2X2 _1199_ (
    .A(_421_),
    .B(_425_),
    .Y(_426_)
);

FILL FILL_2__1413_ (
);

FILL FILL_0__1659_ (
);

FILL FILL_0__1239_ (
);

OAI21X1 _1411_ (
    .A(_619_),
    .B(_615_),
    .C(_618_),
    .Y(_623_)
);

FILL FILL_1__1573_ (
);

FILL FILL_1__1153_ (
);

BUFX2 BUFX2_insert40 (
    .A(Stg[1]),
    .Y(Stg_1_bF$buf2)
);

BUFX2 BUFX2_insert41 (
    .A(Stg[1]),
    .Y(Stg_1_bF$buf1)
);

BUFX2 BUFX2_insert42 (
    .A(Stg[1]),
    .Y(Stg_1_bF$buf0)
);

BUFX2 BUFX2_insert43 (
    .A(_183_),
    .Y(_183__bF$buf3)
);

BUFX2 BUFX2_insert44 (
    .A(_183_),
    .Y(_183__bF$buf2)
);

BUFX2 BUFX2_insert45 (
    .A(_183_),
    .Y(_183__bF$buf1)
);

BUFX2 BUFX2_insert46 (
    .A(_183_),
    .Y(_183__bF$buf0)
);

BUFX2 BUFX2_insert47 (
    .A(Ain12b[11]),
    .Y(Ain12b_11_bF$buf4)
);

BUFX2 BUFX2_insert48 (
    .A(Ain12b[11]),
    .Y(Ain12b_11_bF$buf3)
);

BUFX2 BUFX2_insert49 (
    .A(Ain12b[11]),
    .Y(Ain12b_11_bF$buf2)
);

FILL FILL_2__1642_ (
);

FILL FILL_0__1468_ (
);

FILL FILL_0__1048_ (
);

FILL FILL_2__997_ (
);

FILL FILL_1__1629_ (
);

FILL FILL_1__1209_ (
);

AOI21X1 _1640_ (
    .A(_808_),
    .B(_807_),
    .C(_262_),
    .Y(_809_)
);

NOR3X1 _1220_ (
    .A(_434_),
    .B(_445_),
    .C(_430_),
    .Y(_446_)
);

OAI21X1 _971_ (
    .A(Stg_0_bF$buf6),
    .B(_205_),
    .C(_206_),
    .Y(_207_)
);

FILL FILL_1__1382_ (
);

FILL FILL_0__1697_ (
);

FILL FILL_0__1277_ (
);

FILL FILL_1__1438_ (
);

FILL FILL_1__1018_ (
);

FILL FILL_1__1191_ (
);

FILL FILL_2__1260_ (
);

FILL FILL_0__1086_ (
);

NAND3X1 _1505_ (
    .A(_201__bF$buf6),
    .B(_678_),
    .C(_674_),
    .Y(_679_)
);

FILL FILL_1__1667_ (
);

FILL FILL_1__1247_ (
);

FILL FILL_2__1316_ (
);

DFFPOSX1 _1734_ (
    .D(_6_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[4])
);

NAND3X1 _1314_ (
    .A(Stg_0_bF$buf1),
    .B(_183__bF$buf3),
    .C(_164__bF$buf1),
    .Y(_533_)
);

FILL FILL_1__1476_ (
);

FILL FILL_1__1056_ (
);

OAI21X1 _1543_ (
    .A(_164__bF$buf4),
    .B(_714_),
    .C(_715_),
    .Y(_716_)
);

NOR2X1 _1123_ (
    .A(_338_),
    .B(_332_),
    .Y(_353_)
);

FILL FILL_0__871_ (
);

FILL FILL_1__905_ (
);

INVX2 _874_ (
    .A(_116_),
    .Y(_117_)
);

FILL FILL_1__1285_ (
);

FILL FILL_0__927_ (
);

DFFPOSX1 _1772_ (
    .D(_44_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[4])
);

OAI21X1 _1352_ (
    .A(_564_),
    .B(_565_),
    .C(_568_),
    .Y(_569_)
);

FILL FILL_1__1094_ (
);

FILL FILL_0__1812_ (
);

FILL FILL_2__1583_ (
);

FILL FILL_2__1163_ (
);

OAI21X1 _1408_ (
    .A(_619_),
    .B(_615_),
    .C(LoadCtl_6_bF$buf0),
    .Y(_621_)
);

AOI21X1 _1581_ (
    .A(_752_),
    .B(_750_),
    .C(_192_),
    .Y(_753_)
);

OAI21X1 _1161_ (
    .A(_389_),
    .B(_388_),
    .C(_191_),
    .Y(_390_)
);

FILL FILL_1__943_ (
);

FILL FILL_2__1639_ (
);

FILL FILL_0__1621_ (
);

FILL FILL_0__1201_ (
);

FILL FILL_2__1219_ (
);

AOI21X1 _1637_ (
    .A(_805_),
    .B(_802_),
    .C(Yin12b[7]),
    .Y(_806_)
);

NOR2X1 _1217_ (
    .A(_436_),
    .B(_437_),
    .Y(_443_)
);

FILL FILL_0__965_ (
);

OAI21X1 _968_ (
    .A(Stg_0_bF$buf1),
    .B(_202_),
    .C(_203_),
    .Y(_204_)
);

FILL FILL_1__1379_ (
);

INVX1 _1390_ (
    .A(_589_),
    .Y(_604_)
);

FILL FILL_0__1430_ (
);

FILL FILL_0__1010_ (
);

OAI21X1 _1446_ (
    .A(_356_),
    .B(_625_),
    .C(_643_),
    .Y(_39_)
);

OAI21X1 _1026_ (
    .A(Stg_0_bF$buf2),
    .B(_200_),
    .C(_259_),
    .Y(_260_)
);

FILL FILL_1__1188_ (
);

FILL FILL_1__981_ (
);

FILL FILL_1__1400_ (
);

NOR2X1 _1675_ (
    .A(_827_),
    .B(_824_),
    .Y(_842_)
);

NAND2X1 _1255_ (
    .A(_478_),
    .B(_476_),
    .Y(_479_)
);

FILL FILL_0__1715_ (
);

FILL FILL_2__1486_ (
);

FILL FILL_2__1066_ (
);

OAI21X1 _1484_ (
    .A(_553_),
    .B(_635_),
    .C(_663_),
    .Y(_57_)
);

OR2X2 _1064_ (
    .A(_296_),
    .B(_295_),
    .Y(_297_)
);

FILL FILL_0__1524_ (
);

FILL FILL_0__1104_ (
);

FILL FILL_0__868_ (
);

NAND2X1 _1293_ (
    .A(_512_),
    .B(_505_),
    .Y(_514_)
);

FILL FILL_0__1333_ (
);

DFFPOSX1 _1769_ (
    .D(_41_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[9])
);

NOR2X1 _1349_ (
    .A(_564_),
    .B(_565_),
    .Y(_566_)
);

FILL FILL_0__1809_ (
);

FILL FILL_1__884_ (
);

FILL FILL_0__1562_ (
);

FILL FILL_0__1142_ (
);

FILL FILL_1__1723_ (
);

FILL FILL_1__1303_ (
);

NAND2X1 _1578_ (
    .A(_746_),
    .B(_749_),
    .Y(_750_)
);

OAI21X1 _1158_ (
    .A(_331_),
    .B(_383_),
    .C(_386_),
    .Y(_387_)
);

FILL FILL_0__1618_ (
);

FILL FILL_0__1371_ (
);

FILL FILL88350x25350 (
);

FILL FILL_1__1532_ (
);

FILL FILL_1__1112_ (
);

OAI21X1 _1387_ (
    .A(_592_),
    .B(_601_),
    .C(LoadCtl_6_bF$buf0),
    .Y(_602_)
);

FILL FILL_0__1427_ (
);

FILL FILL_0__1007_ (
);

FILL FILL_0__1180_ (
);

OAI21X1 _930_ (
    .A(Stg_0_bF$buf1),
    .B(_165_),
    .C(_166_),
    .Y(_167_)
);

FILL FILL_1__1341_ (
);

NAND3X1 _1196_ (
    .A(_201__bF$buf4),
    .B(_418_),
    .C(_413_),
    .Y(_423_)
);

FILL FILL_1__978_ (
);

FILL FILL_0__1656_ (
);

FILL FILL_0__1236_ (
);

FILL FILL_1__1570_ (
);

FILL FILL_1__1150_ (
);

BUFX2 BUFX2_insert10 (
    .A(_188_),
    .Y(_188__bF$buf1)
);

BUFX2 BUFX2_insert11 (
    .A(_188_),
    .Y(_188__bF$buf0)
);

FILL FILL_0__1465_ (
);

FILL FILL_0__1045_ (
);

FILL FILL_2__994_ (
);

FILL FILL_1__1626_ (
);

FILL FILL_1__1206_ (
);

FILL FILL_0__1694_ (
);

FILL FILL_0__1274_ (
);

FILL FILL_1__1435_ (
);

FILL FILL_1__1015_ (
);

FILL FILL_0__1083_ (
);

MUX2X1 _1502_ (
    .A(_675_),
    .B(_196_),
    .S(Stg_1_bF$buf3),
    .Y(_676_)
);

FILL FILL_1__1664_ (
);

FILL FILL_1__1244_ (
);

OAI21X1 _1099_ (
    .A(_188__bF$buf1),
    .B(_330_),
    .C(_307_),
    .Y(_5_)
);

FILL FILL_2__1313_ (
);

FILL FILL_0__1559_ (
);

FILL FILL_0__1139_ (
);

DFFPOSX1 _1731_ (
    .D(_3_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[1])
);

OAI21X1 _1311_ (
    .A(_188__bF$buf0),
    .B(_529_),
    .C(_530_),
    .Y(_17_)
);

FILL FILL_1__1473_ (
);

FILL FILL_1__1053_ (
);

FILL FILL_0__1368_ (
);

FILL FILL_2__897_ (
);

FILL FILL_1__1529_ (
);

FILL FILL_1__1109_ (
);

NAND2X1 _1540_ (
    .A(Stg_0_bF$buf5),
    .B(Xin12b[10]),
    .Y(_713_)
);

NAND2X1 _1120_ (
    .A(_350_),
    .B(_349_),
    .Y(_351_)
);

FILL FILL_1__902_ (
);

OAI21X1 _871_ (
    .A(_110_),
    .B(_113_),
    .C(_111_),
    .Y(_114_)
);

FILL FILL_1__1282_ (
);

FILL FILL_0__1597_ (
);

FILL FILL_0__1177_ (
);

FILL FILL_0__924_ (
);

INVX8 _927_ (
    .A(Stg_1_bF$buf0),
    .Y(_164_)
);

FILL FILL_1__1338_ (
);

FILL FILL_1__1091_ (
);

FILL FILL_2__1580_ (
);

FILL FILL_2__1160_ (
);

NAND2X1 _1405_ (
    .A(Ain12b[10]),
    .B(_201__bF$buf0),
    .Y(_618_)
);

FILL FILL_1__1567_ (
);

FILL FILL_1__1147_ (
);

FILL FILL_1__940_ (
);

FILL FILL_2__1636_ (
);

FILL FILL_2__1216_ (
);

INVX1 _1634_ (
    .A(_801_),
    .Y(_803_)
);

NAND3X1 _1214_ (
    .A(Xin12b[9]),
    .B(_438_),
    .C(_439_),
    .Y(_440_)
);

FILL FILL_0__962_ (
);

INVX8 _965_ (
    .A(Ain12b_11_bF$buf0),
    .Y(_201_)
);

FILL FILL_1__1376_ (
);

NAND2X1 _1443_ (
    .A(Yin[0]),
    .B(_625_),
    .Y(_642_)
);

NAND2X1 _1023_ (
    .A(Stg_0_bF$buf2),
    .B(Yin12b[4]),
    .Y(_257_)
);

FILL FILL_1__1185_ (
);

AOI22X1 _1672_ (
    .A(_817_),
    .B(_188__bF$buf2),
    .C(_839_),
    .D(_815_),
    .Y(_69_)
);

OAI21X1 _1252_ (
    .A(Ain12b_11_bF$buf3),
    .B(_459_),
    .C(_475_),
    .Y(_476_)
);

FILL FILL_0__1712_ (
);

FILL FILL_2__1483_ (
);

FILL FILL_2__1063_ (
);

DFFPOSX1 _1728_ (
    .D(_0_),
    .CLK(clk_bF$buf5),
    .Q(Ycalc[0])
);

NAND3X1 _1308_ (
    .A(_527_),
    .B(_524_),
    .C(_516_),
    .Y(_528_)
);

NAND2X1 _1481_ (
    .A(Ain[0]),
    .B(_635_),
    .Y(_662_)
);

NAND2X1 _1061_ (
    .A(_291_),
    .B(_293_),
    .Y(_294_)
);

FILL FILL_0__1521_ (
);

FILL FILL_2__1539_ (
);

FILL FILL_2__1119_ (
);

FILL FILL_0__1101_ (
);

OAI21X1 _1537_ (
    .A(_699_),
    .B(_673_),
    .C(_700_),
    .Y(_710_)
);

INVX1 _1117_ (
    .A(_347_),
    .Y(_348_)
);

FILL FILL_0__865_ (
);

NAND2X1 _868_ (
    .A(LoadCtl[2]),
    .B(Acalc[4]),
    .Y(_111_)
);

FILL FILL_1__1699_ (
);

FILL FILL_1__1279_ (
);

NAND2X1 _1290_ (
    .A(_509_),
    .B(_510_),
    .Y(_511_)
);

FILL FILL_0__1330_ (
);

DFFPOSX1 _1766_ (
    .D(_38_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[10])
);

OAI21X1 _1346_ (
    .A(Stg_2_bF$buf2),
    .B(_485_),
    .C(_191_),
    .Y(_563_)
);

FILL FILL_1__1088_ (
);

FILL FILL_1__881_ (
);

FILL FILL_1__1720_ (
);

FILL FILL_1_CLKBUF1_insert12 (
);

FILL FILL_1__1300_ (
);

FILL FILL_1_CLKBUF1_insert13 (
);

FILL FILL_1_CLKBUF1_insert14 (
);

FILL FILL_1_CLKBUF1_insert15 (
);

FILL FILL_1_CLKBUF1_insert16 (
);

FILL FILL_1_CLKBUF1_insert17 (
);

FILL FILL_1_CLKBUF1_insert18 (
);

FILL FILL_1_CLKBUF1_insert19 (
);

INVX1 _1575_ (
    .A(_742_),
    .Y(_747_)
);

INVX1 _1155_ (
    .A(_343_),
    .Y(_384_)
);

FILL FILL_1__937_ (
);

FILL FILL_0__1615_ (
);

FILL FILL_2__1386_ (
);

FILL FILL_0__959_ (
);

OAI21X1 _1384_ (
    .A(_598_),
    .B(_542_),
    .C(_597_),
    .Y(_599_)
);

FILL FILL_0__1424_ (
);

FILL FILL_0__1004_ (
);

FILL FILL88350x46950 (
);

NAND2X1 _1193_ (
    .A(_418_),
    .B(_419_),
    .Y(_420_)
);

FILL FILL_1__975_ (
);

FILL FILL_0__1653_ (
);

FILL FILL_0__1233_ (
);

FILL FILL_1__1814_ (
);

AND2X2 _1669_ (
    .A(_823_),
    .B(_836_),
    .Y(_837_)
);

NAND2X1 _1249_ (
    .A(Xin12b[11]),
    .B(_356_),
    .Y(_473_)
);

FILL FILL_0__997_ (
);

FILL FILL_0__1709_ (
);

FILL FILL_0__1462_ (
);

FILL FILL_0__1042_ (
);

FILL FILL_2__991_ (
);

FILL FILL_1__1623_ (
);

FILL FILL_1__1203_ (
);

INVX1 _1478_ (
    .A(Ain[1]),
    .Y(_660_)
);

NAND2X1 _1058_ (
    .A(_246_),
    .B(_290_),
    .Y(_291_)
);

FILL FILL_0__1518_ (
);

FILL FILL_0__1691_ (
);

FILL FILL_0__1271_ (
);

FILL FILL_1__1432_ (
);

FILL FILL_1__1012_ (
);

OAI21X1 _1287_ (
    .A(Stg_2_bF$buf0),
    .B(_506_),
    .C(_507_),
    .Y(_508_)
);

FILL FILL_0__1327_ (
);

FILL FILL_1_BUFX2_insert40 (
);

FILL FILL_1_BUFX2_insert41 (
);

FILL FILL_1_BUFX2_insert42 (
);

FILL FILL_1_BUFX2_insert43 (
);

FILL FILL_1_BUFX2_insert44 (
);

FILL FILL_1_BUFX2_insert45 (
);

FILL FILL_1_BUFX2_insert46 (
);

FILL FILL_1_BUFX2_insert47 (
);

FILL FILL_1_BUFX2_insert48 (
);

FILL FILL_1_BUFX2_insert49 (
);

FILL FILL_0__1080_ (
);

FILL FILL_1__1661_ (
);

FILL FILL_1__1241_ (
);

OR2X2 _1096_ (
    .A(_327_),
    .B(_309_),
    .Y(_328_)
);

FILL FILL_1__878_ (
);

FILL FILL_0__1556_ (
);

FILL FILL_0__1136_ (
);

FILL FILL_1__1717_ (
);

FILL FILL_1__1470_ (
);

FILL FILL_1__1050_ (
);

FILL FILL_0__1365_ (
);

FILL FILL_2__894_ (
);

FILL FILL_1__1526_ (
);

FILL FILL_1__1106_ (
);

FILL FILL_0__1594_ (
);

FILL FILL_0__1174_ (
);

FILL FILL_0__921_ (
);

OAI21X1 _924_ (
    .A(_117_),
    .B(_160_),
    .C(_161_),
    .Y(_861_[1])
);

FILL FILL_1__1335_ (
);

FILL FILL88650x54150 (
);

AOI21X1 _1402_ (
    .A(_599_),
    .B(_614_),
    .C(_612_),
    .Y(_615_)
);

FILL FILL_1__1564_ (
);

FILL FILL_1__1144_ (
);

FILL FILL_2__1633_ (
);

FILL FILL_2__1213_ (
);

FILL FILL_0__1459_ (
);

FILL FILL_0__1039_ (
);

FILL FILL_2__988_ (
);

NOR2X1 _1631_ (
    .A(_183__bF$buf2),
    .B(_471_),
    .Y(_800_)
);

OAI21X1 _1211_ (
    .A(_416_),
    .B(_413_),
    .C(_201__bF$buf4),
    .Y(_437_)
);

MUX2X1 _962_ (
    .A(_197_),
    .B(_196_),
    .S(_164__bF$buf0),
    .Y(_198_)
);

FILL FILL_1__1373_ (
);

FILL FILL_0__1688_ (
);

FILL FILL_0__1268_ (
);

FILL FILL_1__1429_ (
);

FILL FILL_1__1009_ (
);

OAI21X1 _1440_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_168_),
    .C(_640_),
    .Y(_36_)
);

NAND2X1 _1020_ (
    .A(Xcalc[1]),
    .B(_188__bF$buf0),
    .Y(_254_)
);

FILL FILL_1__1182_ (
);

FILL FILL_0__1497_ (
);

FILL FILL_0__1077_ (
);

FILL FILL_1__1658_ (
);

FILL FILL_1__1238_ (
);

FILL FILL_2__1480_ (
);

FILL FILL_2__1060_ (
);

OAI21X1 _1725_ (
    .A(_100_),
    .B(_103_),
    .C(_191_),
    .Y(_104_)
);

INVX1 _1305_ (
    .A(_524_),
    .Y(_525_)
);

FILL FILL_1__1467_ (
);

FILL FILL_1__1047_ (
);

FILL FILL_2__1536_ (
);

FILL FILL_2__1116_ (
);

OAI21X1 _1534_ (
    .A(_707_),
    .B(_706_),
    .C(_672_),
    .Y(_63_)
);

NAND2X1 _1114_ (
    .A(_338_),
    .B(_344_),
    .Y(_345_)
);

OAI21X1 _865_ (
    .A(LoadCtl[4]),
    .B(_106_),
    .C(_107_),
    .Y(_108_)
);

FILL FILL_1__1696_ (
);

FILL FILL_1__1276_ (
);

FILL FILL_0__918_ (
);

DFFPOSX1 _1763_ (
    .D(_35_),
    .CLK(clk_bF$buf2),
    .Q(Xin1[1])
);

NOR2X1 _1343_ (
    .A(_541_),
    .B(_555_),
    .Y(_560_)
);

FILL FILL_1__1085_ (
);

INVX1 _1572_ (
    .A(_741_),
    .Y(_744_)
);

NAND3X1 _1152_ (
    .A(_172_),
    .B(_378_),
    .C(_377_),
    .Y(_381_)
);

FILL FILL_1__934_ (
);

FILL FILL_0__1612_ (
);

FILL FILL_2__1383_ (
);

OAI21X1 _1628_ (
    .A(_793_),
    .B(_752_),
    .C(_796_),
    .Y(_797_)
);

INVX1 _1208_ (
    .A(_421_),
    .Y(_434_)
);

FILL FILL_0__956_ (
);

MUX2X1 _959_ (
    .A(_194_),
    .B(_193_),
    .S(_164__bF$buf2),
    .Y(_195_)
);

INVX1 _1381_ (
    .A(_595_),
    .Y(_596_)
);

FILL FILL_0__1421_ (
);

FILL FILL_0__1001_ (
);

NAND2X1 _1437_ (
    .A(Xin[1]),
    .B(_119_),
    .Y(_639_)
);

OAI21X1 _1017_ (
    .A(_183__bF$buf3),
    .B(_251_),
    .C(_240_),
    .Y(_252_)
);

FILL FILL_1__1599_ (
);

FILL FILL_1__1179_ (
);

NAND3X1 _1190_ (
    .A(_201__bF$buf4),
    .B(_416_),
    .C(_413_),
    .Y(_417_)
);

FILL FILL_1__972_ (
);

FILL FILL_0__1650_ (
);

FILL FILL_0__1230_ (
);

FILL FILL_1__1811_ (
);

NAND2X1 _1666_ (
    .A(_827_),
    .B(_833_),
    .Y(_834_)
);

AOI22X1 _1246_ (
    .A(_146_),
    .B(_188__bF$buf3),
    .C(_470_),
    .D(_186_),
    .Y(_12_)
);

FILL FILL_0__994_ (
);

OAI21X1 _997_ (
    .A(_188__bF$buf1),
    .B(_232_),
    .C(_189_),
    .Y(_1_)
);

FILL FILL_0__1706_ (
);

FILL FILL_2__1477_ (
);

FILL FILL_2__1057_ (
);

FILL FILL88050x79350 (
);

FILL FILL_1__1620_ (
);

FILL FILL_1__1200_ (
);

OAI21X1 _1475_ (
    .A(_606_),
    .B(_629_),
    .C(_658_),
    .Y(_53_)
);

OAI21X1 _1055_ (
    .A(_164__bF$buf4),
    .B(_286_),
    .C(_287_),
    .Y(_288_)
);

FILL FILL_0__1515_ (
);

OAI21X1 _1284_ (
    .A(_504_),
    .B(_496_),
    .C(_501_),
    .Y(_505_)
);

FILL FILL_0__1324_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

INVX1 _1093_ (
    .A(_324_),
    .Y(_325_)
);

FILL FILL_1__875_ (
);

FILL FILL_0__1553_ (
);

FILL FILL_0__1133_ (
);

FILL FILL_1__1714_ (
);

OAI21X1 _1569_ (
    .A(Stg_2_bF$buf3),
    .B(_178_),
    .C(_740_),
    .Y(_741_)
);

OAI21X1 _1149_ (
    .A(Ain12b_11_bF$buf3),
    .B(_371_),
    .C(_375_),
    .Y(_378_)
);

FILL FILL_0__897_ (
);

FILL FILL_0__1609_ (
);

FILL FILL_0__1362_ (
);

FILL FILL_2__891_ (
);

FILL FILL_1__1523_ (
);

FILL FILL_1__1103_ (
);

DFFPOSX1 _1798_ (
    .D(_63_),
    .CLK(clk_bF$buf5),
    .Q(Ycalc[2])
);

INVX1 _1378_ (
    .A(_592_),
    .Y(_593_)
);

FILL FILL_0__1418_ (
);

FILL FILL_2__947_ (
);

FILL FILL_0__1591_ (
);

FILL FILL_0__1171_ (
);

OAI22X1 _921_ (
    .A(_112_),
    .B(_158_),
    .C(_157_),
    .D(_113_),
    .Y(_159_)
);

FILL FILL_1__1332_ (
);

INVX1 _1187_ (
    .A(_336_),
    .Y(_414_)
);

FILL FILL_1__969_ (
);

FILL FILL_0__1647_ (
);

FILL FILL_0__1227_ (
);

FILL FILL_1__1808_ (
);

FILL FILL_1__1561_ (
);

FILL FILL_1__1141_ (
);

FILL FILL88650x75750 (
);

FILL FILL_2__1630_ (
);

FILL FILL_2__1210_ (
);

FILL FILL_0__1456_ (
);

FILL FILL_0__1036_ (
);

FILL FILL_1__1617_ (
);

FILL FILL_1__1370_ (
);

FILL FILL_0__1685_ (
);

FILL FILL_0__1265_ (
);

FILL FILL_1__1426_ (
);

FILL FILL_1__1006_ (
);

FILL FILL_0__1494_ (
);

FILL FILL_0__1074_ (
);

FILL FILL_1__1655_ (
);

FILL FILL_1__1235_ (
);

INVX1 _1722_ (
    .A(_100_),
    .Y(_101_)
);

OAI21X1 _1302_ (
    .A(_492_),
    .B(_521_),
    .C(_520_),
    .Y(_522_)
);

FILL FILL_1__1464_ (
);

FILL FILL_1__1044_ (
);

FILL FILL_2__1533_ (
);

FILL FILL_2__1113_ (
);

FILL FILL_0__1359_ (
);

FILL FILL_2__888_ (
);

OAI21X1 _1531_ (
    .A(_699_),
    .B(_701_),
    .C(_673_),
    .Y(_705_)
);

AOI21X1 _1111_ (
    .A(_332_),
    .B(_201__bF$buf1),
    .C(_339_),
    .Y(_342_)
);

FILL FILL_1__1693_ (
);

FILL FILL_1__1273_ (
);

FILL FILL88350x7350 (
);

FILL FILL_0__1588_ (
);

FILL FILL_0__1168_ (
);

FILL FILL_0__915_ (
);

OAI21X1 _918_ (
    .A(LoadCtl[4]),
    .B(_154_),
    .C(_155_),
    .Y(_156_)
);

FILL FILL_1__1329_ (
);

DFFPOSX1 _1760_ (
    .D(_32_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[4])
);

NAND2X1 _1340_ (
    .A(_556_),
    .B(_545_),
    .Y(_558_)
);

FILL FILL_1__1082_ (
);

FILL FILL_0__1397_ (
);

FILL FILL_1__1558_ (
);

FILL FILL_1__1138_ (
);

FILL FILL_1__931_ (
);

FILL FILL_2__1380_ (
);

INVX1 _1625_ (
    .A(_749_),
    .Y(_794_)
);

NAND2X1 _1205_ (
    .A(_186_),
    .B(_431_),
    .Y(_432_)
);

FILL FILL_0__953_ (
);

INVX2 _956_ (
    .A(_191_),
    .Y(_192_)
);

FILL FILL_1__1367_ (
);

FILL FILL_2__1436_ (
);

FILL FILL_2__1016_ (
);

OAI21X1 _1434_ (
    .A(_212_),
    .B(_635_),
    .C(_637_),
    .Y(_33_)
);

AND2X2 _1014_ (
    .A(_240_),
    .B(_248_),
    .Y(_249_)
);

FILL FILL_1__1596_ (
);

FILL FILL_1__1176_ (
);

AOI21X1 _1663_ (
    .A(_824_),
    .B(_201__bF$buf2),
    .C(_828_),
    .Y(_831_)
);

NOR2X1 _1243_ (
    .A(_463_),
    .B(_465_),
    .Y(_468_)
);

FILL FILL_0__991_ (
);

OAI21X1 _994_ (
    .A(Yin0[0]),
    .B(_199_),
    .C(_229_),
    .Y(_230_)
);

FILL FILL_0__1703_ (
);

NAND2X1 _1719_ (
    .A(_475_),
    .B(_97_),
    .Y(_98_)
);

NAND2X1 _1472_ (
    .A(Ain[0]),
    .B(_629_),
    .Y(_657_)
);

NAND2X1 _1052_ (
    .A(Stg_0_bF$buf0),
    .B(_284_),
    .Y(_285_)
);

FILL FILL_0__1512_ (
);

FILL FILL_2__1283_ (
);

OR2X2 _1528_ (
    .A(_701_),
    .B(_699_),
    .Y(_702_)
);

INVX1 _1108_ (
    .A(_338_),
    .Y(_339_)
);

OAI21X1 _1281_ (
    .A(_500_),
    .B(_502_),
    .C(_491_),
    .Y(_15_)
);

FILL FILL_0__1321_ (
);

DFFPOSX1 _1757_ (
    .D(_29_),
    .CLK(clk_bF$buf4),
    .Q(Xin12b[9])
);

NAND2X1 _1337_ (
    .A(_554_),
    .B(_552_),
    .Y(_555_)
);

FILL FILL_1__1499_ (
);

FILL FILL_1__1079_ (
);

INVX1 _1090_ (
    .A(_319_),
    .Y(_322_)
);

FILL FILL_1__872_ (
);

FILL FILL_0__1550_ (
);

FILL FILL_0__1130_ (
);

FILL FILL_1__1711_ (
);

NAND2X1 _1566_ (
    .A(Stg_1_bF$buf3),
    .B(_737_),
    .Y(_738_)
);

OAI21X1 _1146_ (
    .A(_183__bF$buf2),
    .B(_373_),
    .C(_374_),
    .Y(_375_)
);

FILL FILL_0__894_ (
);

FILL FILL_1__928_ (
);

INVX1 _897_ (
    .A(LoadCtl[4]),
    .Y(_137_)
);

FILL FILL_0__1606_ (
);

FILL FILL_2__1377_ (
);

FILL FILL_1__1520_ (
);

FILL FILL_1__1100_ (
);

FILL FILL_2_BUFX2_insert31 (
);

FILL FILL_2_BUFX2_insert33 (
);

FILL FILL_2_BUFX2_insert36 (
);

FILL FILL_2_BUFX2_insert39 (
);

DFFPOSX1 _1795_ (
    .D(LoadCtl[4]),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[5])
);

INVX1 _1375_ (
    .A(Ain12b[8]),
    .Y(_590_)
);

FILL FILL_0__1415_ (
);

FILL FILL_2__944_ (
);

NAND3X1 _1184_ (
    .A(_382_),
    .B(_387_),
    .C(_405_),
    .Y(_411_)
);

FILL FILL_1__966_ (
);

FILL FILL_0__1644_ (
);

FILL FILL_0__1224_ (
);

FILL FILL_0__988_ (
);

FILL FILL88650x150 (
);

FILL FILL_0__1453_ (
);

FILL FILL_0__1033_ (
);

FILL FILL_1__1614_ (
);

OAI21X1 _1469_ (
    .A(_616_),
    .B(_625_),
    .C(_655_),
    .Y(_50_)
);

AOI21X1 _1049_ (
    .A(_255_),
    .B(_275_),
    .C(_273_),
    .Y(_282_)
);

FILL FILL_0__1509_ (
);

FILL FILL_0__1682_ (
);

FILL FILL_0__1262_ (
);

FILL FILL_1__1423_ (
);

FILL FILL_1__1003_ (
);

INVX1 _1698_ (
    .A(_77_),
    .Y(_78_)
);

NOR2X1 _1278_ (
    .A(_487_),
    .B(_499_),
    .Y(_500_)
);

FILL FILL_0__1318_ (
);

FILL FILL_0__1491_ (
);

FILL FILL_0__1071_ (
);

FILL FILL_1__1652_ (
);

FILL FILL_1__1232_ (
);

AOI21X1 _1087_ (
    .A(_315_),
    .B(Stg_2_bF$buf1),
    .C(_318_),
    .Y(_319_)
);

FILL FILL_1__869_ (
);

FILL FILL_0__1547_ (
);

FILL FILL_0__1127_ (
);

FILL FILL_1__1708_ (
);

FILL FILL_1__1461_ (
);

FILL FILL_1__1041_ (
);

FILL FILL_2__1530_ (
);

FILL FILL_2__1110_ (
);

FILL FILL_0__1356_ (
);

FILL FILL_2__885_ (
);

FILL FILL_1__1517_ (
);

FILL FILL_1__1690_ (
);

FILL FILL_1__1270_ (
);

FILL FILL_0__1585_ (
);

FILL FILL_0__1165_ (
);

FILL FILL_0__912_ (
);

OAI21X1 _915_ (
    .A(_117_),
    .B(_152_),
    .C(_153_),
    .Y(_861_[0])
);

FILL FILL_1__1326_ (
);

FILL FILL88650x61350 (
);

FILL FILL_0__1394_ (
);

BUFX2 _1813_ (
    .A(_861_[1]),
    .Y(Xout[1])
);

FILL FILL_1__1555_ (
);

FILL FILL_1__1135_ (
);

INVX1 _1622_ (
    .A(_785_),
    .Y(_791_)
);

INVX1 _1202_ (
    .A(_426_),
    .Y(_429_)
);

FILL FILL_0__950_ (
);

NAND2X1 _953_ (
    .A(Ycalc[1]),
    .B(_188__bF$buf2),
    .Y(_189_)
);

FILL FILL_1__1364_ (
);

FILL FILL_2__1433_ (
);

FILL FILL_2__1013_ (
);

FILL FILL_0__1679_ (
);

FILL FILL_0__1259_ (
);

NAND2X1 _1431_ (
    .A(Xin[0]),
    .B(_635_),
    .Y(_636_)
);

OAI21X1 _1011_ (
    .A(Stg_0_bF$buf0),
    .B(_244_),
    .C(_245_),
    .Y(_246_)
);

FILL FILL_1__1593_ (
);

FILL FILL_1__1173_ (
);

FILL FILL_0__1488_ (
);

FILL FILL_0__1068_ (
);

FILL FILL87750x86550 (
);

FILL FILL_1__1649_ (
);

FILL FILL_1__1229_ (
);

INVX1 _1660_ (
    .A(_827_),
    .Y(_828_)
);

AOI21X1 _1240_ (
    .A(_410_),
    .B(_411_),
    .C(_464_),
    .Y(_465_)
);

INVX1 _991_ (
    .A(_226_),
    .Y(_227_)
);

FILL FILL_0__1700_ (
);

FILL FILL_0__1297_ (
);

NAND2X1 _1716_ (
    .A(Ycalc[11]),
    .B(_188__bF$buf2),
    .Y(_95_)
);

FILL FILL_1__1458_ (
);

FILL FILL_1__1038_ (
);

FILL FILL_2__1107_ (
);

FILL FILL_2__1280_ (
);

AOI21X1 _1525_ (
    .A(_698_),
    .B(_679_),
    .C(Yin1[0]),
    .Y(_699_)
);

OAI21X1 _1105_ (
    .A(Stg_1_bF$buf3),
    .B(_286_),
    .C(_335_),
    .Y(_336_)
);

FILL FILL_1__1687_ (
);

FILL FILL_1__1267_ (
);

FILL FILL_2__1336_ (
);

FILL FILL_0__909_ (
);

DFFPOSX1 _1754_ (
    .D(_26_),
    .CLK(clk_bF$buf4),
    .Q(Xin12b[10])
);

INVX1 _1334_ (
    .A(_551_),
    .Y(_552_)
);

FILL FILL_1__1496_ (
);

FILL FILL_1__1076_ (
);

NAND3X1 _1563_ (
    .A(_678_),
    .B(_726_),
    .C(_696_),
    .Y(_735_)
);

INVX1 _1143_ (
    .A(_371_),
    .Y(_372_)
);

FILL FILL_0__891_ (
);

FILL FILL_1__925_ (
);

AOI21X1 _894_ (
    .A(_109_),
    .B(_131_),
    .C(_134_),
    .Y(_135_)
);

FILL FILL_0__1603_ (
);

AOI21X1 _1619_ (
    .A(_788_),
    .B(_786_),
    .C(_192_),
    .Y(_789_)
);

FILL FILL_0__947_ (
);

DFFPOSX1 _1792_ (
    .D(LoadCtl[1]),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[2])
);

NAND2X1 _1372_ (
    .A(_521_),
    .B(_586_),
    .Y(_587_)
);

FILL FILL_0__1412_ (
);

FILL FILL_2__941_ (
);

FILL FILL_2__1183_ (
);

NAND2X1 _1428_ (
    .A(Xin[1]),
    .B(_632_),
    .Y(_634_)
);

OAI21X1 _1008_ (
    .A(Stg_0_bF$buf0),
    .B(_241_),
    .C(_242_),
    .Y(_243_)
);

NAND2X1 _1181_ (
    .A(Xcalc[8]),
    .B(_188__bF$buf3),
    .Y(_408_)
);

FILL FILL_1__963_ (
);

FILL FILL_0__1641_ (
);

FILL FILL_0__1221_ (
);

INVX1 _1657_ (
    .A(_739_),
    .Y(_825_)
);

AND2X2 _1237_ (
    .A(_457_),
    .B(_461_),
    .Y(_462_)
);

FILL FILL_0__985_ (
);

MUX2X1 _988_ (
    .A(_223_),
    .B(_220_),
    .S(Stg_2_bF$buf1),
    .Y(_224_)
);

FILL FILL_1__1399_ (
);

FILL FILL88050x86550 (
);

FILL FILL_0__1450_ (
);

FILL FILL_0__1030_ (
);

FILL FILL_1__1611_ (
);

NAND2X1 _1466_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Yin[1]),
    .Y(_654_)
);

AOI21X1 _1046_ (
    .A(_279_),
    .B(_276_),
    .C(_192_),
    .Y(_280_)
);

FILL FILL_0__1506_ (
);

FILL FILL_2__1697_ (
);

FILL FILL_2__1277_ (
);

FILL FILL_1__1420_ (
);

FILL FILL_1__1000_ (
);

OR2X2 _1695_ (
    .A(_74_),
    .B(_73_),
    .Y(_75_)
);

OR2X2 _1275_ (
    .A(_496_),
    .B(Ain0[1]),
    .Y(_497_)
);

FILL FILL_0__1315_ (
);

NAND2X1 _1084_ (
    .A(_267_),
    .B(_290_),
    .Y(_316_)
);

FILL FILL_1__866_ (
);

FILL FILL_0__1544_ (
);

FILL FILL_0__1124_ (
);

FILL FILL_1__1705_ (
);

FILL FILL_0__888_ (
);

FILL FILL_0__1353_ (
);

FILL FILL_1__1514_ (
);

DFFPOSX1 _1789_ (
    .D(_61_),
    .CLK(clk_bF$buf7),
    .Q(Ain0[1])
);

AOI22X1 _1369_ (
    .A(_124_),
    .B(_188__bF$buf3),
    .C(_583_),
    .D(_584_),
    .Y(_21_)
);

FILL FILL_0__1409_ (
);

FILL FILL_2__938_ (
);

FILL FILL_0__1582_ (
);

FILL FILL_0__1162_ (
);

OAI22X1 _912_ (
    .A(_112_),
    .B(_150_),
    .C(_149_),
    .D(_113_),
    .Y(_151_)
);

FILL FILL_1__1323_ (
);

AND2X2 _1598_ (
    .A(_766_),
    .B(_768_),
    .Y(_769_)
);

OR2X2 _1178_ (
    .A(_393_),
    .B(_405_),
    .Y(_406_)
);

FILL FILL_0__1638_ (
);

FILL FILL_0__1218_ (
);

FILL FILL88650x82950 (
);

FILL FILL_0__1391_ (
);

BUFX2 _1810_ (
    .A(_860_),
    .Y(ISout)
);

FILL FILL_1__1552_ (
);

FILL FILL_1__1132_ (
);

FILL FILL87450x64950 (
);

FILL FILL_0__1447_ (
);

FILL FILL_0__1027_ (
);

FILL FILL_1__1608_ (
);

OAI21X1 _950_ (
    .A(_180_),
    .B(_182_),
    .C(_186_),
    .Y(_187_)
);

FILL FILL_1__1361_ (
);

FILL FILL_1__998_ (
);

FILL FILL_2__1430_ (
);

FILL FILL_2__1010_ (
);

FILL FILL_0__1676_ (
);

FILL FILL_0__1256_ (
);

FILL FILL_1__1417_ (
);

FILL FILL_1__1590_ (
);

FILL FILL_1__1170_ (
);

FILL FILL_0__1485_ (
);

FILL FILL_0__1065_ (
);

FILL FILL_1__1646_ (
);

FILL FILL_1__1226_ (
);

FILL FILL_0__1294_ (
);

OAI21X1 _1713_ (
    .A(_87_),
    .B(_92_),
    .C(_191_),
    .Y(_93_)
);

FILL FILL_1__1455_ (
);

FILL FILL_1__1035_ (
);

FILL FILL88650x14550 (
);

AOI22X1 _1522_ (
    .A(_684_),
    .B(_689_),
    .C(_692_),
    .D(_695_),
    .Y(_696_)
);

NAND2X1 _1102_ (
    .A(Stg_0_bF$buf5),
    .B(Yin12b[11]),
    .Y(_333_)
);

FILL FILL_1__1684_ (
);

FILL FILL_1__1264_ (
);

FILL FILL_2__1333_ (
);

FILL FILL_0__1579_ (
);

FILL FILL_0__1159_ (
);

FILL FILL_0__906_ (
);

OAI21X1 _909_ (
    .A(LoadCtl[4]),
    .B(_146_),
    .C(_147_),
    .Y(_148_)
);

DFFPOSX1 _1751_ (
    .D(_23_),
    .CLK(clk_bF$buf7),
    .Q(Acalc[9])
);

NOR2X1 _1331_ (
    .A(_201__bF$buf0),
    .B(_548_),
    .Y(_549_)
);

FILL FILL_1__1493_ (
);

FILL FILL_1__1073_ (
);

FILL FILL_0__1388_ (
);

DFFPOSX1 _1807_ (
    .D(_72_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[11])
);

FILL FILL88650x3750 (
);

FILL FILL_1__1549_ (
);

FILL FILL_1__1129_ (
);

AOI21X1 _1560_ (
    .A(_732_),
    .B(_711_),
    .C(_192_),
    .Y(_733_)
);

OAI21X1 _1140_ (
    .A(_368_),
    .B(_352_),
    .C(_186_),
    .Y(_370_)
);

FILL FILL_1__922_ (
);

INVX1 _891_ (
    .A(Ycalc[6]),
    .Y(_132_)
);

FILL FILL_0__1600_ (
);

FILL FILL_0__1197_ (
);

NAND2X1 _1616_ (
    .A(_782_),
    .B(_785_),
    .Y(_786_)
);

FILL FILL_0__944_ (
);

NAND2X1 _947_ (
    .A(_183__bF$buf1),
    .B(_164__bF$buf2),
    .Y(_184_)
);

FILL FILL_1__1358_ (
);

FILL FILL87750x72150 (
);

FILL FILL_2__1427_ (
);

FILL FILL_2__1007_ (
);

FILL FILL87750x39750 (
);

FILL FILL_2__1180_ (
);

NOR2X1 _1425_ (
    .A(_113_),
    .B(_117_),
    .Y(_632_)
);

NAND2X1 _1005_ (
    .A(_183__bF$buf3),
    .B(_239_),
    .Y(_240_)
);

FILL FILL_1__1587_ (
);

FILL FILL_1__1167_ (
);

FILL FILL_1__960_ (
);

NAND3X1 _1654_ (
    .A(_818_),
    .B(_821_),
    .C(_820_),
    .Y(_822_)
);

NOR2X1 _1234_ (
    .A(_449_),
    .B(_455_),
    .Y(_459_)
);

FILL FILL_0__982_ (
);

MUX2X1 _985_ (
    .A(Xin12b[8]),
    .B(Xin12b[7]),
    .S(Stg_0_bF$buf3),
    .Y(_221_)
);

FILL FILL_1__1396_ (
);

OAI21X1 _1463_ (
    .A(_256_),
    .B(_119_),
    .C(_652_),
    .Y(_47_)
);

INVX1 _1043_ (
    .A(_255_),
    .Y(_277_)
);

FILL FILL_0__1503_ (
);

FILL FILL_2__1694_ (
);

FILL FILL_2__1274_ (
);

NAND2X1 _1519_ (
    .A(_164__bF$buf0),
    .B(_214_),
    .Y(_693_)
);

OAI21X1 _1692_ (
    .A(Stg_2_bF$buf3),
    .B(_775_),
    .C(_826_),
    .Y(_858_)
);

OAI21X1 _1272_ (
    .A(Stg_2_bF$buf2),
    .B(_492_),
    .C(_493_),
    .Y(_494_)
);

FILL FILL_0__1312_ (
);

DFFPOSX1 _1748_ (
    .D(_20_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[6])
);

OAI21X1 _1328_ (
    .A(_190_),
    .B(_292_),
    .C(_201__bF$buf3),
    .Y(_546_)
);

OAI21X1 _1081_ (
    .A(Stg_0_bF$buf5),
    .B(Yin12b[9]),
    .C(_312_),
    .Y(_313_)
);

FILL FILL_1__863_ (
);

FILL FILL_0__1541_ (
);

FILL FILL_0__1121_ (
);

FILL FILL_1__1702_ (
);

NOR2X1 _1557_ (
    .A(Yin1[1]),
    .B(_728_),
    .Y(_730_)
);

NAND2X1 _1137_ (
    .A(_363_),
    .B(_366_),
    .Y(_367_)
);

FILL FILL_0__885_ (
);

FILL FILL_1__919_ (
);

INVX1 _888_ (
    .A(Ycalc[10]),
    .Y(_129_)
);

FILL FILL_1__1299_ (
);

FILL FILL_0__1350_ (
);

FILL FILL_1__1511_ (
);

DFFPOSX1 _1786_ (
    .D(_58_),
    .CLK(clk_bF$buf7),
    .Q(Ain1[0])
);

INVX1 _1366_ (
    .A(_581_),
    .Y(_582_)
);

FILL FILL_0__1406_ (
);

FILL FILL_2__1597_ (
);

FILL FILL_2__1177_ (
);

FILL FILL88050x72150 (
);

FILL FILL_1__1320_ (
);

FILL FILL88050x39750 (
);

NAND3X1 _1595_ (
    .A(_265_),
    .B(_765_),
    .C(_764_),
    .Y(_766_)
);

NAND2X1 _1175_ (
    .A(_401_),
    .B(_402_),
    .Y(_403_)
);

FILL FILL_1__957_ (
);

FILL FILL_0__1635_ (
);

FILL FILL_0__1215_ (
);

FILL FILL_0__979_ (
);

FILL FILL_0__1444_ (
);

FILL FILL_0__1024_ (
);

FILL FILL_1__1605_ (
);

FILL FILL_1__995_ (
);

FILL FILL_0__1673_ (
);

FILL FILL_0__1253_ (
);

FILL FILL_1__1414_ (
);

OAI21X1 _1689_ (
    .A(_854_),
    .B(_841_),
    .C(_191_),
    .Y(_856_)
);

NAND2X1 _1269_ (
    .A(Acalc[1]),
    .B(_188__bF$buf0),
    .Y(_491_)
);

FILL FILL_0__1309_ (
);

FILL FILL_0__1482_ (
);

FILL FILL_0__1062_ (
);

FILL FILL_1__1643_ (
);

FILL FILL_1__1223_ (
);

NAND2X1 _1498_ (
    .A(Ycalc[2]),
    .B(_188__bF$buf1),
    .Y(_672_)
);

NAND2X1 _1078_ (
    .A(_295_),
    .B(_298_),
    .Y(_310_)
);

FILL FILL_0__1538_ (
);

FILL FILL_0__1118_ (
);

FILL FILL_0__1291_ (
);

AOI21X1 _1710_ (
    .A(_89_),
    .B(_797_),
    .C(_88_),
    .Y(_90_)
);

FILL FILL_1__1452_ (
);

FILL FILL_1__1032_ (
);

FILL FILL_0__1347_ (
);

FILL FILL_1__1508_ (
);

FILL FILL_1__1681_ (
);

FILL FILL_1__1261_ (
);

FILL FILL_1__898_ (
);

FILL FILL_2__1330_ (
);

FILL FILL_0__1576_ (
);

FILL FILL_0__1156_ (
);

FILL FILL_0__903_ (
);

OAI21X1 _906_ (
    .A(_117_),
    .B(_144_),
    .C(_145_),
    .Y(_862_[1])
);

FILL FILL_1__1317_ (
);

FILL FILL_1__1490_ (
);

FILL FILL_1__1070_ (
);

FILL FILL_0__1385_ (
);

DFFPOSX1 _1804_ (
    .D(_69_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[8])
);

FILL FILL_1__1546_ (
);

FILL FILL_1__1126_ (
);

FILL FILL_0__1194_ (
);

NAND3X1 _1613_ (
    .A(_201__bF$buf5),
    .B(_780_),
    .C(_774_),
    .Y(_783_)
);

FILL FILL_0__941_ (
);

NAND2X1 _944_ (
    .A(_163_),
    .B(_179_),
    .Y(_181_)
);

FILL FILL_1__1355_ (
);

FILL FILL_2__1004_ (
);

OAI21X1 _1422_ (
    .A(_422_),
    .B(_629_),
    .C(_630_),
    .Y(_28_)
);

NAND2X1 _1002_ (
    .A(Stg_0_bF$buf2),
    .B(Yin0[1]),
    .Y(_237_)
);

FILL FILL_1__1584_ (
);

FILL FILL_1__1164_ (
);

FILL FILL_2__1653_ (
);

FILL FILL_2__1233_ (
);

FILL FILL_0__1479_ (
);

FILL FILL_0__1059_ (
);

AOI21X1 _1651_ (
    .A(_791_),
    .B(_818_),
    .C(_809_),
    .Y(_819_)
);

NOR2X1 _1231_ (
    .A(_454_),
    .B(_455_),
    .Y(_456_)
);

MUX2X1 _982_ (
    .A(Xin12b[4]),
    .B(Xin1[1]),
    .S(Stg_0_bF$buf1),
    .Y(_218_)
);

FILL FILL_1__1393_ (
);

FILL FILL_0__1288_ (
);

AND2X2 _1707_ (
    .A(_79_),
    .B(_81_),
    .Y(_87_)
);

FILL FILL_1__1449_ (
);

FILL FILL_1__1029_ (
);

NAND2X1 _1460_ (
    .A(Yin[0]),
    .B(_119_),
    .Y(_651_)
);

INVX1 _1040_ (
    .A(_273_),
    .Y(_274_)
);

FILL FILL_0__1500_ (
);

FILL FILL_0__1097_ (
);

NAND2X1 _1516_ (
    .A(Stg_1_bF$buf2),
    .B(_204_),
    .Y(_690_)
);

FILL FILL_1__1678_ (
);

FILL FILL_1__1258_ (
);

FILL FILL_2__1327_ (
);

FILL FILL_2__1080_ (
);

DFFPOSX1 _1745_ (
    .D(_17_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[3])
);

OAI21X1 _1325_ (
    .A(_540_),
    .B(_543_),
    .C(_531_),
    .Y(_18_)
);

FILL FILL_1__1487_ (
);

FILL FILL_1__1067_ (
);

OAI21X1 _1554_ (
    .A(Ain12b_11_bF$buf1),
    .B(_721_),
    .C(_726_),
    .Y(_727_)
);

NAND3X1 _1134_ (
    .A(_201__bF$buf1),
    .B(_361_),
    .C(_354_),
    .Y(_364_)
);

FILL FILL_0__882_ (
);

FILL FILL_1__916_ (
);

AOI21X1 _885_ (
    .A(_109_),
    .B(_123_),
    .C(_126_),
    .Y(_127_)
);

FILL FILL_1__1296_ (
);

FILL FILL_0__938_ (
);

DFFPOSX1 _1783_ (
    .D(_55_),
    .CLK(clk_bF$buf7),
    .Q(Ain12b[7])
);

INVX1 _1363_ (
    .A(_578_),
    .Y(_579_)
);

FILL FILL_0__1403_ (
);

FILL FILL_2__1594_ (
);

FILL FILL_2__1174_ (
);

NOR2X1 _1419_ (
    .A(_137_),
    .B(_117_),
    .Y(_628_)
);

NOR2X1 _1592_ (
    .A(_761_),
    .B(_762_),
    .Y(_763_)
);

OAI21X1 _1172_ (
    .A(_399_),
    .B(_398_),
    .C(Xin12b[7]),
    .Y(_400_)
);

FILL FILL_1__954_ (
);

FILL FILL_0__1632_ (
);

FILL FILL_0__1212_ (
);

OAI21X1 _1648_ (
    .A(_141_),
    .B(LoadCtl_6_bF$buf3),
    .C(_816_),
    .Y(_68_)
);

NOR2X1 _1228_ (
    .A(_449_),
    .B(_452_),
    .Y(_453_)
);

FILL FILL_0__976_ (
);

MUX2X1 _979_ (
    .A(_214_),
    .B(_211_),
    .S(_164__bF$buf0),
    .Y(_215_)
);

FILL FILL_0__1441_ (
);

FILL FILL_0__1021_ (
);

FILL FILL_1__1602_ (
);

OAI21X1 _1457_ (
    .A(_244_),
    .B(_635_),
    .C(_649_),
    .Y(_44_)
);

INVX1 _1037_ (
    .A(_269_),
    .Y(_271_)
);

FILL FILL_1__1199_ (
);

FILL FILL_1__992_ (
);

FILL FILL_0__1670_ (
);

FILL FILL_0__1250_ (
);

FILL FILL_1__1411_ (
);

OAI21X1 _1686_ (
    .A(_850_),
    .B(_852_),
    .C(Yin12b[9]),
    .Y(_853_)
);

OR2X2 _1266_ (
    .A(_488_),
    .B(_487_),
    .Y(_489_)
);

FILL FILL_0__1726_ (
);

FILL FILL_0__1306_ (
);

FILL FILL_2__1497_ (
);

FILL FILL_2__1077_ (
);

FILL FILL_1__1640_ (
);

FILL FILL_1__1220_ (
);

INVX1 _1495_ (
    .A(_860_),
    .Y(_670_)
);

NAND2X1 _1075_ (
    .A(Xcalc[3]),
    .B(_188__bF$buf4),
    .Y(_307_)
);

FILL FILL_0__1535_ (
);

FILL FILL_0__1115_ (
);

FILL FILL_0__879_ (
);

FILL FILL_0__1344_ (
);

FILL FILL_1__1505_ (
);

FILL FILL88050x25350 (
);

FILL FILL_1__895_ (
);

FILL FILL_0__1573_ (
);

FILL FILL_0__1153_ (
);

FILL FILL_0__900_ (
);

OAI22X1 _903_ (
    .A(_112_),
    .B(_142_),
    .C(_141_),
    .D(_113_),
    .Y(_143_)
);

FILL FILL_1__1314_ (
);

OAI21X1 _1589_ (
    .A(_183__bF$buf0),
    .B(_758_),
    .C(_759_),
    .Y(_760_)
);

NAND3X1 _1169_ (
    .A(_201__bF$buf4),
    .B(_396_),
    .C(_394_),
    .Y(_397_)
);

FILL FILL_0__1629_ (
);

FILL FILL_0__1209_ (
);

FILL FILL_0__1382_ (
);

DFFPOSX1 _1801_ (
    .D(_66_),
    .CLK(clk_bF$buf1),
    .Q(Ycalc[5])
);

FILL FILL_1__1543_ (
);

FILL FILL_1__1123_ (
);

OAI21X1 _1398_ (
    .A(_611_),
    .B(_610_),
    .C(_603_),
    .Y(_23_)
);

FILL FILL_0__1438_ (
);

FILL FILL_0__1018_ (
);

FILL FILL_0__1191_ (
);

INVX1 _1610_ (
    .A(_777_),
    .Y(_780_)
);

MUX2X1 _941_ (
    .A(_177_),
    .B(_174_),
    .S(_164__bF$buf0),
    .Y(_178_)
);

FILL FILL_1__1352_ (
);

FILL FILL_1__989_ (
);

FILL FILL_0__1667_ (
);

FILL FILL_0__1247_ (
);

FILL FILL_1__1408_ (
);

FILL FILL_1__1581_ (
);

FILL FILL_1__1161_ (
);

FILL FILL_2__1650_ (
);

FILL FILL_2__1230_ (
);

FILL FILL_0__1476_ (
);

FILL FILL_0__1056_ (
);

FILL FILL_1__1637_ (
);

FILL FILL_1__1217_ (
);

FILL FILL_1__1390_ (
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_2__1706_ (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert2 (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_0_BUFX2_insert4 (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_0__1285_ (
);

AOI21X1 _1704_ (
    .A(_840_),
    .B(_849_),
    .C(_83_),
    .Y(_84_)
);

FILL FILL_1__1446_ (
);

FILL FILL_1__1026_ (
);

FILL FILL88650x21750 (
);

FILL FILL_0__1094_ (
);

NAND3X1 _1513_ (
    .A(_164__bF$buf2),
    .B(_686_),
    .C(_685_),
    .Y(_687_)
);

FILL FILL_1__1675_ (
);

FILL FILL_1__1255_ (
);

FILL FILL_2__1324_ (
);

DFFPOSX1 _1742_ (
    .D(_14_),
    .CLK(clk_bF$buf0),
    .Q(Acalc[0])
);

NAND2X1 _1322_ (
    .A(_538_),
    .B(_536_),
    .Y(_541_)
);

FILL FILL_1__1484_ (
);

FILL FILL_1__1064_ (
);

FILL FILL_2__1553_ (
);

FILL FILL_0__1379_ (
);

NAND2X1 _1551_ (
    .A(_164__bF$buf0),
    .B(_211_),
    .Y(_724_)
);

INVX1 _1131_ (
    .A(_359_),
    .Y(_361_)
);

FILL FILL_1__913_ (
);

INVX1 _882_ (
    .A(Acalc[7]),
    .Y(_124_)
);

FILL FILL_1__1293_ (
);

FILL FILL_2_BUFX2_insert0 (
);

FILL FILL_2_BUFX2_insert3 (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_0__1188_ (
);

OAI21X1 _1607_ (
    .A(_183__bF$buf0),
    .B(_775_),
    .C(_776_),
    .Y(_777_)
);

FILL FILL_0__935_ (
);

FILL FILL87750x46950 (
);

INVX1 _938_ (
    .A(Xin12b[4]),
    .Y(_175_)
);

FILL FILL_1__1349_ (
);

DFFPOSX1 _1780_ (
    .D(_52_),
    .CLK(clk_bF$buf3),
    .Q(Ain12b[8])
);

NAND2X1 _1360_ (
    .A(_575_),
    .B(_574_),
    .Y(_576_)
);

FILL FILL_0__1400_ (
);

FILL FILL_2__1171_ (
);

OAI21X1 _1416_ (
    .A(_458_),
    .B(_625_),
    .C(_626_),
    .Y(_26_)
);

FILL FILL_1__1578_ (
);

FILL FILL_1__1158_ (
);

FILL FILL_1__951_ (
);

FILL FILL_2__1647_ (
);

FILL FILL_2__1227_ (
);

OAI21X1 _1645_ (
    .A(_201__bF$buf6),
    .B(_191_),
    .C(LoadCtl_6_bF$buf3),
    .Y(_814_)
);

OR2X2 _1225_ (
    .A(_413_),
    .B(_416_),
    .Y(_450_)
);

FILL FILL_0__973_ (
);

INVX1 _976_ (
    .A(Xin12b[5]),
    .Y(_212_)
);

FILL FILL_1__1387_ (
);

NAND2X1 _1454_ (
    .A(Yin[1]),
    .B(_632_),
    .Y(_648_)
);

MUX2X1 _1034_ (
    .A(_267_),
    .B(_264_),
    .S(_164__bF$buf4),
    .Y(_268_)
);

FILL FILL_1__1196_ (
);

AOI21X1 _1683_ (
    .A(_847_),
    .B(_201__bF$buf2),
    .C(_843_),
    .Y(_850_)
);

OAI21X1 _1263_ (
    .A(_183__bF$buf3),
    .B(_484_),
    .C(_485_),
    .Y(_486_)
);

FILL FILL_0__1723_ (
);

FILL FILL_0__1303_ (
);

FILL FILL_2__1494_ (
);

FILL FILL_2__1074_ (
);

DFFPOSX1 _1739_ (
    .D(_11_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[9])
);

OAI21X1 _1319_ (
    .A(_534_),
    .B(_532_),
    .C(_537_),
    .Y(_538_)
);

OAI21X1 _1492_ (
    .A(LoadCtl_0_bF$buf3),
    .B(_483_),
    .C(_668_),
    .Y(_60_)
);

INVX1 _1072_ (
    .A(_303_),
    .Y(_305_)
);

FILL FILL_0__1532_ (
);

FILL FILL_0__1112_ (
);

INVX1 _1548_ (
    .A(_712_),
    .Y(_721_)
);

OAI21X1 _1128_ (
    .A(_357_),
    .B(_355_),
    .C(Stg_2_bF$buf4),
    .Y(_358_)
);

FILL FILL_0__876_ (
);

INVX1 _879_ (
    .A(Acalc[11]),
    .Y(_121_)
);

FILL FILL_0__1341_ (
);

FILL FILL_1__1502_ (
);

DFFPOSX1 _1777_ (
    .D(_49_),
    .CLK(clk_bF$buf2),
    .Q(Yin0[1])
);

OAI21X1 _1357_ (
    .A(_570_),
    .B(_562_),
    .C(_567_),
    .Y(_573_)
);

FILL FILL_1__1099_ (
);

FILL FILL_1__892_ (
);

FILL FILL88050x46950 (
);

FILL FILL_0__1570_ (
);

FILL FILL_0__1150_ (
);

OAI21X1 _900_ (
    .A(_137_),
    .B(_138_),
    .C(_139_),
    .Y(_140_)
);

FILL FILL_1__1311_ (
);

FILL FILL88050x3750 (
);

NOR2X1 _1586_ (
    .A(_164__bF$buf3),
    .B(_471_),
    .Y(_757_)
);

NAND3X1 _1166_ (
    .A(_361_),
    .B(_376_),
    .C(_353_),
    .Y(_394_)
);

FILL FILL_1__948_ (
);

FILL FILL_0__1626_ (
);

FILL FILL_0__1206_ (
);

FILL FILL_2__1397_ (
);

FILL FILL_1__1540_ (
);

FILL FILL_1__1120_ (
);

NAND2X1 _1395_ (
    .A(_607_),
    .B(_608_),
    .Y(_609_)
);

FILL FILL_0__1435_ (
);

FILL FILL_0__1015_ (
);

FILL FILL_1__986_ (
);

FILL FILL_0__1664_ (
);

FILL FILL_0__1244_ (
);

FILL FILL_1__1405_ (
);

FILL FILL_0__1473_ (
);

FILL FILL_0__1053_ (
);

FILL FILL_1__1634_ (
);

FILL FILL_1__1214_ (
);

OAI21X1 _1489_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_118_),
    .C(Ain1[1]),
    .Y(_667_)
);

AOI21X1 _1069_ (
    .A(_297_),
    .B(_299_),
    .C(Xin1[0]),
    .Y(_302_)
);

FILL FILL_2__1703_ (
);

FILL FILL_0__1529_ (
);

FILL FILL_0__1109_ (
);

FILL FILL_0__1282_ (
);

OAI21X1 _1701_ (
    .A(_77_),
    .B(_80_),
    .C(Yin12b[10]),
    .Y(_81_)
);

FILL FILL_1__1443_ (
);

FILL FILL_1__1023_ (
);

INVX1 _1298_ (
    .A(Ain1[1]),
    .Y(_518_)
);

FILL FILL_0__1338_ (
);

FILL FILL_0__1091_ (
);

NAND3X1 _1510_ (
    .A(_183__bF$buf1),
    .B(_682_),
    .C(_683_),
    .Y(_684_)
);

FILL FILL_1__1672_ (
);

FILL FILL_1__1252_ (
);

FILL FILL_1__889_ (
);

FILL FILL_0__1567_ (
);

FILL FILL_0__1147_ (
);

FILL FILL_1__1308_ (
);

FILL FILL_0_BUFX2_insert50 (
);

FILL FILL_0_BUFX2_insert51 (
);

FILL FILL_0_BUFX2_insert52 (
);

FILL FILL_0_BUFX2_insert53 (
);

FILL FILL_0_BUFX2_insert54 (
);

FILL FILL_0_BUFX2_insert55 (
);

FILL FILL_0_BUFX2_insert56 (
);

FILL FILL_0_BUFX2_insert57 (
);

FILL FILL_0_BUFX2_insert58 (
);

FILL FILL_1__1481_ (
);

FILL FILL_1__1061_ (
);

FILL FILL_2__1550_ (
);

FILL FILL_2__1130_ (
);

FILL FILL88350x54150 (
);

FILL FILL_0__1376_ (
);

FILL FILL_1__1537_ (
);

FILL FILL_1__1117_ (
);

FILL FILL_1__910_ (
);

FILL FILL_1__1290_ (
);

FILL FILL_0__1185_ (
);

NAND3X1 _1604_ (
    .A(_744_),
    .B(_761_),
    .C(_743_),
    .Y(_774_)
);

FILL FILL_0__932_ (
);

INVX1 _935_ (
    .A(Xin12b[6]),
    .Y(_172_)
);

FILL FILL_1__1346_ (
);

NAND3X1 _1413_ (
    .A(LoadCtl[5]),
    .B(_137_),
    .C(_109_),
    .Y(_624_)
);

FILL FILL_1__1575_ (
);

FILL FILL_1__1155_ (
);

FILL FILL_2__1644_ (
);

FILL FILL_2__1224_ (
);

NOR2X1 _1642_ (
    .A(_810_),
    .B(_798_),
    .Y(_811_)
);

OAI21X1 _1222_ (
    .A(_446_),
    .B(_447_),
    .C(_186_),
    .Y(_448_)
);

FILL FILL_0__970_ (
);

INVX1 _973_ (
    .A(Xin12b[7]),
    .Y(_209_)
);

FILL FILL_1__1384_ (
);

FILL FILL_0__1699_ (
);

FILL FILL_0__1279_ (
);

OAI21X1 _1451_ (
    .A(_284_),
    .B(_629_),
    .C(_646_),
    .Y(_41_)
);

INVX1 _1031_ (
    .A(Yin12b[5]),
    .Y(_265_)
);

FILL FILL_1__1193_ (
);

FILL FILL_0__1088_ (
);

NAND2X1 _1507_ (
    .A(Stg_0_bF$buf1),
    .B(_202_),
    .Y(_681_)
);

FILL FILL_1__1669_ (
);

FILL FILL_1__1249_ (
);

NAND3X1 _1680_ (
    .A(_801_),
    .B(_828_),
    .C(_846_),
    .Y(_847_)
);

INVX1 _1260_ (
    .A(Ain0[0]),
    .Y(_483_)
);

FILL FILL_0__1720_ (
);

FILL FILL_0__1300_ (
);

FILL FILL_2__1491_ (
);

FILL FILL_2__1071_ (
);

DFFPOSX1 _1736_ (
    .D(_8_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[6])
);

NOR2X1 _1316_ (
    .A(_534_),
    .B(_532_),
    .Y(_535_)
);

FILL FILL_1__1478_ (
);

FILL FILL_1__1058_ (
);

FILL FILL_2__1547_ (
);

FILL FILL_2__1127_ (
);

INVX1 _1545_ (
    .A(_717_),
    .Y(_718_)
);

NOR2X1 _1125_ (
    .A(Stg_1_bF$buf0),
    .B(_313_),
    .Y(_355_)
);

FILL FILL_0__873_ (
);

FILL FILL_1__907_ (
);

NOR2X1 _876_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_118_),
    .Y(_119_)
);

FILL FILL_1__1287_ (
);

FILL FILL_0__929_ (
);

DFFPOSX1 _1774_ (
    .D(_46_),
    .CLK(clk_bF$buf2),
    .Q(Yin1[0])
);

AND2X2 _1354_ (
    .A(_562_),
    .B(_570_),
    .Y(_571_)
);

FILL FILL_1__1096_ (
);

FILL FILL_0__1814_ (
);

AOI22X1 _1583_ (
    .A(_133_),
    .B(_188__bF$buf2),
    .C(_754_),
    .D(_709_),
    .Y(_65_)
);

OAI21X1 _1163_ (
    .A(_149_),
    .B(LoadCtl_6_bF$buf1),
    .C(_391_),
    .Y(_8_)
);

FILL FILL_1__945_ (
);

FILL FILL_0__1623_ (
);

FILL FILL_0__1203_ (
);

FILL FILL_2__1394_ (
);

NAND2X1 _1639_ (
    .A(_801_),
    .B(_804_),
    .Y(_808_)
);

NAND2X1 _1219_ (
    .A(_444_),
    .B(_440_),
    .Y(_445_)
);

FILL FILL_0__967_ (
);

INVX1 _1392_ (
    .A(Ain12b[9]),
    .Y(_606_)
);

FILL FILL_0__1432_ (
);

FILL FILL_0__1012_ (
);

FILL FILL_2__961_ (
);

NAND2X1 _1448_ (
    .A(Yin[0]),
    .B(_629_),
    .Y(_645_)
);

INVX1 _1028_ (
    .A(Yin12b[7]),
    .Y(_262_)
);

FILL FILL_1__983_ (
);

endmodule
