VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic_element
  CLASS BLOCK ;
  FOREIGN cordic_element ;
  ORIGIN 6.000 6.000 ;
  SIZE 903.000 BY 915.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 900.300 900.300 902.700 ;
        RECT 891.300 830.700 900.300 900.300 ;
        RECT 0.600 828.300 900.300 830.700 ;
        RECT 891.300 758.700 900.300 828.300 ;
        RECT 0.600 756.300 900.300 758.700 ;
        RECT 891.300 686.700 900.300 756.300 ;
        RECT 0.600 684.300 900.300 686.700 ;
        RECT 891.300 614.700 900.300 684.300 ;
        RECT 0.600 612.300 900.300 614.700 ;
        RECT 891.300 542.700 900.300 612.300 ;
        RECT 0.600 540.300 900.300 542.700 ;
        RECT 891.300 470.700 900.300 540.300 ;
        RECT 0.600 468.300 900.300 470.700 ;
        RECT 891.300 398.700 900.300 468.300 ;
        RECT 0.600 396.300 900.300 398.700 ;
        RECT 891.300 326.700 900.300 396.300 ;
        RECT 0.600 324.300 900.300 326.700 ;
        RECT 891.300 254.700 900.300 324.300 ;
        RECT 0.600 252.300 900.300 254.700 ;
        RECT 891.300 182.700 900.300 252.300 ;
        RECT 0.600 180.300 900.300 182.700 ;
        RECT 891.300 110.700 900.300 180.300 ;
        RECT 0.600 108.300 900.300 110.700 ;
        RECT 891.300 38.700 900.300 108.300 ;
        RECT 0.600 36.300 900.300 38.700 ;
        RECT 891.300 0.300 900.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 866.700 -0.300 902.700 ;
        RECT -9.300 864.300 890.400 866.700 ;
        RECT -9.300 794.700 -0.300 864.300 ;
        RECT -9.300 792.300 890.400 794.700 ;
        RECT -9.300 722.700 -0.300 792.300 ;
        RECT -9.300 720.300 890.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT -9.300 648.300 890.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT -9.300 576.300 890.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT -9.300 504.300 890.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT -9.300 432.300 890.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT -9.300 360.300 890.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT -9.300 288.300 890.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT -9.300 216.300 890.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT -9.300 144.300 890.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT -9.300 72.300 890.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT -9.300 0.300 890.400 2.700 ;
    END
  END vdd
  PIN Ain[1]
    PORT
      LAYER metal2 ;
        RECT 292.950 666.450 295.050 667.050 ;
        RECT 290.400 665.400 295.050 666.450 ;
        RECT 290.400 661.050 291.450 665.400 ;
        RECT 292.950 664.950 295.050 665.400 ;
        RECT 427.950 664.950 430.050 667.050 ;
        RECT 428.400 661.050 429.450 664.950 ;
        RECT 289.950 658.950 292.050 661.050 ;
        RECT 427.950 658.950 430.050 661.050 ;
        RECT 517.950 658.950 520.050 661.050 ;
        RECT 1.950 637.950 4.050 640.050 ;
        RECT 2.400 586.050 3.450 637.950 ;
        RECT 290.400 586.050 291.450 658.950 ;
        RECT 1.950 583.950 4.050 586.050 ;
        RECT 214.950 583.950 217.050 586.050 ;
        RECT 289.950 583.950 292.050 586.050 ;
        RECT 215.400 562.050 216.450 583.950 ;
        RECT 214.950 559.950 217.050 562.050 ;
        RECT 518.400 508.050 519.450 658.950 ;
        RECT 799.950 520.950 802.050 523.050 ;
        RECT 800.400 517.050 801.450 520.950 ;
        RECT 694.950 514.950 697.050 517.050 ;
        RECT 799.950 514.950 802.050 517.050 ;
        RECT 695.400 508.050 696.450 514.950 ;
        RECT 517.950 505.950 520.050 508.050 ;
        RECT 694.950 505.950 697.050 508.050 ;
        RECT 691.950 480.450 694.050 481.050 ;
        RECT 695.400 480.450 696.450 505.950 ;
        RECT 691.950 479.400 696.450 480.450 ;
        RECT 691.950 478.950 694.050 479.400 ;
      LAYER metal3 ;
        RECT 289.950 660.600 292.050 661.050 ;
        RECT 427.950 660.600 430.050 661.050 ;
        RECT 517.950 660.600 520.050 661.050 ;
        RECT 289.950 659.400 520.050 660.600 ;
        RECT 289.950 658.950 292.050 659.400 ;
        RECT 427.950 658.950 430.050 659.400 ;
        RECT 517.950 658.950 520.050 659.400 ;
        RECT 1.950 639.600 4.050 640.050 ;
        RECT -3.600 638.400 4.050 639.600 ;
        RECT 1.950 637.950 4.050 638.400 ;
        RECT 1.950 585.600 4.050 586.050 ;
        RECT 214.950 585.600 217.050 586.050 ;
        RECT 289.950 585.600 292.050 586.050 ;
        RECT 1.950 584.400 292.050 585.600 ;
        RECT 1.950 583.950 4.050 584.400 ;
        RECT 214.950 583.950 217.050 584.400 ;
        RECT 289.950 583.950 292.050 584.400 ;
        RECT 694.950 516.600 697.050 517.050 ;
        RECT 799.950 516.600 802.050 517.050 ;
        RECT 694.950 515.400 802.050 516.600 ;
        RECT 694.950 514.950 697.050 515.400 ;
        RECT 799.950 514.950 802.050 515.400 ;
        RECT 517.950 507.600 520.050 508.050 ;
        RECT 694.950 507.600 697.050 508.050 ;
        RECT 517.950 506.400 697.050 507.600 ;
        RECT 517.950 505.950 520.050 506.400 ;
        RECT 694.950 505.950 697.050 506.400 ;
    END
  END Ain[1]
  PIN Ain[0]
    PORT
      LAYER metal2 ;
        RECT 397.950 703.950 400.050 706.050 ;
        RECT 415.950 703.950 418.050 706.050 ;
        RECT 538.950 705.450 541.050 706.050 ;
        RECT 538.950 704.400 543.450 705.450 ;
        RECT 538.950 703.950 541.050 704.400 ;
        RECT 398.400 688.050 399.450 703.950 ;
        RECT 542.400 688.050 543.450 704.400 ;
        RECT 397.950 685.950 400.050 688.050 ;
        RECT 541.950 685.950 544.050 688.050 ;
        RECT 595.950 685.950 598.050 688.050 ;
        RECT 398.400 678.450 399.450 685.950 ;
        RECT 395.400 677.400 399.450 678.450 ;
        RECT 370.950 634.950 373.050 637.050 ;
        RECT 371.400 634.050 372.450 634.950 ;
        RECT 395.400 634.050 396.450 677.400 ;
        RECT 596.400 637.050 597.450 685.950 ;
        RECT 595.950 634.950 598.050 637.050 ;
        RECT 658.950 634.950 661.050 637.050 ;
        RECT 757.950 634.950 760.050 637.050 ;
        RECT 659.400 634.050 660.450 634.950 ;
        RECT 370.950 631.950 373.050 634.050 ;
        RECT 394.950 631.950 397.050 634.050 ;
        RECT 397.950 631.950 400.050 634.050 ;
        RECT 658.950 631.950 661.050 634.050 ;
        RECT 398.400 595.050 399.450 631.950 ;
        RECT 758.400 604.050 759.450 634.950 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 397.950 592.950 400.050 595.050 ;
        RECT 409.950 592.950 412.050 595.050 ;
      LAYER metal3 ;
        RECT 397.950 705.600 400.050 706.050 ;
        RECT 415.950 705.600 418.050 706.050 ;
        RECT 397.950 704.400 418.050 705.600 ;
        RECT 397.950 703.950 400.050 704.400 ;
        RECT 415.950 703.950 418.050 704.400 ;
        RECT 397.950 687.600 400.050 688.050 ;
        RECT 541.950 687.600 544.050 688.050 ;
        RECT 595.950 687.600 598.050 688.050 ;
        RECT 397.950 686.400 598.050 687.600 ;
        RECT 397.950 685.950 400.050 686.400 ;
        RECT 541.950 685.950 544.050 686.400 ;
        RECT 595.950 685.950 598.050 686.400 ;
        RECT 370.950 636.600 373.050 637.050 ;
        RECT -3.600 635.400 373.050 636.600 ;
        RECT -3.600 632.400 -2.400 635.400 ;
        RECT 370.950 634.950 373.050 635.400 ;
        RECT 595.950 636.600 598.050 637.050 ;
        RECT 658.950 636.600 661.050 637.050 ;
        RECT 757.950 636.600 760.050 637.050 ;
        RECT 595.950 635.400 760.050 636.600 ;
        RECT 595.950 634.950 598.050 635.400 ;
        RECT 658.950 634.950 661.050 635.400 ;
        RECT 757.950 634.950 760.050 635.400 ;
        RECT 370.950 633.600 373.050 634.050 ;
        RECT 394.950 633.600 397.050 634.050 ;
        RECT 397.950 633.600 400.050 634.050 ;
        RECT 370.950 632.400 400.050 633.600 ;
        RECT 370.950 631.950 373.050 632.400 ;
        RECT 394.950 631.950 397.050 632.400 ;
        RECT 397.950 631.950 400.050 632.400 ;
        RECT 397.950 594.600 400.050 595.050 ;
        RECT 409.950 594.600 412.050 595.050 ;
        RECT 397.950 593.400 412.050 594.600 ;
        RECT 397.950 592.950 400.050 593.400 ;
        RECT 409.950 592.950 412.050 593.400 ;
    END
  END Ain[0]
  PIN Aout[1]
    PORT
      LAYER metal2 ;
        RECT 812.400 889.050 813.450 909.450 ;
        RECT 811.950 886.950 814.050 889.050 ;
    END
  END Aout[1]
  PIN Aout[0]
    PORT
      LAYER metal2 ;
        RECT 758.400 889.050 759.450 909.450 ;
        RECT 757.950 886.950 760.050 889.050 ;
    END
  END Aout[0]
  PIN ISin
    PORT
      LAYER metal2 ;
        RECT 1.950 880.950 4.050 883.050 ;
        RECT 121.950 880.950 124.050 883.050 ;
        RECT 2.400 877.050 3.450 880.950 ;
        RECT 122.400 877.050 123.450 880.950 ;
        RECT 1.950 874.950 4.050 877.050 ;
        RECT 121.950 874.950 124.050 877.050 ;
      LAYER metal3 ;
        RECT 1.950 882.600 4.050 883.050 ;
        RECT -3.600 881.400 4.050 882.600 ;
        RECT 1.950 880.950 4.050 881.400 ;
        RECT 1.950 876.600 4.050 877.050 ;
        RECT 121.950 876.600 124.050 877.050 ;
        RECT 1.950 875.400 124.050 876.600 ;
        RECT 1.950 874.950 4.050 875.400 ;
        RECT 121.950 874.950 124.050 875.400 ;
    END
  END ISin
  PIN ISout
    PORT
      LAYER metal2 ;
        RECT 671.400 904.050 672.450 909.450 ;
        RECT 346.950 901.950 349.050 904.050 ;
        RECT 670.950 901.950 673.050 904.050 ;
        RECT 347.400 889.050 348.450 901.950 ;
        RECT 346.950 886.950 349.050 889.050 ;
      LAYER metal3 ;
        RECT 346.950 903.600 349.050 904.050 ;
        RECT 670.950 903.600 673.050 904.050 ;
        RECT 346.950 902.400 673.050 903.600 ;
        RECT 346.950 901.950 349.050 902.400 ;
        RECT 670.950 901.950 673.050 902.400 ;
    END
  END ISout
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 31.950 481.950 34.050 484.050 ;
      LAYER metal3 ;
        RECT -3.600 485.400 33.600 486.600 ;
        RECT 32.400 484.050 33.600 485.400 ;
        RECT 31.950 481.950 34.050 484.050 ;
    END
  END Rdy
  PIN Stg[2]
    PORT
      LAYER metal2 ;
        RECT 286.950 339.450 289.050 340.050 ;
        RECT 286.950 338.400 291.450 339.450 ;
        RECT 286.950 337.950 289.050 338.400 ;
        RECT 290.400 265.050 291.450 338.400 ;
        RECT 472.950 337.950 475.050 340.050 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 473.400 334.050 474.450 337.950 ;
        RECT 454.950 331.950 457.050 334.050 ;
        RECT 472.950 331.950 475.050 334.050 ;
        RECT 424.950 265.950 427.050 268.050 ;
        RECT 425.400 265.050 426.450 265.950 ;
        RECT 455.400 265.050 456.450 331.950 ;
        RECT 695.400 331.050 696.450 337.950 ;
        RECT 694.950 328.950 697.050 331.050 ;
        RECT 289.950 262.950 292.050 265.050 ;
        RECT 298.950 262.950 301.050 265.050 ;
        RECT 424.950 262.950 427.050 265.050 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 299.400 196.050 300.450 262.950 ;
        RECT 289.950 193.950 292.050 196.050 ;
        RECT 298.950 193.950 301.050 196.050 ;
        RECT 290.400 133.050 291.450 193.950 ;
        RECT 277.950 130.950 280.050 133.050 ;
        RECT 289.950 130.950 292.050 133.050 ;
        RECT 278.400 42.450 279.450 130.950 ;
        RECT 275.400 41.400 279.450 42.450 ;
        RECT 275.400 4.050 276.450 41.400 ;
        RECT 274.950 1.950 277.050 4.050 ;
        RECT 280.950 1.950 283.050 4.050 ;
        RECT 281.400 -3.600 282.450 1.950 ;
      LAYER metal3 ;
        RECT 454.950 333.600 457.050 334.050 ;
        RECT 472.950 333.600 475.050 334.050 ;
        RECT 454.950 332.400 663.600 333.600 ;
        RECT 454.950 331.950 457.050 332.400 ;
        RECT 472.950 331.950 475.050 332.400 ;
        RECT 662.400 330.600 663.600 332.400 ;
        RECT 694.950 330.600 697.050 331.050 ;
        RECT 662.400 329.400 697.050 330.600 ;
        RECT 694.950 328.950 697.050 329.400 ;
        RECT 289.950 264.600 292.050 265.050 ;
        RECT 298.950 264.600 301.050 265.050 ;
        RECT 424.950 264.600 427.050 265.050 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 289.950 263.400 457.050 264.600 ;
        RECT 289.950 262.950 292.050 263.400 ;
        RECT 298.950 262.950 301.050 263.400 ;
        RECT 424.950 262.950 427.050 263.400 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 289.950 195.600 292.050 196.050 ;
        RECT 298.950 195.600 301.050 196.050 ;
        RECT 289.950 194.400 301.050 195.600 ;
        RECT 289.950 193.950 292.050 194.400 ;
        RECT 298.950 193.950 301.050 194.400 ;
        RECT 277.950 132.600 280.050 133.050 ;
        RECT 289.950 132.600 292.050 133.050 ;
        RECT 277.950 131.400 292.050 132.600 ;
        RECT 277.950 130.950 280.050 131.400 ;
        RECT 289.950 130.950 292.050 131.400 ;
        RECT 274.950 3.600 277.050 4.050 ;
        RECT 280.950 3.600 283.050 4.050 ;
        RECT 274.950 2.400 283.050 3.600 ;
        RECT 274.950 1.950 277.050 2.400 ;
        RECT 280.950 1.950 283.050 2.400 ;
    END
  END Stg[2]
  PIN Stg[1]
    PORT
      LAYER metal2 ;
        RECT 205.950 337.950 208.050 340.050 ;
        RECT 364.950 337.950 367.050 340.050 ;
        RECT 538.950 339.450 541.050 340.050 ;
        RECT 536.400 338.400 541.050 339.450 ;
        RECT 206.400 295.050 207.450 337.950 ;
        RECT 365.400 336.450 366.450 337.950 ;
        RECT 365.400 335.400 369.450 336.450 ;
        RECT 368.400 295.050 369.450 335.400 ;
        RECT 536.400 295.050 537.450 338.400 ;
        RECT 538.950 337.950 541.050 338.400 ;
        RECT 205.950 292.950 208.050 295.050 ;
        RECT 325.950 292.950 328.050 295.050 ;
        RECT 367.950 292.950 370.050 295.050 ;
        RECT 535.950 292.950 538.050 295.050 ;
        RECT 206.400 267.450 207.450 292.950 ;
        RECT 208.950 267.450 211.050 268.050 ;
        RECT 206.400 266.400 211.050 267.450 ;
        RECT 208.950 265.950 211.050 266.400 ;
        RECT 326.400 208.050 327.450 292.950 ;
        RECT 319.950 205.950 322.050 208.050 ;
        RECT 325.950 205.950 328.050 208.050 ;
        RECT 320.400 60.450 321.450 205.950 ;
        RECT 320.400 59.400 324.450 60.450 ;
        RECT 323.400 27.450 324.450 59.400 ;
        RECT 320.400 26.400 324.450 27.450 ;
        RECT 320.400 7.050 321.450 26.400 ;
        RECT 259.950 4.950 262.050 7.050 ;
        RECT 319.950 4.950 322.050 7.050 ;
        RECT 260.400 -3.600 261.450 4.950 ;
      LAYER metal3 ;
        RECT 205.950 294.600 208.050 295.050 ;
        RECT 325.950 294.600 328.050 295.050 ;
        RECT 367.950 294.600 370.050 295.050 ;
        RECT 535.950 294.600 538.050 295.050 ;
        RECT 205.950 293.400 538.050 294.600 ;
        RECT 205.950 292.950 208.050 293.400 ;
        RECT 325.950 292.950 328.050 293.400 ;
        RECT 367.950 292.950 370.050 293.400 ;
        RECT 535.950 292.950 538.050 293.400 ;
        RECT 319.950 207.600 322.050 208.050 ;
        RECT 325.950 207.600 328.050 208.050 ;
        RECT 319.950 206.400 328.050 207.600 ;
        RECT 319.950 205.950 322.050 206.400 ;
        RECT 325.950 205.950 328.050 206.400 ;
        RECT 259.950 6.600 262.050 7.050 ;
        RECT 319.950 6.600 322.050 7.050 ;
        RECT 259.950 5.400 322.050 6.600 ;
        RECT 259.950 4.950 262.050 5.400 ;
        RECT 319.950 4.950 322.050 5.400 ;
    END
  END Stg[1]
  PIN Stg[0]
    PORT
      LAYER metal2 ;
        RECT 157.950 463.950 160.050 466.050 ;
        RECT 274.950 463.950 277.050 466.050 ;
        RECT 158.400 457.050 159.450 463.950 ;
        RECT 275.400 457.050 276.450 463.950 ;
        RECT 157.950 456.450 160.050 457.050 ;
        RECT 155.400 455.400 160.050 456.450 ;
        RECT 151.950 411.450 154.050 412.050 ;
        RECT 155.400 411.450 156.450 455.400 ;
        RECT 157.950 454.950 160.050 455.400 ;
        RECT 274.950 456.450 277.050 457.050 ;
        RECT 274.950 455.400 279.450 456.450 ;
        RECT 274.950 454.950 277.050 455.400 ;
        RECT 278.400 436.050 279.450 455.400 ;
        RECT 277.950 433.950 280.050 436.050 ;
        RECT 490.950 433.950 493.050 436.050 ;
        RECT 151.950 410.400 156.450 411.450 ;
        RECT 491.400 411.450 492.450 433.950 ;
        RECT 493.950 411.450 496.050 412.050 ;
        RECT 491.400 410.400 496.050 411.450 ;
        RECT 151.950 409.950 154.050 410.400 ;
        RECT 493.950 409.950 496.050 410.400 ;
        RECT 494.400 385.050 495.450 409.950 ;
        RECT 493.950 382.950 496.050 385.050 ;
        RECT 502.950 382.950 505.050 385.050 ;
        RECT 494.400 358.050 495.450 382.950 ;
        RECT 481.950 355.950 484.050 358.050 ;
        RECT 493.950 355.950 496.050 358.050 ;
        RECT 482.400 301.050 483.450 355.950 ;
        RECT 481.950 298.950 484.050 301.050 ;
        RECT 490.950 298.950 493.050 301.050 ;
        RECT 491.400 240.450 492.450 298.950 ;
        RECT 493.950 240.450 496.050 241.050 ;
        RECT 491.400 239.400 496.050 240.450 ;
        RECT 491.400 226.050 492.450 239.400 ;
        RECT 493.950 238.950 496.050 239.400 ;
        RECT 277.950 223.950 280.050 226.050 ;
        RECT 490.950 223.950 493.050 226.050 ;
        RECT 278.400 172.050 279.450 223.950 ;
        RECT 241.950 169.950 244.050 172.050 ;
        RECT 256.950 169.950 259.050 172.050 ;
        RECT 277.950 169.950 280.050 172.050 ;
        RECT 242.400 58.050 243.450 169.950 ;
        RECT 257.400 169.050 258.450 169.950 ;
        RECT 256.950 166.950 259.050 169.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 248.400 27.450 249.450 55.950 ;
        RECT 245.400 26.400 249.450 27.450 ;
        RECT 245.400 4.050 246.450 26.400 ;
        RECT 244.950 1.950 247.050 4.050 ;
        RECT 253.950 1.950 256.050 4.050 ;
        RECT 254.400 -3.600 255.450 1.950 ;
      LAYER metal3 ;
        RECT 157.950 465.600 160.050 466.050 ;
        RECT 274.950 465.600 277.050 466.050 ;
        RECT 157.950 464.400 277.050 465.600 ;
        RECT 157.950 463.950 160.050 464.400 ;
        RECT 274.950 463.950 277.050 464.400 ;
        RECT 277.950 435.600 280.050 436.050 ;
        RECT 490.950 435.600 493.050 436.050 ;
        RECT 277.950 434.400 493.050 435.600 ;
        RECT 277.950 433.950 280.050 434.400 ;
        RECT 490.950 433.950 493.050 434.400 ;
        RECT 493.950 384.600 496.050 385.050 ;
        RECT 502.950 384.600 505.050 385.050 ;
        RECT 493.950 383.400 505.050 384.600 ;
        RECT 493.950 382.950 496.050 383.400 ;
        RECT 502.950 382.950 505.050 383.400 ;
        RECT 481.950 357.600 484.050 358.050 ;
        RECT 493.950 357.600 496.050 358.050 ;
        RECT 481.950 356.400 496.050 357.600 ;
        RECT 481.950 355.950 484.050 356.400 ;
        RECT 493.950 355.950 496.050 356.400 ;
        RECT 481.950 300.600 484.050 301.050 ;
        RECT 490.950 300.600 493.050 301.050 ;
        RECT 481.950 299.400 493.050 300.600 ;
        RECT 481.950 298.950 484.050 299.400 ;
        RECT 490.950 298.950 493.050 299.400 ;
        RECT 277.950 225.600 280.050 226.050 ;
        RECT 490.950 225.600 493.050 226.050 ;
        RECT 277.950 224.400 493.050 225.600 ;
        RECT 277.950 223.950 280.050 224.400 ;
        RECT 490.950 223.950 493.050 224.400 ;
        RECT 241.950 171.600 244.050 172.050 ;
        RECT 256.950 171.600 259.050 172.050 ;
        RECT 277.950 171.600 280.050 172.050 ;
        RECT 241.950 170.400 280.050 171.600 ;
        RECT 241.950 169.950 244.050 170.400 ;
        RECT 256.950 169.950 259.050 170.400 ;
        RECT 277.950 169.950 280.050 170.400 ;
        RECT 241.950 57.600 244.050 58.050 ;
        RECT 247.950 57.600 250.050 58.050 ;
        RECT 241.950 56.400 250.050 57.600 ;
        RECT 241.950 55.950 244.050 56.400 ;
        RECT 247.950 55.950 250.050 56.400 ;
        RECT 244.950 3.600 247.050 4.050 ;
        RECT 253.950 3.600 256.050 4.050 ;
        RECT 244.950 2.400 256.050 3.600 ;
        RECT 244.950 1.950 247.050 2.400 ;
        RECT 253.950 1.950 256.050 2.400 ;
    END
  END Stg[0]
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 665.400 908.400 669.450 909.450 ;
        RECT 668.400 889.050 669.450 908.400 ;
        RECT 667.950 886.950 670.050 889.050 ;
    END
  END Vld
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 649.950 375.450 652.050 376.050 ;
        RECT 655.950 375.450 658.050 376.050 ;
        RECT 649.950 374.550 658.050 375.450 ;
        RECT 649.950 373.950 652.050 374.550 ;
        RECT 655.950 373.950 658.050 374.550 ;
      LAYER metal2 ;
        RECT 286.950 592.950 289.050 595.050 ;
        RECT 287.400 591.450 288.450 592.950 ;
        RECT 284.400 590.400 288.450 591.450 ;
        RECT 284.400 577.050 285.450 590.400 ;
        RECT 283.950 574.950 286.050 577.050 ;
        RECT 427.950 574.950 430.050 577.050 ;
        RECT 649.950 574.950 652.050 577.050 ;
        RECT 211.950 520.950 214.050 523.050 ;
        RECT 212.400 511.050 213.450 520.950 ;
        RECT 284.400 511.050 285.450 574.950 ;
        RECT 428.400 562.050 429.450 574.950 ;
        RECT 427.950 559.950 430.050 562.050 ;
        RECT 28.950 508.950 31.050 511.050 ;
        RECT 211.950 508.950 214.050 511.050 ;
        RECT 283.950 508.950 286.050 511.050 ;
        RECT 29.400 471.450 30.450 508.950 ;
        RECT 26.400 470.400 30.450 471.450 ;
        RECT 16.950 376.950 19.050 379.050 ;
        RECT 17.400 355.050 18.450 376.950 ;
        RECT 26.400 355.050 27.450 470.400 ;
        RECT 650.400 376.050 651.450 574.950 ;
        RECT 655.950 376.950 658.050 379.050 ;
        RECT 656.400 376.050 657.450 376.950 ;
        RECT 649.950 373.950 652.050 376.050 ;
        RECT 655.950 373.950 658.050 376.050 ;
        RECT 16.950 352.950 19.050 355.050 ;
        RECT 25.950 352.950 28.050 355.050 ;
        RECT 26.400 232.050 27.450 352.950 ;
        RECT 656.400 274.050 657.450 373.950 ;
        RECT 631.950 271.950 634.050 274.050 ;
        RECT 655.950 271.950 658.050 274.050 ;
        RECT 16.950 229.950 19.050 232.050 ;
        RECT 25.950 229.950 28.050 232.050 ;
        RECT 17.400 202.050 18.450 229.950 ;
        RECT 16.950 199.950 19.050 202.050 ;
        RECT 632.400 129.450 633.450 271.950 ;
        RECT 629.400 128.400 633.450 129.450 ;
        RECT 629.400 103.050 630.450 128.400 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 701.400 -2.550 702.450 100.950 ;
        RECT 698.400 -3.600 702.450 -2.550 ;
      LAYER metal3 ;
        RECT 283.950 576.600 286.050 577.050 ;
        RECT 427.950 576.600 430.050 577.050 ;
        RECT 649.950 576.600 652.050 577.050 ;
        RECT 283.950 575.400 652.050 576.600 ;
        RECT 283.950 574.950 286.050 575.400 ;
        RECT 427.950 574.950 430.050 575.400 ;
        RECT 649.950 574.950 652.050 575.400 ;
        RECT 28.950 510.600 31.050 511.050 ;
        RECT 211.950 510.600 214.050 511.050 ;
        RECT 283.950 510.600 286.050 511.050 ;
        RECT 28.950 509.400 286.050 510.600 ;
        RECT 28.950 508.950 31.050 509.400 ;
        RECT 211.950 508.950 214.050 509.400 ;
        RECT 283.950 508.950 286.050 509.400 ;
        RECT 16.950 354.600 19.050 355.050 ;
        RECT 25.950 354.600 28.050 355.050 ;
        RECT 16.950 353.400 28.050 354.600 ;
        RECT 16.950 352.950 19.050 353.400 ;
        RECT 25.950 352.950 28.050 353.400 ;
        RECT 631.950 273.600 634.050 274.050 ;
        RECT 655.950 273.600 658.050 274.050 ;
        RECT 631.950 272.400 658.050 273.600 ;
        RECT 631.950 271.950 634.050 272.400 ;
        RECT 655.950 271.950 658.050 272.400 ;
        RECT 16.950 231.600 19.050 232.050 ;
        RECT 25.950 231.600 28.050 232.050 ;
        RECT 16.950 230.400 28.050 231.600 ;
        RECT 16.950 229.950 19.050 230.400 ;
        RECT 25.950 229.950 28.050 230.400 ;
        RECT 628.950 102.600 631.050 103.050 ;
        RECT 700.950 102.600 703.050 103.050 ;
        RECT 628.950 101.400 703.050 102.600 ;
        RECT 628.950 100.950 631.050 101.400 ;
        RECT 700.950 100.950 703.050 101.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 76.950 522.450 79.050 523.050 ;
        RECT 76.950 521.400 81.450 522.450 ;
        RECT 76.950 520.950 79.050 521.400 ;
        RECT 80.400 448.050 81.450 521.400 ;
        RECT 415.950 502.950 418.050 505.050 ;
        RECT 607.950 502.950 610.050 505.050 ;
        RECT 416.400 502.050 417.450 502.950 ;
        RECT 343.950 499.950 346.050 502.050 ;
        RECT 415.950 499.950 418.050 502.050 ;
        RECT 340.950 489.450 343.050 490.050 ;
        RECT 344.400 489.450 345.450 499.950 ;
        RECT 416.400 490.050 417.450 499.950 ;
        RECT 340.950 488.400 345.450 489.450 ;
        RECT 340.950 487.950 343.050 488.400 ;
        RECT 344.400 481.050 345.450 488.400 ;
        RECT 415.950 487.950 418.050 490.050 ;
        RECT 295.950 478.950 298.050 481.050 ;
        RECT 343.950 478.950 346.050 481.050 ;
        RECT 127.950 448.950 130.050 451.050 ;
        RECT 229.950 448.950 232.050 451.050 ;
        RECT 128.400 448.050 129.450 448.950 ;
        RECT 230.400 448.050 231.450 448.950 ;
        RECT 296.400 448.050 297.450 478.950 ;
        RECT 79.950 445.950 82.050 448.050 ;
        RECT 127.950 445.950 130.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 295.950 445.950 298.050 448.050 ;
        RECT 608.400 445.050 609.450 502.950 ;
        RECT 607.950 442.950 610.050 445.050 ;
        RECT 700.950 442.950 703.050 445.050 ;
        RECT 701.400 418.050 702.450 442.950 ;
        RECT 700.950 417.450 703.050 418.050 ;
        RECT 698.400 416.400 703.050 417.450 ;
        RECT 698.400 241.050 699.450 416.400 ;
        RECT 700.950 415.950 703.050 416.400 ;
        RECT 691.950 238.950 694.050 241.050 ;
        RECT 697.950 238.950 700.050 241.050 ;
        RECT 692.400 139.050 693.450 238.950 ;
        RECT 679.950 136.950 682.050 139.050 ;
        RECT 691.950 136.950 694.050 139.050 ;
        RECT 680.400 4.050 681.450 136.950 ;
        RECT 679.950 1.950 682.050 4.050 ;
        RECT 691.950 1.950 694.050 4.050 ;
        RECT 692.400 -3.600 693.450 1.950 ;
      LAYER metal3 ;
        RECT 415.950 504.600 418.050 505.050 ;
        RECT 607.950 504.600 610.050 505.050 ;
        RECT 415.950 503.400 610.050 504.600 ;
        RECT 415.950 502.950 418.050 503.400 ;
        RECT 607.950 502.950 610.050 503.400 ;
        RECT 343.950 501.600 346.050 502.050 ;
        RECT 415.950 501.600 418.050 502.050 ;
        RECT 343.950 500.400 418.050 501.600 ;
        RECT 343.950 499.950 346.050 500.400 ;
        RECT 415.950 499.950 418.050 500.400 ;
        RECT 295.950 480.600 298.050 481.050 ;
        RECT 343.950 480.600 346.050 481.050 ;
        RECT 295.950 479.400 346.050 480.600 ;
        RECT 295.950 478.950 298.050 479.400 ;
        RECT 343.950 478.950 346.050 479.400 ;
        RECT 79.950 447.600 82.050 448.050 ;
        RECT 127.950 447.600 130.050 448.050 ;
        RECT 229.950 447.600 232.050 448.050 ;
        RECT 295.950 447.600 298.050 448.050 ;
        RECT 79.950 446.400 298.050 447.600 ;
        RECT 79.950 445.950 82.050 446.400 ;
        RECT 127.950 445.950 130.050 446.400 ;
        RECT 229.950 445.950 232.050 446.400 ;
        RECT 295.950 445.950 298.050 446.400 ;
        RECT 607.950 444.600 610.050 445.050 ;
        RECT 700.950 444.600 703.050 445.050 ;
        RECT 607.950 443.400 703.050 444.600 ;
        RECT 607.950 442.950 610.050 443.400 ;
        RECT 700.950 442.950 703.050 443.400 ;
        RECT 691.950 240.600 694.050 241.050 ;
        RECT 697.950 240.600 700.050 241.050 ;
        RECT 691.950 239.400 700.050 240.600 ;
        RECT 691.950 238.950 694.050 239.400 ;
        RECT 697.950 238.950 700.050 239.400 ;
        RECT 679.950 138.600 682.050 139.050 ;
        RECT 691.950 138.600 694.050 139.050 ;
        RECT 679.950 137.400 694.050 138.600 ;
        RECT 679.950 136.950 682.050 137.400 ;
        RECT 691.950 136.950 694.050 137.400 ;
        RECT 679.950 3.600 682.050 4.050 ;
        RECT 691.950 3.600 694.050 4.050 ;
        RECT 679.950 2.400 694.050 3.600 ;
        RECT 679.950 1.950 682.050 2.400 ;
        RECT 691.950 1.950 694.050 2.400 ;
    END
  END Xin[0]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 889.950 886.950 892.050 889.050 ;
        RECT 890.400 838.050 891.450 886.950 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 857.400 817.050 858.450 835.950 ;
        RECT 856.950 814.950 859.050 817.050 ;
      LAYER metal3 ;
        RECT 889.950 888.600 892.050 889.050 ;
        RECT 889.950 887.400 897.600 888.600 ;
        RECT 889.950 886.950 892.050 887.400 ;
        RECT 856.950 837.600 859.050 838.050 ;
        RECT 889.950 837.600 892.050 838.050 ;
        RECT 856.950 836.400 892.050 837.600 ;
        RECT 856.950 835.950 859.050 836.400 ;
        RECT 889.950 835.950 892.050 836.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 868.950 888.450 871.050 889.050 ;
        RECT 868.950 887.400 873.450 888.450 ;
        RECT 868.950 886.950 871.050 887.400 ;
        RECT 872.400 883.050 873.450 887.400 ;
        RECT 871.950 880.950 874.050 883.050 ;
      LAYER metal3 ;
        RECT 871.950 882.600 874.050 883.050 ;
        RECT 871.950 881.400 897.600 882.600 ;
        RECT 871.950 880.950 874.050 881.400 ;
    END
  END Xout[0]
  PIN Yin[1]
    PORT
      LAYER metal1 ;
        RECT 436.950 204.450 439.050 205.050 ;
        RECT 442.950 204.450 445.050 205.050 ;
        RECT 436.950 203.550 445.050 204.450 ;
        RECT 436.950 202.950 439.050 203.550 ;
        RECT 442.950 202.950 445.050 203.550 ;
      LAYER metal2 ;
        RECT 436.950 202.950 439.050 205.050 ;
        RECT 442.950 202.950 445.050 205.050 ;
        RECT 437.400 184.050 438.450 202.950 ;
        RECT 443.400 202.050 444.450 202.950 ;
        RECT 442.950 199.950 445.050 202.050 ;
        RECT 601.950 201.450 604.050 202.050 ;
        RECT 599.400 200.400 604.050 201.450 ;
        RECT 599.400 184.050 600.450 200.400 ;
        RECT 601.950 199.950 604.050 200.400 ;
        RECT 643.950 199.950 646.050 202.050 ;
        RECT 694.950 199.950 697.050 202.050 ;
        RECT 436.950 181.950 439.050 184.050 ;
        RECT 598.950 181.950 601.050 184.050 ;
        RECT 79.950 160.950 82.050 163.050 ;
        RECT 80.400 136.050 81.450 160.950 ;
        RECT 437.400 151.050 438.450 181.950 ;
        RECT 301.950 148.950 304.050 151.050 ;
        RECT 436.950 148.950 439.050 151.050 ;
        RECT 302.400 136.050 303.450 148.950 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 146.400 130.050 147.450 133.950 ;
        RECT 145.950 127.950 148.050 130.050 ;
        RECT 302.400 27.450 303.450 133.950 ;
        RECT 302.400 26.400 306.450 27.450 ;
        RECT 305.400 -3.600 306.450 26.400 ;
      LAYER metal3 ;
        RECT 601.950 201.600 604.050 202.050 ;
        RECT 643.950 201.600 646.050 202.050 ;
        RECT 694.950 201.600 697.050 202.050 ;
        RECT 601.950 200.400 697.050 201.600 ;
        RECT 601.950 199.950 604.050 200.400 ;
        RECT 643.950 199.950 646.050 200.400 ;
        RECT 694.950 199.950 697.050 200.400 ;
        RECT 436.950 183.600 439.050 184.050 ;
        RECT 598.950 183.600 601.050 184.050 ;
        RECT 436.950 182.400 601.050 183.600 ;
        RECT 436.950 181.950 439.050 182.400 ;
        RECT 598.950 181.950 601.050 182.400 ;
        RECT 301.950 150.600 304.050 151.050 ;
        RECT 436.950 150.600 439.050 151.050 ;
        RECT 301.950 149.400 439.050 150.600 ;
        RECT 301.950 148.950 304.050 149.400 ;
        RECT 436.950 148.950 439.050 149.400 ;
        RECT 79.950 135.600 82.050 136.050 ;
        RECT 145.950 135.600 148.050 136.050 ;
        RECT 301.950 135.600 304.050 136.050 ;
        RECT 79.950 134.400 304.050 135.600 ;
        RECT 79.950 133.950 82.050 134.400 ;
        RECT 145.950 133.950 148.050 134.400 ;
        RECT 301.950 133.950 304.050 134.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 520.950 232.950 523.050 235.050 ;
        RECT 682.950 232.950 685.050 235.050 ;
        RECT 694.950 232.950 697.050 235.050 ;
        RECT 521.400 220.050 522.450 232.950 ;
        RECT 683.400 220.050 684.450 232.950 ;
        RECT 695.400 220.050 696.450 232.950 ;
        RECT 313.950 217.950 316.050 220.050 ;
        RECT 520.950 217.950 523.050 220.050 ;
        RECT 682.950 217.950 685.050 220.050 ;
        RECT 694.950 217.950 697.050 220.050 ;
        RECT 310.950 201.450 313.050 202.050 ;
        RECT 314.400 201.450 315.450 217.950 ;
        RECT 310.950 200.400 315.450 201.450 ;
        RECT 310.950 199.950 313.050 200.400 ;
        RECT 40.950 160.950 43.050 163.050 ;
        RECT 41.400 133.050 42.450 160.950 ;
        RECT 314.400 157.050 315.450 200.400 ;
        RECT 163.950 154.950 166.050 157.050 ;
        RECT 298.950 154.950 301.050 157.050 ;
        RECT 313.950 154.950 316.050 157.050 ;
        RECT 164.400 133.050 165.450 154.950 ;
        RECT 40.950 130.950 43.050 133.050 ;
        RECT 163.950 130.950 166.050 133.050 ;
        RECT 164.400 130.050 165.450 130.950 ;
        RECT 163.950 127.950 166.050 130.050 ;
        RECT 299.400 33.450 300.450 154.950 ;
        RECT 296.400 32.400 300.450 33.450 ;
        RECT 296.400 -2.550 297.450 32.400 ;
        RECT 296.400 -3.600 300.450 -2.550 ;
      LAYER metal3 ;
        RECT 313.950 219.600 316.050 220.050 ;
        RECT 520.950 219.600 523.050 220.050 ;
        RECT 682.950 219.600 685.050 220.050 ;
        RECT 694.950 219.600 697.050 220.050 ;
        RECT 313.950 218.400 697.050 219.600 ;
        RECT 313.950 217.950 316.050 218.400 ;
        RECT 520.950 217.950 523.050 218.400 ;
        RECT 682.950 217.950 685.050 218.400 ;
        RECT 694.950 217.950 697.050 218.400 ;
        RECT 163.950 156.600 166.050 157.050 ;
        RECT 298.950 156.600 301.050 157.050 ;
        RECT 313.950 156.600 316.050 157.050 ;
        RECT 163.950 155.400 316.050 156.600 ;
        RECT 163.950 154.950 166.050 155.400 ;
        RECT 298.950 154.950 301.050 155.400 ;
        RECT 313.950 154.950 316.050 155.400 ;
        RECT 40.950 132.600 43.050 133.050 ;
        RECT 163.950 132.600 166.050 133.050 ;
        RECT 40.950 131.400 166.050 132.600 ;
        RECT 40.950 130.950 43.050 131.400 ;
        RECT 163.950 130.950 166.050 131.400 ;
    END
  END Yin[0]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 880.950 337.950 883.050 340.050 ;
      LAYER metal3 ;
        RECT 880.950 339.600 883.050 340.050 ;
        RECT 896.400 339.600 897.600 342.600 ;
        RECT 880.950 338.400 897.600 339.600 ;
        RECT 880.950 337.950 883.050 338.400 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 883.950 312.450 886.050 313.050 ;
        RECT 883.950 311.400 888.450 312.450 ;
        RECT 883.950 310.950 886.050 311.400 ;
        RECT 887.400 307.050 888.450 311.400 ;
        RECT 886.950 304.950 889.050 307.050 ;
      LAYER metal3 ;
        RECT 886.950 306.600 889.050 307.050 ;
        RECT 886.950 305.400 897.600 306.600 ;
        RECT 886.950 304.950 889.050 305.400 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 334.950 774.450 337.050 775.050 ;
        RECT 874.950 774.450 877.050 775.050 ;
        RECT 334.950 773.400 339.450 774.450 ;
        RECT 334.950 772.950 337.050 773.400 ;
        RECT 338.400 730.050 339.450 773.400 ;
        RECT 874.950 773.400 879.450 774.450 ;
        RECT 874.950 772.950 877.050 773.400 ;
        RECT 878.400 742.050 879.450 773.400 ;
        RECT 871.950 739.950 874.050 742.050 ;
        RECT 877.950 739.950 880.050 742.050 ;
        RECT 886.950 739.950 889.050 742.050 ;
        RECT 184.950 727.950 187.050 730.050 ;
        RECT 337.950 727.950 340.050 730.050 ;
        RECT 103.950 595.950 106.050 598.050 ;
        RECT 104.400 580.050 105.450 595.950 ;
        RECT 185.400 580.050 186.450 727.950 ;
        RECT 1.950 577.950 4.050 580.050 ;
        RECT 103.950 577.950 106.050 580.050 ;
        RECT 184.950 577.950 187.050 580.050 ;
        RECT 2.400 202.050 3.450 577.950 ;
        RECT 887.400 316.050 888.450 739.950 ;
        RECT 871.950 313.950 874.050 316.050 ;
        RECT 886.950 313.950 889.050 316.050 ;
        RECT 872.400 292.050 873.450 313.950 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 871.950 289.950 874.050 292.050 ;
        RECT 470.400 271.050 471.450 289.950 ;
        RECT 469.950 270.450 472.050 271.050 ;
        RECT 467.400 269.400 472.050 270.450 ;
        RECT 872.400 270.450 873.450 289.950 ;
        RECT 874.950 270.450 877.050 271.050 ;
        RECT 872.400 269.400 879.450 270.450 ;
        RECT 467.400 205.050 468.450 269.400 ;
        RECT 469.950 268.950 472.050 269.400 ;
        RECT 874.950 268.950 877.050 269.400 ;
        RECT 49.950 202.950 52.050 205.050 ;
        RECT 466.950 202.950 469.050 205.050 ;
        RECT 50.400 202.050 51.450 202.950 ;
        RECT 1.950 199.950 4.050 202.050 ;
        RECT 49.950 199.950 52.050 202.050 ;
        RECT 50.400 199.050 51.450 199.950 ;
        RECT 878.400 199.050 879.450 269.400 ;
        RECT 49.950 196.950 52.050 199.050 ;
        RECT 877.950 196.950 880.050 199.050 ;
      LAYER metal3 ;
        RECT 871.950 741.600 874.050 742.050 ;
        RECT 877.950 741.600 880.050 742.050 ;
        RECT 886.950 741.600 889.050 742.050 ;
        RECT 871.950 740.400 889.050 741.600 ;
        RECT 871.950 739.950 874.050 740.400 ;
        RECT 877.950 739.950 880.050 740.400 ;
        RECT 886.950 739.950 889.050 740.400 ;
        RECT 184.950 729.600 187.050 730.050 ;
        RECT 337.950 729.600 340.050 730.050 ;
        RECT 184.950 728.400 340.050 729.600 ;
        RECT 184.950 727.950 187.050 728.400 ;
        RECT 337.950 727.950 340.050 728.400 ;
        RECT 1.950 579.600 4.050 580.050 ;
        RECT 103.950 579.600 106.050 580.050 ;
        RECT 184.950 579.600 187.050 580.050 ;
        RECT 1.950 578.400 187.050 579.600 ;
        RECT 1.950 577.950 4.050 578.400 ;
        RECT 103.950 577.950 106.050 578.400 ;
        RECT 184.950 577.950 187.050 578.400 ;
        RECT 871.950 315.600 874.050 316.050 ;
        RECT 886.950 315.600 889.050 316.050 ;
        RECT 871.950 314.400 889.050 315.600 ;
        RECT 871.950 313.950 874.050 314.400 ;
        RECT 886.950 313.950 889.050 314.400 ;
        RECT 469.950 291.600 472.050 292.050 ;
        RECT 871.950 291.600 874.050 292.050 ;
        RECT 469.950 290.400 874.050 291.600 ;
        RECT 469.950 289.950 472.050 290.400 ;
        RECT 871.950 289.950 874.050 290.400 ;
        RECT 49.950 204.600 52.050 205.050 ;
        RECT 466.950 204.600 469.050 205.050 ;
        RECT 49.950 203.400 469.050 204.600 ;
        RECT 49.950 202.950 52.050 203.400 ;
        RECT 466.950 202.950 469.050 203.400 ;
        RECT 1.950 201.600 4.050 202.050 ;
        RECT 49.950 201.600 52.050 202.050 ;
        RECT -3.600 200.400 52.050 201.600 ;
        RECT 1.950 199.950 4.050 200.400 ;
        RECT 49.950 199.950 52.050 200.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 10.650 896.400 12.450 899.250 ;
        RECT 13.650 896.400 15.450 899.250 ;
        RECT 11.400 888.150 12.600 896.400 ;
        RECT 29.850 892.200 31.650 899.250 ;
        RECT 34.350 893.400 36.150 899.250 ;
        RECT 44.550 894.300 46.350 899.250 ;
        RECT 47.550 895.200 49.350 899.250 ;
        RECT 50.550 894.300 52.350 899.250 ;
        RECT 44.550 892.950 52.350 894.300 ;
        RECT 53.550 893.400 55.350 899.250 ;
        RECT 60.150 893.400 61.950 899.250 ;
        RECT 63.150 896.400 64.950 899.250 ;
        RECT 67.950 897.300 69.750 899.250 ;
        RECT 66.000 896.400 69.750 897.300 ;
        RECT 72.450 896.400 74.250 899.250 ;
        RECT 75.750 896.400 77.550 899.250 ;
        RECT 79.650 896.400 81.450 899.250 ;
        RECT 83.850 896.400 85.650 899.250 ;
        RECT 88.350 896.400 90.150 899.250 ;
        RECT 66.000 895.500 67.050 896.400 ;
        RECT 64.950 893.400 67.050 895.500 ;
        RECT 75.750 894.600 76.800 896.400 ;
        RECT 29.850 891.300 33.450 892.200 ;
        RECT 53.550 891.300 54.750 893.400 ;
        RECT 10.950 886.050 13.050 888.150 ;
        RECT 13.950 887.850 16.050 889.950 ;
        RECT 14.100 886.050 15.900 887.850 ;
        RECT 11.400 873.600 12.600 886.050 ;
        RECT 29.100 885.150 30.900 886.950 ;
        RECT 28.950 883.050 31.050 885.150 ;
        RECT 32.250 883.950 33.450 891.300 ;
        RECT 51.000 890.250 54.750 891.300 ;
        RECT 47.100 888.150 48.900 889.950 ;
        RECT 35.100 885.150 36.900 886.950 ;
        RECT 31.950 881.850 34.050 883.950 ;
        RECT 34.950 883.050 37.050 885.150 ;
        RECT 43.950 884.850 46.050 886.950 ;
        RECT 46.950 886.050 49.050 888.150 ;
        RECT 50.850 886.950 52.050 890.250 ;
        RECT 49.950 884.850 52.050 886.950 ;
        RECT 44.100 883.050 45.900 884.850 ;
        RECT 32.250 873.600 33.450 881.850 ;
        RECT 49.950 879.600 51.150 884.850 ;
        RECT 52.950 881.850 55.050 883.950 ;
        RECT 52.950 880.050 54.750 881.850 ;
        RECT 60.150 880.800 61.050 893.400 ;
        RECT 68.550 892.800 70.350 894.600 ;
        RECT 71.850 893.550 76.800 894.600 ;
        RECT 84.300 895.500 85.350 896.400 ;
        RECT 84.300 894.300 88.050 895.500 ;
        RECT 71.850 892.800 73.650 893.550 ;
        RECT 68.850 891.900 69.900 892.800 ;
        RECT 79.050 892.200 80.850 894.000 ;
        RECT 85.950 893.400 88.050 894.300 ;
        RECT 91.650 893.400 93.450 899.250 ;
        RECT 101.850 893.400 103.650 899.250 ;
        RECT 79.050 891.900 79.950 892.200 ;
        RECT 68.850 891.000 79.950 891.900 ;
        RECT 92.250 891.150 93.450 893.400 ;
        RECT 106.350 892.200 108.150 899.250 ;
        RECT 68.850 889.800 69.900 891.000 ;
        RECT 63.000 888.600 69.900 889.800 ;
        RECT 63.000 887.850 63.900 888.600 ;
        RECT 68.100 888.000 69.900 888.600 ;
        RECT 62.100 886.050 63.900 887.850 ;
        RECT 65.100 886.950 66.900 887.700 ;
        RECT 79.050 886.950 79.950 891.000 ;
        RECT 88.950 889.050 93.450 891.150 ;
        RECT 87.150 887.250 91.050 889.050 ;
        RECT 88.950 886.950 91.050 887.250 ;
        RECT 65.100 885.900 73.050 886.950 ;
        RECT 70.950 884.850 73.050 885.900 ;
        RECT 76.950 884.850 79.950 886.950 ;
        RECT 69.450 881.100 71.250 881.400 ;
        RECT 69.450 880.800 77.850 881.100 ;
        RECT 60.150 880.200 77.850 880.800 ;
        RECT 60.150 879.600 71.250 880.200 ;
        RECT 10.650 867.750 12.450 873.600 ;
        RECT 13.650 867.750 15.450 873.600 ;
        RECT 28.650 867.750 30.450 873.600 ;
        RECT 31.650 867.750 33.450 873.600 ;
        RECT 34.650 867.750 36.450 873.600 ;
        RECT 45.300 867.750 47.100 879.600 ;
        RECT 49.500 867.750 51.300 879.600 ;
        RECT 52.800 867.750 54.600 873.600 ;
        RECT 60.150 867.750 61.950 879.600 ;
        RECT 74.250 878.700 76.050 879.300 ;
        RECT 68.550 877.500 76.050 878.700 ;
        RECT 76.950 878.100 77.850 880.200 ;
        RECT 79.050 880.200 79.950 884.850 ;
        RECT 89.250 881.400 91.050 883.200 ;
        RECT 85.950 880.200 90.150 881.400 ;
        RECT 79.050 879.300 85.050 880.200 ;
        RECT 85.950 879.300 88.050 880.200 ;
        RECT 92.250 879.600 93.450 889.050 ;
        RECT 104.550 891.300 108.150 892.200 ;
        RECT 122.850 892.200 124.650 899.250 ;
        RECT 127.350 893.400 129.150 899.250 ;
        RECT 132.150 893.400 133.950 899.250 ;
        RECT 135.150 896.400 136.950 899.250 ;
        RECT 139.950 897.300 141.750 899.250 ;
        RECT 138.000 896.400 141.750 897.300 ;
        RECT 144.450 896.400 146.250 899.250 ;
        RECT 147.750 896.400 149.550 899.250 ;
        RECT 151.650 896.400 153.450 899.250 ;
        RECT 155.850 896.400 157.650 899.250 ;
        RECT 160.350 896.400 162.150 899.250 ;
        RECT 138.000 895.500 139.050 896.400 ;
        RECT 136.950 893.400 139.050 895.500 ;
        RECT 147.750 894.600 148.800 896.400 ;
        RECT 122.850 891.300 126.450 892.200 ;
        RECT 101.100 885.150 102.900 886.950 ;
        RECT 100.950 883.050 103.050 885.150 ;
        RECT 104.550 883.950 105.750 891.300 ;
        RECT 107.100 885.150 108.900 886.950 ;
        RECT 122.100 885.150 123.900 886.950 ;
        RECT 103.950 881.850 106.050 883.950 ;
        RECT 106.950 883.050 109.050 885.150 ;
        RECT 121.950 883.050 124.050 885.150 ;
        RECT 125.250 883.950 126.450 891.300 ;
        RECT 128.100 885.150 129.900 886.950 ;
        RECT 124.950 881.850 127.050 883.950 ;
        RECT 127.950 883.050 130.050 885.150 ;
        RECT 84.150 878.400 85.050 879.300 ;
        RECT 81.450 878.100 83.250 878.400 ;
        RECT 68.550 876.600 69.750 877.500 ;
        RECT 76.950 877.200 83.250 878.100 ;
        RECT 81.450 876.600 83.250 877.200 ;
        RECT 84.150 876.600 86.850 878.400 ;
        RECT 64.950 874.500 69.750 876.600 ;
        RECT 72.150 874.500 79.050 876.300 ;
        RECT 68.550 873.600 69.750 874.500 ;
        RECT 63.150 867.750 64.950 873.600 ;
        RECT 68.250 867.750 70.050 873.600 ;
        RECT 73.050 867.750 74.850 873.600 ;
        RECT 76.050 867.750 77.850 874.500 ;
        RECT 84.150 873.600 88.050 875.700 ;
        RECT 79.950 867.750 81.750 873.600 ;
        RECT 84.150 867.750 85.950 873.600 ;
        RECT 88.650 867.750 90.450 870.600 ;
        RECT 91.650 867.750 93.450 879.600 ;
        RECT 104.550 873.600 105.750 881.850 ;
        RECT 125.250 873.600 126.450 881.850 ;
        RECT 132.150 880.800 133.050 893.400 ;
        RECT 140.550 892.800 142.350 894.600 ;
        RECT 143.850 893.550 148.800 894.600 ;
        RECT 156.300 895.500 157.350 896.400 ;
        RECT 156.300 894.300 160.050 895.500 ;
        RECT 143.850 892.800 145.650 893.550 ;
        RECT 140.850 891.900 141.900 892.800 ;
        RECT 151.050 892.200 152.850 894.000 ;
        RECT 157.950 893.400 160.050 894.300 ;
        RECT 163.650 893.400 165.450 899.250 ;
        RECT 176.550 896.400 178.350 899.250 ;
        RECT 179.550 896.400 181.350 899.250 ;
        RECT 151.050 891.900 151.950 892.200 ;
        RECT 140.850 891.000 151.950 891.900 ;
        RECT 164.250 891.150 165.450 893.400 ;
        RECT 140.850 889.800 141.900 891.000 ;
        RECT 135.000 888.600 141.900 889.800 ;
        RECT 135.000 887.850 135.900 888.600 ;
        RECT 140.100 888.000 141.900 888.600 ;
        RECT 134.100 886.050 135.900 887.850 ;
        RECT 137.100 886.950 138.900 887.700 ;
        RECT 151.050 886.950 151.950 891.000 ;
        RECT 160.950 889.050 165.450 891.150 ;
        RECT 159.150 887.250 163.050 889.050 ;
        RECT 160.950 886.950 163.050 887.250 ;
        RECT 137.100 885.900 145.050 886.950 ;
        RECT 142.950 884.850 145.050 885.900 ;
        RECT 148.950 884.850 151.950 886.950 ;
        RECT 141.450 881.100 143.250 881.400 ;
        RECT 141.450 880.800 149.850 881.100 ;
        RECT 132.150 880.200 149.850 880.800 ;
        RECT 132.150 879.600 143.250 880.200 ;
        RECT 101.550 867.750 103.350 873.600 ;
        RECT 104.550 867.750 106.350 873.600 ;
        RECT 107.550 867.750 109.350 873.600 ;
        RECT 121.650 867.750 123.450 873.600 ;
        RECT 124.650 867.750 126.450 873.600 ;
        RECT 127.650 867.750 129.450 873.600 ;
        RECT 132.150 867.750 133.950 879.600 ;
        RECT 146.250 878.700 148.050 879.300 ;
        RECT 140.550 877.500 148.050 878.700 ;
        RECT 148.950 878.100 149.850 880.200 ;
        RECT 151.050 880.200 151.950 884.850 ;
        RECT 161.250 881.400 163.050 883.200 ;
        RECT 157.950 880.200 162.150 881.400 ;
        RECT 151.050 879.300 157.050 880.200 ;
        RECT 157.950 879.300 160.050 880.200 ;
        RECT 164.250 879.600 165.450 889.050 ;
        RECT 175.950 887.850 178.050 889.950 ;
        RECT 179.400 888.150 180.600 896.400 ;
        RECT 197.850 892.200 199.650 899.250 ;
        RECT 202.350 893.400 204.150 899.250 ;
        RECT 207.150 893.400 208.950 899.250 ;
        RECT 210.150 896.400 211.950 899.250 ;
        RECT 214.950 897.300 216.750 899.250 ;
        RECT 213.000 896.400 216.750 897.300 ;
        RECT 219.450 896.400 221.250 899.250 ;
        RECT 222.750 896.400 224.550 899.250 ;
        RECT 226.650 896.400 228.450 899.250 ;
        RECT 230.850 896.400 232.650 899.250 ;
        RECT 235.350 896.400 237.150 899.250 ;
        RECT 213.000 895.500 214.050 896.400 ;
        RECT 211.950 893.400 214.050 895.500 ;
        RECT 222.750 894.600 223.800 896.400 ;
        RECT 197.850 891.300 201.450 892.200 ;
        RECT 176.100 886.050 177.900 887.850 ;
        RECT 178.950 886.050 181.050 888.150 ;
        RECT 156.150 878.400 157.050 879.300 ;
        RECT 153.450 878.100 155.250 878.400 ;
        RECT 140.550 876.600 141.750 877.500 ;
        RECT 148.950 877.200 155.250 878.100 ;
        RECT 153.450 876.600 155.250 877.200 ;
        RECT 156.150 876.600 158.850 878.400 ;
        RECT 136.950 874.500 141.750 876.600 ;
        RECT 144.150 874.500 151.050 876.300 ;
        RECT 140.550 873.600 141.750 874.500 ;
        RECT 135.150 867.750 136.950 873.600 ;
        RECT 140.250 867.750 142.050 873.600 ;
        RECT 145.050 867.750 146.850 873.600 ;
        RECT 148.050 867.750 149.850 874.500 ;
        RECT 156.150 873.600 160.050 875.700 ;
        RECT 151.950 867.750 153.750 873.600 ;
        RECT 156.150 867.750 157.950 873.600 ;
        RECT 160.650 867.750 162.450 870.600 ;
        RECT 163.650 867.750 165.450 879.600 ;
        RECT 179.400 873.600 180.600 886.050 ;
        RECT 197.100 885.150 198.900 886.950 ;
        RECT 196.950 883.050 199.050 885.150 ;
        RECT 200.250 883.950 201.450 891.300 ;
        RECT 203.100 885.150 204.900 886.950 ;
        RECT 199.950 881.850 202.050 883.950 ;
        RECT 202.950 883.050 205.050 885.150 ;
        RECT 200.250 873.600 201.450 881.850 ;
        RECT 207.150 880.800 208.050 893.400 ;
        RECT 215.550 892.800 217.350 894.600 ;
        RECT 218.850 893.550 223.800 894.600 ;
        RECT 231.300 895.500 232.350 896.400 ;
        RECT 231.300 894.300 235.050 895.500 ;
        RECT 218.850 892.800 220.650 893.550 ;
        RECT 215.850 891.900 216.900 892.800 ;
        RECT 226.050 892.200 227.850 894.000 ;
        RECT 232.950 893.400 235.050 894.300 ;
        RECT 238.650 893.400 240.450 899.250 ;
        RECT 251.550 896.400 253.350 899.250 ;
        RECT 254.550 896.400 256.350 899.250 ;
        RECT 226.050 891.900 226.950 892.200 ;
        RECT 215.850 891.000 226.950 891.900 ;
        RECT 239.250 891.150 240.450 893.400 ;
        RECT 215.850 889.800 216.900 891.000 ;
        RECT 210.000 888.600 216.900 889.800 ;
        RECT 210.000 887.850 210.900 888.600 ;
        RECT 215.100 888.000 216.900 888.600 ;
        RECT 209.100 886.050 210.900 887.850 ;
        RECT 212.100 886.950 213.900 887.700 ;
        RECT 226.050 886.950 226.950 891.000 ;
        RECT 235.950 889.050 240.450 891.150 ;
        RECT 234.150 887.250 238.050 889.050 ;
        RECT 235.950 886.950 238.050 887.250 ;
        RECT 212.100 885.900 220.050 886.950 ;
        RECT 217.950 884.850 220.050 885.900 ;
        RECT 223.950 884.850 226.950 886.950 ;
        RECT 216.450 881.100 218.250 881.400 ;
        RECT 216.450 880.800 224.850 881.100 ;
        RECT 207.150 880.200 224.850 880.800 ;
        RECT 207.150 879.600 218.250 880.200 ;
        RECT 176.550 867.750 178.350 873.600 ;
        RECT 179.550 867.750 181.350 873.600 ;
        RECT 196.650 867.750 198.450 873.600 ;
        RECT 199.650 867.750 201.450 873.600 ;
        RECT 202.650 867.750 204.450 873.600 ;
        RECT 207.150 867.750 208.950 879.600 ;
        RECT 221.250 878.700 223.050 879.300 ;
        RECT 215.550 877.500 223.050 878.700 ;
        RECT 223.950 878.100 224.850 880.200 ;
        RECT 226.050 880.200 226.950 884.850 ;
        RECT 236.250 881.400 238.050 883.200 ;
        RECT 232.950 880.200 237.150 881.400 ;
        RECT 226.050 879.300 232.050 880.200 ;
        RECT 232.950 879.300 235.050 880.200 ;
        RECT 239.250 879.600 240.450 889.050 ;
        RECT 250.950 887.850 253.050 889.950 ;
        RECT 254.400 888.150 255.600 896.400 ;
        RECT 271.650 893.400 273.450 899.250 ;
        RECT 272.250 891.300 273.450 893.400 ;
        RECT 274.650 894.300 276.450 899.250 ;
        RECT 277.650 895.200 279.450 899.250 ;
        RECT 280.650 894.300 282.450 899.250 ;
        RECT 274.650 892.950 282.450 894.300 ;
        RECT 285.150 893.400 286.950 899.250 ;
        RECT 288.150 896.400 289.950 899.250 ;
        RECT 292.950 897.300 294.750 899.250 ;
        RECT 291.000 896.400 294.750 897.300 ;
        RECT 297.450 896.400 299.250 899.250 ;
        RECT 300.750 896.400 302.550 899.250 ;
        RECT 304.650 896.400 306.450 899.250 ;
        RECT 308.850 896.400 310.650 899.250 ;
        RECT 313.350 896.400 315.150 899.250 ;
        RECT 291.000 895.500 292.050 896.400 ;
        RECT 289.950 893.400 292.050 895.500 ;
        RECT 300.750 894.600 301.800 896.400 ;
        RECT 272.250 890.250 276.000 891.300 ;
        RECT 251.100 886.050 252.900 887.850 ;
        RECT 253.950 886.050 256.050 888.150 ;
        RECT 274.950 886.950 276.150 890.250 ;
        RECT 278.100 888.150 279.900 889.950 ;
        RECT 231.150 878.400 232.050 879.300 ;
        RECT 228.450 878.100 230.250 878.400 ;
        RECT 215.550 876.600 216.750 877.500 ;
        RECT 223.950 877.200 230.250 878.100 ;
        RECT 228.450 876.600 230.250 877.200 ;
        RECT 231.150 876.600 233.850 878.400 ;
        RECT 211.950 874.500 216.750 876.600 ;
        RECT 219.150 874.500 226.050 876.300 ;
        RECT 215.550 873.600 216.750 874.500 ;
        RECT 210.150 867.750 211.950 873.600 ;
        RECT 215.250 867.750 217.050 873.600 ;
        RECT 220.050 867.750 221.850 873.600 ;
        RECT 223.050 867.750 224.850 874.500 ;
        RECT 231.150 873.600 235.050 875.700 ;
        RECT 226.950 867.750 228.750 873.600 ;
        RECT 231.150 867.750 232.950 873.600 ;
        RECT 235.650 867.750 237.450 870.600 ;
        RECT 238.650 867.750 240.450 879.600 ;
        RECT 254.400 873.600 255.600 886.050 ;
        RECT 274.950 884.850 277.050 886.950 ;
        RECT 277.950 886.050 280.050 888.150 ;
        RECT 280.950 884.850 283.050 886.950 ;
        RECT 271.950 881.850 274.050 883.950 ;
        RECT 272.250 880.050 274.050 881.850 ;
        RECT 275.850 879.600 277.050 884.850 ;
        RECT 281.100 883.050 282.900 884.850 ;
        RECT 285.150 880.800 286.050 893.400 ;
        RECT 293.550 892.800 295.350 894.600 ;
        RECT 296.850 893.550 301.800 894.600 ;
        RECT 309.300 895.500 310.350 896.400 ;
        RECT 309.300 894.300 313.050 895.500 ;
        RECT 296.850 892.800 298.650 893.550 ;
        RECT 293.850 891.900 294.900 892.800 ;
        RECT 304.050 892.200 305.850 894.000 ;
        RECT 310.950 893.400 313.050 894.300 ;
        RECT 316.650 893.400 318.450 899.250 ;
        RECT 326.550 896.400 328.350 899.250 ;
        RECT 329.550 896.400 331.350 899.250 ;
        RECT 341.550 896.400 343.350 899.250 ;
        RECT 304.050 891.900 304.950 892.200 ;
        RECT 293.850 891.000 304.950 891.900 ;
        RECT 317.250 891.150 318.450 893.400 ;
        RECT 293.850 889.800 294.900 891.000 ;
        RECT 288.000 888.600 294.900 889.800 ;
        RECT 288.000 887.850 288.900 888.600 ;
        RECT 293.100 888.000 294.900 888.600 ;
        RECT 287.100 886.050 288.900 887.850 ;
        RECT 290.100 886.950 291.900 887.700 ;
        RECT 304.050 886.950 304.950 891.000 ;
        RECT 313.950 889.050 318.450 891.150 ;
        RECT 312.150 887.250 316.050 889.050 ;
        RECT 313.950 886.950 316.050 887.250 ;
        RECT 290.100 885.900 298.050 886.950 ;
        RECT 295.950 884.850 298.050 885.900 ;
        RECT 301.950 884.850 304.950 886.950 ;
        RECT 294.450 881.100 296.250 881.400 ;
        RECT 294.450 880.800 302.850 881.100 ;
        RECT 285.150 880.200 302.850 880.800 ;
        RECT 285.150 879.600 296.250 880.200 ;
        RECT 251.550 867.750 253.350 873.600 ;
        RECT 254.550 867.750 256.350 873.600 ;
        RECT 272.400 867.750 274.200 873.600 ;
        RECT 275.700 867.750 277.500 879.600 ;
        RECT 279.900 867.750 281.700 879.600 ;
        RECT 285.150 867.750 286.950 879.600 ;
        RECT 299.250 878.700 301.050 879.300 ;
        RECT 293.550 877.500 301.050 878.700 ;
        RECT 301.950 878.100 302.850 880.200 ;
        RECT 304.050 880.200 304.950 884.850 ;
        RECT 314.250 881.400 316.050 883.200 ;
        RECT 310.950 880.200 315.150 881.400 ;
        RECT 304.050 879.300 310.050 880.200 ;
        RECT 310.950 879.300 313.050 880.200 ;
        RECT 317.250 879.600 318.450 889.050 ;
        RECT 325.950 887.850 328.050 889.950 ;
        RECT 329.400 888.150 330.600 896.400 ;
        RECT 342.150 892.500 343.350 896.400 ;
        RECT 344.850 893.400 346.650 899.250 ;
        RECT 347.850 893.400 349.650 899.250 ;
        RECT 342.150 891.600 347.250 892.500 ;
        RECT 345.000 890.700 347.250 891.600 ;
        RECT 326.100 886.050 327.900 887.850 ;
        RECT 328.950 886.050 331.050 888.150 ;
        RECT 309.150 878.400 310.050 879.300 ;
        RECT 306.450 878.100 308.250 878.400 ;
        RECT 293.550 876.600 294.750 877.500 ;
        RECT 301.950 877.200 308.250 878.100 ;
        RECT 306.450 876.600 308.250 877.200 ;
        RECT 309.150 876.600 311.850 878.400 ;
        RECT 289.950 874.500 294.750 876.600 ;
        RECT 297.150 874.500 304.050 876.300 ;
        RECT 293.550 873.600 294.750 874.500 ;
        RECT 288.150 867.750 289.950 873.600 ;
        RECT 293.250 867.750 295.050 873.600 ;
        RECT 298.050 867.750 299.850 873.600 ;
        RECT 301.050 867.750 302.850 874.500 ;
        RECT 309.150 873.600 313.050 875.700 ;
        RECT 304.950 867.750 306.750 873.600 ;
        RECT 309.150 867.750 310.950 873.600 ;
        RECT 313.650 867.750 315.450 870.600 ;
        RECT 316.650 867.750 318.450 879.600 ;
        RECT 329.400 873.600 330.600 886.050 ;
        RECT 340.950 884.850 343.050 886.950 ;
        RECT 341.100 883.050 342.900 884.850 ;
        RECT 345.000 882.300 346.050 890.700 ;
        RECT 348.150 886.950 349.350 893.400 ;
        RECT 365.850 892.200 367.650 899.250 ;
        RECT 370.350 893.400 372.150 899.250 ;
        RECT 380.550 896.400 382.350 899.250 ;
        RECT 383.550 896.400 385.350 899.250 ;
        RECT 386.550 896.400 388.350 899.250 ;
        RECT 365.850 891.300 369.450 892.200 ;
        RECT 346.950 884.850 349.350 886.950 ;
        RECT 365.100 885.150 366.900 886.950 ;
        RECT 345.000 881.400 347.250 882.300 ;
        RECT 341.550 880.500 347.250 881.400 ;
        RECT 341.550 873.600 342.750 880.500 ;
        RECT 348.150 879.600 349.350 884.850 ;
        RECT 364.950 883.050 367.050 885.150 ;
        RECT 368.250 883.950 369.450 891.300 ;
        RECT 384.000 889.950 385.050 896.400 ;
        RECT 398.550 894.300 400.350 899.250 ;
        RECT 401.550 895.200 403.350 899.250 ;
        RECT 404.550 894.300 406.350 899.250 ;
        RECT 398.550 892.950 406.350 894.300 ;
        RECT 407.550 893.400 409.350 899.250 ;
        RECT 414.150 893.400 415.950 899.250 ;
        RECT 417.150 896.400 418.950 899.250 ;
        RECT 421.950 897.300 423.750 899.250 ;
        RECT 420.000 896.400 423.750 897.300 ;
        RECT 426.450 896.400 428.250 899.250 ;
        RECT 429.750 896.400 431.550 899.250 ;
        RECT 433.650 896.400 435.450 899.250 ;
        RECT 437.850 896.400 439.650 899.250 ;
        RECT 442.350 896.400 444.150 899.250 ;
        RECT 420.000 895.500 421.050 896.400 ;
        RECT 418.950 893.400 421.050 895.500 ;
        RECT 429.750 894.600 430.800 896.400 ;
        RECT 407.550 891.300 408.750 893.400 ;
        RECT 405.000 890.250 408.750 891.300 ;
        RECT 382.950 887.850 385.050 889.950 ;
        RECT 401.100 888.150 402.900 889.950 ;
        RECT 371.100 885.150 372.900 886.950 ;
        RECT 367.950 881.850 370.050 883.950 ;
        RECT 370.950 883.050 373.050 885.150 ;
        RECT 379.950 884.850 382.050 886.950 ;
        RECT 380.100 883.050 381.900 884.850 ;
        RECT 326.550 867.750 328.350 873.600 ;
        RECT 329.550 867.750 331.350 873.600 ;
        RECT 341.550 867.750 343.350 873.600 ;
        RECT 344.850 867.750 346.650 879.600 ;
        RECT 347.850 867.750 349.650 879.600 ;
        RECT 368.250 873.600 369.450 881.850 ;
        RECT 384.000 880.650 385.050 887.850 ;
        RECT 385.950 884.850 388.050 886.950 ;
        RECT 397.950 884.850 400.050 886.950 ;
        RECT 400.950 886.050 403.050 888.150 ;
        RECT 404.850 886.950 406.050 890.250 ;
        RECT 403.950 884.850 406.050 886.950 ;
        RECT 386.100 883.050 387.900 884.850 ;
        RECT 398.100 883.050 399.900 884.850 ;
        RECT 370.950 879.450 373.050 880.050 ;
        RECT 376.950 879.450 379.050 880.050 ;
        RECT 384.000 879.600 386.550 880.650 ;
        RECT 403.950 879.600 405.150 884.850 ;
        RECT 406.950 881.850 409.050 883.950 ;
        RECT 406.950 880.050 408.750 881.850 ;
        RECT 414.150 880.800 415.050 893.400 ;
        RECT 422.550 892.800 424.350 894.600 ;
        RECT 425.850 893.550 430.800 894.600 ;
        RECT 438.300 895.500 439.350 896.400 ;
        RECT 438.300 894.300 442.050 895.500 ;
        RECT 425.850 892.800 427.650 893.550 ;
        RECT 422.850 891.900 423.900 892.800 ;
        RECT 433.050 892.200 434.850 894.000 ;
        RECT 439.950 893.400 442.050 894.300 ;
        RECT 445.650 893.400 447.450 899.250 ;
        RECT 455.850 893.400 457.650 899.250 ;
        RECT 433.050 891.900 433.950 892.200 ;
        RECT 422.850 891.000 433.950 891.900 ;
        RECT 446.250 891.150 447.450 893.400 ;
        RECT 460.350 892.200 462.150 899.250 ;
        RECT 422.850 889.800 423.900 891.000 ;
        RECT 417.000 888.600 423.900 889.800 ;
        RECT 417.000 887.850 417.900 888.600 ;
        RECT 422.100 888.000 423.900 888.600 ;
        RECT 416.100 886.050 417.900 887.850 ;
        RECT 419.100 886.950 420.900 887.700 ;
        RECT 433.050 886.950 433.950 891.000 ;
        RECT 442.950 889.050 447.450 891.150 ;
        RECT 441.150 887.250 445.050 889.050 ;
        RECT 442.950 886.950 445.050 887.250 ;
        RECT 419.100 885.900 427.050 886.950 ;
        RECT 424.950 884.850 427.050 885.900 ;
        RECT 430.950 884.850 433.950 886.950 ;
        RECT 423.450 881.100 425.250 881.400 ;
        RECT 423.450 880.800 431.850 881.100 ;
        RECT 414.150 880.200 431.850 880.800 ;
        RECT 414.150 879.600 425.250 880.200 ;
        RECT 370.950 878.550 379.050 879.450 ;
        RECT 370.950 877.950 373.050 878.550 ;
        RECT 376.950 877.950 379.050 878.550 ;
        RECT 364.650 867.750 366.450 873.600 ;
        RECT 367.650 867.750 369.450 873.600 ;
        RECT 370.650 867.750 372.450 873.600 ;
        RECT 380.550 867.750 382.350 879.600 ;
        RECT 384.750 867.750 386.550 879.600 ;
        RECT 399.300 867.750 401.100 879.600 ;
        RECT 403.500 867.750 405.300 879.600 ;
        RECT 406.800 867.750 408.600 873.600 ;
        RECT 414.150 867.750 415.950 879.600 ;
        RECT 428.250 878.700 430.050 879.300 ;
        RECT 422.550 877.500 430.050 878.700 ;
        RECT 430.950 878.100 431.850 880.200 ;
        RECT 433.050 880.200 433.950 884.850 ;
        RECT 443.250 881.400 445.050 883.200 ;
        RECT 439.950 880.200 444.150 881.400 ;
        RECT 433.050 879.300 439.050 880.200 ;
        RECT 439.950 879.300 442.050 880.200 ;
        RECT 446.250 879.600 447.450 889.050 ;
        RECT 458.550 891.300 462.150 892.200 ;
        RECT 468.150 893.400 469.950 899.250 ;
        RECT 471.150 896.400 472.950 899.250 ;
        RECT 475.950 897.300 477.750 899.250 ;
        RECT 474.000 896.400 477.750 897.300 ;
        RECT 480.450 896.400 482.250 899.250 ;
        RECT 483.750 896.400 485.550 899.250 ;
        RECT 487.650 896.400 489.450 899.250 ;
        RECT 491.850 896.400 493.650 899.250 ;
        RECT 496.350 896.400 498.150 899.250 ;
        RECT 474.000 895.500 475.050 896.400 ;
        RECT 472.950 893.400 475.050 895.500 ;
        RECT 483.750 894.600 484.800 896.400 ;
        RECT 455.100 885.150 456.900 886.950 ;
        RECT 454.950 883.050 457.050 885.150 ;
        RECT 458.550 883.950 459.750 891.300 ;
        RECT 461.100 885.150 462.900 886.950 ;
        RECT 457.950 881.850 460.050 883.950 ;
        RECT 460.950 883.050 463.050 885.150 ;
        RECT 438.150 878.400 439.050 879.300 ;
        RECT 435.450 878.100 437.250 878.400 ;
        RECT 422.550 876.600 423.750 877.500 ;
        RECT 430.950 877.200 437.250 878.100 ;
        RECT 435.450 876.600 437.250 877.200 ;
        RECT 438.150 876.600 440.850 878.400 ;
        RECT 418.950 874.500 423.750 876.600 ;
        RECT 426.150 874.500 433.050 876.300 ;
        RECT 422.550 873.600 423.750 874.500 ;
        RECT 417.150 867.750 418.950 873.600 ;
        RECT 422.250 867.750 424.050 873.600 ;
        RECT 427.050 867.750 428.850 873.600 ;
        RECT 430.050 867.750 431.850 874.500 ;
        RECT 438.150 873.600 442.050 875.700 ;
        RECT 433.950 867.750 435.750 873.600 ;
        RECT 438.150 867.750 439.950 873.600 ;
        RECT 442.650 867.750 444.450 870.600 ;
        RECT 445.650 867.750 447.450 879.600 ;
        RECT 458.550 873.600 459.750 881.850 ;
        RECT 468.150 880.800 469.050 893.400 ;
        RECT 476.550 892.800 478.350 894.600 ;
        RECT 479.850 893.550 484.800 894.600 ;
        RECT 492.300 895.500 493.350 896.400 ;
        RECT 492.300 894.300 496.050 895.500 ;
        RECT 479.850 892.800 481.650 893.550 ;
        RECT 476.850 891.900 477.900 892.800 ;
        RECT 487.050 892.200 488.850 894.000 ;
        RECT 493.950 893.400 496.050 894.300 ;
        RECT 499.650 893.400 501.450 899.250 ;
        RECT 509.550 896.400 511.350 899.250 ;
        RECT 512.550 896.400 514.350 899.250 ;
        RECT 524.550 896.400 526.350 899.250 ;
        RECT 527.550 896.400 529.350 899.250 ;
        RECT 545.700 896.400 547.500 899.250 ;
        RECT 487.050 891.900 487.950 892.200 ;
        RECT 476.850 891.000 487.950 891.900 ;
        RECT 500.250 891.150 501.450 893.400 ;
        RECT 476.850 889.800 477.900 891.000 ;
        RECT 471.000 888.600 477.900 889.800 ;
        RECT 471.000 887.850 471.900 888.600 ;
        RECT 476.100 888.000 477.900 888.600 ;
        RECT 470.100 886.050 471.900 887.850 ;
        RECT 473.100 886.950 474.900 887.700 ;
        RECT 487.050 886.950 487.950 891.000 ;
        RECT 496.950 889.050 501.450 891.150 ;
        RECT 495.150 887.250 499.050 889.050 ;
        RECT 496.950 886.950 499.050 887.250 ;
        RECT 473.100 885.900 481.050 886.950 ;
        RECT 478.950 884.850 481.050 885.900 ;
        RECT 484.950 884.850 487.950 886.950 ;
        RECT 477.450 881.100 479.250 881.400 ;
        RECT 477.450 880.800 485.850 881.100 ;
        RECT 468.150 880.200 485.850 880.800 ;
        RECT 468.150 879.600 479.250 880.200 ;
        RECT 455.550 867.750 457.350 873.600 ;
        RECT 458.550 867.750 460.350 873.600 ;
        RECT 461.550 867.750 463.350 873.600 ;
        RECT 468.150 867.750 469.950 879.600 ;
        RECT 482.250 878.700 484.050 879.300 ;
        RECT 476.550 877.500 484.050 878.700 ;
        RECT 484.950 878.100 485.850 880.200 ;
        RECT 487.050 880.200 487.950 884.850 ;
        RECT 497.250 881.400 499.050 883.200 ;
        RECT 493.950 880.200 498.150 881.400 ;
        RECT 487.050 879.300 493.050 880.200 ;
        RECT 493.950 879.300 496.050 880.200 ;
        RECT 500.250 879.600 501.450 889.050 ;
        RECT 508.950 887.850 511.050 889.950 ;
        RECT 512.400 888.150 513.600 896.400 ;
        RECT 509.100 886.050 510.900 887.850 ;
        RECT 511.950 886.050 514.050 888.150 ;
        RECT 523.950 887.850 526.050 889.950 ;
        RECT 527.400 888.150 528.600 896.400 ;
        RECT 549.000 895.050 550.800 899.250 ;
        RECT 545.100 893.400 550.800 895.050 ;
        RECT 553.200 893.400 555.000 899.250 ;
        RECT 565.650 896.400 567.450 899.250 ;
        RECT 568.650 896.400 570.450 899.250 ;
        RECT 578.550 896.400 580.350 899.250 ;
        RECT 581.550 896.400 583.350 899.250 ;
        RECT 584.550 896.400 586.350 899.250 ;
        RECT 599.550 896.400 601.350 899.250 ;
        RECT 602.550 896.400 604.350 899.250 ;
        RECT 524.100 886.050 525.900 887.850 ;
        RECT 526.950 886.050 529.050 888.150 ;
        RECT 545.100 886.950 546.300 893.400 ;
        RECT 548.100 888.150 549.900 889.950 ;
        RECT 492.150 878.400 493.050 879.300 ;
        RECT 489.450 878.100 491.250 878.400 ;
        RECT 476.550 876.600 477.750 877.500 ;
        RECT 484.950 877.200 491.250 878.100 ;
        RECT 489.450 876.600 491.250 877.200 ;
        RECT 492.150 876.600 494.850 878.400 ;
        RECT 472.950 874.500 477.750 876.600 ;
        RECT 480.150 874.500 487.050 876.300 ;
        RECT 476.550 873.600 477.750 874.500 ;
        RECT 471.150 867.750 472.950 873.600 ;
        RECT 476.250 867.750 478.050 873.600 ;
        RECT 481.050 867.750 482.850 873.600 ;
        RECT 484.050 867.750 485.850 874.500 ;
        RECT 492.150 873.600 496.050 875.700 ;
        RECT 487.950 867.750 489.750 873.600 ;
        RECT 492.150 867.750 493.950 873.600 ;
        RECT 496.650 867.750 498.450 870.600 ;
        RECT 499.650 867.750 501.450 879.600 ;
        RECT 512.400 873.600 513.600 886.050 ;
        RECT 527.400 873.600 528.600 886.050 ;
        RECT 544.950 884.850 547.050 886.950 ;
        RECT 547.950 886.050 550.050 888.150 ;
        RECT 550.950 887.850 553.050 889.950 ;
        RECT 554.100 888.150 555.900 889.950 ;
        RECT 566.400 888.150 567.600 896.400 ;
        RECT 582.000 889.950 583.050 896.400 ;
        RECT 551.100 886.050 552.900 887.850 ;
        RECT 553.950 886.050 556.050 888.150 ;
        RECT 565.950 886.050 568.050 888.150 ;
        RECT 568.950 887.850 571.050 889.950 ;
        RECT 580.950 887.850 583.050 889.950 ;
        RECT 598.950 887.850 601.050 889.950 ;
        RECT 602.400 888.150 603.600 896.400 ;
        RECT 614.550 894.300 616.350 899.250 ;
        RECT 617.550 895.200 619.350 899.250 ;
        RECT 620.550 894.300 622.350 899.250 ;
        RECT 614.550 892.950 622.350 894.300 ;
        RECT 623.550 893.400 625.350 899.250 ;
        RECT 638.550 894.300 640.350 899.250 ;
        RECT 641.550 895.200 643.350 899.250 ;
        RECT 644.550 894.300 646.350 899.250 ;
        RECT 607.950 891.450 610.050 892.050 ;
        RECT 613.950 891.450 616.050 892.050 ;
        RECT 607.950 890.550 616.050 891.450 ;
        RECT 623.550 891.300 624.750 893.400 ;
        RECT 638.550 892.950 646.350 894.300 ;
        RECT 647.550 893.400 649.350 899.250 ;
        RECT 662.550 896.400 664.350 899.250 ;
        RECT 647.550 891.300 648.750 893.400 ;
        RECT 663.150 892.500 664.350 896.400 ;
        RECT 665.850 893.400 667.650 899.250 ;
        RECT 668.850 893.400 670.650 899.250 ;
        RECT 675.150 893.400 676.950 899.250 ;
        RECT 678.150 896.400 679.950 899.250 ;
        RECT 682.950 897.300 684.750 899.250 ;
        RECT 681.000 896.400 684.750 897.300 ;
        RECT 687.450 896.400 689.250 899.250 ;
        RECT 690.750 896.400 692.550 899.250 ;
        RECT 694.650 896.400 696.450 899.250 ;
        RECT 698.850 896.400 700.650 899.250 ;
        RECT 703.350 896.400 705.150 899.250 ;
        RECT 681.000 895.500 682.050 896.400 ;
        RECT 679.950 893.400 682.050 895.500 ;
        RECT 690.750 894.600 691.800 896.400 ;
        RECT 663.150 891.600 668.250 892.500 ;
        RECT 607.950 889.950 610.050 890.550 ;
        RECT 613.950 889.950 616.050 890.550 ;
        RECT 621.000 890.250 624.750 891.300 ;
        RECT 645.000 890.250 648.750 891.300 ;
        RECT 666.000 890.700 668.250 891.600 ;
        RECT 617.100 888.150 618.900 889.950 ;
        RECT 569.100 886.050 570.900 887.850 ;
        RECT 545.100 879.600 546.300 884.850 ;
        RECT 509.550 867.750 511.350 873.600 ;
        RECT 512.550 867.750 514.350 873.600 ;
        RECT 524.550 867.750 526.350 873.600 ;
        RECT 527.550 867.750 529.350 873.600 ;
        RECT 544.650 867.750 546.450 879.600 ;
        RECT 547.650 878.700 555.450 879.600 ;
        RECT 547.650 867.750 549.450 878.700 ;
        RECT 550.650 867.750 552.450 877.800 ;
        RECT 553.650 867.750 555.450 878.700 ;
        RECT 566.400 873.600 567.600 886.050 ;
        RECT 577.950 884.850 580.050 886.950 ;
        RECT 578.100 883.050 579.900 884.850 ;
        RECT 582.000 880.650 583.050 887.850 ;
        RECT 583.950 884.850 586.050 886.950 ;
        RECT 599.100 886.050 600.900 887.850 ;
        RECT 601.950 886.050 604.050 888.150 ;
        RECT 584.100 883.050 585.900 884.850 ;
        RECT 582.000 879.600 584.550 880.650 ;
        RECT 565.650 867.750 567.450 873.600 ;
        RECT 568.650 867.750 570.450 873.600 ;
        RECT 578.550 867.750 580.350 879.600 ;
        RECT 582.750 867.750 584.550 879.600 ;
        RECT 602.400 873.600 603.600 886.050 ;
        RECT 613.950 884.850 616.050 886.950 ;
        RECT 616.950 886.050 619.050 888.150 ;
        RECT 620.850 886.950 622.050 890.250 ;
        RECT 641.100 888.150 642.900 889.950 ;
        RECT 619.950 884.850 622.050 886.950 ;
        RECT 637.950 884.850 640.050 886.950 ;
        RECT 640.950 886.050 643.050 888.150 ;
        RECT 644.850 886.950 646.050 890.250 ;
        RECT 643.950 884.850 646.050 886.950 ;
        RECT 661.950 884.850 664.050 886.950 ;
        RECT 614.100 883.050 615.900 884.850 ;
        RECT 619.950 879.600 621.150 884.850 ;
        RECT 622.950 881.850 625.050 883.950 ;
        RECT 638.100 883.050 639.900 884.850 ;
        RECT 622.950 880.050 624.750 881.850 ;
        RECT 643.950 879.600 645.150 884.850 ;
        RECT 646.950 881.850 649.050 883.950 ;
        RECT 662.100 883.050 663.900 884.850 ;
        RECT 666.000 882.300 667.050 890.700 ;
        RECT 669.150 886.950 670.350 893.400 ;
        RECT 667.950 884.850 670.350 886.950 ;
        RECT 646.950 880.050 648.750 881.850 ;
        RECT 666.000 881.400 668.250 882.300 ;
        RECT 662.550 880.500 668.250 881.400 ;
        RECT 599.550 867.750 601.350 873.600 ;
        RECT 602.550 867.750 604.350 873.600 ;
        RECT 615.300 867.750 617.100 879.600 ;
        RECT 619.500 867.750 621.300 879.600 ;
        RECT 622.800 867.750 624.600 873.600 ;
        RECT 639.300 867.750 641.100 879.600 ;
        RECT 643.500 867.750 645.300 879.600 ;
        RECT 662.550 873.600 663.750 880.500 ;
        RECT 669.150 879.600 670.350 884.850 ;
        RECT 675.150 880.800 676.050 893.400 ;
        RECT 683.550 892.800 685.350 894.600 ;
        RECT 686.850 893.550 691.800 894.600 ;
        RECT 699.300 895.500 700.350 896.400 ;
        RECT 699.300 894.300 703.050 895.500 ;
        RECT 686.850 892.800 688.650 893.550 ;
        RECT 683.850 891.900 684.900 892.800 ;
        RECT 694.050 892.200 695.850 894.000 ;
        RECT 700.950 893.400 703.050 894.300 ;
        RECT 706.650 893.400 708.450 899.250 ;
        RECT 716.850 893.400 718.650 899.250 ;
        RECT 694.050 891.900 694.950 892.200 ;
        RECT 683.850 891.000 694.950 891.900 ;
        RECT 707.250 891.150 708.450 893.400 ;
        RECT 721.350 892.200 723.150 899.250 ;
        RECT 683.850 889.800 684.900 891.000 ;
        RECT 678.000 888.600 684.900 889.800 ;
        RECT 678.000 887.850 678.900 888.600 ;
        RECT 683.100 888.000 684.900 888.600 ;
        RECT 677.100 886.050 678.900 887.850 ;
        RECT 680.100 886.950 681.900 887.700 ;
        RECT 694.050 886.950 694.950 891.000 ;
        RECT 703.950 889.050 708.450 891.150 ;
        RECT 702.150 887.250 706.050 889.050 ;
        RECT 703.950 886.950 706.050 887.250 ;
        RECT 680.100 885.900 688.050 886.950 ;
        RECT 685.950 884.850 688.050 885.900 ;
        RECT 691.950 884.850 694.950 886.950 ;
        RECT 684.450 881.100 686.250 881.400 ;
        RECT 684.450 880.800 692.850 881.100 ;
        RECT 675.150 880.200 692.850 880.800 ;
        RECT 675.150 879.600 686.250 880.200 ;
        RECT 646.800 867.750 648.600 873.600 ;
        RECT 662.550 867.750 664.350 873.600 ;
        RECT 665.850 867.750 667.650 879.600 ;
        RECT 668.850 867.750 670.650 879.600 ;
        RECT 675.150 867.750 676.950 879.600 ;
        RECT 689.250 878.700 691.050 879.300 ;
        RECT 683.550 877.500 691.050 878.700 ;
        RECT 691.950 878.100 692.850 880.200 ;
        RECT 694.050 880.200 694.950 884.850 ;
        RECT 704.250 881.400 706.050 883.200 ;
        RECT 700.950 880.200 705.150 881.400 ;
        RECT 694.050 879.300 700.050 880.200 ;
        RECT 700.950 879.300 703.050 880.200 ;
        RECT 707.250 879.600 708.450 889.050 ;
        RECT 719.550 891.300 723.150 892.200 ;
        RECT 737.850 892.200 739.650 899.250 ;
        RECT 742.350 893.400 744.150 899.250 ;
        RECT 757.350 893.400 759.150 899.250 ;
        RECT 760.350 893.400 762.150 899.250 ;
        RECT 763.650 896.400 765.450 899.250 ;
        RECT 737.850 891.300 741.450 892.200 ;
        RECT 716.100 885.150 717.900 886.950 ;
        RECT 715.950 883.050 718.050 885.150 ;
        RECT 719.550 883.950 720.750 891.300 ;
        RECT 722.100 885.150 723.900 886.950 ;
        RECT 737.100 885.150 738.900 886.950 ;
        RECT 718.950 881.850 721.050 883.950 ;
        RECT 721.950 883.050 724.050 885.150 ;
        RECT 736.950 883.050 739.050 885.150 ;
        RECT 740.250 883.950 741.450 891.300 ;
        RECT 757.650 886.950 758.850 893.400 ;
        RECT 763.650 892.500 764.850 896.400 ;
        RECT 759.750 891.600 764.850 892.500 ;
        RECT 767.550 893.400 769.350 899.250 ;
        RECT 770.850 896.400 772.650 899.250 ;
        RECT 775.350 896.400 777.150 899.250 ;
        RECT 779.550 896.400 781.350 899.250 ;
        RECT 783.450 896.400 785.250 899.250 ;
        RECT 786.750 896.400 788.550 899.250 ;
        RECT 791.250 897.300 793.050 899.250 ;
        RECT 791.250 896.400 795.000 897.300 ;
        RECT 796.050 896.400 797.850 899.250 ;
        RECT 775.650 895.500 776.700 896.400 ;
        RECT 772.950 894.300 776.700 895.500 ;
        RECT 784.200 894.600 785.250 896.400 ;
        RECT 793.950 895.500 795.000 896.400 ;
        RECT 772.950 893.400 775.050 894.300 ;
        RECT 759.750 890.700 762.000 891.600 ;
        RECT 743.100 885.150 744.900 886.950 ;
        RECT 739.950 881.850 742.050 883.950 ;
        RECT 742.950 883.050 745.050 885.150 ;
        RECT 757.650 884.850 760.050 886.950 ;
        RECT 699.150 878.400 700.050 879.300 ;
        RECT 696.450 878.100 698.250 878.400 ;
        RECT 683.550 876.600 684.750 877.500 ;
        RECT 691.950 877.200 698.250 878.100 ;
        RECT 696.450 876.600 698.250 877.200 ;
        RECT 699.150 876.600 701.850 878.400 ;
        RECT 679.950 874.500 684.750 876.600 ;
        RECT 687.150 874.500 694.050 876.300 ;
        RECT 683.550 873.600 684.750 874.500 ;
        RECT 678.150 867.750 679.950 873.600 ;
        RECT 683.250 867.750 685.050 873.600 ;
        RECT 688.050 867.750 689.850 873.600 ;
        RECT 691.050 867.750 692.850 874.500 ;
        RECT 699.150 873.600 703.050 875.700 ;
        RECT 694.950 867.750 696.750 873.600 ;
        RECT 699.150 867.750 700.950 873.600 ;
        RECT 703.650 867.750 705.450 870.600 ;
        RECT 706.650 867.750 708.450 879.600 ;
        RECT 719.550 873.600 720.750 881.850 ;
        RECT 740.250 873.600 741.450 881.850 ;
        RECT 757.650 879.600 758.850 884.850 ;
        RECT 760.950 882.300 762.000 890.700 ;
        RECT 767.550 891.150 768.750 893.400 ;
        RECT 780.150 892.200 781.950 894.000 ;
        RECT 784.200 893.550 789.150 894.600 ;
        RECT 787.350 892.800 789.150 893.550 ;
        RECT 790.650 892.800 792.450 894.600 ;
        RECT 793.950 893.400 796.050 895.500 ;
        RECT 799.050 893.400 800.850 899.250 ;
        RECT 811.350 893.400 813.150 899.250 ;
        RECT 814.350 893.400 816.150 899.250 ;
        RECT 817.650 896.400 819.450 899.250 ;
        RECT 832.650 896.400 834.450 899.250 ;
        RECT 835.650 896.400 837.450 899.250 ;
        RECT 781.050 891.900 781.950 892.200 ;
        RECT 791.100 891.900 792.150 892.800 ;
        RECT 767.550 889.050 772.050 891.150 ;
        RECT 781.050 891.000 792.150 891.900 ;
        RECT 763.950 884.850 766.050 886.950 ;
        RECT 764.100 883.050 765.900 884.850 ;
        RECT 759.750 881.400 762.000 882.300 ;
        RECT 759.750 880.500 765.450 881.400 ;
        RECT 716.550 867.750 718.350 873.600 ;
        RECT 719.550 867.750 721.350 873.600 ;
        RECT 722.550 867.750 724.350 873.600 ;
        RECT 736.650 867.750 738.450 873.600 ;
        RECT 739.650 867.750 741.450 873.600 ;
        RECT 742.650 867.750 744.450 873.600 ;
        RECT 757.350 867.750 759.150 879.600 ;
        RECT 760.350 867.750 762.150 879.600 ;
        RECT 764.250 873.600 765.450 880.500 ;
        RECT 763.650 867.750 765.450 873.600 ;
        RECT 767.550 879.600 768.750 889.050 ;
        RECT 769.950 887.250 773.850 889.050 ;
        RECT 769.950 886.950 772.050 887.250 ;
        RECT 781.050 886.950 781.950 891.000 ;
        RECT 791.100 889.800 792.150 891.000 ;
        RECT 791.100 888.600 798.000 889.800 ;
        RECT 791.100 888.000 792.900 888.600 ;
        RECT 797.100 887.850 798.000 888.600 ;
        RECT 794.100 886.950 795.900 887.700 ;
        RECT 781.050 884.850 784.050 886.950 ;
        RECT 787.950 885.900 795.900 886.950 ;
        RECT 797.100 886.050 798.900 887.850 ;
        RECT 787.950 884.850 790.050 885.900 ;
        RECT 769.950 881.400 771.750 883.200 ;
        RECT 770.850 880.200 775.050 881.400 ;
        RECT 781.050 880.200 781.950 884.850 ;
        RECT 789.750 881.100 791.550 881.400 ;
        RECT 767.550 867.750 769.350 879.600 ;
        RECT 772.950 879.300 775.050 880.200 ;
        RECT 775.950 879.300 781.950 880.200 ;
        RECT 783.150 880.800 791.550 881.100 ;
        RECT 799.950 880.800 800.850 893.400 ;
        RECT 783.150 880.200 800.850 880.800 ;
        RECT 775.950 878.400 776.850 879.300 ;
        RECT 774.150 876.600 776.850 878.400 ;
        RECT 777.750 878.100 779.550 878.400 ;
        RECT 783.150 878.100 784.050 880.200 ;
        RECT 789.750 879.600 800.850 880.200 ;
        RECT 811.650 886.950 812.850 893.400 ;
        RECT 817.650 892.500 818.850 896.400 ;
        RECT 813.750 891.600 818.850 892.500 ;
        RECT 813.750 890.700 816.000 891.600 ;
        RECT 811.650 884.850 814.050 886.950 ;
        RECT 811.650 879.600 812.850 884.850 ;
        RECT 814.950 882.300 816.000 890.700 ;
        RECT 833.400 888.150 834.600 896.400 ;
        RECT 845.850 893.400 847.650 899.250 ;
        RECT 850.350 892.200 852.150 899.250 ;
        RECT 863.550 896.400 865.350 899.250 ;
        RECT 848.550 891.300 852.150 892.200 ;
        RECT 864.150 892.500 865.350 896.400 ;
        RECT 866.850 893.400 868.650 899.250 ;
        RECT 869.850 893.400 871.650 899.250 ;
        RECT 864.150 891.600 869.250 892.500 ;
        RECT 817.950 884.850 820.050 886.950 ;
        RECT 832.950 886.050 835.050 888.150 ;
        RECT 835.950 887.850 838.050 889.950 ;
        RECT 836.100 886.050 837.900 887.850 ;
        RECT 818.100 883.050 819.900 884.850 ;
        RECT 813.750 881.400 816.000 882.300 ;
        RECT 813.750 880.500 819.450 881.400 ;
        RECT 777.750 877.200 784.050 878.100 ;
        RECT 784.950 878.700 786.750 879.300 ;
        RECT 784.950 877.500 792.450 878.700 ;
        RECT 777.750 876.600 779.550 877.200 ;
        RECT 791.250 876.600 792.450 877.500 ;
        RECT 772.950 873.600 776.850 875.700 ;
        RECT 781.950 874.500 788.850 876.300 ;
        RECT 791.250 874.500 796.050 876.600 ;
        RECT 770.550 867.750 772.350 870.600 ;
        RECT 775.050 867.750 776.850 873.600 ;
        RECT 779.250 867.750 781.050 873.600 ;
        RECT 783.150 867.750 784.950 874.500 ;
        RECT 791.250 873.600 792.450 874.500 ;
        RECT 786.150 867.750 787.950 873.600 ;
        RECT 790.950 867.750 792.750 873.600 ;
        RECT 796.050 867.750 797.850 873.600 ;
        RECT 799.050 867.750 800.850 879.600 ;
        RECT 811.350 867.750 813.150 879.600 ;
        RECT 814.350 867.750 816.150 879.600 ;
        RECT 818.250 873.600 819.450 880.500 ;
        RECT 833.400 873.600 834.600 886.050 ;
        RECT 845.100 885.150 846.900 886.950 ;
        RECT 844.950 883.050 847.050 885.150 ;
        RECT 848.550 883.950 849.750 891.300 ;
        RECT 867.000 890.700 869.250 891.600 ;
        RECT 851.100 885.150 852.900 886.950 ;
        RECT 847.950 881.850 850.050 883.950 ;
        RECT 850.950 883.050 853.050 885.150 ;
        RECT 862.950 884.850 865.050 886.950 ;
        RECT 863.100 883.050 864.900 884.850 ;
        RECT 867.000 882.300 868.050 890.700 ;
        RECT 870.150 886.950 871.350 893.400 ;
        RECT 868.950 884.850 871.350 886.950 ;
        RECT 848.550 873.600 849.750 881.850 ;
        RECT 867.000 881.400 869.250 882.300 ;
        RECT 863.550 880.500 869.250 881.400 ;
        RECT 863.550 873.600 864.750 880.500 ;
        RECT 870.150 879.600 871.350 884.850 ;
        RECT 817.650 867.750 819.450 873.600 ;
        RECT 832.650 867.750 834.450 873.600 ;
        RECT 835.650 867.750 837.450 873.600 ;
        RECT 845.550 867.750 847.350 873.600 ;
        RECT 848.550 867.750 850.350 873.600 ;
        RECT 851.550 867.750 853.350 873.600 ;
        RECT 863.550 867.750 865.350 873.600 ;
        RECT 866.850 867.750 868.650 879.600 ;
        RECT 869.850 867.750 871.650 879.600 ;
        RECT 13.650 857.400 15.450 863.250 ;
        RECT 16.650 857.400 18.450 863.250 ;
        RECT 14.400 844.950 15.600 857.400 ;
        RECT 26.550 853.500 28.350 863.250 ;
        RECT 29.550 854.400 31.350 863.250 ;
        RECT 32.550 862.500 40.350 863.250 ;
        RECT 32.550 853.500 34.350 862.500 ;
        RECT 26.550 852.600 34.350 853.500 ;
        RECT 35.550 853.800 37.350 861.600 ;
        RECT 38.550 854.700 40.350 862.500 ;
        RECT 42.150 862.500 49.950 863.250 ;
        RECT 42.150 853.800 43.950 862.500 ;
        RECT 35.550 852.900 43.950 853.800 ;
        RECT 45.150 853.800 46.950 861.600 ;
        RECT 45.150 851.400 46.350 853.800 ;
        RECT 48.150 853.200 49.950 862.500 ;
        RECT 60.300 851.400 62.100 863.250 ;
        RECT 64.500 851.400 66.300 863.250 ;
        RECT 67.800 857.400 69.600 863.250 ;
        RECT 80.550 857.400 82.350 863.250 ;
        RECT 83.550 857.400 85.350 863.250 ;
        RECT 98.550 857.400 100.350 863.250 ;
        RECT 101.550 857.400 103.350 863.250 ;
        RECT 104.550 857.400 106.350 863.250 ;
        RECT 118.650 857.400 120.450 863.250 ;
        RECT 121.650 857.400 123.450 863.250 ;
        RECT 124.650 857.400 126.450 863.250 ;
        RECT 42.900 850.200 46.350 851.400 ;
        RECT 29.100 846.150 30.900 847.950 ;
        RECT 38.100 846.150 39.900 847.950 ;
        RECT 13.950 842.850 16.050 844.950 ;
        RECT 17.100 843.150 18.900 844.950 ;
        RECT 28.950 844.050 31.050 846.150 ;
        RECT 14.400 834.600 15.600 842.850 ;
        RECT 16.950 841.050 19.050 843.150 ;
        RECT 34.950 842.850 37.050 844.950 ;
        RECT 37.950 844.050 40.050 846.150 ;
        RECT 42.900 844.950 44.100 850.200 ;
        RECT 59.100 846.150 60.900 847.950 ;
        RECT 64.950 846.150 66.150 851.400 ;
        RECT 67.950 849.150 69.750 850.950 ;
        RECT 67.950 847.050 70.050 849.150 ;
        RECT 42.900 842.850 46.050 844.950 ;
        RECT 58.950 844.050 61.050 846.150 ;
        RECT 61.950 842.850 64.050 844.950 ;
        RECT 64.950 844.050 67.050 846.150 ;
        RECT 83.400 844.950 84.600 857.400 ;
        RECT 101.550 849.150 102.750 857.400 ;
        RECT 122.250 849.150 123.450 857.400 ;
        RECT 129.150 851.400 130.950 863.250 ;
        RECT 132.150 857.400 133.950 863.250 ;
        RECT 137.250 857.400 139.050 863.250 ;
        RECT 142.050 857.400 143.850 863.250 ;
        RECT 137.550 856.500 138.750 857.400 ;
        RECT 145.050 856.500 146.850 863.250 ;
        RECT 148.950 857.400 150.750 863.250 ;
        RECT 153.150 857.400 154.950 863.250 ;
        RECT 157.650 860.400 159.450 863.250 ;
        RECT 133.950 854.400 138.750 856.500 ;
        RECT 141.150 854.700 148.050 856.500 ;
        RECT 153.150 855.300 157.050 857.400 ;
        RECT 137.550 853.500 138.750 854.400 ;
        RECT 150.450 853.800 152.250 854.400 ;
        RECT 137.550 852.300 145.050 853.500 ;
        RECT 143.250 851.700 145.050 852.300 ;
        RECT 145.950 852.900 152.250 853.800 ;
        RECT 129.150 850.800 140.250 851.400 ;
        RECT 145.950 850.800 146.850 852.900 ;
        RECT 150.450 852.600 152.250 852.900 ;
        RECT 153.150 852.600 155.850 854.400 ;
        RECT 153.150 851.700 154.050 852.600 ;
        RECT 129.150 850.200 146.850 850.800 ;
        RECT 97.950 845.850 100.050 847.950 ;
        RECT 100.950 847.050 103.050 849.150 ;
        RECT 35.100 841.050 36.900 842.850 ;
        RECT 42.900 836.400 44.100 842.850 ;
        RECT 62.100 841.050 63.900 842.850 ;
        RECT 65.850 840.750 67.050 844.050 ;
        RECT 80.100 843.150 81.900 844.950 ;
        RECT 79.950 841.050 82.050 843.150 ;
        RECT 82.950 842.850 85.050 844.950 ;
        RECT 98.100 844.050 99.900 845.850 ;
        RECT 66.000 839.700 69.750 840.750 ;
        RECT 33.300 835.500 44.100 836.400 ;
        RECT 59.550 836.700 67.350 838.050 ;
        RECT 33.300 834.600 34.350 835.500 ;
        RECT 39.300 834.600 40.350 835.500 ;
        RECT 13.650 831.750 15.450 834.600 ;
        RECT 16.650 831.750 18.450 834.600 ;
        RECT 29.250 831.750 31.350 834.600 ;
        RECT 32.550 831.750 34.350 834.600 ;
        RECT 35.550 831.750 37.350 834.600 ;
        RECT 38.550 831.750 40.350 834.600 ;
        RECT 59.550 831.750 61.350 836.700 ;
        RECT 62.550 831.750 64.350 835.800 ;
        RECT 65.550 831.750 67.350 836.700 ;
        RECT 68.550 837.600 69.750 839.700 ;
        RECT 68.550 831.750 70.350 837.600 ;
        RECT 83.400 834.600 84.600 842.850 ;
        RECT 101.550 839.700 102.750 847.050 ;
        RECT 103.950 845.850 106.050 847.950 ;
        RECT 118.950 845.850 121.050 847.950 ;
        RECT 121.950 847.050 124.050 849.150 ;
        RECT 104.100 844.050 105.900 845.850 ;
        RECT 119.100 844.050 120.900 845.850 ;
        RECT 122.250 839.700 123.450 847.050 ;
        RECT 124.950 845.850 127.050 847.950 ;
        RECT 125.100 844.050 126.900 845.850 ;
        RECT 101.550 838.800 105.150 839.700 ;
        RECT 80.550 831.750 82.350 834.600 ;
        RECT 83.550 831.750 85.350 834.600 ;
        RECT 98.850 831.750 100.650 837.600 ;
        RECT 103.350 831.750 105.150 838.800 ;
        RECT 119.850 838.800 123.450 839.700 ;
        RECT 119.850 831.750 121.650 838.800 ;
        RECT 129.150 837.600 130.050 850.200 ;
        RECT 138.450 849.900 146.850 850.200 ;
        RECT 148.050 850.800 154.050 851.700 ;
        RECT 154.950 850.800 157.050 851.700 ;
        RECT 160.650 851.400 162.450 863.250 ;
        RECT 173.400 857.400 175.200 863.250 ;
        RECT 176.700 851.400 178.500 863.250 ;
        RECT 180.900 851.400 182.700 863.250 ;
        RECT 186.150 851.400 187.950 863.250 ;
        RECT 189.150 857.400 190.950 863.250 ;
        RECT 194.250 857.400 196.050 863.250 ;
        RECT 199.050 857.400 200.850 863.250 ;
        RECT 194.550 856.500 195.750 857.400 ;
        RECT 202.050 856.500 203.850 863.250 ;
        RECT 205.950 857.400 207.750 863.250 ;
        RECT 210.150 857.400 211.950 863.250 ;
        RECT 214.650 860.400 216.450 863.250 ;
        RECT 190.950 854.400 195.750 856.500 ;
        RECT 198.150 854.700 205.050 856.500 ;
        RECT 210.150 855.300 214.050 857.400 ;
        RECT 194.550 853.500 195.750 854.400 ;
        RECT 207.450 853.800 209.250 854.400 ;
        RECT 194.550 852.300 202.050 853.500 ;
        RECT 200.250 851.700 202.050 852.300 ;
        RECT 202.950 852.900 209.250 853.800 ;
        RECT 138.450 849.600 140.250 849.900 ;
        RECT 148.050 846.150 148.950 850.800 ;
        RECT 154.950 849.600 159.150 850.800 ;
        RECT 158.250 847.800 160.050 849.600 ;
        RECT 139.950 845.100 142.050 846.150 ;
        RECT 131.100 843.150 132.900 844.950 ;
        RECT 134.100 844.050 142.050 845.100 ;
        RECT 145.950 844.050 148.950 846.150 ;
        RECT 134.100 843.300 135.900 844.050 ;
        RECT 132.000 842.400 132.900 843.150 ;
        RECT 137.100 842.400 138.900 843.000 ;
        RECT 132.000 841.200 138.900 842.400 ;
        RECT 137.850 840.000 138.900 841.200 ;
        RECT 148.050 840.000 148.950 844.050 ;
        RECT 157.950 843.750 160.050 844.050 ;
        RECT 156.150 841.950 160.050 843.750 ;
        RECT 161.250 841.950 162.450 851.400 ;
        RECT 173.250 849.150 175.050 850.950 ;
        RECT 172.950 847.050 175.050 849.150 ;
        RECT 176.850 846.150 178.050 851.400 ;
        RECT 186.150 850.800 197.250 851.400 ;
        RECT 202.950 850.800 203.850 852.900 ;
        RECT 207.450 852.600 209.250 852.900 ;
        RECT 210.150 852.600 212.850 854.400 ;
        RECT 210.150 851.700 211.050 852.600 ;
        RECT 186.150 850.200 203.850 850.800 ;
        RECT 182.100 846.150 183.900 847.950 ;
        RECT 137.850 839.100 148.950 840.000 ;
        RECT 157.950 839.850 162.450 841.950 ;
        RECT 175.950 844.050 178.050 846.150 ;
        RECT 175.950 840.750 177.150 844.050 ;
        RECT 178.950 842.850 181.050 844.950 ;
        RECT 181.950 844.050 184.050 846.150 ;
        RECT 179.100 841.050 180.900 842.850 ;
        RECT 137.850 838.200 138.900 839.100 ;
        RECT 148.050 838.800 148.950 839.100 ;
        RECT 124.350 831.750 126.150 837.600 ;
        RECT 129.150 831.750 130.950 837.600 ;
        RECT 133.950 835.500 136.050 837.600 ;
        RECT 137.550 836.400 139.350 838.200 ;
        RECT 140.850 837.450 142.650 838.200 ;
        RECT 140.850 836.400 145.800 837.450 ;
        RECT 148.050 837.000 149.850 838.800 ;
        RECT 161.250 837.600 162.450 839.850 ;
        RECT 173.250 839.700 177.000 840.750 ;
        RECT 173.250 837.600 174.450 839.700 ;
        RECT 154.950 836.700 157.050 837.600 ;
        RECT 135.000 834.600 136.050 835.500 ;
        RECT 144.750 834.600 145.800 836.400 ;
        RECT 153.300 835.500 157.050 836.700 ;
        RECT 153.300 834.600 154.350 835.500 ;
        RECT 132.150 831.750 133.950 834.600 ;
        RECT 135.000 833.700 138.750 834.600 ;
        RECT 136.950 831.750 138.750 833.700 ;
        RECT 141.450 831.750 143.250 834.600 ;
        RECT 144.750 831.750 146.550 834.600 ;
        RECT 148.650 831.750 150.450 834.600 ;
        RECT 152.850 831.750 154.650 834.600 ;
        RECT 157.350 831.750 159.150 834.600 ;
        RECT 160.650 831.750 162.450 837.600 ;
        RECT 172.650 831.750 174.450 837.600 ;
        RECT 175.650 836.700 183.450 838.050 ;
        RECT 175.650 831.750 177.450 836.700 ;
        RECT 178.650 831.750 180.450 835.800 ;
        RECT 181.650 831.750 183.450 836.700 ;
        RECT 186.150 837.600 187.050 850.200 ;
        RECT 195.450 849.900 203.850 850.200 ;
        RECT 205.050 850.800 211.050 851.700 ;
        RECT 211.950 850.800 214.050 851.700 ;
        RECT 217.650 851.400 219.450 863.250 ;
        RECT 229.650 862.500 237.450 863.250 ;
        RECT 229.650 851.400 231.450 862.500 ;
        RECT 232.650 851.400 234.450 861.600 ;
        RECT 235.650 852.600 237.450 862.500 ;
        RECT 238.650 853.500 240.450 863.250 ;
        RECT 241.650 852.600 243.450 863.250 ;
        RECT 235.650 851.700 243.450 852.600 ;
        RECT 246.150 851.400 247.950 863.250 ;
        RECT 249.150 857.400 250.950 863.250 ;
        RECT 254.250 857.400 256.050 863.250 ;
        RECT 259.050 857.400 260.850 863.250 ;
        RECT 254.550 856.500 255.750 857.400 ;
        RECT 262.050 856.500 263.850 863.250 ;
        RECT 265.950 857.400 267.750 863.250 ;
        RECT 270.150 857.400 271.950 863.250 ;
        RECT 274.650 860.400 276.450 863.250 ;
        RECT 250.950 854.400 255.750 856.500 ;
        RECT 258.150 854.700 265.050 856.500 ;
        RECT 270.150 855.300 274.050 857.400 ;
        RECT 254.550 853.500 255.750 854.400 ;
        RECT 267.450 853.800 269.250 854.400 ;
        RECT 254.550 852.300 262.050 853.500 ;
        RECT 260.250 851.700 262.050 852.300 ;
        RECT 262.950 852.900 269.250 853.800 ;
        RECT 195.450 849.600 197.250 849.900 ;
        RECT 205.050 846.150 205.950 850.800 ;
        RECT 211.950 849.600 216.150 850.800 ;
        RECT 215.250 847.800 217.050 849.600 ;
        RECT 196.950 845.100 199.050 846.150 ;
        RECT 188.100 843.150 189.900 844.950 ;
        RECT 191.100 844.050 199.050 845.100 ;
        RECT 202.950 844.050 205.950 846.150 ;
        RECT 191.100 843.300 192.900 844.050 ;
        RECT 189.000 842.400 189.900 843.150 ;
        RECT 194.100 842.400 195.900 843.000 ;
        RECT 189.000 841.200 195.900 842.400 ;
        RECT 194.850 840.000 195.900 841.200 ;
        RECT 205.050 840.000 205.950 844.050 ;
        RECT 214.950 843.750 217.050 844.050 ;
        RECT 213.150 841.950 217.050 843.750 ;
        RECT 218.250 841.950 219.450 851.400 ;
        RECT 232.800 850.500 234.600 851.400 ;
        RECT 246.150 850.800 257.250 851.400 ;
        RECT 262.950 850.800 263.850 852.900 ;
        RECT 267.450 852.600 269.250 852.900 ;
        RECT 270.150 852.600 272.850 854.400 ;
        RECT 270.150 851.700 271.050 852.600 ;
        RECT 232.800 849.600 236.850 850.500 ;
        RECT 230.100 846.150 231.900 847.950 ;
        RECT 235.950 846.150 236.850 849.600 ;
        RECT 246.150 850.200 263.850 850.800 ;
        RECT 241.950 846.150 243.750 847.950 ;
        RECT 229.950 844.050 232.050 846.150 ;
        RECT 232.950 842.850 235.050 844.950 ;
        RECT 235.950 844.050 238.050 846.150 ;
        RECT 194.850 839.100 205.950 840.000 ;
        RECT 214.950 839.850 219.450 841.950 ;
        RECT 233.250 841.050 235.050 842.850 ;
        RECT 194.850 838.200 195.900 839.100 ;
        RECT 205.050 838.800 205.950 839.100 ;
        RECT 186.150 831.750 187.950 837.600 ;
        RECT 190.950 835.500 193.050 837.600 ;
        RECT 194.550 836.400 196.350 838.200 ;
        RECT 197.850 837.450 199.650 838.200 ;
        RECT 197.850 836.400 202.800 837.450 ;
        RECT 205.050 837.000 206.850 838.800 ;
        RECT 218.250 837.600 219.450 839.850 ;
        RECT 237.000 837.600 238.050 844.050 ;
        RECT 238.950 842.850 241.050 844.950 ;
        RECT 241.950 844.050 244.050 846.150 ;
        RECT 238.950 841.050 240.750 842.850 ;
        RECT 246.150 837.600 247.050 850.200 ;
        RECT 255.450 849.900 263.850 850.200 ;
        RECT 265.050 850.800 271.050 851.700 ;
        RECT 271.950 850.800 274.050 851.700 ;
        RECT 277.650 851.400 279.450 863.250 ;
        RECT 288.300 851.400 290.100 863.250 ;
        RECT 292.500 851.400 294.300 863.250 ;
        RECT 295.800 857.400 297.600 863.250 ;
        RECT 303.150 851.400 304.950 863.250 ;
        RECT 306.150 857.400 307.950 863.250 ;
        RECT 311.250 857.400 313.050 863.250 ;
        RECT 316.050 857.400 317.850 863.250 ;
        RECT 311.550 856.500 312.750 857.400 ;
        RECT 319.050 856.500 320.850 863.250 ;
        RECT 322.950 857.400 324.750 863.250 ;
        RECT 327.150 857.400 328.950 863.250 ;
        RECT 331.650 860.400 333.450 863.250 ;
        RECT 307.950 854.400 312.750 856.500 ;
        RECT 315.150 854.700 322.050 856.500 ;
        RECT 327.150 855.300 331.050 857.400 ;
        RECT 311.550 853.500 312.750 854.400 ;
        RECT 324.450 853.800 326.250 854.400 ;
        RECT 311.550 852.300 319.050 853.500 ;
        RECT 317.250 851.700 319.050 852.300 ;
        RECT 319.950 852.900 326.250 853.800 ;
        RECT 255.450 849.600 257.250 849.900 ;
        RECT 265.050 846.150 265.950 850.800 ;
        RECT 271.950 849.600 276.150 850.800 ;
        RECT 275.250 847.800 277.050 849.600 ;
        RECT 256.950 845.100 259.050 846.150 ;
        RECT 248.100 843.150 249.900 844.950 ;
        RECT 251.100 844.050 259.050 845.100 ;
        RECT 262.950 844.050 265.950 846.150 ;
        RECT 251.100 843.300 252.900 844.050 ;
        RECT 249.000 842.400 249.900 843.150 ;
        RECT 254.100 842.400 255.900 843.000 ;
        RECT 249.000 841.200 255.900 842.400 ;
        RECT 254.850 840.000 255.900 841.200 ;
        RECT 265.050 840.000 265.950 844.050 ;
        RECT 274.950 843.750 277.050 844.050 ;
        RECT 273.150 841.950 277.050 843.750 ;
        RECT 278.250 841.950 279.450 851.400 ;
        RECT 287.100 846.150 288.900 847.950 ;
        RECT 292.950 846.150 294.150 851.400 ;
        RECT 295.950 849.150 297.750 850.950 ;
        RECT 303.150 850.800 314.250 851.400 ;
        RECT 319.950 850.800 320.850 852.900 ;
        RECT 324.450 852.600 326.250 852.900 ;
        RECT 327.150 852.600 329.850 854.400 ;
        RECT 327.150 851.700 328.050 852.600 ;
        RECT 303.150 850.200 320.850 850.800 ;
        RECT 295.950 847.050 298.050 849.150 ;
        RECT 286.950 844.050 289.050 846.150 ;
        RECT 289.950 842.850 292.050 844.950 ;
        RECT 292.950 844.050 295.050 846.150 ;
        RECT 254.850 839.100 265.950 840.000 ;
        RECT 274.950 839.850 279.450 841.950 ;
        RECT 290.100 841.050 291.900 842.850 ;
        RECT 293.850 840.750 295.050 844.050 ;
        RECT 254.850 838.200 255.900 839.100 ;
        RECT 265.050 838.800 265.950 839.100 ;
        RECT 211.950 836.700 214.050 837.600 ;
        RECT 192.000 834.600 193.050 835.500 ;
        RECT 201.750 834.600 202.800 836.400 ;
        RECT 210.300 835.500 214.050 836.700 ;
        RECT 210.300 834.600 211.350 835.500 ;
        RECT 189.150 831.750 190.950 834.600 ;
        RECT 192.000 833.700 195.750 834.600 ;
        RECT 193.950 831.750 195.750 833.700 ;
        RECT 198.450 831.750 200.250 834.600 ;
        RECT 201.750 831.750 203.550 834.600 ;
        RECT 205.650 831.750 207.450 834.600 ;
        RECT 209.850 831.750 211.650 834.600 ;
        RECT 214.350 831.750 216.150 834.600 ;
        RECT 217.650 831.750 219.450 837.600 ;
        RECT 232.800 831.750 234.600 837.600 ;
        RECT 237.000 831.750 238.800 837.600 ;
        RECT 241.200 831.750 243.000 837.600 ;
        RECT 246.150 831.750 247.950 837.600 ;
        RECT 250.950 835.500 253.050 837.600 ;
        RECT 254.550 836.400 256.350 838.200 ;
        RECT 257.850 837.450 259.650 838.200 ;
        RECT 257.850 836.400 262.800 837.450 ;
        RECT 265.050 837.000 266.850 838.800 ;
        RECT 278.250 837.600 279.450 839.850 ;
        RECT 294.000 839.700 297.750 840.750 ;
        RECT 271.950 836.700 274.050 837.600 ;
        RECT 252.000 834.600 253.050 835.500 ;
        RECT 261.750 834.600 262.800 836.400 ;
        RECT 270.300 835.500 274.050 836.700 ;
        RECT 270.300 834.600 271.350 835.500 ;
        RECT 249.150 831.750 250.950 834.600 ;
        RECT 252.000 833.700 255.750 834.600 ;
        RECT 253.950 831.750 255.750 833.700 ;
        RECT 258.450 831.750 260.250 834.600 ;
        RECT 261.750 831.750 263.550 834.600 ;
        RECT 265.650 831.750 267.450 834.600 ;
        RECT 269.850 831.750 271.650 834.600 ;
        RECT 274.350 831.750 276.150 834.600 ;
        RECT 277.650 831.750 279.450 837.600 ;
        RECT 287.550 836.700 295.350 838.050 ;
        RECT 287.550 831.750 289.350 836.700 ;
        RECT 290.550 831.750 292.350 835.800 ;
        RECT 293.550 831.750 295.350 836.700 ;
        RECT 296.550 837.600 297.750 839.700 ;
        RECT 303.150 837.600 304.050 850.200 ;
        RECT 312.450 849.900 320.850 850.200 ;
        RECT 322.050 850.800 328.050 851.700 ;
        RECT 328.950 850.800 331.050 851.700 ;
        RECT 334.650 851.400 336.450 863.250 ;
        RECT 349.650 862.500 357.450 863.250 ;
        RECT 349.650 851.400 351.450 862.500 ;
        RECT 352.650 851.400 354.450 861.600 ;
        RECT 355.650 852.600 357.450 862.500 ;
        RECT 358.650 853.500 360.450 863.250 ;
        RECT 361.650 852.600 363.450 863.250 ;
        RECT 371.550 857.400 373.350 863.250 ;
        RECT 374.550 857.400 376.350 863.250 ;
        RECT 377.550 857.400 379.350 863.250 ;
        RECT 355.650 851.700 363.450 852.600 ;
        RECT 312.450 849.600 314.250 849.900 ;
        RECT 322.050 846.150 322.950 850.800 ;
        RECT 328.950 849.600 333.150 850.800 ;
        RECT 332.250 847.800 334.050 849.600 ;
        RECT 313.950 845.100 316.050 846.150 ;
        RECT 305.100 843.150 306.900 844.950 ;
        RECT 308.100 844.050 316.050 845.100 ;
        RECT 319.950 844.050 322.950 846.150 ;
        RECT 308.100 843.300 309.900 844.050 ;
        RECT 306.000 842.400 306.900 843.150 ;
        RECT 311.100 842.400 312.900 843.000 ;
        RECT 306.000 841.200 312.900 842.400 ;
        RECT 311.850 840.000 312.900 841.200 ;
        RECT 322.050 840.000 322.950 844.050 ;
        RECT 331.950 843.750 334.050 844.050 ;
        RECT 330.150 841.950 334.050 843.750 ;
        RECT 335.250 841.950 336.450 851.400 ;
        RECT 352.800 850.500 354.600 851.400 ;
        RECT 352.800 849.600 356.850 850.500 ;
        RECT 350.100 846.150 351.900 847.950 ;
        RECT 355.950 846.150 356.850 849.600 ;
        RECT 374.550 849.150 375.750 857.400 ;
        RECT 384.150 851.400 385.950 863.250 ;
        RECT 387.150 857.400 388.950 863.250 ;
        RECT 392.250 857.400 394.050 863.250 ;
        RECT 397.050 857.400 398.850 863.250 ;
        RECT 392.550 856.500 393.750 857.400 ;
        RECT 400.050 856.500 401.850 863.250 ;
        RECT 403.950 857.400 405.750 863.250 ;
        RECT 408.150 857.400 409.950 863.250 ;
        RECT 412.650 860.400 414.450 863.250 ;
        RECT 388.950 854.400 393.750 856.500 ;
        RECT 396.150 854.700 403.050 856.500 ;
        RECT 408.150 855.300 412.050 857.400 ;
        RECT 392.550 853.500 393.750 854.400 ;
        RECT 405.450 853.800 407.250 854.400 ;
        RECT 392.550 852.300 400.050 853.500 ;
        RECT 398.250 851.700 400.050 852.300 ;
        RECT 400.950 852.900 407.250 853.800 ;
        RECT 384.150 850.800 395.250 851.400 ;
        RECT 400.950 850.800 401.850 852.900 ;
        RECT 405.450 852.600 407.250 852.900 ;
        RECT 408.150 852.600 410.850 854.400 ;
        RECT 408.150 851.700 409.050 852.600 ;
        RECT 384.150 850.200 401.850 850.800 ;
        RECT 361.950 846.150 363.750 847.950 ;
        RECT 349.950 844.050 352.050 846.150 ;
        RECT 352.950 842.850 355.050 844.950 ;
        RECT 355.950 844.050 358.050 846.150 ;
        RECT 311.850 839.100 322.950 840.000 ;
        RECT 331.950 839.850 336.450 841.950 ;
        RECT 353.250 841.050 355.050 842.850 ;
        RECT 311.850 838.200 312.900 839.100 ;
        RECT 322.050 838.800 322.950 839.100 ;
        RECT 296.550 831.750 298.350 837.600 ;
        RECT 303.150 831.750 304.950 837.600 ;
        RECT 307.950 835.500 310.050 837.600 ;
        RECT 311.550 836.400 313.350 838.200 ;
        RECT 314.850 837.450 316.650 838.200 ;
        RECT 314.850 836.400 319.800 837.450 ;
        RECT 322.050 837.000 323.850 838.800 ;
        RECT 335.250 837.600 336.450 839.850 ;
        RECT 357.000 837.600 358.050 844.050 ;
        RECT 358.950 842.850 361.050 844.950 ;
        RECT 361.950 844.050 364.050 846.150 ;
        RECT 370.950 845.850 373.050 847.950 ;
        RECT 373.950 847.050 376.050 849.150 ;
        RECT 371.100 844.050 372.900 845.850 ;
        RECT 358.950 841.050 360.750 842.850 ;
        RECT 374.550 839.700 375.750 847.050 ;
        RECT 376.950 845.850 379.050 847.950 ;
        RECT 377.100 844.050 378.900 845.850 ;
        RECT 374.550 838.800 378.150 839.700 ;
        RECT 328.950 836.700 331.050 837.600 ;
        RECT 309.000 834.600 310.050 835.500 ;
        RECT 318.750 834.600 319.800 836.400 ;
        RECT 327.300 835.500 331.050 836.700 ;
        RECT 327.300 834.600 328.350 835.500 ;
        RECT 306.150 831.750 307.950 834.600 ;
        RECT 309.000 833.700 312.750 834.600 ;
        RECT 310.950 831.750 312.750 833.700 ;
        RECT 315.450 831.750 317.250 834.600 ;
        RECT 318.750 831.750 320.550 834.600 ;
        RECT 322.650 831.750 324.450 834.600 ;
        RECT 326.850 831.750 328.650 834.600 ;
        RECT 331.350 831.750 333.150 834.600 ;
        RECT 334.650 831.750 336.450 837.600 ;
        RECT 352.800 831.750 354.600 837.600 ;
        RECT 357.000 831.750 358.800 837.600 ;
        RECT 361.200 831.750 363.000 837.600 ;
        RECT 371.850 831.750 373.650 837.600 ;
        RECT 376.350 831.750 378.150 838.800 ;
        RECT 384.150 837.600 385.050 850.200 ;
        RECT 393.450 849.900 401.850 850.200 ;
        RECT 403.050 850.800 409.050 851.700 ;
        RECT 409.950 850.800 412.050 851.700 ;
        RECT 415.650 851.400 417.450 863.250 ;
        RECT 425.550 857.400 427.350 863.250 ;
        RECT 428.550 857.400 430.350 863.250 ;
        RECT 393.450 849.600 395.250 849.900 ;
        RECT 403.050 846.150 403.950 850.800 ;
        RECT 409.950 849.600 414.150 850.800 ;
        RECT 413.250 847.800 415.050 849.600 ;
        RECT 394.950 845.100 397.050 846.150 ;
        RECT 386.100 843.150 387.900 844.950 ;
        RECT 389.100 844.050 397.050 845.100 ;
        RECT 400.950 844.050 403.950 846.150 ;
        RECT 389.100 843.300 390.900 844.050 ;
        RECT 387.000 842.400 387.900 843.150 ;
        RECT 392.100 842.400 393.900 843.000 ;
        RECT 387.000 841.200 393.900 842.400 ;
        RECT 392.850 840.000 393.900 841.200 ;
        RECT 403.050 840.000 403.950 844.050 ;
        RECT 412.950 843.750 415.050 844.050 ;
        RECT 411.150 841.950 415.050 843.750 ;
        RECT 416.250 841.950 417.450 851.400 ;
        RECT 428.400 844.950 429.600 857.400 ;
        RECT 435.150 851.400 436.950 863.250 ;
        RECT 438.150 857.400 439.950 863.250 ;
        RECT 443.250 857.400 445.050 863.250 ;
        RECT 448.050 857.400 449.850 863.250 ;
        RECT 443.550 856.500 444.750 857.400 ;
        RECT 451.050 856.500 452.850 863.250 ;
        RECT 454.950 857.400 456.750 863.250 ;
        RECT 459.150 857.400 460.950 863.250 ;
        RECT 463.650 860.400 465.450 863.250 ;
        RECT 439.950 854.400 444.750 856.500 ;
        RECT 447.150 854.700 454.050 856.500 ;
        RECT 459.150 855.300 463.050 857.400 ;
        RECT 443.550 853.500 444.750 854.400 ;
        RECT 456.450 853.800 458.250 854.400 ;
        RECT 443.550 852.300 451.050 853.500 ;
        RECT 449.250 851.700 451.050 852.300 ;
        RECT 451.950 852.900 458.250 853.800 ;
        RECT 435.150 850.800 446.250 851.400 ;
        RECT 451.950 850.800 452.850 852.900 ;
        RECT 456.450 852.600 458.250 852.900 ;
        RECT 459.150 852.600 461.850 854.400 ;
        RECT 459.150 851.700 460.050 852.600 ;
        RECT 435.150 850.200 452.850 850.800 ;
        RECT 425.100 843.150 426.900 844.950 ;
        RECT 392.850 839.100 403.950 840.000 ;
        RECT 412.950 839.850 417.450 841.950 ;
        RECT 424.950 841.050 427.050 843.150 ;
        RECT 427.950 842.850 430.050 844.950 ;
        RECT 392.850 838.200 393.900 839.100 ;
        RECT 403.050 838.800 403.950 839.100 ;
        RECT 384.150 831.750 385.950 837.600 ;
        RECT 388.950 835.500 391.050 837.600 ;
        RECT 392.550 836.400 394.350 838.200 ;
        RECT 395.850 837.450 397.650 838.200 ;
        RECT 395.850 836.400 400.800 837.450 ;
        RECT 403.050 837.000 404.850 838.800 ;
        RECT 416.250 837.600 417.450 839.850 ;
        RECT 409.950 836.700 412.050 837.600 ;
        RECT 390.000 834.600 391.050 835.500 ;
        RECT 399.750 834.600 400.800 836.400 ;
        RECT 408.300 835.500 412.050 836.700 ;
        RECT 408.300 834.600 409.350 835.500 ;
        RECT 387.150 831.750 388.950 834.600 ;
        RECT 390.000 833.700 393.750 834.600 ;
        RECT 391.950 831.750 393.750 833.700 ;
        RECT 396.450 831.750 398.250 834.600 ;
        RECT 399.750 831.750 401.550 834.600 ;
        RECT 403.650 831.750 405.450 834.600 ;
        RECT 407.850 831.750 409.650 834.600 ;
        RECT 412.350 831.750 414.150 834.600 ;
        RECT 415.650 831.750 417.450 837.600 ;
        RECT 428.400 834.600 429.600 842.850 ;
        RECT 435.150 837.600 436.050 850.200 ;
        RECT 444.450 849.900 452.850 850.200 ;
        RECT 454.050 850.800 460.050 851.700 ;
        RECT 460.950 850.800 463.050 851.700 ;
        RECT 466.650 851.400 468.450 863.250 ;
        RECT 478.650 851.400 480.450 863.250 ;
        RECT 481.650 852.300 483.450 863.250 ;
        RECT 484.650 853.200 486.450 863.250 ;
        RECT 487.650 852.300 489.450 863.250 ;
        RECT 481.650 851.400 489.450 852.300 ;
        RECT 497.550 851.400 499.350 863.250 ;
        RECT 502.050 851.550 503.850 863.250 ;
        RECT 505.050 852.900 506.850 863.250 ;
        RECT 523.650 862.500 531.450 863.250 ;
        RECT 505.050 851.550 507.450 852.900 ;
        RECT 444.450 849.600 446.250 849.900 ;
        RECT 454.050 846.150 454.950 850.800 ;
        RECT 460.950 849.600 465.150 850.800 ;
        RECT 464.250 847.800 466.050 849.600 ;
        RECT 445.950 845.100 448.050 846.150 ;
        RECT 437.100 843.150 438.900 844.950 ;
        RECT 440.100 844.050 448.050 845.100 ;
        RECT 451.950 844.050 454.950 846.150 ;
        RECT 440.100 843.300 441.900 844.050 ;
        RECT 438.000 842.400 438.900 843.150 ;
        RECT 443.100 842.400 444.900 843.000 ;
        RECT 438.000 841.200 444.900 842.400 ;
        RECT 443.850 840.000 444.900 841.200 ;
        RECT 454.050 840.000 454.950 844.050 ;
        RECT 463.950 843.750 466.050 844.050 ;
        RECT 462.150 841.950 466.050 843.750 ;
        RECT 467.250 841.950 468.450 851.400 ;
        RECT 479.100 846.150 480.300 851.400 ;
        RECT 497.550 850.200 498.750 851.400 ;
        RECT 502.950 850.200 504.750 850.650 ;
        RECT 497.550 849.000 504.750 850.200 ;
        RECT 502.950 848.850 504.750 849.000 ;
        RECT 500.100 846.150 501.900 847.950 ;
        RECT 478.950 844.050 481.050 846.150 ;
        RECT 443.850 839.100 454.950 840.000 ;
        RECT 463.950 839.850 468.450 841.950 ;
        RECT 443.850 838.200 444.900 839.100 ;
        RECT 454.050 838.800 454.950 839.100 ;
        RECT 425.550 831.750 427.350 834.600 ;
        RECT 428.550 831.750 430.350 834.600 ;
        RECT 435.150 831.750 436.950 837.600 ;
        RECT 439.950 835.500 442.050 837.600 ;
        RECT 443.550 836.400 445.350 838.200 ;
        RECT 446.850 837.450 448.650 838.200 ;
        RECT 446.850 836.400 451.800 837.450 ;
        RECT 454.050 837.000 455.850 838.800 ;
        RECT 467.250 837.600 468.450 839.850 ;
        RECT 460.950 836.700 463.050 837.600 ;
        RECT 441.000 834.600 442.050 835.500 ;
        RECT 450.750 834.600 451.800 836.400 ;
        RECT 459.300 835.500 463.050 836.700 ;
        RECT 459.300 834.600 460.350 835.500 ;
        RECT 438.150 831.750 439.950 834.600 ;
        RECT 441.000 833.700 444.750 834.600 ;
        RECT 442.950 831.750 444.750 833.700 ;
        RECT 447.450 831.750 449.250 834.600 ;
        RECT 450.750 831.750 452.550 834.600 ;
        RECT 454.650 831.750 456.450 834.600 ;
        RECT 458.850 831.750 460.650 834.600 ;
        RECT 463.350 831.750 465.150 834.600 ;
        RECT 466.650 831.750 468.450 837.600 ;
        RECT 479.100 837.600 480.300 844.050 ;
        RECT 481.950 842.850 484.050 844.950 ;
        RECT 485.100 843.150 486.900 844.950 ;
        RECT 482.100 841.050 483.900 842.850 ;
        RECT 484.950 841.050 487.050 843.150 ;
        RECT 487.950 842.850 490.050 844.950 ;
        RECT 497.100 843.150 498.900 844.950 ;
        RECT 499.950 844.050 502.050 846.150 ;
        RECT 488.100 841.050 489.900 842.850 ;
        RECT 496.950 841.050 499.050 843.150 ;
        RECT 503.700 840.600 504.600 848.850 ;
        RECT 506.100 844.950 507.450 851.550 ;
        RECT 523.650 851.400 525.450 862.500 ;
        RECT 526.650 851.400 528.450 861.600 ;
        RECT 529.650 852.600 531.450 862.500 ;
        RECT 532.650 853.500 534.450 863.250 ;
        RECT 535.650 852.600 537.450 863.250 ;
        RECT 529.650 851.700 537.450 852.600 ;
        RECT 546.300 851.400 548.100 863.250 ;
        RECT 550.500 851.400 552.300 863.250 ;
        RECT 553.800 857.400 555.600 863.250 ;
        RECT 569.550 857.400 571.350 863.250 ;
        RECT 572.550 857.400 574.350 863.250 ;
        RECT 575.550 857.400 577.350 863.250 ;
        RECT 592.650 857.400 594.450 863.250 ;
        RECT 595.650 857.400 597.450 863.250 ;
        RECT 598.650 857.400 600.450 863.250 ;
        RECT 610.650 857.400 612.450 863.250 ;
        RECT 613.650 857.400 615.450 863.250 ;
        RECT 526.800 850.500 528.600 851.400 ;
        RECT 526.800 849.600 530.850 850.500 ;
        RECT 524.100 846.150 525.900 847.950 ;
        RECT 529.950 846.150 530.850 849.600 ;
        RECT 535.950 846.150 537.750 847.950 ;
        RECT 545.100 846.150 546.900 847.950 ;
        RECT 550.950 846.150 552.150 851.400 ;
        RECT 553.950 849.150 555.750 850.950 ;
        RECT 572.550 849.150 573.750 857.400 ;
        RECT 596.250 849.150 597.450 857.400 ;
        RECT 553.950 847.050 556.050 849.150 ;
        RECT 505.950 842.850 508.050 844.950 ;
        RECT 523.950 844.050 526.050 846.150 ;
        RECT 526.950 842.850 529.050 844.950 ;
        RECT 529.950 844.050 532.050 846.150 ;
        RECT 502.950 839.700 504.750 840.600 ;
        RECT 501.450 838.800 504.750 839.700 ;
        RECT 479.100 835.950 484.800 837.600 ;
        RECT 479.700 831.750 481.500 834.600 ;
        RECT 483.000 831.750 484.800 835.950 ;
        RECT 487.200 831.750 489.000 837.600 ;
        RECT 501.450 834.600 502.350 838.800 ;
        RECT 507.000 837.600 508.050 842.850 ;
        RECT 527.250 841.050 529.050 842.850 ;
        RECT 531.000 837.600 532.050 844.050 ;
        RECT 532.950 842.850 535.050 844.950 ;
        RECT 535.950 844.050 538.050 846.150 ;
        RECT 544.950 844.050 547.050 846.150 ;
        RECT 547.950 842.850 550.050 844.950 ;
        RECT 550.950 844.050 553.050 846.150 ;
        RECT 568.950 845.850 571.050 847.950 ;
        RECT 571.950 847.050 574.050 849.150 ;
        RECT 569.100 844.050 570.900 845.850 ;
        RECT 532.950 841.050 534.750 842.850 ;
        RECT 548.100 841.050 549.900 842.850 ;
        RECT 551.850 840.750 553.050 844.050 ;
        RECT 552.000 839.700 555.750 840.750 ;
        RECT 497.550 831.750 499.350 834.600 ;
        RECT 500.550 831.750 502.350 834.600 ;
        RECT 503.550 831.750 505.350 834.600 ;
        RECT 506.550 831.750 508.350 837.600 ;
        RECT 526.800 831.750 528.600 837.600 ;
        RECT 531.000 831.750 532.800 837.600 ;
        RECT 535.200 831.750 537.000 837.600 ;
        RECT 545.550 836.700 553.350 838.050 ;
        RECT 545.550 831.750 547.350 836.700 ;
        RECT 548.550 831.750 550.350 835.800 ;
        RECT 551.550 831.750 553.350 836.700 ;
        RECT 554.550 837.600 555.750 839.700 ;
        RECT 572.550 839.700 573.750 847.050 ;
        RECT 574.950 845.850 577.050 847.950 ;
        RECT 592.950 845.850 595.050 847.950 ;
        RECT 595.950 847.050 598.050 849.150 ;
        RECT 575.100 844.050 576.900 845.850 ;
        RECT 593.100 844.050 594.900 845.850 ;
        RECT 596.250 839.700 597.450 847.050 ;
        RECT 598.950 845.850 601.050 847.950 ;
        RECT 599.100 844.050 600.900 845.850 ;
        RECT 611.400 844.950 612.600 857.400 ;
        RECT 626.550 851.400 628.350 863.250 ;
        RECT 631.050 851.550 632.850 863.250 ;
        RECT 634.050 852.900 635.850 863.250 ;
        RECT 647.550 857.400 649.350 863.250 ;
        RECT 650.550 857.400 652.350 863.250 ;
        RECT 634.050 851.550 636.450 852.900 ;
        RECT 626.550 850.200 627.750 851.400 ;
        RECT 631.950 850.200 633.750 850.650 ;
        RECT 626.550 849.000 633.750 850.200 ;
        RECT 631.950 848.850 633.750 849.000 ;
        RECT 629.100 846.150 630.900 847.950 ;
        RECT 610.950 842.850 613.050 844.950 ;
        RECT 614.100 843.150 615.900 844.950 ;
        RECT 626.100 843.150 627.900 844.950 ;
        RECT 628.950 844.050 631.050 846.150 ;
        RECT 572.550 838.800 576.150 839.700 ;
        RECT 554.550 831.750 556.350 837.600 ;
        RECT 569.850 831.750 571.650 837.600 ;
        RECT 574.350 831.750 576.150 838.800 ;
        RECT 593.850 838.800 597.450 839.700 ;
        RECT 593.850 831.750 595.650 838.800 ;
        RECT 598.350 831.750 600.150 837.600 ;
        RECT 611.400 834.600 612.600 842.850 ;
        RECT 613.950 841.050 616.050 843.150 ;
        RECT 625.950 841.050 628.050 843.150 ;
        RECT 632.700 840.600 633.600 848.850 ;
        RECT 635.100 844.950 636.450 851.550 ;
        RECT 647.100 846.150 648.900 847.950 ;
        RECT 634.950 842.850 637.050 844.950 ;
        RECT 646.950 844.050 649.050 846.150 ;
        RECT 631.950 839.700 633.750 840.600 ;
        RECT 630.450 838.800 633.750 839.700 ;
        RECT 630.450 834.600 631.350 838.800 ;
        RECT 636.000 837.600 637.050 842.850 ;
        RECT 650.700 840.300 651.900 857.400 ;
        RECT 654.150 851.400 655.950 863.250 ;
        RECT 657.150 851.400 658.950 863.250 ;
        RECT 672.300 851.400 674.100 863.250 ;
        RECT 676.500 851.400 678.300 863.250 ;
        RECT 679.800 857.400 681.600 863.250 ;
        RECT 693.300 851.400 695.100 863.250 ;
        RECT 697.500 851.400 699.300 863.250 ;
        RECT 700.800 857.400 702.600 863.250 ;
        RECT 715.650 857.400 717.450 863.250 ;
        RECT 718.650 857.400 720.450 863.250 ;
        RECT 721.650 857.400 723.450 863.250 ;
        RECT 652.950 845.850 655.050 847.950 ;
        RECT 657.150 846.150 658.350 851.400 ;
        RECT 671.100 846.150 672.900 847.950 ;
        RECT 676.950 846.150 678.150 851.400 ;
        RECT 679.950 849.150 681.750 850.950 ;
        RECT 679.950 847.050 682.050 849.150 ;
        RECT 692.100 846.150 693.900 847.950 ;
        RECT 697.950 846.150 699.150 851.400 ;
        RECT 700.950 849.150 702.750 850.950 ;
        RECT 719.250 849.150 720.450 857.400 ;
        RECT 726.150 851.400 727.950 863.250 ;
        RECT 729.150 857.400 730.950 863.250 ;
        RECT 734.250 857.400 736.050 863.250 ;
        RECT 739.050 857.400 740.850 863.250 ;
        RECT 734.550 856.500 735.750 857.400 ;
        RECT 742.050 856.500 743.850 863.250 ;
        RECT 745.950 857.400 747.750 863.250 ;
        RECT 750.150 857.400 751.950 863.250 ;
        RECT 754.650 860.400 756.450 863.250 ;
        RECT 730.950 854.400 735.750 856.500 ;
        RECT 738.150 854.700 745.050 856.500 ;
        RECT 750.150 855.300 754.050 857.400 ;
        RECT 734.550 853.500 735.750 854.400 ;
        RECT 747.450 853.800 749.250 854.400 ;
        RECT 734.550 852.300 742.050 853.500 ;
        RECT 740.250 851.700 742.050 852.300 ;
        RECT 742.950 852.900 749.250 853.800 ;
        RECT 726.150 850.800 737.250 851.400 ;
        RECT 742.950 850.800 743.850 852.900 ;
        RECT 747.450 852.600 749.250 852.900 ;
        RECT 750.150 852.600 752.850 854.400 ;
        RECT 750.150 851.700 751.050 852.600 ;
        RECT 726.150 850.200 743.850 850.800 ;
        RECT 700.950 847.050 703.050 849.150 ;
        RECT 653.100 844.050 654.900 845.850 ;
        RECT 655.950 844.050 658.350 846.150 ;
        RECT 670.950 844.050 673.050 846.150 ;
        RECT 647.550 839.100 655.050 840.300 ;
        RECT 610.650 831.750 612.450 834.600 ;
        RECT 613.650 831.750 615.450 834.600 ;
        RECT 626.550 831.750 628.350 834.600 ;
        RECT 629.550 831.750 631.350 834.600 ;
        RECT 632.550 831.750 634.350 834.600 ;
        RECT 635.550 831.750 637.350 837.600 ;
        RECT 647.550 831.750 649.350 839.100 ;
        RECT 653.250 838.500 655.050 839.100 ;
        RECT 657.150 837.600 658.350 844.050 ;
        RECT 673.950 842.850 676.050 844.950 ;
        RECT 676.950 844.050 679.050 846.150 ;
        RECT 691.950 844.050 694.050 846.150 ;
        RECT 674.100 841.050 675.900 842.850 ;
        RECT 677.850 840.750 679.050 844.050 ;
        RECT 694.950 842.850 697.050 844.950 ;
        RECT 697.950 844.050 700.050 846.150 ;
        RECT 715.950 845.850 718.050 847.950 ;
        RECT 718.950 847.050 721.050 849.150 ;
        RECT 716.100 844.050 717.900 845.850 ;
        RECT 695.100 841.050 696.900 842.850 ;
        RECT 698.850 840.750 700.050 844.050 ;
        RECT 678.000 839.700 681.750 840.750 ;
        RECT 699.000 839.700 702.750 840.750 ;
        RECT 719.250 839.700 720.450 847.050 ;
        RECT 721.950 845.850 724.050 847.950 ;
        RECT 722.100 844.050 723.900 845.850 ;
        RECT 652.050 831.750 653.850 837.600 ;
        RECT 655.050 836.100 658.350 837.600 ;
        RECT 671.550 836.700 679.350 838.050 ;
        RECT 655.050 831.750 656.850 836.100 ;
        RECT 671.550 831.750 673.350 836.700 ;
        RECT 674.550 831.750 676.350 835.800 ;
        RECT 677.550 831.750 679.350 836.700 ;
        RECT 680.550 837.600 681.750 839.700 ;
        RECT 680.550 831.750 682.350 837.600 ;
        RECT 692.550 836.700 700.350 838.050 ;
        RECT 692.550 831.750 694.350 836.700 ;
        RECT 695.550 831.750 697.350 835.800 ;
        RECT 698.550 831.750 700.350 836.700 ;
        RECT 701.550 837.600 702.750 839.700 ;
        RECT 716.850 838.800 720.450 839.700 ;
        RECT 701.550 831.750 703.350 837.600 ;
        RECT 716.850 831.750 718.650 838.800 ;
        RECT 726.150 837.600 727.050 850.200 ;
        RECT 735.450 849.900 743.850 850.200 ;
        RECT 745.050 850.800 751.050 851.700 ;
        RECT 751.950 850.800 754.050 851.700 ;
        RECT 757.650 851.400 759.450 863.250 ;
        RECT 772.650 857.400 774.450 863.250 ;
        RECT 775.650 857.400 777.450 863.250 ;
        RECT 778.650 857.400 780.450 863.250 ;
        RECT 791.400 857.400 793.200 863.250 ;
        RECT 735.450 849.600 737.250 849.900 ;
        RECT 745.050 846.150 745.950 850.800 ;
        RECT 751.950 849.600 756.150 850.800 ;
        RECT 755.250 847.800 757.050 849.600 ;
        RECT 736.950 845.100 739.050 846.150 ;
        RECT 728.100 843.150 729.900 844.950 ;
        RECT 731.100 844.050 739.050 845.100 ;
        RECT 742.950 844.050 745.950 846.150 ;
        RECT 731.100 843.300 732.900 844.050 ;
        RECT 729.000 842.400 729.900 843.150 ;
        RECT 734.100 842.400 735.900 843.000 ;
        RECT 729.000 841.200 735.900 842.400 ;
        RECT 734.850 840.000 735.900 841.200 ;
        RECT 745.050 840.000 745.950 844.050 ;
        RECT 754.950 843.750 757.050 844.050 ;
        RECT 753.150 841.950 757.050 843.750 ;
        RECT 758.250 841.950 759.450 851.400 ;
        RECT 776.250 849.150 777.450 857.400 ;
        RECT 794.700 851.400 796.500 863.250 ;
        RECT 798.900 851.400 800.700 863.250 ;
        RECT 812.550 852.300 814.350 863.250 ;
        RECT 815.550 853.200 817.350 863.250 ;
        RECT 818.550 852.300 820.350 863.250 ;
        RECT 812.550 851.400 820.350 852.300 ;
        RECT 821.550 851.400 823.350 863.250 ;
        RECT 836.400 857.400 838.200 863.250 ;
        RECT 839.700 851.400 841.500 863.250 ;
        RECT 843.900 851.400 845.700 863.250 ;
        RECT 848.550 851.400 850.350 863.250 ;
        RECT 851.550 860.400 853.350 863.250 ;
        RECT 856.050 857.400 857.850 863.250 ;
        RECT 860.250 857.400 862.050 863.250 ;
        RECT 853.950 855.300 857.850 857.400 ;
        RECT 864.150 856.500 865.950 863.250 ;
        RECT 867.150 857.400 868.950 863.250 ;
        RECT 871.950 857.400 873.750 863.250 ;
        RECT 877.050 857.400 878.850 863.250 ;
        RECT 872.250 856.500 873.450 857.400 ;
        RECT 862.950 854.700 869.850 856.500 ;
        RECT 872.250 854.400 877.050 856.500 ;
        RECT 855.150 852.600 857.850 854.400 ;
        RECT 858.750 853.800 860.550 854.400 ;
        RECT 858.750 852.900 865.050 853.800 ;
        RECT 872.250 853.500 873.450 854.400 ;
        RECT 858.750 852.600 860.550 852.900 ;
        RECT 856.950 851.700 857.850 852.600 ;
        RECT 791.250 849.150 793.050 850.950 ;
        RECT 772.950 845.850 775.050 847.950 ;
        RECT 775.950 847.050 778.050 849.150 ;
        RECT 773.100 844.050 774.900 845.850 ;
        RECT 734.850 839.100 745.950 840.000 ;
        RECT 754.950 839.850 759.450 841.950 ;
        RECT 734.850 838.200 735.900 839.100 ;
        RECT 745.050 838.800 745.950 839.100 ;
        RECT 721.350 831.750 723.150 837.600 ;
        RECT 726.150 831.750 727.950 837.600 ;
        RECT 730.950 835.500 733.050 837.600 ;
        RECT 734.550 836.400 736.350 838.200 ;
        RECT 737.850 837.450 739.650 838.200 ;
        RECT 737.850 836.400 742.800 837.450 ;
        RECT 745.050 837.000 746.850 838.800 ;
        RECT 758.250 837.600 759.450 839.850 ;
        RECT 776.250 839.700 777.450 847.050 ;
        RECT 778.950 845.850 781.050 847.950 ;
        RECT 790.950 847.050 793.050 849.150 ;
        RECT 794.850 846.150 796.050 851.400 ;
        RECT 800.100 846.150 801.900 847.950 ;
        RECT 821.700 846.150 822.900 851.400 ;
        RECT 836.250 849.150 838.050 850.950 ;
        RECT 835.950 847.050 838.050 849.150 ;
        RECT 839.850 846.150 841.050 851.400 ;
        RECT 845.100 846.150 846.900 847.950 ;
        RECT 779.100 844.050 780.900 845.850 ;
        RECT 793.950 844.050 796.050 846.150 ;
        RECT 793.950 840.750 795.150 844.050 ;
        RECT 796.950 842.850 799.050 844.950 ;
        RECT 799.950 844.050 802.050 846.150 ;
        RECT 811.950 842.850 814.050 844.950 ;
        RECT 815.100 843.150 816.900 844.950 ;
        RECT 797.100 841.050 798.900 842.850 ;
        RECT 812.100 841.050 813.900 842.850 ;
        RECT 814.950 841.050 817.050 843.150 ;
        RECT 817.950 842.850 820.050 844.950 ;
        RECT 820.950 844.050 823.050 846.150 ;
        RECT 838.950 844.050 841.050 846.150 ;
        RECT 818.100 841.050 819.900 842.850 ;
        RECT 751.950 836.700 754.050 837.600 ;
        RECT 732.000 834.600 733.050 835.500 ;
        RECT 741.750 834.600 742.800 836.400 ;
        RECT 750.300 835.500 754.050 836.700 ;
        RECT 750.300 834.600 751.350 835.500 ;
        RECT 729.150 831.750 730.950 834.600 ;
        RECT 732.000 833.700 735.750 834.600 ;
        RECT 733.950 831.750 735.750 833.700 ;
        RECT 738.450 831.750 740.250 834.600 ;
        RECT 741.750 831.750 743.550 834.600 ;
        RECT 745.650 831.750 747.450 834.600 ;
        RECT 749.850 831.750 751.650 834.600 ;
        RECT 754.350 831.750 756.150 834.600 ;
        RECT 757.650 831.750 759.450 837.600 ;
        RECT 773.850 838.800 777.450 839.700 ;
        RECT 791.250 839.700 795.000 840.750 ;
        RECT 773.850 831.750 775.650 838.800 ;
        RECT 791.250 837.600 792.450 839.700 ;
        RECT 778.350 831.750 780.150 837.600 ;
        RECT 790.650 831.750 792.450 837.600 ;
        RECT 793.650 836.700 801.450 838.050 ;
        RECT 821.700 837.600 822.900 844.050 ;
        RECT 838.950 840.750 840.150 844.050 ;
        RECT 841.950 842.850 844.050 844.950 ;
        RECT 844.950 844.050 847.050 846.150 ;
        RECT 842.100 841.050 843.900 842.850 ;
        RECT 848.550 841.950 849.750 851.400 ;
        RECT 853.950 850.800 856.050 851.700 ;
        RECT 856.950 850.800 862.950 851.700 ;
        RECT 851.850 849.600 856.050 850.800 ;
        RECT 850.950 847.800 852.750 849.600 ;
        RECT 862.050 846.150 862.950 850.800 ;
        RECT 864.150 850.800 865.050 852.900 ;
        RECT 865.950 852.300 873.450 853.500 ;
        RECT 865.950 851.700 867.750 852.300 ;
        RECT 880.050 851.400 881.850 863.250 ;
        RECT 870.750 850.800 881.850 851.400 ;
        RECT 864.150 850.200 881.850 850.800 ;
        RECT 864.150 849.900 872.550 850.200 ;
        RECT 870.750 849.600 872.550 849.900 ;
        RECT 862.050 844.050 865.050 846.150 ;
        RECT 868.950 845.100 871.050 846.150 ;
        RECT 868.950 844.050 876.900 845.100 ;
        RECT 850.950 843.750 853.050 844.050 ;
        RECT 850.950 841.950 854.850 843.750 ;
        RECT 836.250 839.700 840.000 840.750 ;
        RECT 848.550 839.850 853.050 841.950 ;
        RECT 862.050 840.000 862.950 844.050 ;
        RECT 875.100 843.300 876.900 844.050 ;
        RECT 878.100 843.150 879.900 844.950 ;
        RECT 872.100 842.400 873.900 843.000 ;
        RECT 878.100 842.400 879.000 843.150 ;
        RECT 872.100 841.200 879.000 842.400 ;
        RECT 872.100 840.000 873.150 841.200 ;
        RECT 836.250 837.600 837.450 839.700 ;
        RECT 793.650 831.750 795.450 836.700 ;
        RECT 796.650 831.750 798.450 835.800 ;
        RECT 799.650 831.750 801.450 836.700 ;
        RECT 813.000 831.750 814.800 837.600 ;
        RECT 817.200 835.950 822.900 837.600 ;
        RECT 817.200 831.750 819.000 835.950 ;
        RECT 820.500 831.750 822.300 834.600 ;
        RECT 835.650 831.750 837.450 837.600 ;
        RECT 838.650 836.700 846.450 838.050 ;
        RECT 838.650 831.750 840.450 836.700 ;
        RECT 841.650 831.750 843.450 835.800 ;
        RECT 844.650 831.750 846.450 836.700 ;
        RECT 848.550 837.600 849.750 839.850 ;
        RECT 862.050 839.100 873.150 840.000 ;
        RECT 862.050 838.800 862.950 839.100 ;
        RECT 848.550 831.750 850.350 837.600 ;
        RECT 853.950 836.700 856.050 837.600 ;
        RECT 861.150 837.000 862.950 838.800 ;
        RECT 872.100 838.200 873.150 839.100 ;
        RECT 868.350 837.450 870.150 838.200 ;
        RECT 853.950 835.500 857.700 836.700 ;
        RECT 856.650 834.600 857.700 835.500 ;
        RECT 865.200 836.400 870.150 837.450 ;
        RECT 871.650 836.400 873.450 838.200 ;
        RECT 880.950 837.600 881.850 850.200 ;
        RECT 865.200 834.600 866.250 836.400 ;
        RECT 874.950 835.500 877.050 837.600 ;
        RECT 874.950 834.600 876.000 835.500 ;
        RECT 851.850 831.750 853.650 834.600 ;
        RECT 856.350 831.750 858.150 834.600 ;
        RECT 860.550 831.750 862.350 834.600 ;
        RECT 864.450 831.750 866.250 834.600 ;
        RECT 867.750 831.750 869.550 834.600 ;
        RECT 872.250 833.700 876.000 834.600 ;
        RECT 872.250 831.750 874.050 833.700 ;
        RECT 877.050 831.750 878.850 834.600 ;
        RECT 880.050 831.750 881.850 837.600 ;
        RECT 13.650 821.400 15.450 827.250 ;
        RECT 14.250 819.300 15.450 821.400 ;
        RECT 16.650 822.300 18.450 827.250 ;
        RECT 19.650 823.200 21.450 827.250 ;
        RECT 22.650 822.300 24.450 827.250 ;
        RECT 16.650 820.950 24.450 822.300 ;
        RECT 36.000 821.400 37.800 827.250 ;
        RECT 40.200 821.400 42.000 827.250 ;
        RECT 44.400 821.400 46.200 827.250 ;
        RECT 59.550 824.400 61.350 827.250 ;
        RECT 62.550 824.400 64.350 827.250 ;
        RECT 14.250 818.250 18.000 819.300 ;
        RECT 16.950 814.950 18.150 818.250 ;
        RECT 20.100 816.150 21.900 817.950 ;
        RECT 38.250 816.150 40.050 817.950 ;
        RECT 16.950 812.850 19.050 814.950 ;
        RECT 19.950 814.050 22.050 816.150 ;
        RECT 22.950 812.850 25.050 814.950 ;
        RECT 34.950 812.850 37.050 814.950 ;
        RECT 37.950 814.050 40.050 816.150 ;
        RECT 40.950 814.950 42.000 821.400 ;
        RECT 43.950 816.150 45.750 817.950 ;
        RECT 40.950 812.850 43.050 814.950 ;
        RECT 43.950 814.050 46.050 816.150 ;
        RECT 58.950 815.850 61.050 817.950 ;
        RECT 62.400 816.150 63.600 824.400 ;
        RECT 79.650 821.400 81.450 827.250 ;
        RECT 80.250 819.300 81.450 821.400 ;
        RECT 82.650 822.300 84.450 827.250 ;
        RECT 85.650 823.200 87.450 827.250 ;
        RECT 88.650 822.300 90.450 827.250 ;
        RECT 98.550 824.400 100.350 827.250 ;
        RECT 101.550 824.400 103.350 827.250 ;
        RECT 104.550 824.400 106.350 827.250 ;
        RECT 82.650 820.950 90.450 822.300 ;
        RECT 80.250 818.250 84.000 819.300 ;
        RECT 46.950 812.850 49.050 814.950 ;
        RECT 59.100 814.050 60.900 815.850 ;
        RECT 61.950 814.050 64.050 816.150 ;
        RECT 82.950 814.950 84.150 818.250 ;
        RECT 102.000 817.950 103.050 824.400 ;
        RECT 122.850 820.200 124.650 827.250 ;
        RECT 127.350 821.400 129.150 827.250 ;
        RECT 139.650 826.500 147.450 827.250 ;
        RECT 139.650 821.400 141.450 826.500 ;
        RECT 142.650 821.400 144.450 825.600 ;
        RECT 145.650 822.000 147.450 826.500 ;
        RECT 148.650 822.900 150.450 827.250 ;
        RECT 151.650 822.000 153.450 827.250 ;
        RECT 122.850 819.300 126.450 820.200 ;
        RECT 86.100 816.150 87.900 817.950 ;
        RECT 13.950 809.850 16.050 811.950 ;
        RECT 14.250 808.050 16.050 809.850 ;
        RECT 17.850 807.600 19.050 812.850 ;
        RECT 23.100 811.050 24.900 812.850 ;
        RECT 35.250 811.050 37.050 812.850 ;
        RECT 42.150 809.400 43.050 812.850 ;
        RECT 47.100 811.050 48.900 812.850 ;
        RECT 42.150 808.500 46.200 809.400 ;
        RECT 44.400 807.600 46.200 808.500 ;
        RECT 14.400 795.750 16.200 801.600 ;
        RECT 17.700 795.750 19.500 807.600 ;
        RECT 21.900 795.750 23.700 807.600 ;
        RECT 35.550 806.400 43.350 807.300 ;
        RECT 35.550 795.750 37.350 806.400 ;
        RECT 38.550 795.750 40.350 805.500 ;
        RECT 41.550 796.500 43.350 806.400 ;
        RECT 44.550 797.400 46.350 807.600 ;
        RECT 47.550 796.500 49.350 807.600 ;
        RECT 62.400 801.600 63.600 814.050 ;
        RECT 82.950 812.850 85.050 814.950 ;
        RECT 85.950 814.050 88.050 816.150 ;
        RECT 100.950 815.850 103.050 817.950 ;
        RECT 88.950 812.850 91.050 814.950 ;
        RECT 97.950 812.850 100.050 814.950 ;
        RECT 79.950 809.850 82.050 811.950 ;
        RECT 80.250 808.050 82.050 809.850 ;
        RECT 83.850 807.600 85.050 812.850 ;
        RECT 89.100 811.050 90.900 812.850 ;
        RECT 98.100 811.050 99.900 812.850 ;
        RECT 102.000 808.650 103.050 815.850 ;
        RECT 103.950 812.850 106.050 814.950 ;
        RECT 122.100 813.150 123.900 814.950 ;
        RECT 104.100 811.050 105.900 812.850 ;
        RECT 121.950 811.050 124.050 813.150 ;
        RECT 125.250 811.950 126.450 819.300 ;
        RECT 143.250 819.900 144.150 821.400 ;
        RECT 145.650 821.100 153.450 822.000 ;
        RECT 169.800 821.400 171.600 827.250 ;
        RECT 174.000 821.400 175.800 827.250 ;
        RECT 178.200 821.400 180.000 827.250 ;
        RECT 191.550 824.400 193.350 827.250 ;
        RECT 194.550 824.400 196.350 827.250 ;
        RECT 208.650 824.400 210.450 827.250 ;
        RECT 211.650 824.400 213.450 827.250 ;
        RECT 143.250 818.850 147.600 819.900 ;
        RECT 143.700 816.150 145.500 817.950 ;
        RECT 128.100 813.150 129.900 814.950 ;
        RECT 124.950 809.850 127.050 811.950 ;
        RECT 127.950 811.050 130.050 813.150 ;
        RECT 139.950 812.850 142.050 814.950 ;
        RECT 142.950 814.050 145.050 816.150 ;
        RECT 146.400 814.950 147.600 818.850 ;
        RECT 149.100 816.150 150.900 817.950 ;
        RECT 170.250 816.150 172.050 817.950 ;
        RECT 145.950 812.850 148.050 814.950 ;
        RECT 148.950 814.050 151.050 816.150 ;
        RECT 151.950 812.850 154.050 814.950 ;
        RECT 166.950 812.850 169.050 814.950 ;
        RECT 169.950 814.050 172.050 816.150 ;
        RECT 174.000 814.950 175.050 821.400 ;
        RECT 172.950 812.850 175.050 814.950 ;
        RECT 175.950 816.150 177.750 817.950 ;
        RECT 175.950 814.050 178.050 816.150 ;
        RECT 190.950 815.850 193.050 817.950 ;
        RECT 194.400 816.150 195.600 824.400 ;
        RECT 209.400 816.150 210.600 824.400 ;
        RECT 224.850 820.200 226.650 827.250 ;
        RECT 229.350 821.400 231.150 827.250 ;
        RECT 244.650 821.400 246.450 827.250 ;
        RECT 224.850 819.300 228.450 820.200 ;
        RECT 178.950 812.850 181.050 814.950 ;
        RECT 191.100 814.050 192.900 815.850 ;
        RECT 193.950 814.050 196.050 816.150 ;
        RECT 208.950 814.050 211.050 816.150 ;
        RECT 211.950 815.850 214.050 817.950 ;
        RECT 212.100 814.050 213.900 815.850 ;
        RECT 140.250 811.050 142.050 812.850 ;
        RECT 102.000 807.600 104.550 808.650 ;
        RECT 41.550 795.750 49.350 796.500 ;
        RECT 59.550 795.750 61.350 801.600 ;
        RECT 62.550 795.750 64.350 801.600 ;
        RECT 80.400 795.750 82.200 801.600 ;
        RECT 83.700 795.750 85.500 807.600 ;
        RECT 87.900 795.750 89.700 807.600 ;
        RECT 98.550 795.750 100.350 807.600 ;
        RECT 102.750 795.750 104.550 807.600 ;
        RECT 125.250 801.600 126.450 809.850 ;
        RECT 146.250 807.600 147.450 812.850 ;
        RECT 152.100 811.050 153.900 812.850 ;
        RECT 167.100 811.050 168.900 812.850 ;
        RECT 172.950 809.400 173.850 812.850 ;
        RECT 178.950 811.050 180.750 812.850 ;
        RECT 169.800 808.500 173.850 809.400 ;
        RECT 169.800 807.600 171.600 808.500 ;
        RECT 121.650 795.750 123.450 801.600 ;
        RECT 124.650 795.750 126.450 801.600 ;
        RECT 127.650 795.750 129.450 801.600 ;
        RECT 141.150 795.750 142.950 807.600 ;
        RECT 145.650 795.750 148.950 807.600 ;
        RECT 151.650 795.750 153.450 807.600 ;
        RECT 166.650 796.500 168.450 807.600 ;
        RECT 169.650 797.400 171.450 807.600 ;
        RECT 172.650 806.400 180.450 807.300 ;
        RECT 172.650 796.500 174.450 806.400 ;
        RECT 166.650 795.750 174.450 796.500 ;
        RECT 175.650 795.750 177.450 805.500 ;
        RECT 178.650 795.750 180.450 806.400 ;
        RECT 194.400 801.600 195.600 814.050 ;
        RECT 209.400 801.600 210.600 814.050 ;
        RECT 224.100 813.150 225.900 814.950 ;
        RECT 223.950 811.050 226.050 813.150 ;
        RECT 227.250 811.950 228.450 819.300 ;
        RECT 245.250 819.300 246.450 821.400 ;
        RECT 247.650 822.300 249.450 827.250 ;
        RECT 250.650 823.200 252.450 827.250 ;
        RECT 253.650 822.300 255.450 827.250 ;
        RECT 247.650 820.950 255.450 822.300 ;
        RECT 263.550 822.300 265.350 827.250 ;
        RECT 266.550 823.200 268.350 827.250 ;
        RECT 269.550 822.300 271.350 827.250 ;
        RECT 263.550 820.950 271.350 822.300 ;
        RECT 272.550 821.400 274.350 827.250 ;
        RECT 284.550 824.400 286.350 827.250 ;
        RECT 287.550 824.400 289.350 827.250 ;
        RECT 304.650 826.500 312.450 827.250 ;
        RECT 272.550 819.300 273.750 821.400 ;
        RECT 245.250 818.250 249.000 819.300 ;
        RECT 270.000 818.250 273.750 819.300 ;
        RECT 247.950 814.950 249.150 818.250 ;
        RECT 251.100 816.150 252.900 817.950 ;
        RECT 266.100 816.150 267.900 817.950 ;
        RECT 230.100 813.150 231.900 814.950 ;
        RECT 226.950 809.850 229.050 811.950 ;
        RECT 229.950 811.050 232.050 813.150 ;
        RECT 247.950 812.850 250.050 814.950 ;
        RECT 250.950 814.050 253.050 816.150 ;
        RECT 253.950 812.850 256.050 814.950 ;
        RECT 262.950 812.850 265.050 814.950 ;
        RECT 265.950 814.050 268.050 816.150 ;
        RECT 269.850 814.950 271.050 818.250 ;
        RECT 283.950 815.850 286.050 817.950 ;
        RECT 287.400 816.150 288.600 824.400 ;
        RECT 304.650 821.400 306.450 826.500 ;
        RECT 307.650 821.400 309.450 825.600 ;
        RECT 310.650 822.000 312.450 826.500 ;
        RECT 313.650 822.900 315.450 827.250 ;
        RECT 316.650 822.000 318.450 827.250 ;
        RECT 328.650 824.400 330.450 827.250 ;
        RECT 331.650 824.400 333.450 827.250 ;
        RECT 343.650 826.500 351.450 827.250 ;
        RECT 308.250 819.900 309.150 821.400 ;
        RECT 310.650 821.100 318.450 822.000 ;
        RECT 308.250 818.850 312.600 819.900 ;
        RECT 308.700 816.150 310.500 817.950 ;
        RECT 268.950 812.850 271.050 814.950 ;
        RECT 284.100 814.050 285.900 815.850 ;
        RECT 286.950 814.050 289.050 816.150 ;
        RECT 244.950 809.850 247.050 811.950 ;
        RECT 227.250 801.600 228.450 809.850 ;
        RECT 245.250 808.050 247.050 809.850 ;
        RECT 248.850 807.600 250.050 812.850 ;
        RECT 254.100 811.050 255.900 812.850 ;
        RECT 263.100 811.050 264.900 812.850 ;
        RECT 268.950 807.600 270.150 812.850 ;
        RECT 271.950 809.850 274.050 811.950 ;
        RECT 271.950 808.050 273.750 809.850 ;
        RECT 191.550 795.750 193.350 801.600 ;
        RECT 194.550 795.750 196.350 801.600 ;
        RECT 208.650 795.750 210.450 801.600 ;
        RECT 211.650 795.750 213.450 801.600 ;
        RECT 223.650 795.750 225.450 801.600 ;
        RECT 226.650 795.750 228.450 801.600 ;
        RECT 229.650 795.750 231.450 801.600 ;
        RECT 245.400 795.750 247.200 801.600 ;
        RECT 248.700 795.750 250.500 807.600 ;
        RECT 252.900 795.750 254.700 807.600 ;
        RECT 264.300 795.750 266.100 807.600 ;
        RECT 268.500 795.750 270.300 807.600 ;
        RECT 287.400 801.600 288.600 814.050 ;
        RECT 304.950 812.850 307.050 814.950 ;
        RECT 307.950 814.050 310.050 816.150 ;
        RECT 311.400 814.950 312.600 818.850 ;
        RECT 314.100 816.150 315.900 817.950 ;
        RECT 329.400 816.150 330.600 824.400 ;
        RECT 343.650 821.400 345.450 826.500 ;
        RECT 346.650 821.400 348.450 825.600 ;
        RECT 349.650 822.000 351.450 826.500 ;
        RECT 352.650 822.900 354.450 827.250 ;
        RECT 355.650 822.000 357.450 827.250 ;
        RECT 347.250 819.900 348.150 821.400 ;
        RECT 349.650 821.100 357.450 822.000 ;
        RECT 367.650 826.500 375.450 827.250 ;
        RECT 367.650 821.400 369.450 826.500 ;
        RECT 370.650 821.400 372.450 825.600 ;
        RECT 373.650 822.000 375.450 826.500 ;
        RECT 376.650 822.900 378.450 827.250 ;
        RECT 379.650 822.000 381.450 827.250 ;
        RECT 395.700 824.400 397.500 827.250 ;
        RECT 399.000 823.050 400.800 827.250 ;
        RECT 371.250 819.900 372.150 821.400 ;
        RECT 373.650 821.100 381.450 822.000 ;
        RECT 395.100 821.400 400.800 823.050 ;
        RECT 403.200 821.400 405.000 827.250 ;
        RECT 417.000 821.400 418.800 827.250 ;
        RECT 421.200 823.050 423.000 827.250 ;
        RECT 424.500 824.400 426.300 827.250 ;
        RECT 439.650 824.400 441.450 827.250 ;
        RECT 442.650 824.400 444.450 827.250 ;
        RECT 421.200 821.400 426.900 823.050 ;
        RECT 347.250 818.850 351.600 819.900 ;
        RECT 371.250 818.850 375.600 819.900 ;
        RECT 310.950 812.850 313.050 814.950 ;
        RECT 313.950 814.050 316.050 816.150 ;
        RECT 316.950 812.850 319.050 814.950 ;
        RECT 328.950 814.050 331.050 816.150 ;
        RECT 331.950 815.850 334.050 817.950 ;
        RECT 347.700 816.150 349.500 817.950 ;
        RECT 332.100 814.050 333.900 815.850 ;
        RECT 305.250 811.050 307.050 812.850 ;
        RECT 311.250 807.600 312.450 812.850 ;
        RECT 317.100 811.050 318.900 812.850 ;
        RECT 271.800 795.750 273.600 801.600 ;
        RECT 284.550 795.750 286.350 801.600 ;
        RECT 287.550 795.750 289.350 801.600 ;
        RECT 306.150 795.750 307.950 807.600 ;
        RECT 310.650 795.750 313.950 807.600 ;
        RECT 316.650 795.750 318.450 807.600 ;
        RECT 329.400 801.600 330.600 814.050 ;
        RECT 343.950 812.850 346.050 814.950 ;
        RECT 346.950 814.050 349.050 816.150 ;
        RECT 350.400 814.950 351.600 818.850 ;
        RECT 353.100 816.150 354.900 817.950 ;
        RECT 371.700 816.150 373.500 817.950 ;
        RECT 349.950 812.850 352.050 814.950 ;
        RECT 352.950 814.050 355.050 816.150 ;
        RECT 355.950 812.850 358.050 814.950 ;
        RECT 367.950 812.850 370.050 814.950 ;
        RECT 370.950 814.050 373.050 816.150 ;
        RECT 374.400 814.950 375.600 818.850 ;
        RECT 377.100 816.150 378.900 817.950 ;
        RECT 373.950 812.850 376.050 814.950 ;
        RECT 376.950 814.050 379.050 816.150 ;
        RECT 395.100 814.950 396.300 821.400 ;
        RECT 398.100 816.150 399.900 817.950 ;
        RECT 379.950 812.850 382.050 814.950 ;
        RECT 394.950 812.850 397.050 814.950 ;
        RECT 397.950 814.050 400.050 816.150 ;
        RECT 400.950 815.850 403.050 817.950 ;
        RECT 404.100 816.150 405.900 817.950 ;
        RECT 416.100 816.150 417.900 817.950 ;
        RECT 401.100 814.050 402.900 815.850 ;
        RECT 403.950 814.050 406.050 816.150 ;
        RECT 415.950 814.050 418.050 816.150 ;
        RECT 418.950 815.850 421.050 817.950 ;
        RECT 422.100 816.150 423.900 817.950 ;
        RECT 419.100 814.050 420.900 815.850 ;
        RECT 421.950 814.050 424.050 816.150 ;
        RECT 425.700 814.950 426.900 821.400 ;
        RECT 440.400 816.150 441.600 824.400 ;
        RECT 458.850 820.200 460.650 827.250 ;
        RECT 463.350 821.400 465.150 827.250 ;
        RECT 476.850 820.200 478.650 827.250 ;
        RECT 481.350 821.400 483.150 827.250 ;
        RECT 491.850 821.400 493.650 827.250 ;
        RECT 496.350 820.200 498.150 827.250 ;
        RECT 511.650 821.400 513.450 827.250 ;
        RECT 458.850 819.300 462.450 820.200 ;
        RECT 476.850 819.300 480.450 820.200 ;
        RECT 424.950 812.850 427.050 814.950 ;
        RECT 439.950 814.050 442.050 816.150 ;
        RECT 442.950 815.850 445.050 817.950 ;
        RECT 443.100 814.050 444.900 815.850 ;
        RECT 344.250 811.050 346.050 812.850 ;
        RECT 350.250 807.600 351.450 812.850 ;
        RECT 356.100 811.050 357.900 812.850 ;
        RECT 368.250 811.050 370.050 812.850 ;
        RECT 374.250 807.600 375.450 812.850 ;
        RECT 380.100 811.050 381.900 812.850 ;
        RECT 395.100 807.600 396.300 812.850 ;
        RECT 425.700 807.600 426.900 812.850 ;
        RECT 328.650 795.750 330.450 801.600 ;
        RECT 331.650 795.750 333.450 801.600 ;
        RECT 345.150 795.750 346.950 807.600 ;
        RECT 349.650 795.750 352.950 807.600 ;
        RECT 355.650 795.750 357.450 807.600 ;
        RECT 369.150 795.750 370.950 807.600 ;
        RECT 373.650 795.750 376.950 807.600 ;
        RECT 379.650 795.750 381.450 807.600 ;
        RECT 394.650 795.750 396.450 807.600 ;
        RECT 397.650 806.700 405.450 807.600 ;
        RECT 397.650 795.750 399.450 806.700 ;
        RECT 400.650 795.750 402.450 805.800 ;
        RECT 403.650 795.750 405.450 806.700 ;
        RECT 416.550 806.700 424.350 807.600 ;
        RECT 416.550 795.750 418.350 806.700 ;
        RECT 419.550 795.750 421.350 805.800 ;
        RECT 422.550 795.750 424.350 806.700 ;
        RECT 425.550 795.750 427.350 807.600 ;
        RECT 440.400 801.600 441.600 814.050 ;
        RECT 458.100 813.150 459.900 814.950 ;
        RECT 457.950 811.050 460.050 813.150 ;
        RECT 461.250 811.950 462.450 819.300 ;
        RECT 464.100 813.150 465.900 814.950 ;
        RECT 476.100 813.150 477.900 814.950 ;
        RECT 460.950 809.850 463.050 811.950 ;
        RECT 463.950 811.050 466.050 813.150 ;
        RECT 475.950 811.050 478.050 813.150 ;
        RECT 479.250 811.950 480.450 819.300 ;
        RECT 494.550 819.300 498.150 820.200 ;
        RECT 512.250 819.300 513.450 821.400 ;
        RECT 514.650 822.300 516.450 827.250 ;
        RECT 517.650 823.200 519.450 827.250 ;
        RECT 520.650 822.300 522.450 827.250 ;
        RECT 514.650 820.950 522.450 822.300 ;
        RECT 536.850 820.200 538.650 827.250 ;
        RECT 541.350 821.400 543.150 827.250 ;
        RECT 554.850 820.200 556.650 827.250 ;
        RECT 559.350 821.400 561.150 827.250 ;
        RECT 572.850 820.200 574.650 827.250 ;
        RECT 577.350 821.400 579.150 827.250 ;
        RECT 591.000 821.400 592.800 827.250 ;
        RECT 595.200 823.050 597.000 827.250 ;
        RECT 598.500 824.400 600.300 827.250 ;
        RECT 595.200 821.400 600.900 823.050 ;
        RECT 616.650 821.400 618.450 827.250 ;
        RECT 536.850 819.300 540.450 820.200 ;
        RECT 554.850 819.300 558.450 820.200 ;
        RECT 572.850 819.300 576.450 820.200 ;
        RECT 482.100 813.150 483.900 814.950 ;
        RECT 491.100 813.150 492.900 814.950 ;
        RECT 478.950 809.850 481.050 811.950 ;
        RECT 481.950 811.050 484.050 813.150 ;
        RECT 490.950 811.050 493.050 813.150 ;
        RECT 494.550 811.950 495.750 819.300 ;
        RECT 512.250 818.250 516.000 819.300 ;
        RECT 514.950 814.950 516.150 818.250 ;
        RECT 518.100 816.150 519.900 817.950 ;
        RECT 497.100 813.150 498.900 814.950 ;
        RECT 493.950 809.850 496.050 811.950 ;
        RECT 496.950 811.050 499.050 813.150 ;
        RECT 514.950 812.850 517.050 814.950 ;
        RECT 517.950 814.050 520.050 816.150 ;
        RECT 520.950 812.850 523.050 814.950 ;
        RECT 536.100 813.150 537.900 814.950 ;
        RECT 511.950 809.850 514.050 811.950 ;
        RECT 461.250 801.600 462.450 809.850 ;
        RECT 479.250 801.600 480.450 809.850 ;
        RECT 494.550 801.600 495.750 809.850 ;
        RECT 512.250 808.050 514.050 809.850 ;
        RECT 515.850 807.600 517.050 812.850 ;
        RECT 521.100 811.050 522.900 812.850 ;
        RECT 535.950 811.050 538.050 813.150 ;
        RECT 539.250 811.950 540.450 819.300 ;
        RECT 542.100 813.150 543.900 814.950 ;
        RECT 554.100 813.150 555.900 814.950 ;
        RECT 538.950 809.850 541.050 811.950 ;
        RECT 541.950 811.050 544.050 813.150 ;
        RECT 553.950 811.050 556.050 813.150 ;
        RECT 557.250 811.950 558.450 819.300 ;
        RECT 560.100 813.150 561.900 814.950 ;
        RECT 572.100 813.150 573.900 814.950 ;
        RECT 556.950 809.850 559.050 811.950 ;
        RECT 559.950 811.050 562.050 813.150 ;
        RECT 571.950 811.050 574.050 813.150 ;
        RECT 575.250 811.950 576.450 819.300 ;
        RECT 590.100 816.150 591.900 817.950 ;
        RECT 578.100 813.150 579.900 814.950 ;
        RECT 589.950 814.050 592.050 816.150 ;
        RECT 592.950 815.850 595.050 817.950 ;
        RECT 596.100 816.150 597.900 817.950 ;
        RECT 593.100 814.050 594.900 815.850 ;
        RECT 595.950 814.050 598.050 816.150 ;
        RECT 599.700 814.950 600.900 821.400 ;
        RECT 617.250 819.300 618.450 821.400 ;
        RECT 619.650 822.300 621.450 827.250 ;
        RECT 622.650 823.200 624.450 827.250 ;
        RECT 625.650 822.300 627.450 827.250 ;
        RECT 619.650 820.950 627.450 822.300 ;
        RECT 625.950 819.450 628.050 820.050 ;
        RECT 631.950 819.450 634.050 820.050 ;
        RECT 617.250 818.250 621.000 819.300 ;
        RECT 625.950 818.550 634.050 819.450 ;
        RECT 635.550 819.900 637.350 827.250 ;
        RECT 640.050 821.400 641.850 827.250 ;
        RECT 643.050 822.900 644.850 827.250 ;
        RECT 643.050 821.400 646.350 822.900 ;
        RECT 641.250 819.900 643.050 820.500 ;
        RECT 635.550 818.700 643.050 819.900 ;
        RECT 619.950 814.950 621.150 818.250 ;
        RECT 625.950 817.950 628.050 818.550 ;
        RECT 631.950 817.950 634.050 818.550 ;
        RECT 623.100 816.150 624.900 817.950 ;
        RECT 574.950 809.850 577.050 811.950 ;
        RECT 577.950 811.050 580.050 813.150 ;
        RECT 598.950 812.850 601.050 814.950 ;
        RECT 619.950 812.850 622.050 814.950 ;
        RECT 622.950 814.050 625.050 816.150 ;
        RECT 625.950 812.850 628.050 814.950 ;
        RECT 634.950 812.850 637.050 814.950 ;
        RECT 439.650 795.750 441.450 801.600 ;
        RECT 442.650 795.750 444.450 801.600 ;
        RECT 457.650 795.750 459.450 801.600 ;
        RECT 460.650 795.750 462.450 801.600 ;
        RECT 463.650 795.750 465.450 801.600 ;
        RECT 475.650 795.750 477.450 801.600 ;
        RECT 478.650 795.750 480.450 801.600 ;
        RECT 481.650 795.750 483.450 801.600 ;
        RECT 491.550 795.750 493.350 801.600 ;
        RECT 494.550 795.750 496.350 801.600 ;
        RECT 497.550 795.750 499.350 801.600 ;
        RECT 512.400 795.750 514.200 801.600 ;
        RECT 515.700 795.750 517.500 807.600 ;
        RECT 519.900 795.750 521.700 807.600 ;
        RECT 539.250 801.600 540.450 809.850 ;
        RECT 557.250 801.600 558.450 809.850 ;
        RECT 575.250 801.600 576.450 809.850 ;
        RECT 599.700 807.600 600.900 812.850 ;
        RECT 616.950 809.850 619.050 811.950 ;
        RECT 617.250 808.050 619.050 809.850 ;
        RECT 620.850 807.600 622.050 812.850 ;
        RECT 626.100 811.050 627.900 812.850 ;
        RECT 635.100 811.050 636.900 812.850 ;
        RECT 590.550 806.700 598.350 807.600 ;
        RECT 535.650 795.750 537.450 801.600 ;
        RECT 538.650 795.750 540.450 801.600 ;
        RECT 541.650 795.750 543.450 801.600 ;
        RECT 553.650 795.750 555.450 801.600 ;
        RECT 556.650 795.750 558.450 801.600 ;
        RECT 559.650 795.750 561.450 801.600 ;
        RECT 571.650 795.750 573.450 801.600 ;
        RECT 574.650 795.750 576.450 801.600 ;
        RECT 577.650 795.750 579.450 801.600 ;
        RECT 590.550 795.750 592.350 806.700 ;
        RECT 593.550 795.750 595.350 805.800 ;
        RECT 596.550 795.750 598.350 806.700 ;
        RECT 599.550 795.750 601.350 807.600 ;
        RECT 617.400 795.750 619.200 801.600 ;
        RECT 620.700 795.750 622.500 807.600 ;
        RECT 624.900 795.750 626.700 807.600 ;
        RECT 638.700 801.600 639.900 818.700 ;
        RECT 645.150 814.950 646.350 821.400 ;
        RECT 659.550 822.300 661.350 827.250 ;
        RECT 662.550 823.200 664.350 827.250 ;
        RECT 665.550 822.300 667.350 827.250 ;
        RECT 659.550 820.950 667.350 822.300 ;
        RECT 668.550 821.400 670.350 827.250 ;
        RECT 683.550 822.300 685.350 827.250 ;
        RECT 686.550 823.200 688.350 827.250 ;
        RECT 689.550 822.300 691.350 827.250 ;
        RECT 668.550 819.300 669.750 821.400 ;
        RECT 683.550 820.950 691.350 822.300 ;
        RECT 692.550 821.400 694.350 827.250 ;
        RECT 704.550 822.300 706.350 827.250 ;
        RECT 707.550 823.200 709.350 827.250 ;
        RECT 710.550 822.300 712.350 827.250 ;
        RECT 692.550 819.300 693.750 821.400 ;
        RECT 704.550 820.950 712.350 822.300 ;
        RECT 713.550 821.400 715.350 827.250 ;
        RECT 713.550 819.300 714.750 821.400 ;
        RECT 728.850 820.200 730.650 827.250 ;
        RECT 733.350 821.400 735.150 827.250 ;
        RECT 738.150 821.400 739.950 827.250 ;
        RECT 741.150 824.400 742.950 827.250 ;
        RECT 745.950 825.300 747.750 827.250 ;
        RECT 744.000 824.400 747.750 825.300 ;
        RECT 750.450 824.400 752.250 827.250 ;
        RECT 753.750 824.400 755.550 827.250 ;
        RECT 757.650 824.400 759.450 827.250 ;
        RECT 761.850 824.400 763.650 827.250 ;
        RECT 766.350 824.400 768.150 827.250 ;
        RECT 744.000 823.500 745.050 824.400 ;
        RECT 742.950 821.400 745.050 823.500 ;
        RECT 753.750 822.600 754.800 824.400 ;
        RECT 728.850 819.300 732.450 820.200 ;
        RECT 666.000 818.250 669.750 819.300 ;
        RECT 690.000 818.250 693.750 819.300 ;
        RECT 711.000 818.250 714.750 819.300 ;
        RECT 662.100 816.150 663.900 817.950 ;
        RECT 641.100 813.150 642.900 814.950 ;
        RECT 640.950 811.050 643.050 813.150 ;
        RECT 643.950 812.850 646.350 814.950 ;
        RECT 658.950 812.850 661.050 814.950 ;
        RECT 661.950 814.050 664.050 816.150 ;
        RECT 665.850 814.950 667.050 818.250 ;
        RECT 686.100 816.150 687.900 817.950 ;
        RECT 664.950 812.850 667.050 814.950 ;
        RECT 682.950 812.850 685.050 814.950 ;
        RECT 685.950 814.050 688.050 816.150 ;
        RECT 689.850 814.950 691.050 818.250 ;
        RECT 707.100 816.150 708.900 817.950 ;
        RECT 688.950 812.850 691.050 814.950 ;
        RECT 703.950 812.850 706.050 814.950 ;
        RECT 706.950 814.050 709.050 816.150 ;
        RECT 710.850 814.950 712.050 818.250 ;
        RECT 709.950 812.850 712.050 814.950 ;
        RECT 728.100 813.150 729.900 814.950 ;
        RECT 645.150 807.600 646.350 812.850 ;
        RECT 659.100 811.050 660.900 812.850 ;
        RECT 664.950 807.600 666.150 812.850 ;
        RECT 667.950 809.850 670.050 811.950 ;
        RECT 683.100 811.050 684.900 812.850 ;
        RECT 667.950 808.050 669.750 809.850 ;
        RECT 688.950 807.600 690.150 812.850 ;
        RECT 691.950 809.850 694.050 811.950 ;
        RECT 704.100 811.050 705.900 812.850 ;
        RECT 691.950 808.050 693.750 809.850 ;
        RECT 709.950 807.600 711.150 812.850 ;
        RECT 712.950 809.850 715.050 811.950 ;
        RECT 727.950 811.050 730.050 813.150 ;
        RECT 731.250 811.950 732.450 819.300 ;
        RECT 734.100 813.150 735.900 814.950 ;
        RECT 730.950 809.850 733.050 811.950 ;
        RECT 733.950 811.050 736.050 813.150 ;
        RECT 712.950 808.050 714.750 809.850 ;
        RECT 635.550 795.750 637.350 801.600 ;
        RECT 638.550 795.750 640.350 801.600 ;
        RECT 642.150 795.750 643.950 807.600 ;
        RECT 645.150 795.750 646.950 807.600 ;
        RECT 660.300 795.750 662.100 807.600 ;
        RECT 664.500 795.750 666.300 807.600 ;
        RECT 667.800 795.750 669.600 801.600 ;
        RECT 684.300 795.750 686.100 807.600 ;
        RECT 688.500 795.750 690.300 807.600 ;
        RECT 691.800 795.750 693.600 801.600 ;
        RECT 705.300 795.750 707.100 807.600 ;
        RECT 709.500 795.750 711.300 807.600 ;
        RECT 731.250 801.600 732.450 809.850 ;
        RECT 738.150 808.800 739.050 821.400 ;
        RECT 746.550 820.800 748.350 822.600 ;
        RECT 749.850 821.550 754.800 822.600 ;
        RECT 762.300 823.500 763.350 824.400 ;
        RECT 762.300 822.300 766.050 823.500 ;
        RECT 749.850 820.800 751.650 821.550 ;
        RECT 746.850 819.900 747.900 820.800 ;
        RECT 757.050 820.200 758.850 822.000 ;
        RECT 763.950 821.400 766.050 822.300 ;
        RECT 769.650 821.400 771.450 827.250 ;
        RECT 779.550 824.400 781.350 827.250 ;
        RECT 782.550 824.400 784.350 827.250 ;
        RECT 794.550 824.400 796.350 827.250 ;
        RECT 797.550 824.400 799.350 827.250 ;
        RECT 814.650 824.400 816.450 827.250 ;
        RECT 817.650 824.400 819.450 827.250 ;
        RECT 820.650 824.400 822.450 827.250 ;
        RECT 757.050 819.900 757.950 820.200 ;
        RECT 746.850 819.000 757.950 819.900 ;
        RECT 770.250 819.150 771.450 821.400 ;
        RECT 746.850 817.800 747.900 819.000 ;
        RECT 741.000 816.600 747.900 817.800 ;
        RECT 741.000 815.850 741.900 816.600 ;
        RECT 746.100 816.000 747.900 816.600 ;
        RECT 740.100 814.050 741.900 815.850 ;
        RECT 743.100 814.950 744.900 815.700 ;
        RECT 757.050 814.950 757.950 819.000 ;
        RECT 766.950 817.050 771.450 819.150 ;
        RECT 765.150 815.250 769.050 817.050 ;
        RECT 766.950 814.950 769.050 815.250 ;
        RECT 743.100 813.900 751.050 814.950 ;
        RECT 748.950 812.850 751.050 813.900 ;
        RECT 754.950 812.850 757.950 814.950 ;
        RECT 747.450 809.100 749.250 809.400 ;
        RECT 747.450 808.800 755.850 809.100 ;
        RECT 738.150 808.200 755.850 808.800 ;
        RECT 738.150 807.600 749.250 808.200 ;
        RECT 712.800 795.750 714.600 801.600 ;
        RECT 727.650 795.750 729.450 801.600 ;
        RECT 730.650 795.750 732.450 801.600 ;
        RECT 733.650 795.750 735.450 801.600 ;
        RECT 738.150 795.750 739.950 807.600 ;
        RECT 752.250 806.700 754.050 807.300 ;
        RECT 746.550 805.500 754.050 806.700 ;
        RECT 754.950 806.100 755.850 808.200 ;
        RECT 757.050 808.200 757.950 812.850 ;
        RECT 767.250 809.400 769.050 811.200 ;
        RECT 763.950 808.200 768.150 809.400 ;
        RECT 757.050 807.300 763.050 808.200 ;
        RECT 763.950 807.300 766.050 808.200 ;
        RECT 770.250 807.600 771.450 817.050 ;
        RECT 778.950 815.850 781.050 817.950 ;
        RECT 782.400 816.150 783.600 824.400 ;
        RECT 779.100 814.050 780.900 815.850 ;
        RECT 781.950 814.050 784.050 816.150 ;
        RECT 793.950 815.850 796.050 817.950 ;
        RECT 797.400 816.150 798.600 824.400 ;
        RECT 817.950 817.950 819.000 824.400 ;
        RECT 830.850 821.400 832.650 827.250 ;
        RECT 835.350 820.200 837.150 827.250 ;
        RECT 851.550 824.400 853.350 827.250 ;
        RECT 833.550 819.300 837.150 820.200 ;
        RECT 852.150 820.500 853.350 824.400 ;
        RECT 854.850 821.400 856.650 827.250 ;
        RECT 857.850 821.400 859.650 827.250 ;
        RECT 872.550 821.400 874.350 827.250 ;
        RECT 875.550 821.400 877.350 827.250 ;
        RECT 852.150 819.600 857.250 820.500 ;
        RECT 794.100 814.050 795.900 815.850 ;
        RECT 796.950 814.050 799.050 816.150 ;
        RECT 817.950 815.850 820.050 817.950 ;
        RECT 762.150 806.400 763.050 807.300 ;
        RECT 759.450 806.100 761.250 806.400 ;
        RECT 746.550 804.600 747.750 805.500 ;
        RECT 754.950 805.200 761.250 806.100 ;
        RECT 759.450 804.600 761.250 805.200 ;
        RECT 762.150 804.600 764.850 806.400 ;
        RECT 742.950 802.500 747.750 804.600 ;
        RECT 750.150 802.500 757.050 804.300 ;
        RECT 746.550 801.600 747.750 802.500 ;
        RECT 741.150 795.750 742.950 801.600 ;
        RECT 746.250 795.750 748.050 801.600 ;
        RECT 751.050 795.750 752.850 801.600 ;
        RECT 754.050 795.750 755.850 802.500 ;
        RECT 762.150 801.600 766.050 803.700 ;
        RECT 757.950 795.750 759.750 801.600 ;
        RECT 762.150 795.750 763.950 801.600 ;
        RECT 766.650 795.750 768.450 798.600 ;
        RECT 769.650 795.750 771.450 807.600 ;
        RECT 782.400 801.600 783.600 814.050 ;
        RECT 797.400 801.600 798.600 814.050 ;
        RECT 814.950 812.850 817.050 814.950 ;
        RECT 815.100 811.050 816.900 812.850 ;
        RECT 817.950 808.650 819.000 815.850 ;
        RECT 820.950 812.850 823.050 814.950 ;
        RECT 830.100 813.150 831.900 814.950 ;
        RECT 821.100 811.050 822.900 812.850 ;
        RECT 829.950 811.050 832.050 813.150 ;
        RECT 833.550 811.950 834.750 819.300 ;
        RECT 855.000 818.700 857.250 819.600 ;
        RECT 836.100 813.150 837.900 814.950 ;
        RECT 832.950 809.850 835.050 811.950 ;
        RECT 835.950 811.050 838.050 813.150 ;
        RECT 850.950 812.850 853.050 814.950 ;
        RECT 851.100 811.050 852.900 812.850 ;
        RECT 855.000 810.300 856.050 818.700 ;
        RECT 858.150 814.950 859.350 821.400 ;
        RECT 872.100 816.150 873.900 817.950 ;
        RECT 856.950 812.850 859.350 814.950 ;
        RECT 871.950 814.050 874.050 816.150 ;
        RECT 875.400 814.950 876.600 821.400 ;
        RECT 874.950 812.850 877.050 814.950 ;
        RECT 816.450 807.600 819.000 808.650 ;
        RECT 779.550 795.750 781.350 801.600 ;
        RECT 782.550 795.750 784.350 801.600 ;
        RECT 794.550 795.750 796.350 801.600 ;
        RECT 797.550 795.750 799.350 801.600 ;
        RECT 816.450 795.750 818.250 807.600 ;
        RECT 820.650 795.750 822.450 807.600 ;
        RECT 833.550 801.600 834.750 809.850 ;
        RECT 855.000 809.400 857.250 810.300 ;
        RECT 851.550 808.500 857.250 809.400 ;
        RECT 851.550 801.600 852.750 808.500 ;
        RECT 858.150 807.600 859.350 812.850 ;
        RECT 875.400 807.600 876.600 812.850 ;
        RECT 830.550 795.750 832.350 801.600 ;
        RECT 833.550 795.750 835.350 801.600 ;
        RECT 836.550 795.750 838.350 801.600 ;
        RECT 851.550 795.750 853.350 801.600 ;
        RECT 854.850 795.750 856.650 807.600 ;
        RECT 857.850 795.750 859.650 807.600 ;
        RECT 872.550 795.750 874.350 807.600 ;
        RECT 875.550 795.750 877.350 807.600 ;
        RECT 13.650 785.400 15.450 791.250 ;
        RECT 16.650 785.400 18.450 791.250 ;
        RECT 19.650 785.400 21.450 791.250 ;
        RECT 17.250 777.150 18.450 785.400 ;
        RECT 33.150 780.900 34.950 791.250 ;
        RECT 32.550 779.550 34.950 780.900 ;
        RECT 36.150 779.550 37.950 791.250 ;
        RECT 13.950 773.850 16.050 775.950 ;
        RECT 16.950 775.050 19.050 777.150 ;
        RECT 14.100 772.050 15.900 773.850 ;
        RECT 17.250 767.700 18.450 775.050 ;
        RECT 19.950 773.850 22.050 775.950 ;
        RECT 20.100 772.050 21.900 773.850 ;
        RECT 32.550 772.950 33.900 779.550 ;
        RECT 40.650 779.400 42.450 791.250 ;
        RECT 53.550 785.400 55.350 791.250 ;
        RECT 56.550 785.400 58.350 791.250 ;
        RECT 35.250 778.200 37.050 778.650 ;
        RECT 41.250 778.200 42.450 779.400 ;
        RECT 35.250 777.000 42.450 778.200 ;
        RECT 35.250 776.850 37.050 777.000 ;
        RECT 14.850 766.800 18.450 767.700 ;
        RECT 31.950 770.850 34.050 772.950 ;
        RECT 14.850 759.750 16.650 766.800 ;
        RECT 31.950 765.600 33.000 770.850 ;
        RECT 35.400 768.600 36.300 776.850 ;
        RECT 38.100 774.150 39.900 775.950 ;
        RECT 37.950 772.050 40.050 774.150 ;
        RECT 56.400 772.950 57.600 785.400 ;
        RECT 70.650 779.400 72.450 791.250 ;
        RECT 73.650 780.300 75.450 791.250 ;
        RECT 76.650 781.200 78.450 791.250 ;
        RECT 79.650 780.300 81.450 791.250 ;
        RECT 73.650 779.400 81.450 780.300 ;
        RECT 89.550 780.300 91.350 791.250 ;
        RECT 92.550 781.200 94.350 791.250 ;
        RECT 95.550 780.300 97.350 791.250 ;
        RECT 89.550 779.400 97.350 780.300 ;
        RECT 98.550 779.400 100.350 791.250 ;
        RECT 110.550 785.400 112.350 791.250 ;
        RECT 113.550 785.400 115.350 791.250 ;
        RECT 116.550 786.000 118.350 791.250 ;
        RECT 113.700 785.100 115.350 785.400 ;
        RECT 119.550 785.400 121.350 791.250 ;
        RECT 119.550 785.100 120.750 785.400 ;
        RECT 113.700 784.200 120.750 785.100 ;
        RECT 113.100 780.150 114.900 781.950 ;
        RECT 71.100 774.150 72.300 779.400 ;
        RECT 98.700 774.150 99.900 779.400 ;
        RECT 110.100 777.150 111.900 778.950 ;
        RECT 112.950 778.050 115.050 780.150 ;
        RECT 116.250 777.150 118.050 778.950 ;
        RECT 109.950 775.050 112.050 777.150 ;
        RECT 115.950 775.050 118.050 777.150 ;
        RECT 119.700 775.950 120.750 784.200 ;
        RECT 131.550 779.400 133.350 791.250 ;
        RECT 135.750 779.400 137.550 791.250 ;
        RECT 135.000 778.350 137.550 779.400 ;
        RECT 149.550 779.400 151.350 791.250 ;
        RECT 154.050 779.550 155.850 791.250 ;
        RECT 157.050 780.900 158.850 791.250 ;
        RECT 157.050 779.550 159.450 780.900 ;
        RECT 41.100 771.150 42.900 772.950 ;
        RECT 53.100 771.150 54.900 772.950 ;
        RECT 40.950 769.050 43.050 771.150 ;
        RECT 52.950 769.050 55.050 771.150 ;
        RECT 55.950 770.850 58.050 772.950 ;
        RECT 70.950 772.050 73.050 774.150 ;
        RECT 35.250 767.700 37.050 768.600 ;
        RECT 35.250 766.800 38.550 767.700 ;
        RECT 19.350 759.750 21.150 765.600 ;
        RECT 31.650 759.750 33.450 765.600 ;
        RECT 37.650 762.600 38.550 766.800 ;
        RECT 56.400 762.600 57.600 770.850 ;
        RECT 71.100 765.600 72.300 772.050 ;
        RECT 73.950 770.850 76.050 772.950 ;
        RECT 77.100 771.150 78.900 772.950 ;
        RECT 74.100 769.050 75.900 770.850 ;
        RECT 76.950 769.050 79.050 771.150 ;
        RECT 79.950 770.850 82.050 772.950 ;
        RECT 88.950 770.850 91.050 772.950 ;
        RECT 92.100 771.150 93.900 772.950 ;
        RECT 80.100 769.050 81.900 770.850 ;
        RECT 89.100 769.050 90.900 770.850 ;
        RECT 91.950 769.050 94.050 771.150 ;
        RECT 94.950 770.850 97.050 772.950 ;
        RECT 97.950 772.050 100.050 774.150 ;
        RECT 118.950 773.850 121.050 775.950 ;
        RECT 131.100 774.150 132.900 775.950 ;
        RECT 95.100 769.050 96.900 770.850 ;
        RECT 98.700 765.600 99.900 772.050 ;
        RECT 119.400 769.650 120.600 773.850 ;
        RECT 130.950 772.050 133.050 774.150 ;
        RECT 135.000 771.150 136.050 778.350 ;
        RECT 149.550 778.200 150.750 779.400 ;
        RECT 154.950 778.200 156.750 778.650 ;
        RECT 149.550 777.000 156.750 778.200 ;
        RECT 154.950 776.850 156.750 777.000 ;
        RECT 137.100 774.150 138.900 775.950 ;
        RECT 152.100 774.150 153.900 775.950 ;
        RECT 136.950 772.050 139.050 774.150 ;
        RECT 149.100 771.150 150.900 772.950 ;
        RECT 151.950 772.050 154.050 774.150 ;
        RECT 71.100 763.950 76.800 765.600 ;
        RECT 34.650 759.750 36.450 762.600 ;
        RECT 37.650 759.750 39.450 762.600 ;
        RECT 40.650 759.750 42.450 762.600 ;
        RECT 53.550 759.750 55.350 762.600 ;
        RECT 56.550 759.750 58.350 762.600 ;
        RECT 71.700 759.750 73.500 762.600 ;
        RECT 75.000 759.750 76.800 763.950 ;
        RECT 79.200 759.750 81.000 765.600 ;
        RECT 90.000 759.750 91.800 765.600 ;
        RECT 94.200 763.950 99.900 765.600 ;
        RECT 94.200 759.750 96.000 763.950 ;
        RECT 97.500 759.750 99.300 762.600 ;
        RECT 110.700 759.750 112.500 768.600 ;
        RECT 116.100 768.000 120.600 769.650 ;
        RECT 133.950 769.050 136.050 771.150 ;
        RECT 148.950 769.050 151.050 771.150 ;
        RECT 116.100 759.750 117.900 768.000 ;
        RECT 135.000 762.600 136.050 769.050 ;
        RECT 155.700 768.600 156.600 776.850 ;
        RECT 158.100 772.950 159.450 779.550 ;
        RECT 170.550 780.300 172.350 791.250 ;
        RECT 173.550 781.200 175.350 791.250 ;
        RECT 176.550 780.300 178.350 791.250 ;
        RECT 170.550 779.400 178.350 780.300 ;
        RECT 179.550 779.400 181.350 791.250 ;
        RECT 194.550 779.400 196.350 791.250 ;
        RECT 198.750 779.400 200.550 791.250 ;
        RECT 213.300 779.400 215.100 791.250 ;
        RECT 217.500 779.400 219.300 791.250 ;
        RECT 220.800 785.400 222.600 791.250 ;
        RECT 235.650 785.400 237.450 791.250 ;
        RECT 238.650 785.400 240.450 791.250 ;
        RECT 241.650 785.400 243.450 791.250 ;
        RECT 254.550 785.400 256.350 791.250 ;
        RECT 257.550 785.400 259.350 791.250 ;
        RECT 272.400 785.400 274.200 791.250 ;
        RECT 179.700 774.150 180.900 779.400 ;
        RECT 198.000 778.350 200.550 779.400 ;
        RECT 194.100 774.150 195.900 775.950 ;
        RECT 157.950 770.850 160.050 772.950 ;
        RECT 169.950 770.850 172.050 772.950 ;
        RECT 173.100 771.150 174.900 772.950 ;
        RECT 154.950 767.700 156.750 768.600 ;
        RECT 153.450 766.800 156.750 767.700 ;
        RECT 153.450 762.600 154.350 766.800 ;
        RECT 159.000 765.600 160.050 770.850 ;
        RECT 170.100 769.050 171.900 770.850 ;
        RECT 172.950 769.050 175.050 771.150 ;
        RECT 175.950 770.850 178.050 772.950 ;
        RECT 178.950 772.050 181.050 774.150 ;
        RECT 193.950 772.050 196.050 774.150 ;
        RECT 176.100 769.050 177.900 770.850 ;
        RECT 179.700 765.600 180.900 772.050 ;
        RECT 198.000 771.150 199.050 778.350 ;
        RECT 200.100 774.150 201.900 775.950 ;
        RECT 212.100 774.150 213.900 775.950 ;
        RECT 217.950 774.150 219.150 779.400 ;
        RECT 220.950 777.150 222.750 778.950 ;
        RECT 239.250 777.150 240.450 785.400 ;
        RECT 220.950 775.050 223.050 777.150 ;
        RECT 199.950 772.050 202.050 774.150 ;
        RECT 211.950 772.050 214.050 774.150 ;
        RECT 196.950 769.050 199.050 771.150 ;
        RECT 214.950 770.850 217.050 772.950 ;
        RECT 217.950 772.050 220.050 774.150 ;
        RECT 235.950 773.850 238.050 775.950 ;
        RECT 238.950 775.050 241.050 777.150 ;
        RECT 236.100 772.050 237.900 773.850 ;
        RECT 215.100 769.050 216.900 770.850 ;
        RECT 131.550 759.750 133.350 762.600 ;
        RECT 134.550 759.750 136.350 762.600 ;
        RECT 137.550 759.750 139.350 762.600 ;
        RECT 149.550 759.750 151.350 762.600 ;
        RECT 152.550 759.750 154.350 762.600 ;
        RECT 155.550 759.750 157.350 762.600 ;
        RECT 158.550 759.750 160.350 765.600 ;
        RECT 171.000 759.750 172.800 765.600 ;
        RECT 175.200 763.950 180.900 765.600 ;
        RECT 175.200 759.750 177.000 763.950 ;
        RECT 198.000 762.600 199.050 769.050 ;
        RECT 218.850 768.750 220.050 772.050 ;
        RECT 219.000 767.700 222.750 768.750 ;
        RECT 239.250 767.700 240.450 775.050 ;
        RECT 241.950 773.850 244.050 775.950 ;
        RECT 242.100 772.050 243.900 773.850 ;
        RECT 257.400 772.950 258.600 785.400 ;
        RECT 275.700 779.400 277.500 791.250 ;
        RECT 279.900 779.400 281.700 791.250 ;
        RECT 290.550 785.400 292.350 791.250 ;
        RECT 293.550 785.400 295.350 791.250 ;
        RECT 272.250 777.150 274.050 778.950 ;
        RECT 271.950 775.050 274.050 777.150 ;
        RECT 275.850 774.150 277.050 779.400 ;
        RECT 281.100 774.150 282.900 775.950 ;
        RECT 290.100 774.150 291.900 775.950 ;
        RECT 254.100 771.150 255.900 772.950 ;
        RECT 253.950 769.050 256.050 771.150 ;
        RECT 256.950 770.850 259.050 772.950 ;
        RECT 274.950 772.050 277.050 774.150 ;
        RECT 212.550 764.700 220.350 766.050 ;
        RECT 178.500 759.750 180.300 762.600 ;
        RECT 194.550 759.750 196.350 762.600 ;
        RECT 197.550 759.750 199.350 762.600 ;
        RECT 200.550 759.750 202.350 762.600 ;
        RECT 212.550 759.750 214.350 764.700 ;
        RECT 215.550 759.750 217.350 763.800 ;
        RECT 218.550 759.750 220.350 764.700 ;
        RECT 221.550 765.600 222.750 767.700 ;
        RECT 236.850 766.800 240.450 767.700 ;
        RECT 221.550 759.750 223.350 765.600 ;
        RECT 236.850 759.750 238.650 766.800 ;
        RECT 241.350 759.750 243.150 765.600 ;
        RECT 257.400 762.600 258.600 770.850 ;
        RECT 274.950 768.750 276.150 772.050 ;
        RECT 277.950 770.850 280.050 772.950 ;
        RECT 280.950 772.050 283.050 774.150 ;
        RECT 289.950 772.050 292.050 774.150 ;
        RECT 278.100 769.050 279.900 770.850 ;
        RECT 272.250 767.700 276.000 768.750 ;
        RECT 293.700 768.300 294.900 785.400 ;
        RECT 297.150 779.400 298.950 791.250 ;
        RECT 300.150 779.400 301.950 791.250 ;
        RECT 313.650 779.400 315.450 791.250 ;
        RECT 295.950 773.850 298.050 775.950 ;
        RECT 300.150 774.150 301.350 779.400 ;
        RECT 316.650 778.500 318.450 791.250 ;
        RECT 319.650 779.400 321.450 791.250 ;
        RECT 322.650 778.500 324.450 791.250 ;
        RECT 325.650 779.400 327.450 791.250 ;
        RECT 328.650 778.500 330.450 791.250 ;
        RECT 331.650 779.400 333.450 791.250 ;
        RECT 334.650 778.500 336.450 791.250 ;
        RECT 337.650 779.400 339.450 791.250 ;
        RECT 352.350 779.400 354.150 791.250 ;
        RECT 355.350 779.400 357.150 791.250 ;
        RECT 358.650 785.400 360.450 791.250 ;
        RECT 371.550 785.400 373.350 791.250 ;
        RECT 374.550 785.400 376.350 791.250 ;
        RECT 392.400 785.400 394.200 791.250 ;
        RECT 296.100 772.050 297.900 773.850 ;
        RECT 298.950 772.050 301.350 774.150 ;
        RECT 315.750 777.300 318.450 778.500 ;
        RECT 320.700 777.300 324.450 778.500 ;
        RECT 326.700 777.300 330.450 778.500 ;
        RECT 332.550 777.300 336.450 778.500 ;
        RECT 315.750 772.950 316.800 777.300 ;
        RECT 272.250 765.600 273.450 767.700 ;
        RECT 290.550 767.100 298.050 768.300 ;
        RECT 254.550 759.750 256.350 762.600 ;
        RECT 257.550 759.750 259.350 762.600 ;
        RECT 271.650 759.750 273.450 765.600 ;
        RECT 274.650 764.700 282.450 766.050 ;
        RECT 274.650 759.750 276.450 764.700 ;
        RECT 277.650 759.750 279.450 763.800 ;
        RECT 280.650 759.750 282.450 764.700 ;
        RECT 290.550 759.750 292.350 767.100 ;
        RECT 296.250 766.500 298.050 767.100 ;
        RECT 300.150 765.600 301.350 772.050 ;
        RECT 313.950 770.850 316.800 772.950 ;
        RECT 315.750 767.700 316.800 770.850 ;
        RECT 320.700 770.400 321.900 777.300 ;
        RECT 326.700 770.400 327.900 777.300 ;
        RECT 332.550 770.400 333.750 777.300 ;
        RECT 352.650 774.150 353.850 779.400 ;
        RECT 359.250 778.500 360.450 785.400 ;
        RECT 354.750 777.600 360.450 778.500 ;
        RECT 354.750 776.700 357.000 777.600 ;
        RECT 334.950 770.850 337.050 772.950 ;
        RECT 352.650 772.050 355.050 774.150 ;
        RECT 317.700 768.600 321.900 770.400 ;
        RECT 323.700 768.600 327.900 770.400 ;
        RECT 329.700 768.600 333.750 770.400 ;
        RECT 335.100 769.050 336.900 770.850 ;
        RECT 320.700 767.700 321.900 768.600 ;
        RECT 326.700 767.700 327.900 768.600 ;
        RECT 332.550 767.700 333.750 768.600 ;
        RECT 315.750 766.650 318.600 767.700 ;
        RECT 315.900 766.500 318.600 766.650 ;
        RECT 320.700 766.500 324.600 767.700 ;
        RECT 326.700 766.500 330.450 767.700 ;
        RECT 332.550 766.500 336.600 767.700 ;
        RECT 316.800 765.600 318.600 766.500 ;
        RECT 322.800 765.600 324.600 766.500 ;
        RECT 295.050 759.750 296.850 765.600 ;
        RECT 298.050 764.100 301.350 765.600 ;
        RECT 298.050 759.750 299.850 764.100 ;
        RECT 313.650 759.750 315.450 765.600 ;
        RECT 316.650 759.750 318.450 765.600 ;
        RECT 319.650 759.750 321.450 765.600 ;
        RECT 322.650 759.750 324.450 765.600 ;
        RECT 325.650 759.750 327.450 765.600 ;
        RECT 328.650 759.750 330.450 766.500 ;
        RECT 334.800 765.600 336.600 766.500 ;
        RECT 352.650 765.600 353.850 772.050 ;
        RECT 355.950 768.300 357.000 776.700 ;
        RECT 359.100 774.150 360.900 775.950 ;
        RECT 358.950 772.050 361.050 774.150 ;
        RECT 374.400 772.950 375.600 785.400 ;
        RECT 395.700 779.400 397.500 791.250 ;
        RECT 399.900 779.400 401.700 791.250 ;
        RECT 410.550 779.400 412.350 791.250 ;
        RECT 414.750 779.400 416.550 791.250 ;
        RECT 433.650 785.400 435.450 791.250 ;
        RECT 436.650 785.400 438.450 791.250 ;
        RECT 439.650 785.400 441.450 791.250 ;
        RECT 392.250 777.150 394.050 778.950 ;
        RECT 391.950 775.050 394.050 777.150 ;
        RECT 395.850 774.150 397.050 779.400 ;
        RECT 414.000 778.350 416.550 779.400 ;
        RECT 401.100 774.150 402.900 775.950 ;
        RECT 410.100 774.150 411.900 775.950 ;
        RECT 371.100 771.150 372.900 772.950 ;
        RECT 370.950 769.050 373.050 771.150 ;
        RECT 373.950 770.850 376.050 772.950 ;
        RECT 394.950 772.050 397.050 774.150 ;
        RECT 354.750 767.400 357.000 768.300 ;
        RECT 354.750 766.500 359.850 767.400 ;
        RECT 331.650 759.750 333.450 765.600 ;
        RECT 334.650 759.750 336.450 765.600 ;
        RECT 337.650 759.750 339.450 765.600 ;
        RECT 352.350 759.750 354.150 765.600 ;
        RECT 355.350 759.750 357.150 765.600 ;
        RECT 358.650 762.600 359.850 766.500 ;
        RECT 374.400 762.600 375.600 770.850 ;
        RECT 394.950 768.750 396.150 772.050 ;
        RECT 397.950 770.850 400.050 772.950 ;
        RECT 400.950 772.050 403.050 774.150 ;
        RECT 409.950 772.050 412.050 774.150 ;
        RECT 414.000 771.150 415.050 778.350 ;
        RECT 437.250 777.150 438.450 785.400 ;
        RECT 450.300 779.400 452.100 791.250 ;
        RECT 454.500 779.400 456.300 791.250 ;
        RECT 457.800 785.400 459.600 791.250 ;
        RECT 472.650 785.400 474.450 791.250 ;
        RECT 475.650 785.400 477.450 791.250 ;
        RECT 416.100 774.150 417.900 775.950 ;
        RECT 415.950 772.050 418.050 774.150 ;
        RECT 433.950 773.850 436.050 775.950 ;
        RECT 436.950 775.050 439.050 777.150 ;
        RECT 434.100 772.050 435.900 773.850 ;
        RECT 398.100 769.050 399.900 770.850 ;
        RECT 412.950 769.050 415.050 771.150 ;
        RECT 392.250 767.700 396.000 768.750 ;
        RECT 392.250 765.600 393.450 767.700 ;
        RECT 358.650 759.750 360.450 762.600 ;
        RECT 371.550 759.750 373.350 762.600 ;
        RECT 374.550 759.750 376.350 762.600 ;
        RECT 391.650 759.750 393.450 765.600 ;
        RECT 394.650 764.700 402.450 766.050 ;
        RECT 394.650 759.750 396.450 764.700 ;
        RECT 397.650 759.750 399.450 763.800 ;
        RECT 400.650 759.750 402.450 764.700 ;
        RECT 414.000 762.600 415.050 769.050 ;
        RECT 437.250 767.700 438.450 775.050 ;
        RECT 439.950 773.850 442.050 775.950 ;
        RECT 449.100 774.150 450.900 775.950 ;
        RECT 454.950 774.150 456.150 779.400 ;
        RECT 457.950 777.150 459.750 778.950 ;
        RECT 457.950 775.050 460.050 777.150 ;
        RECT 440.100 772.050 441.900 773.850 ;
        RECT 448.950 772.050 451.050 774.150 ;
        RECT 451.950 770.850 454.050 772.950 ;
        RECT 454.950 772.050 457.050 774.150 ;
        RECT 473.400 772.950 474.600 785.400 ;
        RECT 492.150 780.900 493.950 791.250 ;
        RECT 491.550 779.550 493.950 780.900 ;
        RECT 495.150 779.550 496.950 791.250 ;
        RECT 491.550 772.950 492.900 779.550 ;
        RECT 499.650 779.400 501.450 791.250 ;
        RECT 514.650 785.400 516.450 791.250 ;
        RECT 517.650 785.400 519.450 791.250 ;
        RECT 529.650 785.400 531.450 791.250 ;
        RECT 532.650 785.400 534.450 791.250 ;
        RECT 494.250 778.200 496.050 778.650 ;
        RECT 500.250 778.200 501.450 779.400 ;
        RECT 494.250 777.000 501.450 778.200 ;
        RECT 494.250 776.850 496.050 777.000 ;
        RECT 452.100 769.050 453.900 770.850 ;
        RECT 455.850 768.750 457.050 772.050 ;
        RECT 472.950 770.850 475.050 772.950 ;
        RECT 476.100 771.150 477.900 772.950 ;
        RECT 456.000 767.700 459.750 768.750 ;
        RECT 434.850 766.800 438.450 767.700 ;
        RECT 410.550 759.750 412.350 762.600 ;
        RECT 413.550 759.750 415.350 762.600 ;
        RECT 416.550 759.750 418.350 762.600 ;
        RECT 434.850 759.750 436.650 766.800 ;
        RECT 439.350 759.750 441.150 765.600 ;
        RECT 449.550 764.700 457.350 766.050 ;
        RECT 449.550 759.750 451.350 764.700 ;
        RECT 452.550 759.750 454.350 763.800 ;
        RECT 455.550 759.750 457.350 764.700 ;
        RECT 458.550 765.600 459.750 767.700 ;
        RECT 458.550 759.750 460.350 765.600 ;
        RECT 473.400 762.600 474.600 770.850 ;
        RECT 475.950 769.050 478.050 771.150 ;
        RECT 490.950 770.850 493.050 772.950 ;
        RECT 490.950 765.600 492.000 770.850 ;
        RECT 494.400 768.600 495.300 776.850 ;
        RECT 497.100 774.150 498.900 775.950 ;
        RECT 496.950 772.050 499.050 774.150 ;
        RECT 515.400 772.950 516.600 785.400 ;
        RECT 530.400 772.950 531.600 785.400 ;
        RECT 536.550 779.400 538.350 791.250 ;
        RECT 539.550 788.400 541.350 791.250 ;
        RECT 544.050 785.400 545.850 791.250 ;
        RECT 548.250 785.400 550.050 791.250 ;
        RECT 541.950 783.300 545.850 785.400 ;
        RECT 552.150 784.500 553.950 791.250 ;
        RECT 555.150 785.400 556.950 791.250 ;
        RECT 559.950 785.400 561.750 791.250 ;
        RECT 565.050 785.400 566.850 791.250 ;
        RECT 560.250 784.500 561.450 785.400 ;
        RECT 550.950 782.700 557.850 784.500 ;
        RECT 560.250 782.400 565.050 784.500 ;
        RECT 543.150 780.600 545.850 782.400 ;
        RECT 546.750 781.800 548.550 782.400 ;
        RECT 546.750 780.900 553.050 781.800 ;
        RECT 560.250 781.500 561.450 782.400 ;
        RECT 546.750 780.600 548.550 780.900 ;
        RECT 544.950 779.700 545.850 780.600 ;
        RECT 500.100 771.150 501.900 772.950 ;
        RECT 499.950 769.050 502.050 771.150 ;
        RECT 514.950 770.850 517.050 772.950 ;
        RECT 518.100 771.150 519.900 772.950 ;
        RECT 494.250 767.700 496.050 768.600 ;
        RECT 494.250 766.800 497.550 767.700 ;
        RECT 472.650 759.750 474.450 762.600 ;
        RECT 475.650 759.750 477.450 762.600 ;
        RECT 490.650 759.750 492.450 765.600 ;
        RECT 496.650 762.600 497.550 766.800 ;
        RECT 515.400 762.600 516.600 770.850 ;
        RECT 517.950 769.050 520.050 771.150 ;
        RECT 529.950 770.850 532.050 772.950 ;
        RECT 533.100 771.150 534.900 772.950 ;
        RECT 530.400 762.600 531.600 770.850 ;
        RECT 532.950 769.050 535.050 771.150 ;
        RECT 536.550 769.950 537.750 779.400 ;
        RECT 541.950 778.800 544.050 779.700 ;
        RECT 544.950 778.800 550.950 779.700 ;
        RECT 539.850 777.600 544.050 778.800 ;
        RECT 538.950 775.800 540.750 777.600 ;
        RECT 550.050 774.150 550.950 778.800 ;
        RECT 552.150 778.800 553.050 780.900 ;
        RECT 553.950 780.300 561.450 781.500 ;
        RECT 553.950 779.700 555.750 780.300 ;
        RECT 568.050 779.400 569.850 791.250 ;
        RECT 578.550 785.400 580.350 791.250 ;
        RECT 581.550 785.400 583.350 791.250 ;
        RECT 584.550 785.400 586.350 791.250 ;
        RECT 598.650 785.400 600.450 791.250 ;
        RECT 601.650 785.400 603.450 791.250 ;
        RECT 614.550 785.400 616.350 791.250 ;
        RECT 617.550 785.400 619.350 791.250 ;
        RECT 629.550 785.400 631.350 791.250 ;
        RECT 632.550 785.400 634.350 791.250 ;
        RECT 635.550 785.400 637.350 791.250 ;
        RECT 558.750 778.800 569.850 779.400 ;
        RECT 552.150 778.200 569.850 778.800 ;
        RECT 552.150 777.900 560.550 778.200 ;
        RECT 558.750 777.600 560.550 777.900 ;
        RECT 550.050 772.050 553.050 774.150 ;
        RECT 556.950 773.100 559.050 774.150 ;
        RECT 556.950 772.050 564.900 773.100 ;
        RECT 538.950 771.750 541.050 772.050 ;
        RECT 538.950 769.950 542.850 771.750 ;
        RECT 536.550 767.850 541.050 769.950 ;
        RECT 550.050 768.000 550.950 772.050 ;
        RECT 563.100 771.300 564.900 772.050 ;
        RECT 566.100 771.150 567.900 772.950 ;
        RECT 560.100 770.400 561.900 771.000 ;
        RECT 566.100 770.400 567.000 771.150 ;
        RECT 560.100 769.200 567.000 770.400 ;
        RECT 560.100 768.000 561.150 769.200 ;
        RECT 536.550 765.600 537.750 767.850 ;
        RECT 550.050 767.100 561.150 768.000 ;
        RECT 550.050 766.800 550.950 767.100 ;
        RECT 493.650 759.750 495.450 762.600 ;
        RECT 496.650 759.750 498.450 762.600 ;
        RECT 499.650 759.750 501.450 762.600 ;
        RECT 514.650 759.750 516.450 762.600 ;
        RECT 517.650 759.750 519.450 762.600 ;
        RECT 529.650 759.750 531.450 762.600 ;
        RECT 532.650 759.750 534.450 762.600 ;
        RECT 536.550 759.750 538.350 765.600 ;
        RECT 541.950 764.700 544.050 765.600 ;
        RECT 549.150 765.000 550.950 766.800 ;
        RECT 560.100 766.200 561.150 767.100 ;
        RECT 556.350 765.450 558.150 766.200 ;
        RECT 541.950 763.500 545.700 764.700 ;
        RECT 544.650 762.600 545.700 763.500 ;
        RECT 553.200 764.400 558.150 765.450 ;
        RECT 559.650 764.400 561.450 766.200 ;
        RECT 568.950 765.600 569.850 778.200 ;
        RECT 581.550 777.150 582.750 785.400 ;
        RECT 577.950 773.850 580.050 775.950 ;
        RECT 580.950 775.050 583.050 777.150 ;
        RECT 578.100 772.050 579.900 773.850 ;
        RECT 581.550 767.700 582.750 775.050 ;
        RECT 583.950 773.850 586.050 775.950 ;
        RECT 584.100 772.050 585.900 773.850 ;
        RECT 599.400 772.950 600.600 785.400 ;
        RECT 617.400 772.950 618.600 785.400 ;
        RECT 632.550 777.150 633.750 785.400 ;
        RECT 648.300 779.400 650.100 791.250 ;
        RECT 652.500 779.400 654.300 791.250 ;
        RECT 655.800 785.400 657.600 791.250 ;
        RECT 672.150 779.400 673.950 791.250 ;
        RECT 676.650 779.400 679.950 791.250 ;
        RECT 682.650 779.400 684.450 791.250 ;
        RECT 694.350 779.400 696.150 791.250 ;
        RECT 697.350 779.400 699.150 791.250 ;
        RECT 700.650 785.400 702.450 791.250 ;
        RECT 628.950 773.850 631.050 775.950 ;
        RECT 631.950 775.050 634.050 777.150 ;
        RECT 598.950 770.850 601.050 772.950 ;
        RECT 602.100 771.150 603.900 772.950 ;
        RECT 614.100 771.150 615.900 772.950 ;
        RECT 581.550 766.800 585.150 767.700 ;
        RECT 553.200 762.600 554.250 764.400 ;
        RECT 562.950 763.500 565.050 765.600 ;
        RECT 562.950 762.600 564.000 763.500 ;
        RECT 539.850 759.750 541.650 762.600 ;
        RECT 544.350 759.750 546.150 762.600 ;
        RECT 548.550 759.750 550.350 762.600 ;
        RECT 552.450 759.750 554.250 762.600 ;
        RECT 555.750 759.750 557.550 762.600 ;
        RECT 560.250 761.700 564.000 762.600 ;
        RECT 560.250 759.750 562.050 761.700 ;
        RECT 565.050 759.750 566.850 762.600 ;
        RECT 568.050 759.750 569.850 765.600 ;
        RECT 578.850 759.750 580.650 765.600 ;
        RECT 583.350 759.750 585.150 766.800 ;
        RECT 599.400 762.600 600.600 770.850 ;
        RECT 601.950 769.050 604.050 771.150 ;
        RECT 613.950 769.050 616.050 771.150 ;
        RECT 616.950 770.850 619.050 772.950 ;
        RECT 629.100 772.050 630.900 773.850 ;
        RECT 617.400 762.600 618.600 770.850 ;
        RECT 632.550 767.700 633.750 775.050 ;
        RECT 634.950 773.850 637.050 775.950 ;
        RECT 647.100 774.150 648.900 775.950 ;
        RECT 652.950 774.150 654.150 779.400 ;
        RECT 655.950 777.150 657.750 778.950 ;
        RECT 655.950 775.050 658.050 777.150 ;
        RECT 671.250 774.150 673.050 775.950 ;
        RECT 677.250 774.150 678.450 779.400 ;
        RECT 683.100 774.150 684.900 775.950 ;
        RECT 694.650 774.150 695.850 779.400 ;
        RECT 701.250 778.500 702.450 785.400 ;
        RECT 715.350 779.400 717.150 791.250 ;
        RECT 718.350 779.400 720.150 791.250 ;
        RECT 721.650 785.400 723.450 791.250 ;
        RECT 696.750 777.600 702.450 778.500 ;
        RECT 696.750 776.700 699.000 777.600 ;
        RECT 635.100 772.050 636.900 773.850 ;
        RECT 646.950 772.050 649.050 774.150 ;
        RECT 649.950 770.850 652.050 772.950 ;
        RECT 652.950 772.050 655.050 774.150 ;
        RECT 670.950 772.050 673.050 774.150 ;
        RECT 650.100 769.050 651.900 770.850 ;
        RECT 653.850 768.750 655.050 772.050 ;
        RECT 673.950 770.850 676.050 772.950 ;
        RECT 676.950 772.050 679.050 774.150 ;
        RECT 674.700 769.050 676.500 770.850 ;
        RECT 654.000 767.700 657.750 768.750 ;
        RECT 677.400 768.150 678.600 772.050 ;
        RECT 679.950 770.850 682.050 772.950 ;
        RECT 682.950 772.050 685.050 774.150 ;
        RECT 694.650 772.050 697.050 774.150 ;
        RECT 680.100 769.050 681.900 770.850 ;
        RECT 632.550 766.800 636.150 767.700 ;
        RECT 598.650 759.750 600.450 762.600 ;
        RECT 601.650 759.750 603.450 762.600 ;
        RECT 614.550 759.750 616.350 762.600 ;
        RECT 617.550 759.750 619.350 762.600 ;
        RECT 629.850 759.750 631.650 765.600 ;
        RECT 634.350 759.750 636.150 766.800 ;
        RECT 647.550 764.700 655.350 766.050 ;
        RECT 647.550 759.750 649.350 764.700 ;
        RECT 650.550 759.750 652.350 763.800 ;
        RECT 653.550 759.750 655.350 764.700 ;
        RECT 656.550 765.600 657.750 767.700 ;
        RECT 674.250 767.100 678.600 768.150 ;
        RECT 674.250 765.600 675.150 767.100 ;
        RECT 656.550 759.750 658.350 765.600 ;
        RECT 670.650 760.500 672.450 765.600 ;
        RECT 673.650 761.400 675.450 765.600 ;
        RECT 676.650 765.000 684.450 765.900 ;
        RECT 694.650 765.600 695.850 772.050 ;
        RECT 697.950 768.300 699.000 776.700 ;
        RECT 701.100 774.150 702.900 775.950 ;
        RECT 715.650 774.150 716.850 779.400 ;
        RECT 722.250 778.500 723.450 785.400 ;
        RECT 717.750 777.600 723.450 778.500 ;
        RECT 726.150 779.400 727.950 791.250 ;
        RECT 729.150 785.400 730.950 791.250 ;
        RECT 734.250 785.400 736.050 791.250 ;
        RECT 739.050 785.400 740.850 791.250 ;
        RECT 734.550 784.500 735.750 785.400 ;
        RECT 742.050 784.500 743.850 791.250 ;
        RECT 745.950 785.400 747.750 791.250 ;
        RECT 750.150 785.400 751.950 791.250 ;
        RECT 754.650 788.400 756.450 791.250 ;
        RECT 730.950 782.400 735.750 784.500 ;
        RECT 738.150 782.700 745.050 784.500 ;
        RECT 750.150 783.300 754.050 785.400 ;
        RECT 734.550 781.500 735.750 782.400 ;
        RECT 747.450 781.800 749.250 782.400 ;
        RECT 734.550 780.300 742.050 781.500 ;
        RECT 740.250 779.700 742.050 780.300 ;
        RECT 742.950 780.900 749.250 781.800 ;
        RECT 726.150 778.800 737.250 779.400 ;
        RECT 742.950 778.800 743.850 780.900 ;
        RECT 747.450 780.600 749.250 780.900 ;
        RECT 750.150 780.600 752.850 782.400 ;
        RECT 750.150 779.700 751.050 780.600 ;
        RECT 726.150 778.200 743.850 778.800 ;
        RECT 717.750 776.700 720.000 777.600 ;
        RECT 700.950 772.050 703.050 774.150 ;
        RECT 715.650 772.050 718.050 774.150 ;
        RECT 696.750 767.400 699.000 768.300 ;
        RECT 696.750 766.500 701.850 767.400 ;
        RECT 676.650 760.500 678.450 765.000 ;
        RECT 670.650 759.750 678.450 760.500 ;
        RECT 679.650 759.750 681.450 764.100 ;
        RECT 682.650 759.750 684.450 765.000 ;
        RECT 694.350 759.750 696.150 765.600 ;
        RECT 697.350 759.750 699.150 765.600 ;
        RECT 700.650 762.600 701.850 766.500 ;
        RECT 715.650 765.600 716.850 772.050 ;
        RECT 718.950 768.300 720.000 776.700 ;
        RECT 722.100 774.150 723.900 775.950 ;
        RECT 721.950 772.050 724.050 774.150 ;
        RECT 717.750 767.400 720.000 768.300 ;
        RECT 717.750 766.500 722.850 767.400 ;
        RECT 700.650 759.750 702.450 762.600 ;
        RECT 715.350 759.750 717.150 765.600 ;
        RECT 718.350 759.750 720.150 765.600 ;
        RECT 721.650 762.600 722.850 766.500 ;
        RECT 726.150 765.600 727.050 778.200 ;
        RECT 735.450 777.900 743.850 778.200 ;
        RECT 745.050 778.800 751.050 779.700 ;
        RECT 751.950 778.800 754.050 779.700 ;
        RECT 757.650 779.400 759.450 791.250 ;
        RECT 770.550 785.400 772.350 791.250 ;
        RECT 773.550 785.400 775.350 791.250 ;
        RECT 788.400 785.400 790.200 791.250 ;
        RECT 735.450 777.600 737.250 777.900 ;
        RECT 745.050 774.150 745.950 778.800 ;
        RECT 751.950 777.600 756.150 778.800 ;
        RECT 755.250 775.800 757.050 777.600 ;
        RECT 736.950 773.100 739.050 774.150 ;
        RECT 728.100 771.150 729.900 772.950 ;
        RECT 731.100 772.050 739.050 773.100 ;
        RECT 742.950 772.050 745.950 774.150 ;
        RECT 731.100 771.300 732.900 772.050 ;
        RECT 729.000 770.400 729.900 771.150 ;
        RECT 734.100 770.400 735.900 771.000 ;
        RECT 729.000 769.200 735.900 770.400 ;
        RECT 734.850 768.000 735.900 769.200 ;
        RECT 745.050 768.000 745.950 772.050 ;
        RECT 754.950 771.750 757.050 772.050 ;
        RECT 753.150 769.950 757.050 771.750 ;
        RECT 758.250 769.950 759.450 779.400 ;
        RECT 773.400 772.950 774.600 785.400 ;
        RECT 791.700 779.400 793.500 791.250 ;
        RECT 795.900 779.400 797.700 791.250 ;
        RECT 807.300 779.400 809.100 791.250 ;
        RECT 811.500 779.400 813.300 791.250 ;
        RECT 814.800 785.400 816.600 791.250 ;
        RECT 830.550 780.300 832.350 791.250 ;
        RECT 833.550 781.200 835.350 791.250 ;
        RECT 836.550 780.300 838.350 791.250 ;
        RECT 830.550 779.400 838.350 780.300 ;
        RECT 839.550 779.400 841.350 791.250 ;
        RECT 853.650 779.400 855.450 791.250 ;
        RECT 788.250 777.150 790.050 778.950 ;
        RECT 787.950 775.050 790.050 777.150 ;
        RECT 791.850 774.150 793.050 779.400 ;
        RECT 797.100 774.150 798.900 775.950 ;
        RECT 806.100 774.150 807.900 775.950 ;
        RECT 811.950 774.150 813.150 779.400 ;
        RECT 814.950 777.150 816.750 778.950 ;
        RECT 823.950 777.450 826.050 778.050 ;
        RECT 835.950 777.450 838.050 778.050 ;
        RECT 814.950 775.050 817.050 777.150 ;
        RECT 823.950 776.550 838.050 777.450 ;
        RECT 823.950 775.950 826.050 776.550 ;
        RECT 835.950 775.950 838.050 776.550 ;
        RECT 839.700 774.150 840.900 779.400 ;
        RECT 856.650 778.500 858.450 791.250 ;
        RECT 859.650 779.400 861.450 791.250 ;
        RECT 862.650 778.500 864.450 791.250 ;
        RECT 865.650 779.400 867.450 791.250 ;
        RECT 868.650 778.500 870.450 791.250 ;
        RECT 871.650 779.400 873.450 791.250 ;
        RECT 874.650 778.500 876.450 791.250 ;
        RECT 877.650 779.400 879.450 791.250 ;
        RECT 855.750 777.300 858.450 778.500 ;
        RECT 860.700 777.300 864.450 778.500 ;
        RECT 866.700 777.300 870.450 778.500 ;
        RECT 872.550 777.300 876.450 778.500 ;
        RECT 770.100 771.150 771.900 772.950 ;
        RECT 734.850 767.100 745.950 768.000 ;
        RECT 754.950 767.850 759.450 769.950 ;
        RECT 769.950 769.050 772.050 771.150 ;
        RECT 772.950 770.850 775.050 772.950 ;
        RECT 790.950 772.050 793.050 774.150 ;
        RECT 734.850 766.200 735.900 767.100 ;
        RECT 745.050 766.800 745.950 767.100 ;
        RECT 721.650 759.750 723.450 762.600 ;
        RECT 726.150 759.750 727.950 765.600 ;
        RECT 730.950 763.500 733.050 765.600 ;
        RECT 734.550 764.400 736.350 766.200 ;
        RECT 737.850 765.450 739.650 766.200 ;
        RECT 737.850 764.400 742.800 765.450 ;
        RECT 745.050 765.000 746.850 766.800 ;
        RECT 758.250 765.600 759.450 767.850 ;
        RECT 751.950 764.700 754.050 765.600 ;
        RECT 732.000 762.600 733.050 763.500 ;
        RECT 741.750 762.600 742.800 764.400 ;
        RECT 750.300 763.500 754.050 764.700 ;
        RECT 750.300 762.600 751.350 763.500 ;
        RECT 729.150 759.750 730.950 762.600 ;
        RECT 732.000 761.700 735.750 762.600 ;
        RECT 733.950 759.750 735.750 761.700 ;
        RECT 738.450 759.750 740.250 762.600 ;
        RECT 741.750 759.750 743.550 762.600 ;
        RECT 745.650 759.750 747.450 762.600 ;
        RECT 749.850 759.750 751.650 762.600 ;
        RECT 754.350 759.750 756.150 762.600 ;
        RECT 757.650 759.750 759.450 765.600 ;
        RECT 773.400 762.600 774.600 770.850 ;
        RECT 790.950 768.750 792.150 772.050 ;
        RECT 793.950 770.850 796.050 772.950 ;
        RECT 796.950 772.050 799.050 774.150 ;
        RECT 805.950 772.050 808.050 774.150 ;
        RECT 808.950 770.850 811.050 772.950 ;
        RECT 811.950 772.050 814.050 774.150 ;
        RECT 794.100 769.050 795.900 770.850 ;
        RECT 809.100 769.050 810.900 770.850 ;
        RECT 812.850 768.750 814.050 772.050 ;
        RECT 814.950 771.450 817.050 772.050 ;
        RECT 826.950 771.450 829.050 772.050 ;
        RECT 814.950 770.550 829.050 771.450 ;
        RECT 829.950 770.850 832.050 772.950 ;
        RECT 833.100 771.150 834.900 772.950 ;
        RECT 814.950 769.950 817.050 770.550 ;
        RECT 826.950 769.950 829.050 770.550 ;
        RECT 830.100 769.050 831.900 770.850 ;
        RECT 832.950 769.050 835.050 771.150 ;
        RECT 835.950 770.850 838.050 772.950 ;
        RECT 838.950 772.050 841.050 774.150 ;
        RECT 855.750 772.950 856.800 777.300 ;
        RECT 836.100 769.050 837.900 770.850 ;
        RECT 788.250 767.700 792.000 768.750 ;
        RECT 813.000 767.700 816.750 768.750 ;
        RECT 788.250 765.600 789.450 767.700 ;
        RECT 770.550 759.750 772.350 762.600 ;
        RECT 773.550 759.750 775.350 762.600 ;
        RECT 787.650 759.750 789.450 765.600 ;
        RECT 790.650 764.700 798.450 766.050 ;
        RECT 790.650 759.750 792.450 764.700 ;
        RECT 793.650 759.750 795.450 763.800 ;
        RECT 796.650 759.750 798.450 764.700 ;
        RECT 806.550 764.700 814.350 766.050 ;
        RECT 806.550 759.750 808.350 764.700 ;
        RECT 809.550 759.750 811.350 763.800 ;
        RECT 812.550 759.750 814.350 764.700 ;
        RECT 815.550 765.600 816.750 767.700 ;
        RECT 839.700 765.600 840.900 772.050 ;
        RECT 853.950 770.850 856.800 772.950 ;
        RECT 855.750 767.700 856.800 770.850 ;
        RECT 860.700 770.400 861.900 777.300 ;
        RECT 866.700 770.400 867.900 777.300 ;
        RECT 872.550 770.400 873.750 777.300 ;
        RECT 874.950 770.850 877.050 772.950 ;
        RECT 857.700 768.600 861.900 770.400 ;
        RECT 863.700 768.600 867.900 770.400 ;
        RECT 869.700 768.600 873.750 770.400 ;
        RECT 875.100 769.050 876.900 770.850 ;
        RECT 860.700 767.700 861.900 768.600 ;
        RECT 866.700 767.700 867.900 768.600 ;
        RECT 872.550 767.700 873.750 768.600 ;
        RECT 855.750 766.650 858.600 767.700 ;
        RECT 855.900 766.500 858.600 766.650 ;
        RECT 860.700 766.500 864.600 767.700 ;
        RECT 866.700 766.500 870.450 767.700 ;
        RECT 872.550 766.500 876.600 767.700 ;
        RECT 856.800 765.600 858.600 766.500 ;
        RECT 862.800 765.600 864.600 766.500 ;
        RECT 815.550 759.750 817.350 765.600 ;
        RECT 831.000 759.750 832.800 765.600 ;
        RECT 835.200 763.950 840.900 765.600 ;
        RECT 835.200 759.750 837.000 763.950 ;
        RECT 838.500 759.750 840.300 762.600 ;
        RECT 853.650 759.750 855.450 765.600 ;
        RECT 856.650 759.750 858.450 765.600 ;
        RECT 859.650 759.750 861.450 765.600 ;
        RECT 862.650 759.750 864.450 765.600 ;
        RECT 865.650 759.750 867.450 765.600 ;
        RECT 868.650 759.750 870.450 766.500 ;
        RECT 874.800 765.600 876.600 766.500 ;
        RECT 871.650 759.750 873.450 765.600 ;
        RECT 874.650 759.750 876.450 765.600 ;
        RECT 877.650 759.750 879.450 765.600 ;
        RECT 11.550 747.900 13.350 755.250 ;
        RECT 16.050 749.400 17.850 755.250 ;
        RECT 19.050 750.900 20.850 755.250 ;
        RECT 19.050 749.400 22.350 750.900 ;
        RECT 17.250 747.900 19.050 748.500 ;
        RECT 11.550 746.700 19.050 747.900 ;
        RECT 10.950 740.850 13.050 742.950 ;
        RECT 11.100 739.050 12.900 740.850 ;
        RECT 14.700 729.600 15.900 746.700 ;
        RECT 21.150 742.950 22.350 749.400 ;
        RECT 32.700 746.400 34.500 755.250 ;
        RECT 38.100 747.000 39.900 755.250 ;
        RECT 56.850 749.400 58.650 755.250 ;
        RECT 61.350 748.200 63.150 755.250 ;
        RECT 75.000 749.400 76.800 755.250 ;
        RECT 79.200 751.050 81.000 755.250 ;
        RECT 82.500 752.400 84.300 755.250 ;
        RECT 79.200 749.400 84.900 751.050 ;
        RECT 102.150 750.900 103.950 755.250 ;
        RECT 59.550 747.300 63.150 748.200 ;
        RECT 38.100 745.350 42.600 747.000 ;
        RECT 17.100 741.150 18.900 742.950 ;
        RECT 16.950 739.050 19.050 741.150 ;
        RECT 19.950 740.850 22.350 742.950 ;
        RECT 41.400 741.150 42.600 745.350 ;
        RECT 56.100 741.150 57.900 742.950 ;
        RECT 21.150 735.600 22.350 740.850 ;
        RECT 31.950 737.850 34.050 739.950 ;
        RECT 37.950 737.850 40.050 739.950 ;
        RECT 40.950 739.050 43.050 741.150 ;
        RECT 55.950 739.050 58.050 741.150 ;
        RECT 59.550 739.950 60.750 747.300 ;
        RECT 74.100 744.150 75.900 745.950 ;
        RECT 62.100 741.150 63.900 742.950 ;
        RECT 73.950 742.050 76.050 744.150 ;
        RECT 76.950 743.850 79.050 745.950 ;
        RECT 80.100 744.150 81.900 745.950 ;
        RECT 77.100 742.050 78.900 743.850 ;
        RECT 79.950 742.050 82.050 744.150 ;
        RECT 83.700 742.950 84.900 749.400 ;
        RECT 100.650 749.400 103.950 750.900 ;
        RECT 105.150 749.400 106.950 755.250 ;
        RECT 100.650 742.950 101.850 749.400 ;
        RECT 103.950 747.900 105.750 748.500 ;
        RECT 109.650 747.900 111.450 755.250 ;
        RECT 119.850 749.400 121.650 755.250 ;
        RECT 124.350 748.200 126.150 755.250 ;
        RECT 103.950 746.700 111.450 747.900 ;
        RECT 122.550 747.300 126.150 748.200 ;
        RECT 140.550 747.900 142.350 755.250 ;
        RECT 145.050 749.400 146.850 755.250 ;
        RECT 148.050 750.900 149.850 755.250 ;
        RECT 148.050 749.400 151.350 750.900 ;
        RECT 146.250 747.900 148.050 748.500 ;
        RECT 32.100 736.050 33.900 737.850 ;
        RECT 11.550 723.750 13.350 729.600 ;
        RECT 14.550 723.750 16.350 729.600 ;
        RECT 18.150 723.750 19.950 735.600 ;
        RECT 21.150 723.750 22.950 735.600 ;
        RECT 34.950 734.850 37.050 736.950 ;
        RECT 38.250 736.050 40.050 737.850 ;
        RECT 35.100 733.050 36.900 734.850 ;
        RECT 41.700 730.800 42.750 739.050 ;
        RECT 58.950 737.850 61.050 739.950 ;
        RECT 61.950 739.050 64.050 741.150 ;
        RECT 82.950 740.850 85.050 742.950 ;
        RECT 100.650 740.850 103.050 742.950 ;
        RECT 104.100 741.150 105.900 742.950 ;
        RECT 35.700 729.900 42.750 730.800 ;
        RECT 35.700 729.600 37.350 729.900 ;
        RECT 32.550 723.750 34.350 729.600 ;
        RECT 35.550 723.750 37.350 729.600 ;
        RECT 41.550 729.600 42.750 729.900 ;
        RECT 59.550 729.600 60.750 737.850 ;
        RECT 83.700 735.600 84.900 740.850 ;
        RECT 100.650 735.600 101.850 740.850 ;
        RECT 103.950 739.050 106.050 741.150 ;
        RECT 74.550 734.700 82.350 735.600 ;
        RECT 38.550 723.750 40.350 729.000 ;
        RECT 41.550 723.750 43.350 729.600 ;
        RECT 56.550 723.750 58.350 729.600 ;
        RECT 59.550 723.750 61.350 729.600 ;
        RECT 62.550 723.750 64.350 729.600 ;
        RECT 74.550 723.750 76.350 734.700 ;
        RECT 77.550 723.750 79.350 733.800 ;
        RECT 80.550 723.750 82.350 734.700 ;
        RECT 83.550 723.750 85.350 735.600 ;
        RECT 100.050 723.750 101.850 735.600 ;
        RECT 103.050 723.750 104.850 735.600 ;
        RECT 107.100 729.600 108.300 746.700 ;
        RECT 109.950 740.850 112.050 742.950 ;
        RECT 119.100 741.150 120.900 742.950 ;
        RECT 110.100 739.050 111.900 740.850 ;
        RECT 118.950 739.050 121.050 741.150 ;
        RECT 122.550 739.950 123.750 747.300 ;
        RECT 140.550 746.700 148.050 747.900 ;
        RECT 125.100 741.150 126.900 742.950 ;
        RECT 121.950 737.850 124.050 739.950 ;
        RECT 124.950 739.050 127.050 741.150 ;
        RECT 139.950 740.850 142.050 742.950 ;
        RECT 140.100 739.050 141.900 740.850 ;
        RECT 122.550 729.600 123.750 737.850 ;
        RECT 143.700 729.600 144.900 746.700 ;
        RECT 150.150 742.950 151.350 749.400 ;
        RECT 167.100 747.000 168.900 755.250 ;
        RECT 146.100 741.150 147.900 742.950 ;
        RECT 145.950 739.050 148.050 741.150 ;
        RECT 148.950 740.850 151.350 742.950 ;
        RECT 164.400 745.350 168.900 747.000 ;
        RECT 172.500 746.400 174.300 755.250 ;
        RECT 186.150 750.900 187.950 755.250 ;
        RECT 184.650 749.400 187.950 750.900 ;
        RECT 189.150 749.400 190.950 755.250 ;
        RECT 164.400 741.150 165.600 745.350 ;
        RECT 184.650 742.950 185.850 749.400 ;
        RECT 187.950 747.900 189.750 748.500 ;
        RECT 193.650 747.900 195.450 755.250 ;
        RECT 208.650 749.400 210.450 755.250 ;
        RECT 187.950 746.700 195.450 747.900 ;
        RECT 209.250 747.300 210.450 749.400 ;
        RECT 211.650 750.300 213.450 755.250 ;
        RECT 214.650 751.200 216.450 755.250 ;
        RECT 217.650 750.300 219.450 755.250 ;
        RECT 211.650 748.950 219.450 750.300 ;
        RECT 150.150 735.600 151.350 740.850 ;
        RECT 163.950 739.050 166.050 741.150 ;
        RECT 184.650 740.850 187.050 742.950 ;
        RECT 188.100 741.150 189.900 742.950 ;
        RECT 106.650 723.750 108.450 729.600 ;
        RECT 109.650 723.750 111.450 729.600 ;
        RECT 119.550 723.750 121.350 729.600 ;
        RECT 122.550 723.750 124.350 729.600 ;
        RECT 125.550 723.750 127.350 729.600 ;
        RECT 140.550 723.750 142.350 729.600 ;
        RECT 143.550 723.750 145.350 729.600 ;
        RECT 147.150 723.750 148.950 735.600 ;
        RECT 150.150 723.750 151.950 735.600 ;
        RECT 164.250 730.800 165.300 739.050 ;
        RECT 166.950 737.850 169.050 739.950 ;
        RECT 172.950 737.850 175.050 739.950 ;
        RECT 166.950 736.050 168.750 737.850 ;
        RECT 169.950 734.850 172.050 736.950 ;
        RECT 173.100 736.050 174.900 737.850 ;
        RECT 184.650 735.600 185.850 740.850 ;
        RECT 187.950 739.050 190.050 741.150 ;
        RECT 170.100 733.050 171.900 734.850 ;
        RECT 164.250 729.900 171.300 730.800 ;
        RECT 164.250 729.600 165.450 729.900 ;
        RECT 163.650 723.750 165.450 729.600 ;
        RECT 169.650 729.600 171.300 729.900 ;
        RECT 166.650 723.750 168.450 729.000 ;
        RECT 169.650 723.750 171.450 729.600 ;
        RECT 172.650 723.750 174.450 729.600 ;
        RECT 184.050 723.750 185.850 735.600 ;
        RECT 187.050 723.750 188.850 735.600 ;
        RECT 191.100 729.600 192.300 746.700 ;
        RECT 209.250 746.250 213.000 747.300 ;
        RECT 233.100 747.000 234.900 755.250 ;
        RECT 211.950 742.950 213.150 746.250 ;
        RECT 215.100 744.150 216.900 745.950 ;
        RECT 230.400 745.350 234.900 747.000 ;
        RECT 238.500 746.400 240.300 755.250 ;
        RECT 248.850 749.400 250.650 755.250 ;
        RECT 253.350 748.200 255.150 755.250 ;
        RECT 266.550 752.400 268.350 755.250 ;
        RECT 269.550 752.400 271.350 755.250 ;
        RECT 251.550 747.300 255.150 748.200 ;
        RECT 193.950 740.850 196.050 742.950 ;
        RECT 211.950 740.850 214.050 742.950 ;
        RECT 214.950 742.050 217.050 744.150 ;
        RECT 217.950 740.850 220.050 742.950 ;
        RECT 230.400 741.150 231.600 745.350 ;
        RECT 248.100 741.150 249.900 742.950 ;
        RECT 194.100 739.050 195.900 740.850 ;
        RECT 208.950 737.850 211.050 739.950 ;
        RECT 209.250 736.050 211.050 737.850 ;
        RECT 212.850 735.600 214.050 740.850 ;
        RECT 218.100 739.050 219.900 740.850 ;
        RECT 229.950 739.050 232.050 741.150 ;
        RECT 190.650 723.750 192.450 729.600 ;
        RECT 193.650 723.750 195.450 729.600 ;
        RECT 209.400 723.750 211.200 729.600 ;
        RECT 212.700 723.750 214.500 735.600 ;
        RECT 216.900 723.750 218.700 735.600 ;
        RECT 230.250 730.800 231.300 739.050 ;
        RECT 232.950 737.850 235.050 739.950 ;
        RECT 238.950 737.850 241.050 739.950 ;
        RECT 247.950 739.050 250.050 741.150 ;
        RECT 251.550 739.950 252.750 747.300 ;
        RECT 265.950 743.850 268.050 745.950 ;
        RECT 269.400 744.150 270.600 752.400 ;
        RECT 281.550 750.300 283.350 755.250 ;
        RECT 284.550 751.200 286.350 755.250 ;
        RECT 287.550 750.300 289.350 755.250 ;
        RECT 281.550 748.950 289.350 750.300 ;
        RECT 290.550 749.400 292.350 755.250 ;
        RECT 290.550 747.300 291.750 749.400 ;
        RECT 308.850 748.200 310.650 755.250 ;
        RECT 313.350 749.400 315.150 755.250 ;
        RECT 323.550 752.400 325.350 755.250 ;
        RECT 326.550 752.400 328.350 755.250 ;
        RECT 329.550 752.400 331.350 755.250 ;
        RECT 327.450 748.200 328.350 752.400 ;
        RECT 332.550 749.400 334.350 755.250 ;
        RECT 344.850 749.400 346.650 755.250 ;
        RECT 308.850 747.300 312.450 748.200 ;
        RECT 327.450 747.300 330.750 748.200 ;
        RECT 288.000 746.250 291.750 747.300 ;
        RECT 284.100 744.150 285.900 745.950 ;
        RECT 254.100 741.150 255.900 742.950 ;
        RECT 266.100 742.050 267.900 743.850 ;
        RECT 268.950 742.050 271.050 744.150 ;
        RECT 250.950 737.850 253.050 739.950 ;
        RECT 253.950 739.050 256.050 741.150 ;
        RECT 232.950 736.050 234.750 737.850 ;
        RECT 235.950 734.850 238.050 736.950 ;
        RECT 239.100 736.050 240.900 737.850 ;
        RECT 236.100 733.050 237.900 734.850 ;
        RECT 230.250 729.900 237.300 730.800 ;
        RECT 230.250 729.600 231.450 729.900 ;
        RECT 229.650 723.750 231.450 729.600 ;
        RECT 235.650 729.600 237.300 729.900 ;
        RECT 251.550 729.600 252.750 737.850 ;
        RECT 269.400 729.600 270.600 742.050 ;
        RECT 280.950 740.850 283.050 742.950 ;
        RECT 283.950 742.050 286.050 744.150 ;
        RECT 287.850 742.950 289.050 746.250 ;
        RECT 286.950 740.850 289.050 742.950 ;
        RECT 308.100 741.150 309.900 742.950 ;
        RECT 281.100 739.050 282.900 740.850 ;
        RECT 286.950 735.600 288.150 740.850 ;
        RECT 289.950 737.850 292.050 739.950 ;
        RECT 307.950 739.050 310.050 741.150 ;
        RECT 311.250 739.950 312.450 747.300 ;
        RECT 328.950 746.400 330.750 747.300 ;
        RECT 322.950 743.850 325.050 745.950 ;
        RECT 314.100 741.150 315.900 742.950 ;
        RECT 323.100 742.050 324.900 743.850 ;
        RECT 310.950 737.850 313.050 739.950 ;
        RECT 313.950 739.050 316.050 741.150 ;
        RECT 325.950 740.850 328.050 742.950 ;
        RECT 326.100 739.050 327.900 740.850 ;
        RECT 329.700 738.150 330.600 746.400 ;
        RECT 333.000 744.150 334.050 749.400 ;
        RECT 349.350 748.200 351.150 755.250 ;
        RECT 362.550 752.400 364.350 755.250 ;
        RECT 331.950 742.050 334.050 744.150 ;
        RECT 347.550 747.300 351.150 748.200 ;
        RECT 363.150 748.500 364.350 752.400 ;
        RECT 365.850 749.400 367.650 755.250 ;
        RECT 368.850 749.400 370.650 755.250 ;
        RECT 385.650 749.400 387.450 755.250 ;
        RECT 363.150 747.600 368.250 748.500 ;
        RECT 328.950 738.000 330.750 738.150 ;
        RECT 289.950 736.050 291.750 737.850 ;
        RECT 232.650 723.750 234.450 729.000 ;
        RECT 235.650 723.750 237.450 729.600 ;
        RECT 238.650 723.750 240.450 729.600 ;
        RECT 248.550 723.750 250.350 729.600 ;
        RECT 251.550 723.750 253.350 729.600 ;
        RECT 254.550 723.750 256.350 729.600 ;
        RECT 266.550 723.750 268.350 729.600 ;
        RECT 269.550 723.750 271.350 729.600 ;
        RECT 282.300 723.750 284.100 735.600 ;
        RECT 286.500 723.750 288.300 735.600 ;
        RECT 311.250 729.600 312.450 737.850 ;
        RECT 323.550 736.800 330.750 738.000 ;
        RECT 323.550 735.600 324.750 736.800 ;
        RECT 328.950 736.350 330.750 736.800 ;
        RECT 289.800 723.750 291.600 729.600 ;
        RECT 307.650 723.750 309.450 729.600 ;
        RECT 310.650 723.750 312.450 729.600 ;
        RECT 313.650 723.750 315.450 729.600 ;
        RECT 323.550 723.750 325.350 735.600 ;
        RECT 332.100 735.450 333.450 742.050 ;
        RECT 344.100 741.150 345.900 742.950 ;
        RECT 343.950 739.050 346.050 741.150 ;
        RECT 347.550 739.950 348.750 747.300 ;
        RECT 366.000 746.700 368.250 747.600 ;
        RECT 350.100 741.150 351.900 742.950 ;
        RECT 346.950 737.850 349.050 739.950 ;
        RECT 349.950 739.050 352.050 741.150 ;
        RECT 361.950 740.850 364.050 742.950 ;
        RECT 362.100 739.050 363.900 740.850 ;
        RECT 366.000 738.300 367.050 746.700 ;
        RECT 369.150 742.950 370.350 749.400 ;
        RECT 386.250 747.300 387.450 749.400 ;
        RECT 388.650 750.300 390.450 755.250 ;
        RECT 391.650 751.200 393.450 755.250 ;
        RECT 394.650 750.300 396.450 755.250 ;
        RECT 388.650 748.950 396.450 750.300 ;
        RECT 410.850 748.200 412.650 755.250 ;
        RECT 415.350 749.400 417.150 755.250 ;
        RECT 426.000 749.400 427.800 755.250 ;
        RECT 430.200 751.050 432.000 755.250 ;
        RECT 433.500 752.400 435.300 755.250 ;
        RECT 446.550 752.400 448.350 755.250 ;
        RECT 449.550 752.400 451.350 755.250 ;
        RECT 464.700 752.400 466.500 755.250 ;
        RECT 430.200 749.400 435.900 751.050 ;
        RECT 410.850 747.300 414.450 748.200 ;
        RECT 386.250 746.250 390.000 747.300 ;
        RECT 367.950 740.850 370.350 742.950 ;
        RECT 388.950 742.950 390.150 746.250 ;
        RECT 392.100 744.150 393.900 745.950 ;
        RECT 388.950 740.850 391.050 742.950 ;
        RECT 391.950 742.050 394.050 744.150 ;
        RECT 394.950 740.850 397.050 742.950 ;
        RECT 410.100 741.150 411.900 742.950 ;
        RECT 328.050 723.750 329.850 735.450 ;
        RECT 331.050 734.100 333.450 735.450 ;
        RECT 331.050 723.750 332.850 734.100 ;
        RECT 347.550 729.600 348.750 737.850 ;
        RECT 366.000 737.400 368.250 738.300 ;
        RECT 362.550 736.500 368.250 737.400 ;
        RECT 362.550 729.600 363.750 736.500 ;
        RECT 369.150 735.600 370.350 740.850 ;
        RECT 385.950 737.850 388.050 739.950 ;
        RECT 386.250 736.050 388.050 737.850 ;
        RECT 389.850 735.600 391.050 740.850 ;
        RECT 395.100 739.050 396.900 740.850 ;
        RECT 409.950 739.050 412.050 741.150 ;
        RECT 413.250 739.950 414.450 747.300 ;
        RECT 425.100 744.150 426.900 745.950 ;
        RECT 416.100 741.150 417.900 742.950 ;
        RECT 424.950 742.050 427.050 744.150 ;
        RECT 427.950 743.850 430.050 745.950 ;
        RECT 431.100 744.150 432.900 745.950 ;
        RECT 428.100 742.050 429.900 743.850 ;
        RECT 430.950 742.050 433.050 744.150 ;
        RECT 434.700 742.950 435.900 749.400 ;
        RECT 445.950 743.850 448.050 745.950 ;
        RECT 449.400 744.150 450.600 752.400 ;
        RECT 468.000 751.050 469.800 755.250 ;
        RECT 464.100 749.400 469.800 751.050 ;
        RECT 472.200 749.400 474.000 755.250 ;
        RECT 483.000 749.400 484.800 755.250 ;
        RECT 487.200 751.050 489.000 755.250 ;
        RECT 490.500 752.400 492.300 755.250 ;
        RECT 487.200 749.400 492.900 751.050 ;
        RECT 412.950 737.850 415.050 739.950 ;
        RECT 415.950 739.050 418.050 741.150 ;
        RECT 433.950 740.850 436.050 742.950 ;
        RECT 446.100 742.050 447.900 743.850 ;
        RECT 448.950 742.050 451.050 744.150 ;
        RECT 464.100 742.950 465.300 749.400 ;
        RECT 467.100 744.150 468.900 745.950 ;
        RECT 344.550 723.750 346.350 729.600 ;
        RECT 347.550 723.750 349.350 729.600 ;
        RECT 350.550 723.750 352.350 729.600 ;
        RECT 362.550 723.750 364.350 729.600 ;
        RECT 365.850 723.750 367.650 735.600 ;
        RECT 368.850 723.750 370.650 735.600 ;
        RECT 386.400 723.750 388.200 729.600 ;
        RECT 389.700 723.750 391.500 735.600 ;
        RECT 393.900 723.750 395.700 735.600 ;
        RECT 413.250 729.600 414.450 737.850 ;
        RECT 434.700 735.600 435.900 740.850 ;
        RECT 425.550 734.700 433.350 735.600 ;
        RECT 409.650 723.750 411.450 729.600 ;
        RECT 412.650 723.750 414.450 729.600 ;
        RECT 415.650 723.750 417.450 729.600 ;
        RECT 425.550 723.750 427.350 734.700 ;
        RECT 428.550 723.750 430.350 733.800 ;
        RECT 431.550 723.750 433.350 734.700 ;
        RECT 434.550 723.750 436.350 735.600 ;
        RECT 449.400 729.600 450.600 742.050 ;
        RECT 463.950 740.850 466.050 742.950 ;
        RECT 466.950 742.050 469.050 744.150 ;
        RECT 469.950 743.850 472.050 745.950 ;
        RECT 473.100 744.150 474.900 745.950 ;
        RECT 482.100 744.150 483.900 745.950 ;
        RECT 470.100 742.050 471.900 743.850 ;
        RECT 472.950 742.050 475.050 744.150 ;
        RECT 481.950 742.050 484.050 744.150 ;
        RECT 484.950 743.850 487.050 745.950 ;
        RECT 488.100 744.150 489.900 745.950 ;
        RECT 485.100 742.050 486.900 743.850 ;
        RECT 487.950 742.050 490.050 744.150 ;
        RECT 491.700 742.950 492.900 749.400 ;
        RECT 503.550 750.300 505.350 755.250 ;
        RECT 506.550 751.200 508.350 755.250 ;
        RECT 509.550 750.300 511.350 755.250 ;
        RECT 503.550 748.950 511.350 750.300 ;
        RECT 512.550 749.400 514.350 755.250 ;
        RECT 529.650 749.400 531.450 755.250 ;
        RECT 512.550 747.300 513.750 749.400 ;
        RECT 510.000 746.250 513.750 747.300 ;
        RECT 530.250 747.300 531.450 749.400 ;
        RECT 532.650 750.300 534.450 755.250 ;
        RECT 535.650 751.200 537.450 755.250 ;
        RECT 538.650 750.300 540.450 755.250 ;
        RECT 532.650 748.950 540.450 750.300 ;
        RECT 543.150 749.400 544.950 755.250 ;
        RECT 546.150 752.400 547.950 755.250 ;
        RECT 550.950 753.300 552.750 755.250 ;
        RECT 549.000 752.400 552.750 753.300 ;
        RECT 555.450 752.400 557.250 755.250 ;
        RECT 558.750 752.400 560.550 755.250 ;
        RECT 562.650 752.400 564.450 755.250 ;
        RECT 566.850 752.400 568.650 755.250 ;
        RECT 571.350 752.400 573.150 755.250 ;
        RECT 549.000 751.500 550.050 752.400 ;
        RECT 547.950 749.400 550.050 751.500 ;
        RECT 558.750 750.600 559.800 752.400 ;
        RECT 530.250 746.250 534.000 747.300 ;
        RECT 506.100 744.150 507.900 745.950 ;
        RECT 490.950 740.850 493.050 742.950 ;
        RECT 502.950 740.850 505.050 742.950 ;
        RECT 505.950 742.050 508.050 744.150 ;
        RECT 509.850 742.950 511.050 746.250 ;
        RECT 508.950 740.850 511.050 742.950 ;
        RECT 532.950 742.950 534.150 746.250 ;
        RECT 536.100 744.150 537.900 745.950 ;
        RECT 532.950 740.850 535.050 742.950 ;
        RECT 535.950 742.050 538.050 744.150 ;
        RECT 538.950 740.850 541.050 742.950 ;
        RECT 464.100 735.600 465.300 740.850 ;
        RECT 472.950 738.450 475.050 739.050 ;
        RECT 487.950 738.450 490.050 739.050 ;
        RECT 472.950 737.550 490.050 738.450 ;
        RECT 472.950 736.950 475.050 737.550 ;
        RECT 487.950 736.950 490.050 737.550 ;
        RECT 491.700 735.600 492.900 740.850 ;
        RECT 503.100 739.050 504.900 740.850 ;
        RECT 508.950 735.600 510.150 740.850 ;
        RECT 511.950 737.850 514.050 739.950 ;
        RECT 529.950 737.850 532.050 739.950 ;
        RECT 511.950 736.050 513.750 737.850 ;
        RECT 530.250 736.050 532.050 737.850 ;
        RECT 533.850 735.600 535.050 740.850 ;
        RECT 539.100 739.050 540.900 740.850 ;
        RECT 543.150 736.800 544.050 749.400 ;
        RECT 551.550 748.800 553.350 750.600 ;
        RECT 554.850 749.550 559.800 750.600 ;
        RECT 567.300 751.500 568.350 752.400 ;
        RECT 567.300 750.300 571.050 751.500 ;
        RECT 554.850 748.800 556.650 749.550 ;
        RECT 551.850 747.900 552.900 748.800 ;
        RECT 562.050 748.200 563.850 750.000 ;
        RECT 568.950 749.400 571.050 750.300 ;
        RECT 574.650 749.400 576.450 755.250 ;
        RECT 562.050 747.900 562.950 748.200 ;
        RECT 551.850 747.000 562.950 747.900 ;
        RECT 575.250 747.150 576.450 749.400 ;
        RECT 551.850 745.800 552.900 747.000 ;
        RECT 546.000 744.600 552.900 745.800 ;
        RECT 546.000 743.850 546.900 744.600 ;
        RECT 551.100 744.000 552.900 744.600 ;
        RECT 545.100 742.050 546.900 743.850 ;
        RECT 548.100 742.950 549.900 743.700 ;
        RECT 562.050 742.950 562.950 747.000 ;
        RECT 571.950 745.050 576.450 747.150 ;
        RECT 570.150 743.250 574.050 745.050 ;
        RECT 571.950 742.950 574.050 743.250 ;
        RECT 548.100 741.900 556.050 742.950 ;
        RECT 553.950 740.850 556.050 741.900 ;
        RECT 559.950 740.850 562.950 742.950 ;
        RECT 552.450 737.100 554.250 737.400 ;
        RECT 552.450 736.800 560.850 737.100 ;
        RECT 543.150 736.200 560.850 736.800 ;
        RECT 543.150 735.600 554.250 736.200 ;
        RECT 446.550 723.750 448.350 729.600 ;
        RECT 449.550 723.750 451.350 729.600 ;
        RECT 463.650 723.750 465.450 735.600 ;
        RECT 466.650 734.700 474.450 735.600 ;
        RECT 466.650 723.750 468.450 734.700 ;
        RECT 469.650 723.750 471.450 733.800 ;
        RECT 472.650 723.750 474.450 734.700 ;
        RECT 482.550 734.700 490.350 735.600 ;
        RECT 482.550 723.750 484.350 734.700 ;
        RECT 485.550 723.750 487.350 733.800 ;
        RECT 488.550 723.750 490.350 734.700 ;
        RECT 491.550 723.750 493.350 735.600 ;
        RECT 504.300 723.750 506.100 735.600 ;
        RECT 508.500 723.750 510.300 735.600 ;
        RECT 511.800 723.750 513.600 729.600 ;
        RECT 530.400 723.750 532.200 729.600 ;
        RECT 533.700 723.750 535.500 735.600 ;
        RECT 537.900 723.750 539.700 735.600 ;
        RECT 543.150 723.750 544.950 735.600 ;
        RECT 557.250 734.700 559.050 735.300 ;
        RECT 551.550 733.500 559.050 734.700 ;
        RECT 559.950 734.100 560.850 736.200 ;
        RECT 562.050 736.200 562.950 740.850 ;
        RECT 572.250 737.400 574.050 739.200 ;
        RECT 568.950 736.200 573.150 737.400 ;
        RECT 562.050 735.300 568.050 736.200 ;
        RECT 568.950 735.300 571.050 736.200 ;
        RECT 575.250 735.600 576.450 745.050 ;
        RECT 567.150 734.400 568.050 735.300 ;
        RECT 564.450 734.100 566.250 734.400 ;
        RECT 551.550 732.600 552.750 733.500 ;
        RECT 559.950 733.200 566.250 734.100 ;
        RECT 564.450 732.600 566.250 733.200 ;
        RECT 567.150 732.600 569.850 734.400 ;
        RECT 547.950 730.500 552.750 732.600 ;
        RECT 555.150 730.500 562.050 732.300 ;
        RECT 551.550 729.600 552.750 730.500 ;
        RECT 546.150 723.750 547.950 729.600 ;
        RECT 551.250 723.750 553.050 729.600 ;
        RECT 556.050 723.750 557.850 729.600 ;
        RECT 559.050 723.750 560.850 730.500 ;
        RECT 567.150 729.600 571.050 731.700 ;
        RECT 562.950 723.750 564.750 729.600 ;
        RECT 567.150 723.750 568.950 729.600 ;
        RECT 571.650 723.750 573.450 726.600 ;
        RECT 574.650 723.750 576.450 735.600 ;
        RECT 578.550 749.400 580.350 755.250 ;
        RECT 581.850 752.400 583.650 755.250 ;
        RECT 586.350 752.400 588.150 755.250 ;
        RECT 590.550 752.400 592.350 755.250 ;
        RECT 594.450 752.400 596.250 755.250 ;
        RECT 597.750 752.400 599.550 755.250 ;
        RECT 602.250 753.300 604.050 755.250 ;
        RECT 602.250 752.400 606.000 753.300 ;
        RECT 607.050 752.400 608.850 755.250 ;
        RECT 586.650 751.500 587.700 752.400 ;
        RECT 583.950 750.300 587.700 751.500 ;
        RECT 595.200 750.600 596.250 752.400 ;
        RECT 604.950 751.500 606.000 752.400 ;
        RECT 583.950 749.400 586.050 750.300 ;
        RECT 578.550 747.150 579.750 749.400 ;
        RECT 591.150 748.200 592.950 750.000 ;
        RECT 595.200 749.550 600.150 750.600 ;
        RECT 598.350 748.800 600.150 749.550 ;
        RECT 601.650 748.800 603.450 750.600 ;
        RECT 604.950 749.400 607.050 751.500 ;
        RECT 610.050 749.400 611.850 755.250 ;
        RECT 622.650 749.400 624.450 755.250 ;
        RECT 592.050 747.900 592.950 748.200 ;
        RECT 602.100 747.900 603.150 748.800 ;
        RECT 578.550 745.050 583.050 747.150 ;
        RECT 592.050 747.000 603.150 747.900 ;
        RECT 578.550 735.600 579.750 745.050 ;
        RECT 580.950 743.250 584.850 745.050 ;
        RECT 580.950 742.950 583.050 743.250 ;
        RECT 592.050 742.950 592.950 747.000 ;
        RECT 602.100 745.800 603.150 747.000 ;
        RECT 602.100 744.600 609.000 745.800 ;
        RECT 602.100 744.000 603.900 744.600 ;
        RECT 608.100 743.850 609.000 744.600 ;
        RECT 605.100 742.950 606.900 743.700 ;
        RECT 592.050 740.850 595.050 742.950 ;
        RECT 598.950 741.900 606.900 742.950 ;
        RECT 608.100 742.050 609.900 743.850 ;
        RECT 598.950 740.850 601.050 741.900 ;
        RECT 580.950 737.400 582.750 739.200 ;
        RECT 581.850 736.200 586.050 737.400 ;
        RECT 592.050 736.200 592.950 740.850 ;
        RECT 600.750 737.100 602.550 737.400 ;
        RECT 578.550 723.750 580.350 735.600 ;
        RECT 583.950 735.300 586.050 736.200 ;
        RECT 586.950 735.300 592.950 736.200 ;
        RECT 594.150 736.800 602.550 737.100 ;
        RECT 610.950 736.800 611.850 749.400 ;
        RECT 623.250 747.300 624.450 749.400 ;
        RECT 625.650 750.300 627.450 755.250 ;
        RECT 628.650 751.200 630.450 755.250 ;
        RECT 631.650 750.300 633.450 755.250 ;
        RECT 625.650 748.950 633.450 750.300 ;
        RECT 641.850 749.400 643.650 755.250 ;
        RECT 646.350 748.200 648.150 755.250 ;
        RECT 644.550 747.300 648.150 748.200 ;
        RECT 662.850 748.200 664.650 755.250 ;
        RECT 667.350 749.400 669.150 755.250 ;
        RECT 662.850 747.300 666.450 748.200 ;
        RECT 623.250 746.250 627.000 747.300 ;
        RECT 625.950 742.950 627.150 746.250 ;
        RECT 629.100 744.150 630.900 745.950 ;
        RECT 625.950 740.850 628.050 742.950 ;
        RECT 628.950 742.050 631.050 744.150 ;
        RECT 631.950 740.850 634.050 742.950 ;
        RECT 641.100 741.150 642.900 742.950 ;
        RECT 622.950 737.850 625.050 739.950 ;
        RECT 594.150 736.200 611.850 736.800 ;
        RECT 586.950 734.400 587.850 735.300 ;
        RECT 585.150 732.600 587.850 734.400 ;
        RECT 588.750 734.100 590.550 734.400 ;
        RECT 594.150 734.100 595.050 736.200 ;
        RECT 600.750 735.600 611.850 736.200 ;
        RECT 623.250 736.050 625.050 737.850 ;
        RECT 626.850 735.600 628.050 740.850 ;
        RECT 632.100 739.050 633.900 740.850 ;
        RECT 640.950 739.050 643.050 741.150 ;
        RECT 644.550 739.950 645.750 747.300 ;
        RECT 647.100 741.150 648.900 742.950 ;
        RECT 662.100 741.150 663.900 742.950 ;
        RECT 643.950 737.850 646.050 739.950 ;
        RECT 646.950 739.050 649.050 741.150 ;
        RECT 661.950 739.050 664.050 741.150 ;
        RECT 665.250 739.950 666.450 747.300 ;
        RECT 677.550 747.900 679.350 755.250 ;
        RECT 682.050 749.400 683.850 755.250 ;
        RECT 685.050 750.900 686.850 755.250 ;
        RECT 685.050 749.400 688.350 750.900 ;
        RECT 683.250 747.900 685.050 748.500 ;
        RECT 677.550 746.700 685.050 747.900 ;
        RECT 668.100 741.150 669.900 742.950 ;
        RECT 664.950 737.850 667.050 739.950 ;
        RECT 667.950 739.050 670.050 741.150 ;
        RECT 676.950 740.850 679.050 742.950 ;
        RECT 677.100 739.050 678.900 740.850 ;
        RECT 588.750 733.200 595.050 734.100 ;
        RECT 595.950 734.700 597.750 735.300 ;
        RECT 595.950 733.500 603.450 734.700 ;
        RECT 588.750 732.600 590.550 733.200 ;
        RECT 602.250 732.600 603.450 733.500 ;
        RECT 583.950 729.600 587.850 731.700 ;
        RECT 592.950 730.500 599.850 732.300 ;
        RECT 602.250 730.500 607.050 732.600 ;
        RECT 581.550 723.750 583.350 726.600 ;
        RECT 586.050 723.750 587.850 729.600 ;
        RECT 590.250 723.750 592.050 729.600 ;
        RECT 594.150 723.750 595.950 730.500 ;
        RECT 602.250 729.600 603.450 730.500 ;
        RECT 597.150 723.750 598.950 729.600 ;
        RECT 601.950 723.750 603.750 729.600 ;
        RECT 607.050 723.750 608.850 729.600 ;
        RECT 610.050 723.750 611.850 735.600 ;
        RECT 623.400 723.750 625.200 729.600 ;
        RECT 626.700 723.750 628.500 735.600 ;
        RECT 630.900 723.750 632.700 735.600 ;
        RECT 644.550 729.600 645.750 737.850 ;
        RECT 665.250 729.600 666.450 737.850 ;
        RECT 680.700 729.600 681.900 746.700 ;
        RECT 687.150 742.950 688.350 749.400 ;
        RECT 701.550 750.300 703.350 755.250 ;
        RECT 704.550 751.200 706.350 755.250 ;
        RECT 707.550 750.300 709.350 755.250 ;
        RECT 701.550 748.950 709.350 750.300 ;
        RECT 710.550 749.400 712.350 755.250 ;
        RECT 722.550 752.400 724.350 755.250 ;
        RECT 710.550 747.300 711.750 749.400 ;
        RECT 723.150 748.500 724.350 752.400 ;
        RECT 725.850 749.400 727.650 755.250 ;
        RECT 728.850 749.400 730.650 755.250 ;
        RECT 742.650 754.500 750.450 755.250 ;
        RECT 742.650 749.400 744.450 754.500 ;
        RECT 745.650 749.400 747.450 753.600 ;
        RECT 748.650 750.000 750.450 754.500 ;
        RECT 751.650 750.900 753.450 755.250 ;
        RECT 754.650 750.000 756.450 755.250 ;
        RECT 723.150 747.600 728.250 748.500 ;
        RECT 708.000 746.250 711.750 747.300 ;
        RECT 726.000 746.700 728.250 747.600 ;
        RECT 704.100 744.150 705.900 745.950 ;
        RECT 683.100 741.150 684.900 742.950 ;
        RECT 682.950 739.050 685.050 741.150 ;
        RECT 685.950 740.850 688.350 742.950 ;
        RECT 700.950 740.850 703.050 742.950 ;
        RECT 703.950 742.050 706.050 744.150 ;
        RECT 707.850 742.950 709.050 746.250 ;
        RECT 706.950 740.850 709.050 742.950 ;
        RECT 721.950 740.850 724.050 742.950 ;
        RECT 687.150 735.600 688.350 740.850 ;
        RECT 701.100 739.050 702.900 740.850 ;
        RECT 706.950 735.600 708.150 740.850 ;
        RECT 709.950 737.850 712.050 739.950 ;
        RECT 722.100 739.050 723.900 740.850 ;
        RECT 726.000 738.300 727.050 746.700 ;
        RECT 729.150 742.950 730.350 749.400 ;
        RECT 746.250 747.900 747.150 749.400 ;
        RECT 748.650 749.100 756.450 750.000 ;
        RECT 766.650 749.400 768.450 755.250 ;
        RECT 746.250 746.850 750.600 747.900 ;
        RECT 746.700 744.150 748.500 745.950 ;
        RECT 727.950 740.850 730.350 742.950 ;
        RECT 742.950 740.850 745.050 742.950 ;
        RECT 745.950 742.050 748.050 744.150 ;
        RECT 749.400 742.950 750.600 746.850 ;
        RECT 767.250 747.300 768.450 749.400 ;
        RECT 769.650 750.300 771.450 755.250 ;
        RECT 772.650 751.200 774.450 755.250 ;
        RECT 775.650 750.300 777.450 755.250 ;
        RECT 769.650 748.950 777.450 750.300 ;
        RECT 779.550 749.400 781.350 755.250 ;
        RECT 782.850 752.400 784.650 755.250 ;
        RECT 787.350 752.400 789.150 755.250 ;
        RECT 791.550 752.400 793.350 755.250 ;
        RECT 795.450 752.400 797.250 755.250 ;
        RECT 798.750 752.400 800.550 755.250 ;
        RECT 803.250 753.300 805.050 755.250 ;
        RECT 803.250 752.400 807.000 753.300 ;
        RECT 808.050 752.400 809.850 755.250 ;
        RECT 787.650 751.500 788.700 752.400 ;
        RECT 784.950 750.300 788.700 751.500 ;
        RECT 796.200 750.600 797.250 752.400 ;
        RECT 805.950 751.500 807.000 752.400 ;
        RECT 784.950 749.400 787.050 750.300 ;
        RECT 767.250 746.250 771.000 747.300 ;
        RECT 779.550 747.150 780.750 749.400 ;
        RECT 792.150 748.200 793.950 750.000 ;
        RECT 796.200 749.550 801.150 750.600 ;
        RECT 799.350 748.800 801.150 749.550 ;
        RECT 802.650 748.800 804.450 750.600 ;
        RECT 805.950 749.400 808.050 751.500 ;
        RECT 811.050 749.400 812.850 755.250 ;
        RECT 826.650 749.400 828.450 755.250 ;
        RECT 829.650 749.400 831.450 755.250 ;
        RECT 832.650 749.400 834.450 755.250 ;
        RECT 835.650 749.400 837.450 755.250 ;
        RECT 838.650 749.400 840.450 755.250 ;
        RECT 850.650 749.400 852.450 755.250 ;
        RECT 853.650 749.400 855.450 755.250 ;
        RECT 856.650 749.400 858.450 755.250 ;
        RECT 859.650 749.400 861.450 755.250 ;
        RECT 862.650 749.400 864.450 755.250 ;
        RECT 793.050 747.900 793.950 748.200 ;
        RECT 803.100 747.900 804.150 748.800 ;
        RECT 752.100 744.150 753.900 745.950 ;
        RECT 748.950 740.850 751.050 742.950 ;
        RECT 751.950 742.050 754.050 744.150 ;
        RECT 769.950 742.950 771.150 746.250 ;
        RECT 773.100 744.150 774.900 745.950 ;
        RECT 779.550 745.050 784.050 747.150 ;
        RECT 793.050 747.000 804.150 747.900 ;
        RECT 754.950 740.850 757.050 742.950 ;
        RECT 769.950 740.850 772.050 742.950 ;
        RECT 772.950 742.050 775.050 744.150 ;
        RECT 775.950 740.850 778.050 742.950 ;
        RECT 709.950 736.050 711.750 737.850 ;
        RECT 726.000 737.400 728.250 738.300 ;
        RECT 722.550 736.500 728.250 737.400 ;
        RECT 641.550 723.750 643.350 729.600 ;
        RECT 644.550 723.750 646.350 729.600 ;
        RECT 647.550 723.750 649.350 729.600 ;
        RECT 661.650 723.750 663.450 729.600 ;
        RECT 664.650 723.750 666.450 729.600 ;
        RECT 667.650 723.750 669.450 729.600 ;
        RECT 677.550 723.750 679.350 729.600 ;
        RECT 680.550 723.750 682.350 729.600 ;
        RECT 684.150 723.750 685.950 735.600 ;
        RECT 687.150 723.750 688.950 735.600 ;
        RECT 702.300 723.750 704.100 735.600 ;
        RECT 706.500 723.750 708.300 735.600 ;
        RECT 722.550 729.600 723.750 736.500 ;
        RECT 729.150 735.600 730.350 740.850 ;
        RECT 743.250 739.050 745.050 740.850 ;
        RECT 749.250 735.600 750.450 740.850 ;
        RECT 755.100 739.050 756.900 740.850 ;
        RECT 766.950 737.850 769.050 739.950 ;
        RECT 767.250 736.050 769.050 737.850 ;
        RECT 770.850 735.600 772.050 740.850 ;
        RECT 776.100 739.050 777.900 740.850 ;
        RECT 779.550 735.600 780.750 745.050 ;
        RECT 781.950 743.250 785.850 745.050 ;
        RECT 781.950 742.950 784.050 743.250 ;
        RECT 793.050 742.950 793.950 747.000 ;
        RECT 803.100 745.800 804.150 747.000 ;
        RECT 803.100 744.600 810.000 745.800 ;
        RECT 803.100 744.000 804.900 744.600 ;
        RECT 809.100 743.850 810.000 744.600 ;
        RECT 806.100 742.950 807.900 743.700 ;
        RECT 793.050 740.850 796.050 742.950 ;
        RECT 799.950 741.900 807.900 742.950 ;
        RECT 809.100 742.050 810.900 743.850 ;
        RECT 799.950 740.850 802.050 741.900 ;
        RECT 781.950 737.400 783.750 739.200 ;
        RECT 782.850 736.200 787.050 737.400 ;
        RECT 793.050 736.200 793.950 740.850 ;
        RECT 801.750 737.100 803.550 737.400 ;
        RECT 709.800 723.750 711.600 729.600 ;
        RECT 722.550 723.750 724.350 729.600 ;
        RECT 725.850 723.750 727.650 735.600 ;
        RECT 728.850 723.750 730.650 735.600 ;
        RECT 744.150 723.750 745.950 735.600 ;
        RECT 748.650 723.750 751.950 735.600 ;
        RECT 754.650 723.750 756.450 735.600 ;
        RECT 767.400 723.750 769.200 729.600 ;
        RECT 770.700 723.750 772.500 735.600 ;
        RECT 774.900 723.750 776.700 735.600 ;
        RECT 779.550 723.750 781.350 735.600 ;
        RECT 784.950 735.300 787.050 736.200 ;
        RECT 787.950 735.300 793.950 736.200 ;
        RECT 795.150 736.800 803.550 737.100 ;
        RECT 811.950 736.800 812.850 749.400 ;
        RECT 830.250 748.500 831.450 749.400 ;
        RECT 836.250 748.500 837.450 749.400 ;
        RECT 853.800 748.500 855.600 749.400 ;
        RECT 859.800 748.500 861.600 749.400 ;
        RECT 865.650 748.500 867.450 755.250 ;
        RECT 868.650 749.400 870.450 755.250 ;
        RECT 871.650 749.400 873.450 755.250 ;
        RECT 874.650 749.400 876.450 755.250 ;
        RECT 871.800 748.500 873.600 749.400 ;
        RECT 830.250 747.300 837.450 748.500 ;
        RECT 852.900 748.350 855.600 748.500 ;
        RECT 852.750 747.300 855.600 748.350 ;
        RECT 857.700 747.300 861.600 748.500 ;
        RECT 863.700 747.300 867.450 748.500 ;
        RECT 869.550 747.300 873.600 748.500 ;
        RECT 830.250 742.950 831.450 747.300 ;
        RECT 852.750 744.150 853.800 747.300 ;
        RECT 857.700 746.400 858.900 747.300 ;
        RECT 863.700 746.400 864.900 747.300 ;
        RECT 869.550 746.400 870.750 747.300 ;
        RECT 854.700 744.600 858.900 746.400 ;
        RECT 860.700 744.600 864.900 746.400 ;
        RECT 866.700 744.600 870.750 746.400 ;
        RECT 829.950 740.850 832.050 742.950 ;
        RECT 835.950 740.850 838.050 742.950 ;
        RECT 850.950 742.050 853.800 744.150 ;
        RECT 795.150 736.200 812.850 736.800 ;
        RECT 787.950 734.400 788.850 735.300 ;
        RECT 786.150 732.600 788.850 734.400 ;
        RECT 789.750 734.100 791.550 734.400 ;
        RECT 795.150 734.100 796.050 736.200 ;
        RECT 801.750 735.600 812.850 736.200 ;
        RECT 830.250 737.400 831.450 740.850 ;
        RECT 836.100 739.050 837.900 740.850 ;
        RECT 852.750 737.700 853.800 742.050 ;
        RECT 857.700 737.700 858.900 744.600 ;
        RECT 863.700 737.700 864.900 744.600 ;
        RECT 869.550 737.700 870.750 744.600 ;
        RECT 872.100 744.150 873.900 745.950 ;
        RECT 871.950 742.050 874.050 744.150 ;
        RECT 830.250 736.500 837.450 737.400 ;
        RECT 852.750 736.500 855.450 737.700 ;
        RECT 857.700 736.500 861.450 737.700 ;
        RECT 863.700 736.500 867.450 737.700 ;
        RECT 869.550 736.500 873.450 737.700 ;
        RECT 830.250 735.600 831.450 736.500 ;
        RECT 789.750 733.200 796.050 734.100 ;
        RECT 796.950 734.700 798.750 735.300 ;
        RECT 796.950 733.500 804.450 734.700 ;
        RECT 789.750 732.600 791.550 733.200 ;
        RECT 803.250 732.600 804.450 733.500 ;
        RECT 784.950 729.600 788.850 731.700 ;
        RECT 793.950 730.500 800.850 732.300 ;
        RECT 803.250 730.500 808.050 732.600 ;
        RECT 782.550 723.750 784.350 726.600 ;
        RECT 787.050 723.750 788.850 729.600 ;
        RECT 791.250 723.750 793.050 729.600 ;
        RECT 795.150 723.750 796.950 730.500 ;
        RECT 803.250 729.600 804.450 730.500 ;
        RECT 798.150 723.750 799.950 729.600 ;
        RECT 802.950 723.750 804.750 729.600 ;
        RECT 808.050 723.750 809.850 729.600 ;
        RECT 811.050 723.750 812.850 735.600 ;
        RECT 826.650 723.750 828.450 735.600 ;
        RECT 829.650 723.750 831.450 735.600 ;
        RECT 832.650 723.750 834.450 735.600 ;
        RECT 835.650 723.750 837.450 736.500 ;
        RECT 838.650 723.750 840.450 735.600 ;
        RECT 850.650 723.750 852.450 735.600 ;
        RECT 853.650 723.750 855.450 736.500 ;
        RECT 856.650 723.750 858.450 735.600 ;
        RECT 859.650 723.750 861.450 736.500 ;
        RECT 862.650 723.750 864.450 735.600 ;
        RECT 865.650 723.750 867.450 736.500 ;
        RECT 868.650 723.750 870.450 735.600 ;
        RECT 871.650 723.750 873.450 736.500 ;
        RECT 874.650 723.750 876.450 735.600 ;
        RECT 10.650 713.400 12.450 719.250 ;
        RECT 13.650 713.400 15.450 719.250 ;
        RECT 16.650 713.400 18.450 719.250 ;
        RECT 31.650 713.400 33.450 719.250 ;
        RECT 34.650 714.000 36.450 719.250 ;
        RECT 14.250 705.150 15.450 713.400 ;
        RECT 32.250 713.100 33.450 713.400 ;
        RECT 37.650 713.400 39.450 719.250 ;
        RECT 40.650 713.400 42.450 719.250 ;
        RECT 52.650 713.400 54.450 719.250 ;
        RECT 55.650 713.400 57.450 719.250 ;
        RECT 37.650 713.100 39.300 713.400 ;
        RECT 32.250 712.200 39.300 713.100 ;
        RECT 10.950 701.850 13.050 703.950 ;
        RECT 13.950 703.050 16.050 705.150 ;
        RECT 32.250 703.950 33.300 712.200 ;
        RECT 38.100 708.150 39.900 709.950 ;
        RECT 34.950 705.150 36.750 706.950 ;
        RECT 37.950 706.050 40.050 708.150 ;
        RECT 41.100 705.150 42.900 706.950 ;
        RECT 11.100 700.050 12.900 701.850 ;
        RECT 14.250 695.700 15.450 703.050 ;
        RECT 16.950 701.850 19.050 703.950 ;
        RECT 31.950 701.850 34.050 703.950 ;
        RECT 34.950 703.050 37.050 705.150 ;
        RECT 40.950 703.050 43.050 705.150 ;
        RECT 17.100 700.050 18.900 701.850 ;
        RECT 32.400 697.650 33.600 701.850 ;
        RECT 53.400 700.950 54.600 713.400 ;
        RECT 67.050 707.400 68.850 719.250 ;
        RECT 70.050 707.400 71.850 719.250 ;
        RECT 73.650 713.400 75.450 719.250 ;
        RECT 76.650 713.400 78.450 719.250 ;
        RECT 67.650 702.150 68.850 707.400 ;
        RECT 52.950 698.850 55.050 700.950 ;
        RECT 56.100 699.150 57.900 700.950 ;
        RECT 67.650 700.050 70.050 702.150 ;
        RECT 70.950 701.850 73.050 703.950 ;
        RECT 71.100 700.050 72.900 701.850 ;
        RECT 32.400 696.000 36.900 697.650 ;
        RECT 11.850 694.800 15.450 695.700 ;
        RECT 11.850 687.750 13.650 694.800 ;
        RECT 16.350 687.750 18.150 693.600 ;
        RECT 35.100 687.750 36.900 696.000 ;
        RECT 40.500 687.750 42.300 696.600 ;
        RECT 53.400 690.600 54.600 698.850 ;
        RECT 55.950 697.050 58.050 699.150 ;
        RECT 67.650 693.600 68.850 700.050 ;
        RECT 74.100 696.300 75.300 713.400 ;
        RECT 87.300 707.400 89.100 719.250 ;
        RECT 91.500 707.400 93.300 719.250 ;
        RECT 94.800 713.400 96.600 719.250 ;
        RECT 109.650 707.400 111.450 719.250 ;
        RECT 112.650 708.300 114.450 719.250 ;
        RECT 115.650 709.200 117.450 719.250 ;
        RECT 118.650 708.300 120.450 719.250 ;
        RECT 131.550 713.400 133.350 719.250 ;
        RECT 134.550 713.400 136.350 719.250 ;
        RECT 137.550 714.000 139.350 719.250 ;
        RECT 134.700 713.100 136.350 713.400 ;
        RECT 140.550 713.400 142.350 719.250 ;
        RECT 140.550 713.100 141.750 713.400 ;
        RECT 134.700 712.200 141.750 713.100 ;
        RECT 112.650 707.400 120.450 708.300 ;
        RECT 134.100 708.150 135.900 709.950 ;
        RECT 77.100 702.150 78.900 703.950 ;
        RECT 86.100 702.150 87.900 703.950 ;
        RECT 91.950 702.150 93.150 707.400 ;
        RECT 94.950 705.150 96.750 706.950 ;
        RECT 94.950 703.050 97.050 705.150 ;
        RECT 110.100 702.150 111.300 707.400 ;
        RECT 131.100 705.150 132.900 706.950 ;
        RECT 133.950 706.050 136.050 708.150 ;
        RECT 137.250 705.150 139.050 706.950 ;
        RECT 130.950 703.050 133.050 705.150 ;
        RECT 136.950 703.050 139.050 705.150 ;
        RECT 140.700 703.950 141.750 712.200 ;
        RECT 157.650 707.400 159.450 719.250 ;
        RECT 160.650 707.400 162.450 719.250 ;
        RECT 172.050 707.400 173.850 719.250 ;
        RECT 175.050 707.400 176.850 719.250 ;
        RECT 178.650 713.400 180.450 719.250 ;
        RECT 181.650 713.400 183.450 719.250 ;
        RECT 76.950 700.050 79.050 702.150 ;
        RECT 85.950 700.050 88.050 702.150 ;
        RECT 88.950 698.850 91.050 700.950 ;
        RECT 91.950 700.050 94.050 702.150 ;
        RECT 109.950 700.050 112.050 702.150 ;
        RECT 139.950 701.850 142.050 703.950 ;
        RECT 158.400 702.150 159.600 707.400 ;
        RECT 172.650 702.150 173.850 707.400 ;
        RECT 89.100 697.050 90.900 698.850 ;
        RECT 92.850 696.750 94.050 700.050 ;
        RECT 70.950 695.100 78.450 696.300 ;
        RECT 93.000 695.700 96.750 696.750 ;
        RECT 70.950 694.500 72.750 695.100 ;
        RECT 67.650 692.100 70.950 693.600 ;
        RECT 52.650 687.750 54.450 690.600 ;
        RECT 55.650 687.750 57.450 690.600 ;
        RECT 69.150 687.750 70.950 692.100 ;
        RECT 72.150 687.750 73.950 693.600 ;
        RECT 76.650 687.750 78.450 695.100 ;
        RECT 86.550 692.700 94.350 694.050 ;
        RECT 86.550 687.750 88.350 692.700 ;
        RECT 89.550 687.750 91.350 691.800 ;
        RECT 92.550 687.750 94.350 692.700 ;
        RECT 95.550 693.600 96.750 695.700 ;
        RECT 110.100 693.600 111.300 700.050 ;
        RECT 112.950 698.850 115.050 700.950 ;
        RECT 116.100 699.150 117.900 700.950 ;
        RECT 113.100 697.050 114.900 698.850 ;
        RECT 115.950 697.050 118.050 699.150 ;
        RECT 118.950 698.850 121.050 700.950 ;
        RECT 119.100 697.050 120.900 698.850 ;
        RECT 140.400 697.650 141.600 701.850 ;
        RECT 157.950 700.050 160.050 702.150 ;
        RECT 95.550 687.750 97.350 693.600 ;
        RECT 110.100 691.950 115.800 693.600 ;
        RECT 110.700 687.750 112.500 690.600 ;
        RECT 114.000 687.750 115.800 691.950 ;
        RECT 118.200 687.750 120.000 693.600 ;
        RECT 131.700 687.750 133.500 696.600 ;
        RECT 137.100 696.000 141.600 697.650 ;
        RECT 137.100 687.750 138.900 696.000 ;
        RECT 158.400 693.600 159.600 700.050 ;
        RECT 160.950 698.850 163.050 700.950 ;
        RECT 172.650 700.050 175.050 702.150 ;
        RECT 175.950 701.850 178.050 703.950 ;
        RECT 176.100 700.050 177.900 701.850 ;
        RECT 161.100 697.050 162.900 698.850 ;
        RECT 172.650 693.600 173.850 700.050 ;
        RECT 179.100 696.300 180.300 713.400 ;
        RECT 193.650 707.400 195.450 719.250 ;
        RECT 196.650 708.300 198.450 719.250 ;
        RECT 199.650 709.200 201.450 719.250 ;
        RECT 202.650 708.300 204.450 719.250 ;
        RECT 196.650 707.400 204.450 708.300 ;
        RECT 214.650 707.400 216.450 719.250 ;
        RECT 217.650 708.300 219.450 719.250 ;
        RECT 220.650 709.200 222.450 719.250 ;
        RECT 223.650 708.300 225.450 719.250 ;
        RECT 238.650 713.400 240.450 719.250 ;
        RECT 241.650 713.400 243.450 719.250 ;
        RECT 217.650 707.400 225.450 708.300 ;
        RECT 182.100 702.150 183.900 703.950 ;
        RECT 194.100 702.150 195.300 707.400 ;
        RECT 215.100 702.150 216.300 707.400 ;
        RECT 181.950 700.050 184.050 702.150 ;
        RECT 193.950 700.050 196.050 702.150 ;
        RECT 175.950 695.100 183.450 696.300 ;
        RECT 175.950 694.500 177.750 695.100 ;
        RECT 157.650 687.750 159.450 693.600 ;
        RECT 160.650 687.750 162.450 693.600 ;
        RECT 172.650 692.100 175.950 693.600 ;
        RECT 174.150 687.750 175.950 692.100 ;
        RECT 177.150 687.750 178.950 693.600 ;
        RECT 181.650 687.750 183.450 695.100 ;
        RECT 194.100 693.600 195.300 700.050 ;
        RECT 196.950 698.850 199.050 700.950 ;
        RECT 200.100 699.150 201.900 700.950 ;
        RECT 197.100 697.050 198.900 698.850 ;
        RECT 199.950 697.050 202.050 699.150 ;
        RECT 202.950 698.850 205.050 700.950 ;
        RECT 214.950 700.050 217.050 702.150 ;
        RECT 239.400 700.950 240.600 713.400 ;
        RECT 246.150 707.400 247.950 719.250 ;
        RECT 249.150 713.400 250.950 719.250 ;
        RECT 254.250 713.400 256.050 719.250 ;
        RECT 259.050 713.400 260.850 719.250 ;
        RECT 254.550 712.500 255.750 713.400 ;
        RECT 262.050 712.500 263.850 719.250 ;
        RECT 265.950 713.400 267.750 719.250 ;
        RECT 270.150 713.400 271.950 719.250 ;
        RECT 274.650 716.400 276.450 719.250 ;
        RECT 250.950 710.400 255.750 712.500 ;
        RECT 258.150 710.700 265.050 712.500 ;
        RECT 270.150 711.300 274.050 713.400 ;
        RECT 254.550 709.500 255.750 710.400 ;
        RECT 267.450 709.800 269.250 710.400 ;
        RECT 254.550 708.300 262.050 709.500 ;
        RECT 260.250 707.700 262.050 708.300 ;
        RECT 262.950 708.900 269.250 709.800 ;
        RECT 246.150 706.800 257.250 707.400 ;
        RECT 262.950 706.800 263.850 708.900 ;
        RECT 267.450 708.600 269.250 708.900 ;
        RECT 270.150 708.600 272.850 710.400 ;
        RECT 270.150 707.700 271.050 708.600 ;
        RECT 246.150 706.200 263.850 706.800 ;
        RECT 203.100 697.050 204.900 698.850 ;
        RECT 215.100 693.600 216.300 700.050 ;
        RECT 217.950 698.850 220.050 700.950 ;
        RECT 221.100 699.150 222.900 700.950 ;
        RECT 218.100 697.050 219.900 698.850 ;
        RECT 220.950 697.050 223.050 699.150 ;
        RECT 223.950 698.850 226.050 700.950 ;
        RECT 238.950 698.850 241.050 700.950 ;
        RECT 242.100 699.150 243.900 700.950 ;
        RECT 224.100 697.050 225.900 698.850 ;
        RECT 194.100 691.950 199.800 693.600 ;
        RECT 194.700 687.750 196.500 690.600 ;
        RECT 198.000 687.750 199.800 691.950 ;
        RECT 202.200 687.750 204.000 693.600 ;
        RECT 215.100 691.950 220.800 693.600 ;
        RECT 215.700 687.750 217.500 690.600 ;
        RECT 219.000 687.750 220.800 691.950 ;
        RECT 223.200 687.750 225.000 693.600 ;
        RECT 239.400 690.600 240.600 698.850 ;
        RECT 241.950 697.050 244.050 699.150 ;
        RECT 246.150 693.600 247.050 706.200 ;
        RECT 255.450 705.900 263.850 706.200 ;
        RECT 265.050 706.800 271.050 707.700 ;
        RECT 271.950 706.800 274.050 707.700 ;
        RECT 277.650 707.400 279.450 719.250 ;
        RECT 289.650 713.400 291.450 719.250 ;
        RECT 292.650 713.400 294.450 719.250 ;
        RECT 255.450 705.600 257.250 705.900 ;
        RECT 265.050 702.150 265.950 706.800 ;
        RECT 271.950 705.600 276.150 706.800 ;
        RECT 275.250 703.800 277.050 705.600 ;
        RECT 256.950 701.100 259.050 702.150 ;
        RECT 248.100 699.150 249.900 700.950 ;
        RECT 251.100 700.050 259.050 701.100 ;
        RECT 262.950 700.050 265.950 702.150 ;
        RECT 251.100 699.300 252.900 700.050 ;
        RECT 249.000 698.400 249.900 699.150 ;
        RECT 254.100 698.400 255.900 699.000 ;
        RECT 249.000 697.200 255.900 698.400 ;
        RECT 254.850 696.000 255.900 697.200 ;
        RECT 265.050 696.000 265.950 700.050 ;
        RECT 274.950 699.750 277.050 700.050 ;
        RECT 273.150 697.950 277.050 699.750 ;
        RECT 278.250 697.950 279.450 707.400 ;
        RECT 290.400 700.950 291.600 713.400 ;
        RECT 307.050 707.400 308.850 719.250 ;
        RECT 310.050 707.400 311.850 719.250 ;
        RECT 313.650 713.400 315.450 719.250 ;
        RECT 316.650 713.400 318.450 719.250 ;
        RECT 326.550 713.400 328.350 719.250 ;
        RECT 329.550 713.400 331.350 719.250 ;
        RECT 347.400 713.400 349.200 719.250 ;
        RECT 307.650 702.150 308.850 707.400 ;
        RECT 289.950 698.850 292.050 700.950 ;
        RECT 293.100 699.150 294.900 700.950 ;
        RECT 307.650 700.050 310.050 702.150 ;
        RECT 310.950 701.850 313.050 703.950 ;
        RECT 311.100 700.050 312.900 701.850 ;
        RECT 254.850 695.100 265.950 696.000 ;
        RECT 274.950 695.850 279.450 697.950 ;
        RECT 254.850 694.200 255.900 695.100 ;
        RECT 265.050 694.800 265.950 695.100 ;
        RECT 238.650 687.750 240.450 690.600 ;
        RECT 241.650 687.750 243.450 690.600 ;
        RECT 246.150 687.750 247.950 693.600 ;
        RECT 250.950 691.500 253.050 693.600 ;
        RECT 254.550 692.400 256.350 694.200 ;
        RECT 257.850 693.450 259.650 694.200 ;
        RECT 257.850 692.400 262.800 693.450 ;
        RECT 265.050 693.000 266.850 694.800 ;
        RECT 278.250 693.600 279.450 695.850 ;
        RECT 271.950 692.700 274.050 693.600 ;
        RECT 252.000 690.600 253.050 691.500 ;
        RECT 261.750 690.600 262.800 692.400 ;
        RECT 270.300 691.500 274.050 692.700 ;
        RECT 270.300 690.600 271.350 691.500 ;
        RECT 249.150 687.750 250.950 690.600 ;
        RECT 252.000 689.700 255.750 690.600 ;
        RECT 253.950 687.750 255.750 689.700 ;
        RECT 258.450 687.750 260.250 690.600 ;
        RECT 261.750 687.750 263.550 690.600 ;
        RECT 265.650 687.750 267.450 690.600 ;
        RECT 269.850 687.750 271.650 690.600 ;
        RECT 274.350 687.750 276.150 690.600 ;
        RECT 277.650 687.750 279.450 693.600 ;
        RECT 290.400 690.600 291.600 698.850 ;
        RECT 292.950 697.050 295.050 699.150 ;
        RECT 307.650 693.600 308.850 700.050 ;
        RECT 314.100 696.300 315.300 713.400 ;
        RECT 317.100 702.150 318.900 703.950 ;
        RECT 316.950 700.050 319.050 702.150 ;
        RECT 329.400 700.950 330.600 713.400 ;
        RECT 350.700 707.400 352.500 719.250 ;
        RECT 354.900 707.400 356.700 719.250 ;
        RECT 365.550 713.400 367.350 719.250 ;
        RECT 368.550 713.400 370.350 719.250 ;
        RECT 371.550 713.400 373.350 719.250 ;
        RECT 347.250 705.150 349.050 706.950 ;
        RECT 346.950 703.050 349.050 705.150 ;
        RECT 350.850 702.150 352.050 707.400 ;
        RECT 368.550 705.150 369.750 713.400 ;
        RECT 387.300 707.400 389.100 719.250 ;
        RECT 391.500 707.400 393.300 719.250 ;
        RECT 394.800 713.400 396.600 719.250 ;
        RECT 409.650 713.400 411.450 719.250 ;
        RECT 412.650 713.400 414.450 719.250 ;
        RECT 415.650 713.400 417.450 719.250 ;
        RECT 431.400 713.400 433.200 719.250 ;
        RECT 356.100 702.150 357.900 703.950 ;
        RECT 326.100 699.150 327.900 700.950 ;
        RECT 325.950 697.050 328.050 699.150 ;
        RECT 328.950 698.850 331.050 700.950 ;
        RECT 349.950 700.050 352.050 702.150 ;
        RECT 310.950 695.100 318.450 696.300 ;
        RECT 310.950 694.500 312.750 695.100 ;
        RECT 307.650 692.100 310.950 693.600 ;
        RECT 289.650 687.750 291.450 690.600 ;
        RECT 292.650 687.750 294.450 690.600 ;
        RECT 309.150 687.750 310.950 692.100 ;
        RECT 312.150 687.750 313.950 693.600 ;
        RECT 316.650 687.750 318.450 695.100 ;
        RECT 329.400 690.600 330.600 698.850 ;
        RECT 349.950 696.750 351.150 700.050 ;
        RECT 352.950 698.850 355.050 700.950 ;
        RECT 355.950 700.050 358.050 702.150 ;
        RECT 364.950 701.850 367.050 703.950 ;
        RECT 367.950 703.050 370.050 705.150 ;
        RECT 365.100 700.050 366.900 701.850 ;
        RECT 353.100 697.050 354.900 698.850 ;
        RECT 347.250 695.700 351.000 696.750 ;
        RECT 368.550 695.700 369.750 703.050 ;
        RECT 370.950 701.850 373.050 703.950 ;
        RECT 386.100 702.150 387.900 703.950 ;
        RECT 391.950 702.150 393.150 707.400 ;
        RECT 394.950 705.150 396.750 706.950 ;
        RECT 413.250 705.150 414.450 713.400 ;
        RECT 434.700 707.400 436.500 719.250 ;
        RECT 438.900 707.400 440.700 719.250 ;
        RECT 454.650 713.400 456.450 719.250 ;
        RECT 457.650 713.400 459.450 719.250 ;
        RECT 470.400 713.400 472.200 719.250 ;
        RECT 431.250 705.150 433.050 706.950 ;
        RECT 394.950 703.050 397.050 705.150 ;
        RECT 371.100 700.050 372.900 701.850 ;
        RECT 385.950 700.050 388.050 702.150 ;
        RECT 388.950 698.850 391.050 700.950 ;
        RECT 391.950 700.050 394.050 702.150 ;
        RECT 409.950 701.850 412.050 703.950 ;
        RECT 412.950 703.050 415.050 705.150 ;
        RECT 410.100 700.050 411.900 701.850 ;
        RECT 389.100 697.050 390.900 698.850 ;
        RECT 392.850 696.750 394.050 700.050 ;
        RECT 393.000 695.700 396.750 696.750 ;
        RECT 413.250 695.700 414.450 703.050 ;
        RECT 415.950 701.850 418.050 703.950 ;
        RECT 430.950 703.050 433.050 705.150 ;
        RECT 434.850 702.150 436.050 707.400 ;
        RECT 440.100 702.150 441.900 703.950 ;
        RECT 416.100 700.050 417.900 701.850 ;
        RECT 433.950 700.050 436.050 702.150 ;
        RECT 433.950 696.750 435.150 700.050 ;
        RECT 436.950 698.850 439.050 700.950 ;
        RECT 439.950 700.050 442.050 702.150 ;
        RECT 455.400 700.950 456.600 713.400 ;
        RECT 473.700 707.400 475.500 719.250 ;
        RECT 477.900 707.400 479.700 719.250 ;
        RECT 491.400 713.400 493.200 719.250 ;
        RECT 494.700 707.400 496.500 719.250 ;
        RECT 498.900 707.400 500.700 719.250 ;
        RECT 513.450 707.400 515.250 719.250 ;
        RECT 517.650 707.400 519.450 719.250 ;
        RECT 532.650 713.400 534.450 719.250 ;
        RECT 535.650 713.400 537.450 719.250 ;
        RECT 538.650 713.400 540.450 719.250 ;
        RECT 548.550 713.400 550.350 719.250 ;
        RECT 551.550 713.400 553.350 719.250 ;
        RECT 470.250 705.150 472.050 706.950 ;
        RECT 469.950 703.050 472.050 705.150 ;
        RECT 473.850 702.150 475.050 707.400 ;
        RECT 491.250 705.150 493.050 706.950 ;
        RECT 479.100 702.150 480.900 703.950 ;
        RECT 490.950 703.050 493.050 705.150 ;
        RECT 494.850 702.150 496.050 707.400 ;
        RECT 513.450 706.350 516.000 707.400 ;
        RECT 500.100 702.150 501.900 703.950 ;
        RECT 512.100 702.150 513.900 703.950 ;
        RECT 454.950 698.850 457.050 700.950 ;
        RECT 458.100 699.150 459.900 700.950 ;
        RECT 472.950 700.050 475.050 702.150 ;
        RECT 437.100 697.050 438.900 698.850 ;
        RECT 347.250 693.600 348.450 695.700 ;
        RECT 368.550 694.800 372.150 695.700 ;
        RECT 326.550 687.750 328.350 690.600 ;
        RECT 329.550 687.750 331.350 690.600 ;
        RECT 346.650 687.750 348.450 693.600 ;
        RECT 349.650 692.700 357.450 694.050 ;
        RECT 349.650 687.750 351.450 692.700 ;
        RECT 352.650 687.750 354.450 691.800 ;
        RECT 355.650 687.750 357.450 692.700 ;
        RECT 365.850 687.750 367.650 693.600 ;
        RECT 370.350 687.750 372.150 694.800 ;
        RECT 386.550 692.700 394.350 694.050 ;
        RECT 386.550 687.750 388.350 692.700 ;
        RECT 389.550 687.750 391.350 691.800 ;
        RECT 392.550 687.750 394.350 692.700 ;
        RECT 395.550 693.600 396.750 695.700 ;
        RECT 410.850 694.800 414.450 695.700 ;
        RECT 431.250 695.700 435.000 696.750 ;
        RECT 439.950 696.450 442.050 697.050 ;
        RECT 445.950 696.450 448.050 697.050 ;
        RECT 395.550 687.750 397.350 693.600 ;
        RECT 410.850 687.750 412.650 694.800 ;
        RECT 431.250 693.600 432.450 695.700 ;
        RECT 439.950 695.550 448.050 696.450 ;
        RECT 439.950 694.950 442.050 695.550 ;
        RECT 445.950 694.950 448.050 695.550 ;
        RECT 415.350 687.750 417.150 693.600 ;
        RECT 430.650 687.750 432.450 693.600 ;
        RECT 433.650 692.700 441.450 694.050 ;
        RECT 433.650 687.750 435.450 692.700 ;
        RECT 436.650 687.750 438.450 691.800 ;
        RECT 439.650 687.750 441.450 692.700 ;
        RECT 455.400 690.600 456.600 698.850 ;
        RECT 457.950 697.050 460.050 699.150 ;
        RECT 472.950 696.750 474.150 700.050 ;
        RECT 475.950 698.850 478.050 700.950 ;
        RECT 478.950 700.050 481.050 702.150 ;
        RECT 493.950 700.050 496.050 702.150 ;
        RECT 476.100 697.050 477.900 698.850 ;
        RECT 493.950 696.750 495.150 700.050 ;
        RECT 496.950 698.850 499.050 700.950 ;
        RECT 499.950 700.050 502.050 702.150 ;
        RECT 511.950 700.050 514.050 702.150 ;
        RECT 514.950 699.150 516.000 706.350 ;
        RECT 536.250 705.150 537.450 713.400 ;
        RECT 518.100 702.150 519.900 703.950 ;
        RECT 517.950 700.050 520.050 702.150 ;
        RECT 532.950 701.850 535.050 703.950 ;
        RECT 535.950 703.050 538.050 705.150 ;
        RECT 533.100 700.050 534.900 701.850 ;
        RECT 497.100 697.050 498.900 698.850 ;
        RECT 514.950 697.050 517.050 699.150 ;
        RECT 470.250 695.700 474.000 696.750 ;
        RECT 491.250 695.700 495.000 696.750 ;
        RECT 470.250 693.600 471.450 695.700 ;
        RECT 454.650 687.750 456.450 690.600 ;
        RECT 457.650 687.750 459.450 690.600 ;
        RECT 469.650 687.750 471.450 693.600 ;
        RECT 472.650 692.700 480.450 694.050 ;
        RECT 491.250 693.600 492.450 695.700 ;
        RECT 472.650 687.750 474.450 692.700 ;
        RECT 475.650 687.750 477.450 691.800 ;
        RECT 478.650 687.750 480.450 692.700 ;
        RECT 490.650 687.750 492.450 693.600 ;
        RECT 493.650 692.700 501.450 694.050 ;
        RECT 493.650 687.750 495.450 692.700 ;
        RECT 496.650 687.750 498.450 691.800 ;
        RECT 499.650 687.750 501.450 692.700 ;
        RECT 514.950 690.600 516.000 697.050 ;
        RECT 536.250 695.700 537.450 703.050 ;
        RECT 538.950 701.850 541.050 703.950 ;
        RECT 539.100 700.050 540.900 701.850 ;
        RECT 551.400 700.950 552.600 713.400 ;
        RECT 566.550 707.400 568.350 719.250 ;
        RECT 570.750 707.400 572.550 719.250 ;
        RECT 588.300 707.400 590.100 719.250 ;
        RECT 592.500 707.400 594.300 719.250 ;
        RECT 595.800 713.400 597.600 719.250 ;
        RECT 603.150 707.400 604.950 719.250 ;
        RECT 606.150 713.400 607.950 719.250 ;
        RECT 611.250 713.400 613.050 719.250 ;
        RECT 616.050 713.400 617.850 719.250 ;
        RECT 611.550 712.500 612.750 713.400 ;
        RECT 619.050 712.500 620.850 719.250 ;
        RECT 622.950 713.400 624.750 719.250 ;
        RECT 627.150 713.400 628.950 719.250 ;
        RECT 631.650 716.400 633.450 719.250 ;
        RECT 607.950 710.400 612.750 712.500 ;
        RECT 615.150 710.700 622.050 712.500 ;
        RECT 627.150 711.300 631.050 713.400 ;
        RECT 611.550 709.500 612.750 710.400 ;
        RECT 624.450 709.800 626.250 710.400 ;
        RECT 611.550 708.300 619.050 709.500 ;
        RECT 617.250 707.700 619.050 708.300 ;
        RECT 619.950 708.900 626.250 709.800 ;
        RECT 570.000 706.350 572.550 707.400 ;
        RECT 566.100 702.150 567.900 703.950 ;
        RECT 548.100 699.150 549.900 700.950 ;
        RECT 547.950 697.050 550.050 699.150 ;
        RECT 550.950 698.850 553.050 700.950 ;
        RECT 565.950 700.050 568.050 702.150 ;
        RECT 570.000 699.150 571.050 706.350 ;
        RECT 572.100 702.150 573.900 703.950 ;
        RECT 587.100 702.150 588.900 703.950 ;
        RECT 592.950 702.150 594.150 707.400 ;
        RECT 595.950 705.150 597.750 706.950 ;
        RECT 603.150 706.800 614.250 707.400 ;
        RECT 619.950 706.800 620.850 708.900 ;
        RECT 624.450 708.600 626.250 708.900 ;
        RECT 627.150 708.600 629.850 710.400 ;
        RECT 627.150 707.700 628.050 708.600 ;
        RECT 603.150 706.200 620.850 706.800 ;
        RECT 595.950 703.050 598.050 705.150 ;
        RECT 571.950 700.050 574.050 702.150 ;
        RECT 586.950 700.050 589.050 702.150 ;
        RECT 533.850 694.800 537.450 695.700 ;
        RECT 511.650 687.750 513.450 690.600 ;
        RECT 514.650 687.750 516.450 690.600 ;
        RECT 517.650 687.750 519.450 690.600 ;
        RECT 533.850 687.750 535.650 694.800 ;
        RECT 538.350 687.750 540.150 693.600 ;
        RECT 551.400 690.600 552.600 698.850 ;
        RECT 568.950 697.050 571.050 699.150 ;
        RECT 589.950 698.850 592.050 700.950 ;
        RECT 592.950 700.050 595.050 702.150 ;
        RECT 590.100 697.050 591.900 698.850 ;
        RECT 570.000 690.600 571.050 697.050 ;
        RECT 593.850 696.750 595.050 700.050 ;
        RECT 594.000 695.700 597.750 696.750 ;
        RECT 587.550 692.700 595.350 694.050 ;
        RECT 548.550 687.750 550.350 690.600 ;
        RECT 551.550 687.750 553.350 690.600 ;
        RECT 566.550 687.750 568.350 690.600 ;
        RECT 569.550 687.750 571.350 690.600 ;
        RECT 572.550 687.750 574.350 690.600 ;
        RECT 587.550 687.750 589.350 692.700 ;
        RECT 590.550 687.750 592.350 691.800 ;
        RECT 593.550 687.750 595.350 692.700 ;
        RECT 596.550 693.600 597.750 695.700 ;
        RECT 603.150 693.600 604.050 706.200 ;
        RECT 612.450 705.900 620.850 706.200 ;
        RECT 622.050 706.800 628.050 707.700 ;
        RECT 628.950 706.800 631.050 707.700 ;
        RECT 634.650 707.400 636.450 719.250 ;
        RECT 644.550 713.400 646.350 719.250 ;
        RECT 647.550 713.400 649.350 719.250 ;
        RECT 650.550 713.400 652.350 719.250 ;
        RECT 664.650 713.400 666.450 719.250 ;
        RECT 667.650 713.400 669.450 719.250 ;
        RECT 670.650 713.400 672.450 719.250 ;
        RECT 682.650 718.500 690.450 719.250 ;
        RECT 612.450 705.600 614.250 705.900 ;
        RECT 622.050 702.150 622.950 706.800 ;
        RECT 628.950 705.600 633.150 706.800 ;
        RECT 632.250 703.800 634.050 705.600 ;
        RECT 613.950 701.100 616.050 702.150 ;
        RECT 605.100 699.150 606.900 700.950 ;
        RECT 608.100 700.050 616.050 701.100 ;
        RECT 619.950 700.050 622.950 702.150 ;
        RECT 608.100 699.300 609.900 700.050 ;
        RECT 606.000 698.400 606.900 699.150 ;
        RECT 611.100 698.400 612.900 699.000 ;
        RECT 606.000 697.200 612.900 698.400 ;
        RECT 611.850 696.000 612.900 697.200 ;
        RECT 622.050 696.000 622.950 700.050 ;
        RECT 631.950 699.750 634.050 700.050 ;
        RECT 630.150 697.950 634.050 699.750 ;
        RECT 635.250 697.950 636.450 707.400 ;
        RECT 647.550 705.150 648.750 713.400 ;
        RECT 668.250 705.150 669.450 713.400 ;
        RECT 682.650 707.400 684.450 718.500 ;
        RECT 685.650 707.400 687.450 717.600 ;
        RECT 688.650 708.600 690.450 718.500 ;
        RECT 691.650 709.500 693.450 719.250 ;
        RECT 694.650 708.600 696.450 719.250 ;
        RECT 688.650 707.700 696.450 708.600 ;
        RECT 698.550 707.400 700.350 719.250 ;
        RECT 701.550 716.400 703.350 719.250 ;
        RECT 706.050 713.400 707.850 719.250 ;
        RECT 710.250 713.400 712.050 719.250 ;
        RECT 703.950 711.300 707.850 713.400 ;
        RECT 714.150 712.500 715.950 719.250 ;
        RECT 717.150 713.400 718.950 719.250 ;
        RECT 721.950 713.400 723.750 719.250 ;
        RECT 727.050 713.400 728.850 719.250 ;
        RECT 722.250 712.500 723.450 713.400 ;
        RECT 712.950 710.700 719.850 712.500 ;
        RECT 722.250 710.400 727.050 712.500 ;
        RECT 705.150 708.600 707.850 710.400 ;
        RECT 708.750 709.800 710.550 710.400 ;
        RECT 708.750 708.900 715.050 709.800 ;
        RECT 722.250 709.500 723.450 710.400 ;
        RECT 708.750 708.600 710.550 708.900 ;
        RECT 706.950 707.700 707.850 708.600 ;
        RECT 685.800 706.500 687.600 707.400 ;
        RECT 685.800 705.600 689.850 706.500 ;
        RECT 643.950 701.850 646.050 703.950 ;
        RECT 646.950 703.050 649.050 705.150 ;
        RECT 644.100 700.050 645.900 701.850 ;
        RECT 611.850 695.100 622.950 696.000 ;
        RECT 631.950 695.850 636.450 697.950 ;
        RECT 611.850 694.200 612.900 695.100 ;
        RECT 622.050 694.800 622.950 695.100 ;
        RECT 596.550 687.750 598.350 693.600 ;
        RECT 603.150 687.750 604.950 693.600 ;
        RECT 607.950 691.500 610.050 693.600 ;
        RECT 611.550 692.400 613.350 694.200 ;
        RECT 614.850 693.450 616.650 694.200 ;
        RECT 614.850 692.400 619.800 693.450 ;
        RECT 622.050 693.000 623.850 694.800 ;
        RECT 635.250 693.600 636.450 695.850 ;
        RECT 647.550 695.700 648.750 703.050 ;
        RECT 649.950 701.850 652.050 703.950 ;
        RECT 664.950 701.850 667.050 703.950 ;
        RECT 667.950 703.050 670.050 705.150 ;
        RECT 650.100 700.050 651.900 701.850 ;
        RECT 665.100 700.050 666.900 701.850 ;
        RECT 668.250 695.700 669.450 703.050 ;
        RECT 670.950 701.850 673.050 703.950 ;
        RECT 683.100 702.150 684.900 703.950 ;
        RECT 688.950 702.150 689.850 705.600 ;
        RECT 694.950 702.150 696.750 703.950 ;
        RECT 671.100 700.050 672.900 701.850 ;
        RECT 682.950 700.050 685.050 702.150 ;
        RECT 685.950 698.850 688.050 700.950 ;
        RECT 688.950 700.050 691.050 702.150 ;
        RECT 686.250 697.050 688.050 698.850 ;
        RECT 647.550 694.800 651.150 695.700 ;
        RECT 628.950 692.700 631.050 693.600 ;
        RECT 609.000 690.600 610.050 691.500 ;
        RECT 618.750 690.600 619.800 692.400 ;
        RECT 627.300 691.500 631.050 692.700 ;
        RECT 627.300 690.600 628.350 691.500 ;
        RECT 606.150 687.750 607.950 690.600 ;
        RECT 609.000 689.700 612.750 690.600 ;
        RECT 610.950 687.750 612.750 689.700 ;
        RECT 615.450 687.750 617.250 690.600 ;
        RECT 618.750 687.750 620.550 690.600 ;
        RECT 622.650 687.750 624.450 690.600 ;
        RECT 626.850 687.750 628.650 690.600 ;
        RECT 631.350 687.750 633.150 690.600 ;
        RECT 634.650 687.750 636.450 693.600 ;
        RECT 644.850 687.750 646.650 693.600 ;
        RECT 649.350 687.750 651.150 694.800 ;
        RECT 665.850 694.800 669.450 695.700 ;
        RECT 665.850 687.750 667.650 694.800 ;
        RECT 690.000 693.600 691.050 700.050 ;
        RECT 691.950 698.850 694.050 700.950 ;
        RECT 694.950 700.050 697.050 702.150 ;
        RECT 691.950 697.050 693.750 698.850 ;
        RECT 698.550 697.950 699.750 707.400 ;
        RECT 703.950 706.800 706.050 707.700 ;
        RECT 706.950 706.800 712.950 707.700 ;
        RECT 701.850 705.600 706.050 706.800 ;
        RECT 700.950 703.800 702.750 705.600 ;
        RECT 712.050 702.150 712.950 706.800 ;
        RECT 714.150 706.800 715.050 708.900 ;
        RECT 715.950 708.300 723.450 709.500 ;
        RECT 715.950 707.700 717.750 708.300 ;
        RECT 730.050 707.400 731.850 719.250 ;
        RECT 742.650 713.400 744.450 719.250 ;
        RECT 745.650 713.400 747.450 719.250 ;
        RECT 748.650 713.400 750.450 719.250 ;
        RECT 764.400 713.400 766.200 719.250 ;
        RECT 720.750 706.800 731.850 707.400 ;
        RECT 714.150 706.200 731.850 706.800 ;
        RECT 714.150 705.900 722.550 706.200 ;
        RECT 720.750 705.600 722.550 705.900 ;
        RECT 712.050 700.050 715.050 702.150 ;
        RECT 718.950 701.100 721.050 702.150 ;
        RECT 718.950 700.050 726.900 701.100 ;
        RECT 700.950 699.750 703.050 700.050 ;
        RECT 700.950 697.950 704.850 699.750 ;
        RECT 698.550 695.850 703.050 697.950 ;
        RECT 712.050 696.000 712.950 700.050 ;
        RECT 725.100 699.300 726.900 700.050 ;
        RECT 728.100 699.150 729.900 700.950 ;
        RECT 722.100 698.400 723.900 699.000 ;
        RECT 728.100 698.400 729.000 699.150 ;
        RECT 722.100 697.200 729.000 698.400 ;
        RECT 722.100 696.000 723.150 697.200 ;
        RECT 698.550 693.600 699.750 695.850 ;
        RECT 712.050 695.100 723.150 696.000 ;
        RECT 712.050 694.800 712.950 695.100 ;
        RECT 670.350 687.750 672.150 693.600 ;
        RECT 685.800 687.750 687.600 693.600 ;
        RECT 690.000 687.750 691.800 693.600 ;
        RECT 694.200 687.750 696.000 693.600 ;
        RECT 698.550 687.750 700.350 693.600 ;
        RECT 703.950 692.700 706.050 693.600 ;
        RECT 711.150 693.000 712.950 694.800 ;
        RECT 722.100 694.200 723.150 695.100 ;
        RECT 718.350 693.450 720.150 694.200 ;
        RECT 703.950 691.500 707.700 692.700 ;
        RECT 706.650 690.600 707.700 691.500 ;
        RECT 715.200 692.400 720.150 693.450 ;
        RECT 721.650 692.400 723.450 694.200 ;
        RECT 730.950 693.600 731.850 706.200 ;
        RECT 746.250 705.150 747.450 713.400 ;
        RECT 767.700 707.400 769.500 719.250 ;
        RECT 771.900 707.400 773.700 719.250 ;
        RECT 777.150 707.400 778.950 719.250 ;
        RECT 780.150 713.400 781.950 719.250 ;
        RECT 785.250 713.400 787.050 719.250 ;
        RECT 790.050 713.400 791.850 719.250 ;
        RECT 785.550 712.500 786.750 713.400 ;
        RECT 793.050 712.500 794.850 719.250 ;
        RECT 796.950 713.400 798.750 719.250 ;
        RECT 801.150 713.400 802.950 719.250 ;
        RECT 805.650 716.400 807.450 719.250 ;
        RECT 781.950 710.400 786.750 712.500 ;
        RECT 789.150 710.700 796.050 712.500 ;
        RECT 801.150 711.300 805.050 713.400 ;
        RECT 785.550 709.500 786.750 710.400 ;
        RECT 798.450 709.800 800.250 710.400 ;
        RECT 785.550 708.300 793.050 709.500 ;
        RECT 791.250 707.700 793.050 708.300 ;
        RECT 793.950 708.900 800.250 709.800 ;
        RECT 764.250 705.150 766.050 706.950 ;
        RECT 742.950 701.850 745.050 703.950 ;
        RECT 745.950 703.050 748.050 705.150 ;
        RECT 743.100 700.050 744.900 701.850 ;
        RECT 746.250 695.700 747.450 703.050 ;
        RECT 748.950 701.850 751.050 703.950 ;
        RECT 763.950 703.050 766.050 705.150 ;
        RECT 767.850 702.150 769.050 707.400 ;
        RECT 777.150 706.800 788.250 707.400 ;
        RECT 793.950 706.800 794.850 708.900 ;
        RECT 798.450 708.600 800.250 708.900 ;
        RECT 801.150 708.600 803.850 710.400 ;
        RECT 801.150 707.700 802.050 708.600 ;
        RECT 777.150 706.200 794.850 706.800 ;
        RECT 773.100 702.150 774.900 703.950 ;
        RECT 749.100 700.050 750.900 701.850 ;
        RECT 766.950 700.050 769.050 702.150 ;
        RECT 766.950 696.750 768.150 700.050 ;
        RECT 769.950 698.850 772.050 700.950 ;
        RECT 772.950 700.050 775.050 702.150 ;
        RECT 770.100 697.050 771.900 698.850 ;
        RECT 715.200 690.600 716.250 692.400 ;
        RECT 724.950 691.500 727.050 693.600 ;
        RECT 724.950 690.600 726.000 691.500 ;
        RECT 701.850 687.750 703.650 690.600 ;
        RECT 706.350 687.750 708.150 690.600 ;
        RECT 710.550 687.750 712.350 690.600 ;
        RECT 714.450 687.750 716.250 690.600 ;
        RECT 717.750 687.750 719.550 690.600 ;
        RECT 722.250 689.700 726.000 690.600 ;
        RECT 722.250 687.750 724.050 689.700 ;
        RECT 727.050 687.750 728.850 690.600 ;
        RECT 730.050 687.750 731.850 693.600 ;
        RECT 743.850 694.800 747.450 695.700 ;
        RECT 764.250 695.700 768.000 696.750 ;
        RECT 743.850 687.750 745.650 694.800 ;
        RECT 764.250 693.600 765.450 695.700 ;
        RECT 748.350 687.750 750.150 693.600 ;
        RECT 763.650 687.750 765.450 693.600 ;
        RECT 766.650 692.700 774.450 694.050 ;
        RECT 766.650 687.750 768.450 692.700 ;
        RECT 769.650 687.750 771.450 691.800 ;
        RECT 772.650 687.750 774.450 692.700 ;
        RECT 777.150 693.600 778.050 706.200 ;
        RECT 786.450 705.900 794.850 706.200 ;
        RECT 796.050 706.800 802.050 707.700 ;
        RECT 802.950 706.800 805.050 707.700 ;
        RECT 808.650 707.400 810.450 719.250 ;
        RECT 818.550 708.600 820.350 719.250 ;
        RECT 821.550 709.500 823.350 719.250 ;
        RECT 824.550 718.500 832.350 719.250 ;
        RECT 824.550 708.600 826.350 718.500 ;
        RECT 818.550 707.700 826.350 708.600 ;
        RECT 827.550 707.400 829.350 717.600 ;
        RECT 830.550 707.400 832.350 718.500 ;
        RECT 836.550 707.400 838.350 719.250 ;
        RECT 839.550 716.400 841.350 719.250 ;
        RECT 844.050 713.400 845.850 719.250 ;
        RECT 848.250 713.400 850.050 719.250 ;
        RECT 841.950 711.300 845.850 713.400 ;
        RECT 852.150 712.500 853.950 719.250 ;
        RECT 855.150 713.400 856.950 719.250 ;
        RECT 859.950 713.400 861.750 719.250 ;
        RECT 865.050 713.400 866.850 719.250 ;
        RECT 860.250 712.500 861.450 713.400 ;
        RECT 850.950 710.700 857.850 712.500 ;
        RECT 860.250 710.400 865.050 712.500 ;
        RECT 843.150 708.600 845.850 710.400 ;
        RECT 846.750 709.800 848.550 710.400 ;
        RECT 846.750 708.900 853.050 709.800 ;
        RECT 860.250 709.500 861.450 710.400 ;
        RECT 846.750 708.600 848.550 708.900 ;
        RECT 844.950 707.700 845.850 708.600 ;
        RECT 786.450 705.600 788.250 705.900 ;
        RECT 796.050 702.150 796.950 706.800 ;
        RECT 802.950 705.600 807.150 706.800 ;
        RECT 806.250 703.800 808.050 705.600 ;
        RECT 787.950 701.100 790.050 702.150 ;
        RECT 779.100 699.150 780.900 700.950 ;
        RECT 782.100 700.050 790.050 701.100 ;
        RECT 793.950 700.050 796.950 702.150 ;
        RECT 782.100 699.300 783.900 700.050 ;
        RECT 780.000 698.400 780.900 699.150 ;
        RECT 785.100 698.400 786.900 699.000 ;
        RECT 780.000 697.200 786.900 698.400 ;
        RECT 785.850 696.000 786.900 697.200 ;
        RECT 796.050 696.000 796.950 700.050 ;
        RECT 805.950 699.750 808.050 700.050 ;
        RECT 804.150 697.950 808.050 699.750 ;
        RECT 809.250 697.950 810.450 707.400 ;
        RECT 827.400 706.500 829.200 707.400 ;
        RECT 825.150 705.600 829.200 706.500 ;
        RECT 818.250 702.150 820.050 703.950 ;
        RECT 825.150 702.150 826.050 705.600 ;
        RECT 830.100 702.150 831.900 703.950 ;
        RECT 817.950 700.050 820.050 702.150 ;
        RECT 820.950 698.850 823.050 700.950 ;
        RECT 785.850 695.100 796.950 696.000 ;
        RECT 805.950 695.850 810.450 697.950 ;
        RECT 821.250 697.050 823.050 698.850 ;
        RECT 823.950 700.050 826.050 702.150 ;
        RECT 785.850 694.200 786.900 695.100 ;
        RECT 796.050 694.800 796.950 695.100 ;
        RECT 777.150 687.750 778.950 693.600 ;
        RECT 781.950 691.500 784.050 693.600 ;
        RECT 785.550 692.400 787.350 694.200 ;
        RECT 788.850 693.450 790.650 694.200 ;
        RECT 788.850 692.400 793.800 693.450 ;
        RECT 796.050 693.000 797.850 694.800 ;
        RECT 809.250 693.600 810.450 695.850 ;
        RECT 823.950 693.600 825.000 700.050 ;
        RECT 826.950 698.850 829.050 700.950 ;
        RECT 829.950 700.050 832.050 702.150 ;
        RECT 826.950 697.050 828.750 698.850 ;
        RECT 836.550 697.950 837.750 707.400 ;
        RECT 841.950 706.800 844.050 707.700 ;
        RECT 844.950 706.800 850.950 707.700 ;
        RECT 839.850 705.600 844.050 706.800 ;
        RECT 838.950 703.800 840.750 705.600 ;
        RECT 850.050 702.150 850.950 706.800 ;
        RECT 852.150 706.800 853.050 708.900 ;
        RECT 853.950 708.300 861.450 709.500 ;
        RECT 853.950 707.700 855.750 708.300 ;
        RECT 868.050 707.400 869.850 719.250 ;
        RECT 878.550 707.400 880.350 719.250 ;
        RECT 882.750 707.400 884.550 719.250 ;
        RECT 858.750 706.800 869.850 707.400 ;
        RECT 852.150 706.200 869.850 706.800 ;
        RECT 852.150 705.900 860.550 706.200 ;
        RECT 858.750 705.600 860.550 705.900 ;
        RECT 850.050 700.050 853.050 702.150 ;
        RECT 856.950 701.100 859.050 702.150 ;
        RECT 856.950 700.050 864.900 701.100 ;
        RECT 838.950 699.750 841.050 700.050 ;
        RECT 838.950 697.950 842.850 699.750 ;
        RECT 836.550 695.850 841.050 697.950 ;
        RECT 850.050 696.000 850.950 700.050 ;
        RECT 863.100 699.300 864.900 700.050 ;
        RECT 866.100 699.150 867.900 700.950 ;
        RECT 860.100 698.400 861.900 699.000 ;
        RECT 866.100 698.400 867.000 699.150 ;
        RECT 860.100 697.200 867.000 698.400 ;
        RECT 860.100 696.000 861.150 697.200 ;
        RECT 836.550 693.600 837.750 695.850 ;
        RECT 850.050 695.100 861.150 696.000 ;
        RECT 850.050 694.800 850.950 695.100 ;
        RECT 802.950 692.700 805.050 693.600 ;
        RECT 783.000 690.600 784.050 691.500 ;
        RECT 792.750 690.600 793.800 692.400 ;
        RECT 801.300 691.500 805.050 692.700 ;
        RECT 801.300 690.600 802.350 691.500 ;
        RECT 780.150 687.750 781.950 690.600 ;
        RECT 783.000 689.700 786.750 690.600 ;
        RECT 784.950 687.750 786.750 689.700 ;
        RECT 789.450 687.750 791.250 690.600 ;
        RECT 792.750 687.750 794.550 690.600 ;
        RECT 796.650 687.750 798.450 690.600 ;
        RECT 800.850 687.750 802.650 690.600 ;
        RECT 805.350 687.750 807.150 690.600 ;
        RECT 808.650 687.750 810.450 693.600 ;
        RECT 819.000 687.750 820.800 693.600 ;
        RECT 823.200 687.750 825.000 693.600 ;
        RECT 827.400 687.750 829.200 693.600 ;
        RECT 836.550 687.750 838.350 693.600 ;
        RECT 841.950 692.700 844.050 693.600 ;
        RECT 849.150 693.000 850.950 694.800 ;
        RECT 860.100 694.200 861.150 695.100 ;
        RECT 856.350 693.450 858.150 694.200 ;
        RECT 841.950 691.500 845.700 692.700 ;
        RECT 844.650 690.600 845.700 691.500 ;
        RECT 853.200 692.400 858.150 693.450 ;
        RECT 859.650 692.400 861.450 694.200 ;
        RECT 868.950 693.600 869.850 706.200 ;
        RECT 882.000 706.350 884.550 707.400 ;
        RECT 878.100 702.150 879.900 703.950 ;
        RECT 877.950 700.050 880.050 702.150 ;
        RECT 882.000 699.150 883.050 706.350 ;
        RECT 884.100 702.150 885.900 703.950 ;
        RECT 883.950 700.050 886.050 702.150 ;
        RECT 880.950 697.050 883.050 699.150 ;
        RECT 853.200 690.600 854.250 692.400 ;
        RECT 862.950 691.500 865.050 693.600 ;
        RECT 862.950 690.600 864.000 691.500 ;
        RECT 839.850 687.750 841.650 690.600 ;
        RECT 844.350 687.750 846.150 690.600 ;
        RECT 848.550 687.750 850.350 690.600 ;
        RECT 852.450 687.750 854.250 690.600 ;
        RECT 855.750 687.750 857.550 690.600 ;
        RECT 860.250 689.700 864.000 690.600 ;
        RECT 860.250 687.750 862.050 689.700 ;
        RECT 865.050 687.750 866.850 690.600 ;
        RECT 868.050 687.750 869.850 693.600 ;
        RECT 882.000 690.600 883.050 697.050 ;
        RECT 878.550 687.750 880.350 690.600 ;
        RECT 881.550 687.750 883.350 690.600 ;
        RECT 884.550 687.750 886.350 690.600 ;
        RECT 11.850 676.200 13.650 683.250 ;
        RECT 16.350 677.400 18.150 683.250 ;
        RECT 11.850 675.300 15.450 676.200 ;
        RECT 11.100 669.150 12.900 670.950 ;
        RECT 10.950 667.050 13.050 669.150 ;
        RECT 14.250 667.950 15.450 675.300 ;
        RECT 32.100 675.000 33.900 683.250 ;
        RECT 29.400 673.350 33.900 675.000 ;
        RECT 37.500 674.400 39.300 683.250 ;
        RECT 49.650 677.400 51.450 683.250 ;
        RECT 50.250 675.300 51.450 677.400 ;
        RECT 52.650 678.300 54.450 683.250 ;
        RECT 55.650 679.200 57.450 683.250 ;
        RECT 58.650 678.300 60.450 683.250 ;
        RECT 68.550 680.400 70.350 683.250 ;
        RECT 71.550 680.400 73.350 683.250 ;
        RECT 52.650 676.950 60.450 678.300 ;
        RECT 50.250 674.250 54.000 675.300 ;
        RECT 17.100 669.150 18.900 670.950 ;
        RECT 29.400 669.150 30.600 673.350 ;
        RECT 52.950 670.950 54.150 674.250 ;
        RECT 56.100 672.150 57.900 673.950 ;
        RECT 13.950 665.850 16.050 667.950 ;
        RECT 16.950 667.050 19.050 669.150 ;
        RECT 28.950 667.050 31.050 669.150 ;
        RECT 52.950 668.850 55.050 670.950 ;
        RECT 55.950 670.050 58.050 672.150 ;
        RECT 67.950 671.850 70.050 673.950 ;
        RECT 71.400 672.150 72.600 680.400 ;
        RECT 89.850 676.200 91.650 683.250 ;
        RECT 94.350 677.400 96.150 683.250 ;
        RECT 104.850 677.400 106.650 683.250 ;
        RECT 109.350 676.200 111.150 683.250 ;
        RECT 89.850 675.300 93.450 676.200 ;
        RECT 58.950 668.850 61.050 670.950 ;
        RECT 68.100 670.050 69.900 671.850 ;
        RECT 70.950 670.050 73.050 672.150 ;
        RECT 14.250 657.600 15.450 665.850 ;
        RECT 29.250 658.800 30.300 667.050 ;
        RECT 31.950 665.850 34.050 667.950 ;
        RECT 37.950 665.850 40.050 667.950 ;
        RECT 49.950 665.850 52.050 667.950 ;
        RECT 31.950 664.050 33.750 665.850 ;
        RECT 34.950 662.850 37.050 664.950 ;
        RECT 38.100 664.050 39.900 665.850 ;
        RECT 50.250 664.050 52.050 665.850 ;
        RECT 53.850 663.600 55.050 668.850 ;
        RECT 59.100 667.050 60.900 668.850 ;
        RECT 35.100 661.050 36.900 662.850 ;
        RECT 29.250 657.900 36.300 658.800 ;
        RECT 29.250 657.600 30.450 657.900 ;
        RECT 10.650 651.750 12.450 657.600 ;
        RECT 13.650 651.750 15.450 657.600 ;
        RECT 16.650 651.750 18.450 657.600 ;
        RECT 28.650 651.750 30.450 657.600 ;
        RECT 34.650 657.600 36.300 657.900 ;
        RECT 31.650 651.750 33.450 657.000 ;
        RECT 34.650 651.750 36.450 657.600 ;
        RECT 37.650 651.750 39.450 657.600 ;
        RECT 50.400 651.750 52.200 657.600 ;
        RECT 53.700 651.750 55.500 663.600 ;
        RECT 57.900 651.750 59.700 663.600 ;
        RECT 71.400 657.600 72.600 670.050 ;
        RECT 89.100 669.150 90.900 670.950 ;
        RECT 88.950 667.050 91.050 669.150 ;
        RECT 92.250 667.950 93.450 675.300 ;
        RECT 107.550 675.300 111.150 676.200 ;
        RECT 95.100 669.150 96.900 670.950 ;
        RECT 104.100 669.150 105.900 670.950 ;
        RECT 91.950 665.850 94.050 667.950 ;
        RECT 94.950 667.050 97.050 669.150 ;
        RECT 103.950 667.050 106.050 669.150 ;
        RECT 107.550 667.950 108.750 675.300 ;
        RECT 128.100 675.000 129.900 683.250 ;
        RECT 125.400 673.350 129.900 675.000 ;
        RECT 133.500 674.400 135.300 683.250 ;
        RECT 149.700 680.400 151.500 683.250 ;
        RECT 153.000 679.050 154.800 683.250 ;
        RECT 149.100 677.400 154.800 679.050 ;
        RECT 157.200 677.400 159.000 683.250 ;
        RECT 167.850 677.400 169.650 683.250 ;
        RECT 110.100 669.150 111.900 670.950 ;
        RECT 125.400 669.150 126.600 673.350 ;
        RECT 149.100 670.950 150.300 677.400 ;
        RECT 172.350 676.200 174.150 683.250 ;
        RECT 170.550 675.300 174.150 676.200 ;
        RECT 188.850 676.200 190.650 683.250 ;
        RECT 193.350 677.400 195.150 683.250 ;
        RECT 188.850 675.300 192.450 676.200 ;
        RECT 152.100 672.150 153.900 673.950 ;
        RECT 106.950 665.850 109.050 667.950 ;
        RECT 109.950 667.050 112.050 669.150 ;
        RECT 124.950 667.050 127.050 669.150 ;
        RECT 148.950 668.850 151.050 670.950 ;
        RECT 151.950 670.050 154.050 672.150 ;
        RECT 154.950 671.850 157.050 673.950 ;
        RECT 158.100 672.150 159.900 673.950 ;
        RECT 155.100 670.050 156.900 671.850 ;
        RECT 157.950 670.050 160.050 672.150 ;
        RECT 167.100 669.150 168.900 670.950 ;
        RECT 92.250 657.600 93.450 665.850 ;
        RECT 107.550 657.600 108.750 665.850 ;
        RECT 125.250 658.800 126.300 667.050 ;
        RECT 127.950 665.850 130.050 667.950 ;
        RECT 133.950 665.850 136.050 667.950 ;
        RECT 127.950 664.050 129.750 665.850 ;
        RECT 130.950 662.850 133.050 664.950 ;
        RECT 134.100 664.050 135.900 665.850 ;
        RECT 149.100 663.600 150.300 668.850 ;
        RECT 166.950 667.050 169.050 669.150 ;
        RECT 170.550 667.950 171.750 675.300 ;
        RECT 173.100 669.150 174.900 670.950 ;
        RECT 188.100 669.150 189.900 670.950 ;
        RECT 169.950 665.850 172.050 667.950 ;
        RECT 172.950 667.050 175.050 669.150 ;
        RECT 187.950 667.050 190.050 669.150 ;
        RECT 191.250 667.950 192.450 675.300 ;
        RECT 203.700 674.400 205.500 683.250 ;
        RECT 209.100 675.000 210.900 683.250 ;
        RECT 230.100 675.000 231.900 683.250 ;
        RECT 209.100 673.350 213.600 675.000 ;
        RECT 194.100 669.150 195.900 670.950 ;
        RECT 212.400 669.150 213.600 673.350 ;
        RECT 227.400 673.350 231.900 675.000 ;
        RECT 235.500 674.400 237.300 683.250 ;
        RECT 252.150 678.900 253.950 683.250 ;
        RECT 250.650 677.400 253.950 678.900 ;
        RECT 255.150 677.400 256.950 683.250 ;
        RECT 227.400 669.150 228.600 673.350 ;
        RECT 250.650 670.950 251.850 677.400 ;
        RECT 253.950 675.900 255.750 676.500 ;
        RECT 259.650 675.900 261.450 683.250 ;
        RECT 271.650 677.400 273.450 683.250 ;
        RECT 253.950 674.700 261.450 675.900 ;
        RECT 272.250 675.300 273.450 677.400 ;
        RECT 274.650 678.300 276.450 683.250 ;
        RECT 277.650 679.200 279.450 683.250 ;
        RECT 280.650 678.300 282.450 683.250 ;
        RECT 274.650 676.950 282.450 678.300 ;
        RECT 293.850 677.400 295.650 683.250 ;
        RECT 298.350 676.200 300.150 683.250 ;
        RECT 296.550 675.300 300.150 676.200 ;
        RECT 306.150 677.400 307.950 683.250 ;
        RECT 309.150 680.400 310.950 683.250 ;
        RECT 313.950 681.300 315.750 683.250 ;
        RECT 312.000 680.400 315.750 681.300 ;
        RECT 318.450 680.400 320.250 683.250 ;
        RECT 321.750 680.400 323.550 683.250 ;
        RECT 325.650 680.400 327.450 683.250 ;
        RECT 329.850 680.400 331.650 683.250 ;
        RECT 334.350 680.400 336.150 683.250 ;
        RECT 312.000 679.500 313.050 680.400 ;
        RECT 310.950 677.400 313.050 679.500 ;
        RECT 321.750 678.600 322.800 680.400 ;
        RECT 190.950 665.850 193.050 667.950 ;
        RECT 193.950 667.050 196.050 669.150 ;
        RECT 202.950 665.850 205.050 667.950 ;
        RECT 208.950 665.850 211.050 667.950 ;
        RECT 211.950 667.050 214.050 669.150 ;
        RECT 226.950 667.050 229.050 669.150 ;
        RECT 250.650 668.850 253.050 670.950 ;
        RECT 254.100 669.150 255.900 670.950 ;
        RECT 131.100 661.050 132.900 662.850 ;
        RECT 125.250 657.900 132.300 658.800 ;
        RECT 125.250 657.600 126.450 657.900 ;
        RECT 68.550 651.750 70.350 657.600 ;
        RECT 71.550 651.750 73.350 657.600 ;
        RECT 88.650 651.750 90.450 657.600 ;
        RECT 91.650 651.750 93.450 657.600 ;
        RECT 94.650 651.750 96.450 657.600 ;
        RECT 104.550 651.750 106.350 657.600 ;
        RECT 107.550 651.750 109.350 657.600 ;
        RECT 110.550 651.750 112.350 657.600 ;
        RECT 124.650 651.750 126.450 657.600 ;
        RECT 130.650 657.600 132.300 657.900 ;
        RECT 127.650 651.750 129.450 657.000 ;
        RECT 130.650 651.750 132.450 657.600 ;
        RECT 133.650 651.750 135.450 657.600 ;
        RECT 148.650 651.750 150.450 663.600 ;
        RECT 151.650 662.700 159.450 663.600 ;
        RECT 151.650 651.750 153.450 662.700 ;
        RECT 154.650 651.750 156.450 661.800 ;
        RECT 157.650 651.750 159.450 662.700 ;
        RECT 170.550 657.600 171.750 665.850 ;
        RECT 191.250 657.600 192.450 665.850 ;
        RECT 203.100 664.050 204.900 665.850 ;
        RECT 205.950 662.850 208.050 664.950 ;
        RECT 209.250 664.050 211.050 665.850 ;
        RECT 206.100 661.050 207.900 662.850 ;
        RECT 212.700 658.800 213.750 667.050 ;
        RECT 206.700 657.900 213.750 658.800 ;
        RECT 206.700 657.600 208.350 657.900 ;
        RECT 167.550 651.750 169.350 657.600 ;
        RECT 170.550 651.750 172.350 657.600 ;
        RECT 173.550 651.750 175.350 657.600 ;
        RECT 187.650 651.750 189.450 657.600 ;
        RECT 190.650 651.750 192.450 657.600 ;
        RECT 193.650 651.750 195.450 657.600 ;
        RECT 203.550 651.750 205.350 657.600 ;
        RECT 206.550 651.750 208.350 657.600 ;
        RECT 212.550 657.600 213.750 657.900 ;
        RECT 227.250 658.800 228.300 667.050 ;
        RECT 229.950 665.850 232.050 667.950 ;
        RECT 235.950 665.850 238.050 667.950 ;
        RECT 229.950 664.050 231.750 665.850 ;
        RECT 232.950 662.850 235.050 664.950 ;
        RECT 236.100 664.050 237.900 665.850 ;
        RECT 250.650 663.600 251.850 668.850 ;
        RECT 253.950 667.050 256.050 669.150 ;
        RECT 233.100 661.050 234.900 662.850 ;
        RECT 227.250 657.900 234.300 658.800 ;
        RECT 227.250 657.600 228.450 657.900 ;
        RECT 209.550 651.750 211.350 657.000 ;
        RECT 212.550 651.750 214.350 657.600 ;
        RECT 226.650 651.750 228.450 657.600 ;
        RECT 232.650 657.600 234.300 657.900 ;
        RECT 229.650 651.750 231.450 657.000 ;
        RECT 232.650 651.750 234.450 657.600 ;
        RECT 235.650 651.750 237.450 657.600 ;
        RECT 250.050 651.750 251.850 663.600 ;
        RECT 253.050 651.750 254.850 663.600 ;
        RECT 257.100 657.600 258.300 674.700 ;
        RECT 272.250 674.250 276.000 675.300 ;
        RECT 274.950 670.950 276.150 674.250 ;
        RECT 278.100 672.150 279.900 673.950 ;
        RECT 259.950 668.850 262.050 670.950 ;
        RECT 274.950 668.850 277.050 670.950 ;
        RECT 277.950 670.050 280.050 672.150 ;
        RECT 280.950 668.850 283.050 670.950 ;
        RECT 293.100 669.150 294.900 670.950 ;
        RECT 260.100 667.050 261.900 668.850 ;
        RECT 271.950 665.850 274.050 667.950 ;
        RECT 272.250 664.050 274.050 665.850 ;
        RECT 275.850 663.600 277.050 668.850 ;
        RECT 281.100 667.050 282.900 668.850 ;
        RECT 292.950 667.050 295.050 669.150 ;
        RECT 296.550 667.950 297.750 675.300 ;
        RECT 299.100 669.150 300.900 670.950 ;
        RECT 295.950 665.850 298.050 667.950 ;
        RECT 298.950 667.050 301.050 669.150 ;
        RECT 256.650 651.750 258.450 657.600 ;
        RECT 259.650 651.750 261.450 657.600 ;
        RECT 272.400 651.750 274.200 657.600 ;
        RECT 275.700 651.750 277.500 663.600 ;
        RECT 279.900 651.750 281.700 663.600 ;
        RECT 296.550 657.600 297.750 665.850 ;
        RECT 306.150 664.800 307.050 677.400 ;
        RECT 314.550 676.800 316.350 678.600 ;
        RECT 317.850 677.550 322.800 678.600 ;
        RECT 330.300 679.500 331.350 680.400 ;
        RECT 330.300 678.300 334.050 679.500 ;
        RECT 317.850 676.800 319.650 677.550 ;
        RECT 314.850 675.900 315.900 676.800 ;
        RECT 325.050 676.200 326.850 678.000 ;
        RECT 331.950 677.400 334.050 678.300 ;
        RECT 337.650 677.400 339.450 683.250 ;
        RECT 349.650 680.400 351.450 683.250 ;
        RECT 352.650 680.400 354.450 683.250 ;
        RECT 355.650 680.400 357.450 683.250 ;
        RECT 325.050 675.900 325.950 676.200 ;
        RECT 314.850 675.000 325.950 675.900 ;
        RECT 338.250 675.150 339.450 677.400 ;
        RECT 314.850 673.800 315.900 675.000 ;
        RECT 309.000 672.600 315.900 673.800 ;
        RECT 309.000 671.850 309.900 672.600 ;
        RECT 314.100 672.000 315.900 672.600 ;
        RECT 308.100 670.050 309.900 671.850 ;
        RECT 311.100 670.950 312.900 671.700 ;
        RECT 325.050 670.950 325.950 675.000 ;
        RECT 334.950 673.050 339.450 675.150 ;
        RECT 333.150 671.250 337.050 673.050 ;
        RECT 334.950 670.950 337.050 671.250 ;
        RECT 311.100 669.900 319.050 670.950 ;
        RECT 316.950 668.850 319.050 669.900 ;
        RECT 322.950 668.850 325.950 670.950 ;
        RECT 315.450 665.100 317.250 665.400 ;
        RECT 315.450 664.800 323.850 665.100 ;
        RECT 306.150 664.200 323.850 664.800 ;
        RECT 306.150 663.600 317.250 664.200 ;
        RECT 293.550 651.750 295.350 657.600 ;
        RECT 296.550 651.750 298.350 657.600 ;
        RECT 299.550 651.750 301.350 657.600 ;
        RECT 306.150 651.750 307.950 663.600 ;
        RECT 320.250 662.700 322.050 663.300 ;
        RECT 314.550 661.500 322.050 662.700 ;
        RECT 322.950 662.100 323.850 664.200 ;
        RECT 325.050 664.200 325.950 668.850 ;
        RECT 335.250 665.400 337.050 667.200 ;
        RECT 331.950 664.200 336.150 665.400 ;
        RECT 325.050 663.300 331.050 664.200 ;
        RECT 331.950 663.300 334.050 664.200 ;
        RECT 338.250 663.600 339.450 673.050 ;
        RECT 352.950 673.950 354.000 680.400 ;
        RECT 367.650 677.400 369.450 683.250 ;
        RECT 368.250 675.300 369.450 677.400 ;
        RECT 370.650 678.300 372.450 683.250 ;
        RECT 373.650 679.200 375.450 683.250 ;
        RECT 376.650 678.300 378.450 683.250 ;
        RECT 386.550 680.400 388.350 683.250 ;
        RECT 389.550 680.400 391.350 683.250 ;
        RECT 370.650 676.950 378.450 678.300 ;
        RECT 368.250 674.250 372.000 675.300 ;
        RECT 352.950 671.850 355.050 673.950 ;
        RECT 349.950 668.850 352.050 670.950 ;
        RECT 350.100 667.050 351.900 668.850 ;
        RECT 352.950 664.650 354.000 671.850 ;
        RECT 370.950 670.950 372.150 674.250 ;
        RECT 374.100 672.150 375.900 673.950 ;
        RECT 355.950 668.850 358.050 670.950 ;
        RECT 370.950 668.850 373.050 670.950 ;
        RECT 373.950 670.050 376.050 672.150 ;
        RECT 385.950 671.850 388.050 673.950 ;
        RECT 389.400 672.150 390.600 680.400 ;
        RECT 401.850 677.400 403.650 683.250 ;
        RECT 406.350 676.200 408.150 683.250 ;
        RECT 404.550 675.300 408.150 676.200 ;
        RECT 422.850 676.200 424.650 683.250 ;
        RECT 427.350 677.400 429.150 683.250 ;
        RECT 442.650 677.400 444.450 683.250 ;
        RECT 422.850 675.300 426.450 676.200 ;
        RECT 376.950 668.850 379.050 670.950 ;
        RECT 386.100 670.050 387.900 671.850 ;
        RECT 388.950 670.050 391.050 672.150 ;
        RECT 356.100 667.050 357.900 668.850 ;
        RECT 367.950 665.850 370.050 667.950 ;
        RECT 330.150 662.400 331.050 663.300 ;
        RECT 327.450 662.100 329.250 662.400 ;
        RECT 314.550 660.600 315.750 661.500 ;
        RECT 322.950 661.200 329.250 662.100 ;
        RECT 327.450 660.600 329.250 661.200 ;
        RECT 330.150 660.600 332.850 662.400 ;
        RECT 310.950 658.500 315.750 660.600 ;
        RECT 318.150 658.500 325.050 660.300 ;
        RECT 314.550 657.600 315.750 658.500 ;
        RECT 309.150 651.750 310.950 657.600 ;
        RECT 314.250 651.750 316.050 657.600 ;
        RECT 319.050 651.750 320.850 657.600 ;
        RECT 322.050 651.750 323.850 658.500 ;
        RECT 330.150 657.600 334.050 659.700 ;
        RECT 325.950 651.750 327.750 657.600 ;
        RECT 330.150 651.750 331.950 657.600 ;
        RECT 334.650 651.750 336.450 654.600 ;
        RECT 337.650 651.750 339.450 663.600 ;
        RECT 351.450 663.600 354.000 664.650 ;
        RECT 368.250 664.050 370.050 665.850 ;
        RECT 371.850 663.600 373.050 668.850 ;
        RECT 377.100 667.050 378.900 668.850 ;
        RECT 351.450 651.750 353.250 663.600 ;
        RECT 355.650 651.750 357.450 663.600 ;
        RECT 368.400 651.750 370.200 657.600 ;
        RECT 371.700 651.750 373.500 663.600 ;
        RECT 375.900 651.750 377.700 663.600 ;
        RECT 389.400 657.600 390.600 670.050 ;
        RECT 401.100 669.150 402.900 670.950 ;
        RECT 400.950 667.050 403.050 669.150 ;
        RECT 404.550 667.950 405.750 675.300 ;
        RECT 407.100 669.150 408.900 670.950 ;
        RECT 422.100 669.150 423.900 670.950 ;
        RECT 403.950 665.850 406.050 667.950 ;
        RECT 406.950 667.050 409.050 669.150 ;
        RECT 421.950 667.050 424.050 669.150 ;
        RECT 425.250 667.950 426.450 675.300 ;
        RECT 443.250 675.300 444.450 677.400 ;
        RECT 445.650 678.300 447.450 683.250 ;
        RECT 448.650 679.200 450.450 683.250 ;
        RECT 451.650 678.300 453.450 683.250 ;
        RECT 464.550 680.400 466.350 683.250 ;
        RECT 467.550 680.400 469.350 683.250 ;
        RECT 470.550 680.400 472.350 683.250 ;
        RECT 445.650 676.950 453.450 678.300 ;
        RECT 443.250 674.250 447.000 675.300 ;
        RECT 445.950 670.950 447.150 674.250 ;
        RECT 468.000 673.950 469.050 680.400 ;
        RECT 485.850 676.200 487.650 683.250 ;
        RECT 490.350 677.400 492.150 683.250 ;
        RECT 500.850 677.400 502.650 683.250 ;
        RECT 505.350 676.200 507.150 683.250 ;
        RECT 521.550 680.400 523.350 683.250 ;
        RECT 524.550 680.400 526.350 683.250 ;
        RECT 527.550 680.400 529.350 683.250 ;
        RECT 485.850 675.300 489.450 676.200 ;
        RECT 449.100 672.150 450.900 673.950 ;
        RECT 428.100 669.150 429.900 670.950 ;
        RECT 424.950 665.850 427.050 667.950 ;
        RECT 427.950 667.050 430.050 669.150 ;
        RECT 445.950 668.850 448.050 670.950 ;
        RECT 448.950 670.050 451.050 672.150 ;
        RECT 466.950 671.850 469.050 673.950 ;
        RECT 451.950 668.850 454.050 670.950 ;
        RECT 463.950 668.850 466.050 670.950 ;
        RECT 442.950 665.850 445.050 667.950 ;
        RECT 404.550 657.600 405.750 665.850 ;
        RECT 425.250 657.600 426.450 665.850 ;
        RECT 443.250 664.050 445.050 665.850 ;
        RECT 446.850 663.600 448.050 668.850 ;
        RECT 452.100 667.050 453.900 668.850 ;
        RECT 464.100 667.050 465.900 668.850 ;
        RECT 468.000 664.650 469.050 671.850 ;
        RECT 469.950 668.850 472.050 670.950 ;
        RECT 485.100 669.150 486.900 670.950 ;
        RECT 470.100 667.050 471.900 668.850 ;
        RECT 484.950 667.050 487.050 669.150 ;
        RECT 488.250 667.950 489.450 675.300 ;
        RECT 503.550 675.300 507.150 676.200 ;
        RECT 525.450 676.200 526.350 680.400 ;
        RECT 530.550 677.400 532.350 683.250 ;
        RECT 543.000 677.400 544.800 683.250 ;
        RECT 547.200 679.050 549.000 683.250 ;
        RECT 550.500 680.400 552.300 683.250 ;
        RECT 565.650 680.400 567.450 683.250 ;
        RECT 568.650 680.400 570.450 683.250 ;
        RECT 571.650 680.400 573.450 683.250 ;
        RECT 547.200 677.400 552.900 679.050 ;
        RECT 525.450 675.300 528.750 676.200 ;
        RECT 491.100 669.150 492.900 670.950 ;
        RECT 500.100 669.150 501.900 670.950 ;
        RECT 487.950 665.850 490.050 667.950 ;
        RECT 490.950 667.050 493.050 669.150 ;
        RECT 499.950 667.050 502.050 669.150 ;
        RECT 503.550 667.950 504.750 675.300 ;
        RECT 526.950 674.400 528.750 675.300 ;
        RECT 520.950 671.850 523.050 673.950 ;
        RECT 506.100 669.150 507.900 670.950 ;
        RECT 521.100 670.050 522.900 671.850 ;
        RECT 502.950 665.850 505.050 667.950 ;
        RECT 505.950 667.050 508.050 669.150 ;
        RECT 523.950 668.850 526.050 670.950 ;
        RECT 524.100 667.050 525.900 668.850 ;
        RECT 527.700 666.150 528.600 674.400 ;
        RECT 531.000 672.150 532.050 677.400 ;
        RECT 542.100 672.150 543.900 673.950 ;
        RECT 529.950 670.050 532.050 672.150 ;
        RECT 541.950 670.050 544.050 672.150 ;
        RECT 544.950 671.850 547.050 673.950 ;
        RECT 548.100 672.150 549.900 673.950 ;
        RECT 545.100 670.050 546.900 671.850 ;
        RECT 547.950 670.050 550.050 672.150 ;
        RECT 551.700 670.950 552.900 677.400 ;
        RECT 568.950 673.950 570.000 680.400 ;
        RECT 581.850 677.400 583.650 683.250 ;
        RECT 586.350 676.200 588.150 683.250 ;
        RECT 599.550 680.400 601.350 683.250 ;
        RECT 602.550 680.400 604.350 683.250 ;
        RECT 584.550 675.300 588.150 676.200 ;
        RECT 568.950 671.850 571.050 673.950 ;
        RECT 526.950 666.000 528.750 666.150 ;
        RECT 468.000 663.600 470.550 664.650 ;
        RECT 386.550 651.750 388.350 657.600 ;
        RECT 389.550 651.750 391.350 657.600 ;
        RECT 401.550 651.750 403.350 657.600 ;
        RECT 404.550 651.750 406.350 657.600 ;
        RECT 407.550 651.750 409.350 657.600 ;
        RECT 421.650 651.750 423.450 657.600 ;
        RECT 424.650 651.750 426.450 657.600 ;
        RECT 427.650 651.750 429.450 657.600 ;
        RECT 443.400 651.750 445.200 657.600 ;
        RECT 446.700 651.750 448.500 663.600 ;
        RECT 450.900 651.750 452.700 663.600 ;
        RECT 464.550 651.750 466.350 663.600 ;
        RECT 468.750 651.750 470.550 663.600 ;
        RECT 488.250 657.600 489.450 665.850 ;
        RECT 503.550 657.600 504.750 665.850 ;
        RECT 521.550 664.800 528.750 666.000 ;
        RECT 521.550 663.600 522.750 664.800 ;
        RECT 526.950 664.350 528.750 664.800 ;
        RECT 484.650 651.750 486.450 657.600 ;
        RECT 487.650 651.750 489.450 657.600 ;
        RECT 490.650 651.750 492.450 657.600 ;
        RECT 500.550 651.750 502.350 657.600 ;
        RECT 503.550 651.750 505.350 657.600 ;
        RECT 506.550 651.750 508.350 657.600 ;
        RECT 521.550 651.750 523.350 663.600 ;
        RECT 530.100 663.450 531.450 670.050 ;
        RECT 550.950 668.850 553.050 670.950 ;
        RECT 565.950 668.850 568.050 670.950 ;
        RECT 551.700 663.600 552.900 668.850 ;
        RECT 566.100 667.050 567.900 668.850 ;
        RECT 568.950 664.650 570.000 671.850 ;
        RECT 571.950 668.850 574.050 670.950 ;
        RECT 581.100 669.150 582.900 670.950 ;
        RECT 572.100 667.050 573.900 668.850 ;
        RECT 580.950 667.050 583.050 669.150 ;
        RECT 584.550 667.950 585.750 675.300 ;
        RECT 598.950 671.850 601.050 673.950 ;
        RECT 602.400 672.150 603.600 680.400 ;
        RECT 614.550 678.300 616.350 683.250 ;
        RECT 617.550 679.200 619.350 683.250 ;
        RECT 620.550 678.300 622.350 683.250 ;
        RECT 614.550 676.950 622.350 678.300 ;
        RECT 623.550 677.400 625.350 683.250 ;
        RECT 638.550 680.400 640.350 683.250 ;
        RECT 641.550 680.400 643.350 683.250 ;
        RECT 623.550 675.300 624.750 677.400 ;
        RECT 621.000 674.250 624.750 675.300 ;
        RECT 617.100 672.150 618.900 673.950 ;
        RECT 587.100 669.150 588.900 670.950 ;
        RECT 599.100 670.050 600.900 671.850 ;
        RECT 601.950 670.050 604.050 672.150 ;
        RECT 583.950 665.850 586.050 667.950 ;
        RECT 586.950 667.050 589.050 669.150 ;
        RECT 567.450 663.600 570.000 664.650 ;
        RECT 526.050 651.750 527.850 663.450 ;
        RECT 529.050 662.100 531.450 663.450 ;
        RECT 542.550 662.700 550.350 663.600 ;
        RECT 529.050 651.750 530.850 662.100 ;
        RECT 542.550 651.750 544.350 662.700 ;
        RECT 545.550 651.750 547.350 661.800 ;
        RECT 548.550 651.750 550.350 662.700 ;
        RECT 551.550 651.750 553.350 663.600 ;
        RECT 567.450 651.750 569.250 663.600 ;
        RECT 571.650 651.750 573.450 663.600 ;
        RECT 584.550 657.600 585.750 665.850 ;
        RECT 602.400 657.600 603.600 670.050 ;
        RECT 613.950 668.850 616.050 670.950 ;
        RECT 616.950 670.050 619.050 672.150 ;
        RECT 620.850 670.950 622.050 674.250 ;
        RECT 637.950 671.850 640.050 673.950 ;
        RECT 641.400 672.150 642.600 680.400 ;
        RECT 658.800 677.400 660.600 683.250 ;
        RECT 663.000 677.400 664.800 683.250 ;
        RECT 667.200 677.400 669.000 683.250 ;
        RECT 682.650 677.400 684.450 683.250 ;
        RECT 659.250 672.150 661.050 673.950 ;
        RECT 619.950 668.850 622.050 670.950 ;
        RECT 638.100 670.050 639.900 671.850 ;
        RECT 640.950 670.050 643.050 672.150 ;
        RECT 614.100 667.050 615.900 668.850 ;
        RECT 619.950 663.600 621.150 668.850 ;
        RECT 622.950 665.850 625.050 667.950 ;
        RECT 622.950 664.050 624.750 665.850 ;
        RECT 581.550 651.750 583.350 657.600 ;
        RECT 584.550 651.750 586.350 657.600 ;
        RECT 587.550 651.750 589.350 657.600 ;
        RECT 599.550 651.750 601.350 657.600 ;
        RECT 602.550 651.750 604.350 657.600 ;
        RECT 615.300 651.750 617.100 663.600 ;
        RECT 619.500 651.750 621.300 663.600 ;
        RECT 641.400 657.600 642.600 670.050 ;
        RECT 655.950 668.850 658.050 670.950 ;
        RECT 658.950 670.050 661.050 672.150 ;
        RECT 663.000 670.950 664.050 677.400 ;
        RECT 683.250 675.300 684.450 677.400 ;
        RECT 685.650 678.300 687.450 683.250 ;
        RECT 688.650 679.200 690.450 683.250 ;
        RECT 691.650 678.300 693.450 683.250 ;
        RECT 685.650 676.950 693.450 678.300 ;
        RECT 695.550 677.400 697.350 683.250 ;
        RECT 698.850 680.400 700.650 683.250 ;
        RECT 703.350 680.400 705.150 683.250 ;
        RECT 707.550 680.400 709.350 683.250 ;
        RECT 711.450 680.400 713.250 683.250 ;
        RECT 714.750 680.400 716.550 683.250 ;
        RECT 719.250 681.300 721.050 683.250 ;
        RECT 719.250 680.400 723.000 681.300 ;
        RECT 724.050 680.400 725.850 683.250 ;
        RECT 703.650 679.500 704.700 680.400 ;
        RECT 700.950 678.300 704.700 679.500 ;
        RECT 712.200 678.600 713.250 680.400 ;
        RECT 721.950 679.500 723.000 680.400 ;
        RECT 700.950 677.400 703.050 678.300 ;
        RECT 683.250 674.250 687.000 675.300 ;
        RECT 695.550 675.150 696.750 677.400 ;
        RECT 708.150 676.200 709.950 678.000 ;
        RECT 712.200 677.550 717.150 678.600 ;
        RECT 715.350 676.800 717.150 677.550 ;
        RECT 718.650 676.800 720.450 678.600 ;
        RECT 721.950 677.400 724.050 679.500 ;
        RECT 727.050 677.400 728.850 683.250 ;
        RECT 709.050 675.900 709.950 676.200 ;
        RECT 719.100 675.900 720.150 676.800 ;
        RECT 661.950 668.850 664.050 670.950 ;
        RECT 664.950 672.150 666.750 673.950 ;
        RECT 664.950 670.050 667.050 672.150 ;
        RECT 685.950 670.950 687.150 674.250 ;
        RECT 689.100 672.150 690.900 673.950 ;
        RECT 695.550 673.050 700.050 675.150 ;
        RECT 709.050 675.000 720.150 675.900 ;
        RECT 667.950 668.850 670.050 670.950 ;
        RECT 685.950 668.850 688.050 670.950 ;
        RECT 688.950 670.050 691.050 672.150 ;
        RECT 691.950 668.850 694.050 670.950 ;
        RECT 656.100 667.050 657.900 668.850 ;
        RECT 661.950 665.400 662.850 668.850 ;
        RECT 667.950 667.050 669.750 668.850 ;
        RECT 682.950 665.850 685.050 667.950 ;
        RECT 658.800 664.500 662.850 665.400 ;
        RECT 658.800 663.600 660.600 664.500 ;
        RECT 683.250 664.050 685.050 665.850 ;
        RECT 686.850 663.600 688.050 668.850 ;
        RECT 692.100 667.050 693.900 668.850 ;
        RECT 695.550 663.600 696.750 673.050 ;
        RECT 697.950 671.250 701.850 673.050 ;
        RECT 697.950 670.950 700.050 671.250 ;
        RECT 709.050 670.950 709.950 675.000 ;
        RECT 719.100 673.800 720.150 675.000 ;
        RECT 719.100 672.600 726.000 673.800 ;
        RECT 719.100 672.000 720.900 672.600 ;
        RECT 725.100 671.850 726.000 672.600 ;
        RECT 722.100 670.950 723.900 671.700 ;
        RECT 709.050 668.850 712.050 670.950 ;
        RECT 715.950 669.900 723.900 670.950 ;
        RECT 725.100 670.050 726.900 671.850 ;
        RECT 715.950 668.850 718.050 669.900 ;
        RECT 697.950 665.400 699.750 667.200 ;
        RECT 698.850 664.200 703.050 665.400 ;
        RECT 709.050 664.200 709.950 668.850 ;
        RECT 717.750 665.100 719.550 665.400 ;
        RECT 622.800 651.750 624.600 657.600 ;
        RECT 638.550 651.750 640.350 657.600 ;
        RECT 641.550 651.750 643.350 657.600 ;
        RECT 655.650 652.500 657.450 663.600 ;
        RECT 658.650 653.400 660.450 663.600 ;
        RECT 661.650 662.400 669.450 663.300 ;
        RECT 661.650 652.500 663.450 662.400 ;
        RECT 655.650 651.750 663.450 652.500 ;
        RECT 664.650 651.750 666.450 661.500 ;
        RECT 667.650 651.750 669.450 662.400 ;
        RECT 683.400 651.750 685.200 657.600 ;
        RECT 686.700 651.750 688.500 663.600 ;
        RECT 690.900 651.750 692.700 663.600 ;
        RECT 695.550 651.750 697.350 663.600 ;
        RECT 700.950 663.300 703.050 664.200 ;
        RECT 703.950 663.300 709.950 664.200 ;
        RECT 711.150 664.800 719.550 665.100 ;
        RECT 727.950 664.800 728.850 677.400 ;
        RECT 737.550 678.300 739.350 683.250 ;
        RECT 740.550 679.200 742.350 683.250 ;
        RECT 743.550 678.300 745.350 683.250 ;
        RECT 737.550 676.950 745.350 678.300 ;
        RECT 746.550 677.400 748.350 683.250 ;
        RECT 758.850 677.400 760.650 683.250 ;
        RECT 746.550 675.300 747.750 677.400 ;
        RECT 763.350 676.200 765.150 683.250 ;
        RECT 776.550 678.300 778.350 683.250 ;
        RECT 779.550 679.200 781.350 683.250 ;
        RECT 782.550 678.300 784.350 683.250 ;
        RECT 776.550 676.950 784.350 678.300 ;
        RECT 785.550 677.400 787.350 683.250 ;
        RECT 797.850 677.400 799.650 683.250 ;
        RECT 744.000 674.250 747.750 675.300 ;
        RECT 761.550 675.300 765.150 676.200 ;
        RECT 775.950 675.450 778.050 676.050 ;
        RECT 740.100 672.150 741.900 673.950 ;
        RECT 736.950 668.850 739.050 670.950 ;
        RECT 739.950 670.050 742.050 672.150 ;
        RECT 743.850 670.950 745.050 674.250 ;
        RECT 742.950 668.850 745.050 670.950 ;
        RECT 758.100 669.150 759.900 670.950 ;
        RECT 737.100 667.050 738.900 668.850 ;
        RECT 711.150 664.200 728.850 664.800 ;
        RECT 703.950 662.400 704.850 663.300 ;
        RECT 702.150 660.600 704.850 662.400 ;
        RECT 705.750 662.100 707.550 662.400 ;
        RECT 711.150 662.100 712.050 664.200 ;
        RECT 717.750 663.600 728.850 664.200 ;
        RECT 742.950 663.600 744.150 668.850 ;
        RECT 745.950 665.850 748.050 667.950 ;
        RECT 757.950 667.050 760.050 669.150 ;
        RECT 761.550 667.950 762.750 675.300 ;
        RECT 773.550 674.550 778.050 675.450 ;
        RECT 785.550 675.300 786.750 677.400 ;
        RECT 802.350 676.200 804.150 683.250 ;
        RECT 818.550 680.400 820.350 683.250 ;
        RECT 764.100 669.150 765.900 670.950 ;
        RECT 760.950 665.850 763.050 667.950 ;
        RECT 763.950 667.050 766.050 669.150 ;
        RECT 745.950 664.050 747.750 665.850 ;
        RECT 705.750 661.200 712.050 662.100 ;
        RECT 712.950 662.700 714.750 663.300 ;
        RECT 712.950 661.500 720.450 662.700 ;
        RECT 705.750 660.600 707.550 661.200 ;
        RECT 719.250 660.600 720.450 661.500 ;
        RECT 700.950 657.600 704.850 659.700 ;
        RECT 709.950 658.500 716.850 660.300 ;
        RECT 719.250 658.500 724.050 660.600 ;
        RECT 698.550 651.750 700.350 654.600 ;
        RECT 703.050 651.750 704.850 657.600 ;
        RECT 707.250 651.750 709.050 657.600 ;
        RECT 711.150 651.750 712.950 658.500 ;
        RECT 719.250 657.600 720.450 658.500 ;
        RECT 714.150 651.750 715.950 657.600 ;
        RECT 718.950 651.750 720.750 657.600 ;
        RECT 724.050 651.750 725.850 657.600 ;
        RECT 727.050 651.750 728.850 663.600 ;
        RECT 738.300 651.750 740.100 663.600 ;
        RECT 742.500 651.750 744.300 663.600 ;
        RECT 761.550 657.600 762.750 665.850 ;
        RECT 773.550 664.050 774.450 674.550 ;
        RECT 775.950 673.950 778.050 674.550 ;
        RECT 783.000 674.250 786.750 675.300 ;
        RECT 800.550 675.300 804.150 676.200 ;
        RECT 819.150 676.500 820.350 680.400 ;
        RECT 821.850 677.400 823.650 683.250 ;
        RECT 824.850 677.400 826.650 683.250 ;
        RECT 839.850 677.400 841.650 683.250 ;
        RECT 819.150 675.600 824.250 676.500 ;
        RECT 779.100 672.150 780.900 673.950 ;
        RECT 775.950 668.850 778.050 670.950 ;
        RECT 778.950 670.050 781.050 672.150 ;
        RECT 782.850 670.950 784.050 674.250 ;
        RECT 781.950 668.850 784.050 670.950 ;
        RECT 797.100 669.150 798.900 670.950 ;
        RECT 776.100 667.050 777.900 668.850 ;
        RECT 772.950 661.950 775.050 664.050 ;
        RECT 781.950 663.600 783.150 668.850 ;
        RECT 784.950 665.850 787.050 667.950 ;
        RECT 796.950 667.050 799.050 669.150 ;
        RECT 800.550 667.950 801.750 675.300 ;
        RECT 822.000 674.700 824.250 675.600 ;
        RECT 803.100 669.150 804.900 670.950 ;
        RECT 799.950 665.850 802.050 667.950 ;
        RECT 802.950 667.050 805.050 669.150 ;
        RECT 817.950 668.850 820.050 670.950 ;
        RECT 818.100 667.050 819.900 668.850 ;
        RECT 822.000 666.300 823.050 674.700 ;
        RECT 825.150 670.950 826.350 677.400 ;
        RECT 844.350 676.200 846.150 683.250 ;
        RECT 859.650 677.400 861.450 683.250 ;
        RECT 842.550 675.300 846.150 676.200 ;
        RECT 860.250 675.300 861.450 677.400 ;
        RECT 862.650 678.300 864.450 683.250 ;
        RECT 865.650 679.200 867.450 683.250 ;
        RECT 868.650 678.300 870.450 683.250 ;
        RECT 862.650 676.950 870.450 678.300 ;
        RECT 823.950 668.850 826.350 670.950 ;
        RECT 839.100 669.150 840.900 670.950 ;
        RECT 784.950 664.050 786.750 665.850 ;
        RECT 745.800 651.750 747.600 657.600 ;
        RECT 758.550 651.750 760.350 657.600 ;
        RECT 761.550 651.750 763.350 657.600 ;
        RECT 764.550 651.750 766.350 657.600 ;
        RECT 777.300 651.750 779.100 663.600 ;
        RECT 781.500 651.750 783.300 663.600 ;
        RECT 800.550 657.600 801.750 665.850 ;
        RECT 822.000 665.400 824.250 666.300 ;
        RECT 818.550 664.500 824.250 665.400 ;
        RECT 818.550 657.600 819.750 664.500 ;
        RECT 825.150 663.600 826.350 668.850 ;
        RECT 838.950 667.050 841.050 669.150 ;
        RECT 842.550 667.950 843.750 675.300 ;
        RECT 860.250 674.250 864.000 675.300 ;
        RECT 862.950 670.950 864.150 674.250 ;
        RECT 866.100 672.150 867.900 673.950 ;
        RECT 845.100 669.150 846.900 670.950 ;
        RECT 841.950 665.850 844.050 667.950 ;
        RECT 844.950 667.050 847.050 669.150 ;
        RECT 862.950 668.850 865.050 670.950 ;
        RECT 865.950 670.050 868.050 672.150 ;
        RECT 868.950 668.850 871.050 670.950 ;
        RECT 859.950 665.850 862.050 667.950 ;
        RECT 784.800 651.750 786.600 657.600 ;
        RECT 797.550 651.750 799.350 657.600 ;
        RECT 800.550 651.750 802.350 657.600 ;
        RECT 803.550 651.750 805.350 657.600 ;
        RECT 818.550 651.750 820.350 657.600 ;
        RECT 821.850 651.750 823.650 663.600 ;
        RECT 824.850 651.750 826.650 663.600 ;
        RECT 842.550 657.600 843.750 665.850 ;
        RECT 860.250 664.050 862.050 665.850 ;
        RECT 863.850 663.600 865.050 668.850 ;
        RECT 869.100 667.050 870.900 668.850 ;
        RECT 839.550 651.750 841.350 657.600 ;
        RECT 842.550 651.750 844.350 657.600 ;
        RECT 845.550 651.750 847.350 657.600 ;
        RECT 860.400 651.750 862.200 657.600 ;
        RECT 863.700 651.750 865.500 663.600 ;
        RECT 867.900 651.750 869.700 663.600 ;
        RECT 13.650 641.400 15.450 647.250 ;
        RECT 16.650 641.400 18.450 647.250 ;
        RECT 31.650 641.400 33.450 647.250 ;
        RECT 34.650 642.000 36.450 647.250 ;
        RECT 14.400 628.950 15.600 641.400 ;
        RECT 32.250 641.100 33.450 641.400 ;
        RECT 37.650 641.400 39.450 647.250 ;
        RECT 40.650 641.400 42.450 647.250 ;
        RECT 52.650 641.400 54.450 647.250 ;
        RECT 55.650 642.000 57.450 647.250 ;
        RECT 37.650 641.100 39.300 641.400 ;
        RECT 32.250 640.200 39.300 641.100 ;
        RECT 53.250 641.100 54.450 641.400 ;
        RECT 58.650 641.400 60.450 647.250 ;
        RECT 61.650 641.400 63.450 647.250 ;
        RECT 58.650 641.100 60.300 641.400 ;
        RECT 53.250 640.200 60.300 641.100 ;
        RECT 32.250 631.950 33.300 640.200 ;
        RECT 38.100 636.150 39.900 637.950 ;
        RECT 34.950 633.150 36.750 634.950 ;
        RECT 37.950 634.050 40.050 636.150 ;
        RECT 41.100 633.150 42.900 634.950 ;
        RECT 31.950 629.850 34.050 631.950 ;
        RECT 34.950 631.050 37.050 633.150 ;
        RECT 40.950 631.050 43.050 633.150 ;
        RECT 53.250 631.950 54.300 640.200 ;
        RECT 59.100 636.150 60.900 637.950 ;
        RECT 55.950 633.150 57.750 634.950 ;
        RECT 58.950 634.050 61.050 636.150 ;
        RECT 72.300 635.400 74.100 647.250 ;
        RECT 76.500 635.400 78.300 647.250 ;
        RECT 79.800 641.400 81.600 647.250 ;
        RECT 95.550 641.400 97.350 647.250 ;
        RECT 98.550 641.400 100.350 647.250 ;
        RECT 101.550 642.000 103.350 647.250 ;
        RECT 98.700 641.100 100.350 641.400 ;
        RECT 104.550 641.400 106.350 647.250 ;
        RECT 118.650 641.400 120.450 647.250 ;
        RECT 121.650 642.000 123.450 647.250 ;
        RECT 104.550 641.100 105.750 641.400 ;
        RECT 98.700 640.200 105.750 641.100 ;
        RECT 98.100 636.150 99.900 637.950 ;
        RECT 62.100 633.150 63.900 634.950 ;
        RECT 52.950 629.850 55.050 631.950 ;
        RECT 55.950 631.050 58.050 633.150 ;
        RECT 61.950 631.050 64.050 633.150 ;
        RECT 71.100 630.150 72.900 631.950 ;
        RECT 76.950 630.150 78.150 635.400 ;
        RECT 79.950 633.150 81.750 634.950 ;
        RECT 95.100 633.150 96.900 634.950 ;
        RECT 97.950 634.050 100.050 636.150 ;
        RECT 101.250 633.150 103.050 634.950 ;
        RECT 79.950 631.050 82.050 633.150 ;
        RECT 94.950 631.050 97.050 633.150 ;
        RECT 100.950 631.050 103.050 633.150 ;
        RECT 104.700 631.950 105.750 640.200 ;
        RECT 119.250 641.100 120.450 641.400 ;
        RECT 124.650 641.400 126.450 647.250 ;
        RECT 127.650 641.400 129.450 647.250 ;
        RECT 137.550 641.400 139.350 647.250 ;
        RECT 140.550 641.400 142.350 647.250 ;
        RECT 154.650 641.400 156.450 647.250 ;
        RECT 157.650 641.400 159.450 647.250 ;
        RECT 169.650 641.400 171.450 647.250 ;
        RECT 172.650 642.000 174.450 647.250 ;
        RECT 124.650 641.100 126.300 641.400 ;
        RECT 119.250 640.200 126.300 641.100 ;
        RECT 119.250 631.950 120.300 640.200 ;
        RECT 125.100 636.150 126.900 637.950 ;
        RECT 121.950 633.150 123.750 634.950 ;
        RECT 124.950 634.050 127.050 636.150 ;
        RECT 128.100 633.150 129.900 634.950 ;
        RECT 13.950 626.850 16.050 628.950 ;
        RECT 17.100 627.150 18.900 628.950 ;
        RECT 14.400 618.600 15.600 626.850 ;
        RECT 16.950 625.050 19.050 627.150 ;
        RECT 32.400 625.650 33.600 629.850 ;
        RECT 53.400 625.650 54.600 629.850 ;
        RECT 70.950 628.050 73.050 630.150 ;
        RECT 73.950 626.850 76.050 628.950 ;
        RECT 76.950 628.050 79.050 630.150 ;
        RECT 103.950 629.850 106.050 631.950 ;
        RECT 118.950 629.850 121.050 631.950 ;
        RECT 121.950 631.050 124.050 633.150 ;
        RECT 127.950 631.050 130.050 633.150 ;
        RECT 32.400 624.000 36.900 625.650 ;
        RECT 13.650 615.750 15.450 618.600 ;
        RECT 16.650 615.750 18.450 618.600 ;
        RECT 35.100 615.750 36.900 624.000 ;
        RECT 40.500 615.750 42.300 624.600 ;
        RECT 53.400 624.000 57.900 625.650 ;
        RECT 74.100 625.050 75.900 626.850 ;
        RECT 77.850 624.750 79.050 628.050 ;
        RECT 104.400 625.650 105.600 629.850 ;
        RECT 56.100 615.750 57.900 624.000 ;
        RECT 61.500 615.750 63.300 624.600 ;
        RECT 78.000 623.700 81.750 624.750 ;
        RECT 71.550 620.700 79.350 622.050 ;
        RECT 71.550 615.750 73.350 620.700 ;
        RECT 74.550 615.750 76.350 619.800 ;
        RECT 77.550 615.750 79.350 620.700 ;
        RECT 80.550 621.600 81.750 623.700 ;
        RECT 80.550 615.750 82.350 621.600 ;
        RECT 95.700 615.750 97.500 624.600 ;
        RECT 101.100 624.000 105.600 625.650 ;
        RECT 119.400 625.650 120.600 629.850 ;
        RECT 140.400 628.950 141.600 641.400 ;
        RECT 155.400 628.950 156.600 641.400 ;
        RECT 170.250 641.100 171.450 641.400 ;
        RECT 175.650 641.400 177.450 647.250 ;
        RECT 178.650 641.400 180.450 647.250 ;
        RECT 193.650 641.400 195.450 647.250 ;
        RECT 196.650 642.000 198.450 647.250 ;
        RECT 175.650 641.100 177.300 641.400 ;
        RECT 170.250 640.200 177.300 641.100 ;
        RECT 194.250 641.100 195.450 641.400 ;
        RECT 199.650 641.400 201.450 647.250 ;
        RECT 202.650 641.400 204.450 647.250 ;
        RECT 199.650 641.100 201.300 641.400 ;
        RECT 194.250 640.200 201.300 641.100 ;
        RECT 170.250 631.950 171.300 640.200 ;
        RECT 176.100 636.150 177.900 637.950 ;
        RECT 172.950 633.150 174.750 634.950 ;
        RECT 175.950 634.050 178.050 636.150 ;
        RECT 179.100 633.150 180.900 634.950 ;
        RECT 169.950 629.850 172.050 631.950 ;
        RECT 172.950 631.050 175.050 633.150 ;
        RECT 178.950 631.050 181.050 633.150 ;
        RECT 194.250 631.950 195.300 640.200 ;
        RECT 200.100 636.150 201.900 637.950 ;
        RECT 196.950 633.150 198.750 634.950 ;
        RECT 199.950 634.050 202.050 636.150 ;
        RECT 216.300 635.400 218.100 647.250 ;
        RECT 220.500 635.400 222.300 647.250 ;
        RECT 223.800 641.400 225.600 647.250 ;
        RECT 239.550 641.400 241.350 647.250 ;
        RECT 242.550 641.400 244.350 647.250 ;
        RECT 257.550 641.400 259.350 647.250 ;
        RECT 260.550 641.400 262.350 647.250 ;
        RECT 263.550 642.000 265.350 647.250 ;
        RECT 203.100 633.150 204.900 634.950 ;
        RECT 193.950 629.850 196.050 631.950 ;
        RECT 196.950 631.050 199.050 633.150 ;
        RECT 202.950 631.050 205.050 633.150 ;
        RECT 215.100 630.150 216.900 631.950 ;
        RECT 220.950 630.150 222.150 635.400 ;
        RECT 223.950 633.150 225.750 634.950 ;
        RECT 223.950 631.050 226.050 633.150 ;
        RECT 137.100 627.150 138.900 628.950 ;
        RECT 119.400 624.000 123.900 625.650 ;
        RECT 136.950 625.050 139.050 627.150 ;
        RECT 139.950 626.850 142.050 628.950 ;
        RECT 154.950 626.850 157.050 628.950 ;
        RECT 158.100 627.150 159.900 628.950 ;
        RECT 101.100 615.750 102.900 624.000 ;
        RECT 122.100 615.750 123.900 624.000 ;
        RECT 127.500 615.750 129.300 624.600 ;
        RECT 140.400 618.600 141.600 626.850 ;
        RECT 155.400 618.600 156.600 626.850 ;
        RECT 157.950 625.050 160.050 627.150 ;
        RECT 170.400 625.650 171.600 629.850 ;
        RECT 194.400 625.650 195.600 629.850 ;
        RECT 214.950 628.050 217.050 630.150 ;
        RECT 217.950 626.850 220.050 628.950 ;
        RECT 220.950 628.050 223.050 630.150 ;
        RECT 242.400 628.950 243.600 641.400 ;
        RECT 260.700 641.100 262.350 641.400 ;
        RECT 266.550 641.400 268.350 647.250 ;
        RECT 278.550 641.400 280.350 647.250 ;
        RECT 281.550 641.400 283.350 647.250 ;
        RECT 284.550 642.000 286.350 647.250 ;
        RECT 266.550 641.100 267.750 641.400 ;
        RECT 260.700 640.200 267.750 641.100 ;
        RECT 281.700 641.100 283.350 641.400 ;
        RECT 287.550 641.400 289.350 647.250 ;
        RECT 301.650 641.400 303.450 647.250 ;
        RECT 304.650 641.400 306.450 647.250 ;
        RECT 287.550 641.100 288.750 641.400 ;
        RECT 281.700 640.200 288.750 641.100 ;
        RECT 260.100 636.150 261.900 637.950 ;
        RECT 257.100 633.150 258.900 634.950 ;
        RECT 259.950 634.050 262.050 636.150 ;
        RECT 263.250 633.150 265.050 634.950 ;
        RECT 256.950 631.050 259.050 633.150 ;
        RECT 262.950 631.050 265.050 633.150 ;
        RECT 266.700 631.950 267.750 640.200 ;
        RECT 281.100 636.150 282.900 637.950 ;
        RECT 278.100 633.150 279.900 634.950 ;
        RECT 280.950 634.050 283.050 636.150 ;
        RECT 284.250 633.150 286.050 634.950 ;
        RECT 265.950 629.850 268.050 631.950 ;
        RECT 277.950 631.050 280.050 633.150 ;
        RECT 283.950 631.050 286.050 633.150 ;
        RECT 287.700 631.950 288.750 640.200 ;
        RECT 286.950 629.850 289.050 631.950 ;
        RECT 170.400 624.000 174.900 625.650 ;
        RECT 137.550 615.750 139.350 618.600 ;
        RECT 140.550 615.750 142.350 618.600 ;
        RECT 154.650 615.750 156.450 618.600 ;
        RECT 157.650 615.750 159.450 618.600 ;
        RECT 173.100 615.750 174.900 624.000 ;
        RECT 178.500 615.750 180.300 624.600 ;
        RECT 194.400 624.000 198.900 625.650 ;
        RECT 218.100 625.050 219.900 626.850 ;
        RECT 221.850 624.750 223.050 628.050 ;
        RECT 239.100 627.150 240.900 628.950 ;
        RECT 238.950 625.050 241.050 627.150 ;
        RECT 241.950 626.850 244.050 628.950 ;
        RECT 197.100 615.750 198.900 624.000 ;
        RECT 202.500 615.750 204.300 624.600 ;
        RECT 222.000 623.700 225.750 624.750 ;
        RECT 215.550 620.700 223.350 622.050 ;
        RECT 215.550 615.750 217.350 620.700 ;
        RECT 218.550 615.750 220.350 619.800 ;
        RECT 221.550 615.750 223.350 620.700 ;
        RECT 224.550 621.600 225.750 623.700 ;
        RECT 224.550 615.750 226.350 621.600 ;
        RECT 242.400 618.600 243.600 626.850 ;
        RECT 266.400 625.650 267.600 629.850 ;
        RECT 287.400 625.650 288.600 629.850 ;
        RECT 302.400 628.950 303.600 641.400 ;
        RECT 308.550 635.400 310.350 647.250 ;
        RECT 311.550 644.400 313.350 647.250 ;
        RECT 316.050 641.400 317.850 647.250 ;
        RECT 320.250 641.400 322.050 647.250 ;
        RECT 313.950 639.300 317.850 641.400 ;
        RECT 324.150 640.500 325.950 647.250 ;
        RECT 327.150 641.400 328.950 647.250 ;
        RECT 331.950 641.400 333.750 647.250 ;
        RECT 337.050 641.400 338.850 647.250 ;
        RECT 332.250 640.500 333.450 641.400 ;
        RECT 322.950 638.700 329.850 640.500 ;
        RECT 332.250 638.400 337.050 640.500 ;
        RECT 315.150 636.600 317.850 638.400 ;
        RECT 318.750 637.800 320.550 638.400 ;
        RECT 318.750 636.900 325.050 637.800 ;
        RECT 332.250 637.500 333.450 638.400 ;
        RECT 318.750 636.600 320.550 636.900 ;
        RECT 316.950 635.700 317.850 636.600 ;
        RECT 301.950 626.850 304.050 628.950 ;
        RECT 305.100 627.150 306.900 628.950 ;
        RECT 239.550 615.750 241.350 618.600 ;
        RECT 242.550 615.750 244.350 618.600 ;
        RECT 257.700 615.750 259.500 624.600 ;
        RECT 263.100 624.000 267.600 625.650 ;
        RECT 263.100 615.750 264.900 624.000 ;
        RECT 278.700 615.750 280.500 624.600 ;
        RECT 284.100 624.000 288.600 625.650 ;
        RECT 284.100 615.750 285.900 624.000 ;
        RECT 302.400 618.600 303.600 626.850 ;
        RECT 304.950 625.050 307.050 627.150 ;
        RECT 308.550 625.950 309.750 635.400 ;
        RECT 313.950 634.800 316.050 635.700 ;
        RECT 316.950 634.800 322.950 635.700 ;
        RECT 311.850 633.600 316.050 634.800 ;
        RECT 310.950 631.800 312.750 633.600 ;
        RECT 322.050 630.150 322.950 634.800 ;
        RECT 324.150 634.800 325.050 636.900 ;
        RECT 325.950 636.300 333.450 637.500 ;
        RECT 325.950 635.700 327.750 636.300 ;
        RECT 340.050 635.400 341.850 647.250 ;
        RECT 351.300 635.400 353.100 647.250 ;
        RECT 355.500 635.400 357.300 647.250 ;
        RECT 358.800 641.400 360.600 647.250 ;
        RECT 371.550 641.400 373.350 647.250 ;
        RECT 374.550 641.400 376.350 647.250 ;
        RECT 377.550 641.400 379.350 647.250 ;
        RECT 330.750 634.800 341.850 635.400 ;
        RECT 324.150 634.200 341.850 634.800 ;
        RECT 324.150 633.900 332.550 634.200 ;
        RECT 330.750 633.600 332.550 633.900 ;
        RECT 322.050 628.050 325.050 630.150 ;
        RECT 328.950 629.100 331.050 630.150 ;
        RECT 328.950 628.050 336.900 629.100 ;
        RECT 310.950 627.750 313.050 628.050 ;
        RECT 310.950 625.950 314.850 627.750 ;
        RECT 308.550 623.850 313.050 625.950 ;
        RECT 322.050 624.000 322.950 628.050 ;
        RECT 335.100 627.300 336.900 628.050 ;
        RECT 338.100 627.150 339.900 628.950 ;
        RECT 332.100 626.400 333.900 627.000 ;
        RECT 338.100 626.400 339.000 627.150 ;
        RECT 332.100 625.200 339.000 626.400 ;
        RECT 332.100 624.000 333.150 625.200 ;
        RECT 308.550 621.600 309.750 623.850 ;
        RECT 322.050 623.100 333.150 624.000 ;
        RECT 322.050 622.800 322.950 623.100 ;
        RECT 301.650 615.750 303.450 618.600 ;
        RECT 304.650 615.750 306.450 618.600 ;
        RECT 308.550 615.750 310.350 621.600 ;
        RECT 313.950 620.700 316.050 621.600 ;
        RECT 321.150 621.000 322.950 622.800 ;
        RECT 332.100 622.200 333.150 623.100 ;
        RECT 328.350 621.450 330.150 622.200 ;
        RECT 313.950 619.500 317.700 620.700 ;
        RECT 316.650 618.600 317.700 619.500 ;
        RECT 325.200 620.400 330.150 621.450 ;
        RECT 331.650 620.400 333.450 622.200 ;
        RECT 340.950 621.600 341.850 634.200 ;
        RECT 350.100 630.150 351.900 631.950 ;
        RECT 355.950 630.150 357.150 635.400 ;
        RECT 358.950 633.150 360.750 634.950 ;
        RECT 374.550 633.150 375.750 641.400 ;
        RECT 389.550 635.400 391.350 647.250 ;
        RECT 393.750 635.400 395.550 647.250 ;
        RECT 409.650 635.400 411.450 647.250 ;
        RECT 412.650 636.300 414.450 647.250 ;
        RECT 415.650 637.200 417.450 647.250 ;
        RECT 418.650 636.300 420.450 647.250 ;
        RECT 428.550 641.400 430.350 647.250 ;
        RECT 431.550 641.400 433.350 647.250 ;
        RECT 443.550 641.400 445.350 647.250 ;
        RECT 446.550 641.400 448.350 647.250 ;
        RECT 449.550 641.400 451.350 647.250 ;
        RECT 463.650 641.400 465.450 647.250 ;
        RECT 466.650 641.400 468.450 647.250 ;
        RECT 479.550 641.400 481.350 647.250 ;
        RECT 482.550 641.400 484.350 647.250 ;
        RECT 500.400 641.400 502.200 647.250 ;
        RECT 412.650 635.400 420.450 636.300 ;
        RECT 393.000 634.350 395.550 635.400 ;
        RECT 358.950 631.050 361.050 633.150 ;
        RECT 349.950 628.050 352.050 630.150 ;
        RECT 352.950 626.850 355.050 628.950 ;
        RECT 355.950 628.050 358.050 630.150 ;
        RECT 370.950 629.850 373.050 631.950 ;
        RECT 373.950 631.050 376.050 633.150 ;
        RECT 371.100 628.050 372.900 629.850 ;
        RECT 353.100 625.050 354.900 626.850 ;
        RECT 356.850 624.750 358.050 628.050 ;
        RECT 357.000 623.700 360.750 624.750 ;
        RECT 325.200 618.600 326.250 620.400 ;
        RECT 334.950 619.500 337.050 621.600 ;
        RECT 334.950 618.600 336.000 619.500 ;
        RECT 311.850 615.750 313.650 618.600 ;
        RECT 316.350 615.750 318.150 618.600 ;
        RECT 320.550 615.750 322.350 618.600 ;
        RECT 324.450 615.750 326.250 618.600 ;
        RECT 327.750 615.750 329.550 618.600 ;
        RECT 332.250 617.700 336.000 618.600 ;
        RECT 332.250 615.750 334.050 617.700 ;
        RECT 337.050 615.750 338.850 618.600 ;
        RECT 340.050 615.750 341.850 621.600 ;
        RECT 350.550 620.700 358.350 622.050 ;
        RECT 350.550 615.750 352.350 620.700 ;
        RECT 353.550 615.750 355.350 619.800 ;
        RECT 356.550 615.750 358.350 620.700 ;
        RECT 359.550 621.600 360.750 623.700 ;
        RECT 374.550 623.700 375.750 631.050 ;
        RECT 376.950 629.850 379.050 631.950 ;
        RECT 389.100 630.150 390.900 631.950 ;
        RECT 377.100 628.050 378.900 629.850 ;
        RECT 388.950 628.050 391.050 630.150 ;
        RECT 393.000 627.150 394.050 634.350 ;
        RECT 395.100 630.150 396.900 631.950 ;
        RECT 410.100 630.150 411.300 635.400 ;
        RECT 394.950 628.050 397.050 630.150 ;
        RECT 409.950 628.050 412.050 630.150 ;
        RECT 431.400 628.950 432.600 641.400 ;
        RECT 446.550 633.150 447.750 641.400 ;
        RECT 442.950 629.850 445.050 631.950 ;
        RECT 445.950 631.050 448.050 633.150 ;
        RECT 391.950 625.050 394.050 627.150 ;
        RECT 374.550 622.800 378.150 623.700 ;
        RECT 359.550 615.750 361.350 621.600 ;
        RECT 371.850 615.750 373.650 621.600 ;
        RECT 376.350 615.750 378.150 622.800 ;
        RECT 393.000 618.600 394.050 625.050 ;
        RECT 410.100 621.600 411.300 628.050 ;
        RECT 412.950 626.850 415.050 628.950 ;
        RECT 416.100 627.150 417.900 628.950 ;
        RECT 413.100 625.050 414.900 626.850 ;
        RECT 415.950 625.050 418.050 627.150 ;
        RECT 418.950 626.850 421.050 628.950 ;
        RECT 428.100 627.150 429.900 628.950 ;
        RECT 419.100 625.050 420.900 626.850 ;
        RECT 427.950 625.050 430.050 627.150 ;
        RECT 430.950 626.850 433.050 628.950 ;
        RECT 443.100 628.050 444.900 629.850 ;
        RECT 410.100 619.950 415.800 621.600 ;
        RECT 389.550 615.750 391.350 618.600 ;
        RECT 392.550 615.750 394.350 618.600 ;
        RECT 395.550 615.750 397.350 618.600 ;
        RECT 410.700 615.750 412.500 618.600 ;
        RECT 414.000 615.750 415.800 619.950 ;
        RECT 418.200 615.750 420.000 621.600 ;
        RECT 431.400 618.600 432.600 626.850 ;
        RECT 446.550 623.700 447.750 631.050 ;
        RECT 448.950 629.850 451.050 631.950 ;
        RECT 449.100 628.050 450.900 629.850 ;
        RECT 464.400 628.950 465.600 641.400 ;
        RECT 482.400 628.950 483.600 641.400 ;
        RECT 503.700 635.400 505.500 647.250 ;
        RECT 507.900 635.400 509.700 647.250 ;
        RECT 523.650 641.400 525.450 647.250 ;
        RECT 526.650 641.400 528.450 647.250 ;
        RECT 539.400 641.400 541.200 647.250 ;
        RECT 500.250 633.150 502.050 634.950 ;
        RECT 499.950 631.050 502.050 633.150 ;
        RECT 503.850 630.150 505.050 635.400 ;
        RECT 509.100 630.150 510.900 631.950 ;
        RECT 463.950 626.850 466.050 628.950 ;
        RECT 467.100 627.150 468.900 628.950 ;
        RECT 479.100 627.150 480.900 628.950 ;
        RECT 446.550 622.800 450.150 623.700 ;
        RECT 428.550 615.750 430.350 618.600 ;
        RECT 431.550 615.750 433.350 618.600 ;
        RECT 443.850 615.750 445.650 621.600 ;
        RECT 448.350 615.750 450.150 622.800 ;
        RECT 464.400 618.600 465.600 626.850 ;
        RECT 466.950 625.050 469.050 627.150 ;
        RECT 478.950 625.050 481.050 627.150 ;
        RECT 481.950 626.850 484.050 628.950 ;
        RECT 502.950 628.050 505.050 630.150 ;
        RECT 482.400 618.600 483.600 626.850 ;
        RECT 502.950 624.750 504.150 628.050 ;
        RECT 505.950 626.850 508.050 628.950 ;
        RECT 508.950 628.050 511.050 630.150 ;
        RECT 524.400 628.950 525.600 641.400 ;
        RECT 542.700 635.400 544.500 647.250 ;
        RECT 546.900 635.400 548.700 647.250 ;
        RECT 557.550 635.400 559.350 647.250 ;
        RECT 561.750 635.400 563.550 647.250 ;
        RECT 580.650 641.400 582.450 647.250 ;
        RECT 583.650 641.400 585.450 647.250 ;
        RECT 596.400 641.400 598.200 647.250 ;
        RECT 539.250 633.150 541.050 634.950 ;
        RECT 538.950 631.050 541.050 633.150 ;
        RECT 542.850 630.150 544.050 635.400 ;
        RECT 561.000 634.350 563.550 635.400 ;
        RECT 548.100 630.150 549.900 631.950 ;
        RECT 557.100 630.150 558.900 631.950 ;
        RECT 523.950 626.850 526.050 628.950 ;
        RECT 527.100 627.150 528.900 628.950 ;
        RECT 541.950 628.050 544.050 630.150 ;
        RECT 506.100 625.050 507.900 626.850 ;
        RECT 500.250 623.700 504.000 624.750 ;
        RECT 500.250 621.600 501.450 623.700 ;
        RECT 463.650 615.750 465.450 618.600 ;
        RECT 466.650 615.750 468.450 618.600 ;
        RECT 479.550 615.750 481.350 618.600 ;
        RECT 482.550 615.750 484.350 618.600 ;
        RECT 499.650 615.750 501.450 621.600 ;
        RECT 502.650 620.700 510.450 622.050 ;
        RECT 502.650 615.750 504.450 620.700 ;
        RECT 505.650 615.750 507.450 619.800 ;
        RECT 508.650 615.750 510.450 620.700 ;
        RECT 524.400 618.600 525.600 626.850 ;
        RECT 526.950 625.050 529.050 627.150 ;
        RECT 541.950 624.750 543.150 628.050 ;
        RECT 544.950 626.850 547.050 628.950 ;
        RECT 547.950 628.050 550.050 630.150 ;
        RECT 556.950 628.050 559.050 630.150 ;
        RECT 561.000 627.150 562.050 634.350 ;
        RECT 563.100 630.150 564.900 631.950 ;
        RECT 562.950 628.050 565.050 630.150 ;
        RECT 581.400 628.950 582.600 641.400 ;
        RECT 599.700 635.400 601.500 647.250 ;
        RECT 603.900 635.400 605.700 647.250 ;
        RECT 616.650 641.400 618.450 647.250 ;
        RECT 619.650 641.400 621.450 647.250 ;
        RECT 596.250 633.150 598.050 634.950 ;
        RECT 595.950 631.050 598.050 633.150 ;
        RECT 599.850 630.150 601.050 635.400 ;
        RECT 605.100 630.150 606.900 631.950 ;
        RECT 545.100 625.050 546.900 626.850 ;
        RECT 559.950 625.050 562.050 627.150 ;
        RECT 580.950 626.850 583.050 628.950 ;
        RECT 584.100 627.150 585.900 628.950 ;
        RECT 598.950 628.050 601.050 630.150 ;
        RECT 539.250 623.700 543.000 624.750 ;
        RECT 539.250 621.600 540.450 623.700 ;
        RECT 523.650 615.750 525.450 618.600 ;
        RECT 526.650 615.750 528.450 618.600 ;
        RECT 538.650 615.750 540.450 621.600 ;
        RECT 541.650 620.700 549.450 622.050 ;
        RECT 541.650 615.750 543.450 620.700 ;
        RECT 544.650 615.750 546.450 619.800 ;
        RECT 547.650 615.750 549.450 620.700 ;
        RECT 561.000 618.600 562.050 625.050 ;
        RECT 581.400 618.600 582.600 626.850 ;
        RECT 583.950 625.050 586.050 627.150 ;
        RECT 598.950 624.750 600.150 628.050 ;
        RECT 601.950 626.850 604.050 628.950 ;
        RECT 604.950 628.050 607.050 630.150 ;
        RECT 617.400 628.950 618.600 641.400 ;
        RECT 632.550 636.300 634.350 647.250 ;
        RECT 635.550 637.200 637.350 647.250 ;
        RECT 638.550 636.300 640.350 647.250 ;
        RECT 632.550 635.400 640.350 636.300 ;
        RECT 641.550 635.400 643.350 647.250 ;
        RECT 658.650 641.400 660.450 647.250 ;
        RECT 661.650 641.400 663.450 647.250 ;
        RECT 664.650 641.400 666.450 647.250 ;
        RECT 677.400 641.400 679.200 647.250 ;
        RECT 641.700 630.150 642.900 635.400 ;
        RECT 662.250 633.150 663.450 641.400 ;
        RECT 680.700 635.400 682.500 647.250 ;
        RECT 684.900 635.400 686.700 647.250 ;
        RECT 695.550 641.400 697.350 647.250 ;
        RECT 698.550 641.400 700.350 647.250 ;
        RECT 677.250 633.150 679.050 634.950 ;
        RECT 616.950 626.850 619.050 628.950 ;
        RECT 620.100 627.150 621.900 628.950 ;
        RECT 602.100 625.050 603.900 626.850 ;
        RECT 596.250 623.700 600.000 624.750 ;
        RECT 596.250 621.600 597.450 623.700 ;
        RECT 557.550 615.750 559.350 618.600 ;
        RECT 560.550 615.750 562.350 618.600 ;
        RECT 563.550 615.750 565.350 618.600 ;
        RECT 580.650 615.750 582.450 618.600 ;
        RECT 583.650 615.750 585.450 618.600 ;
        RECT 595.650 615.750 597.450 621.600 ;
        RECT 598.650 620.700 606.450 622.050 ;
        RECT 598.650 615.750 600.450 620.700 ;
        RECT 601.650 615.750 603.450 619.800 ;
        RECT 604.650 615.750 606.450 620.700 ;
        RECT 617.400 618.600 618.600 626.850 ;
        RECT 619.950 625.050 622.050 627.150 ;
        RECT 631.950 626.850 634.050 628.950 ;
        RECT 635.100 627.150 636.900 628.950 ;
        RECT 632.100 625.050 633.900 626.850 ;
        RECT 634.950 625.050 637.050 627.150 ;
        RECT 637.950 626.850 640.050 628.950 ;
        RECT 640.950 628.050 643.050 630.150 ;
        RECT 658.950 629.850 661.050 631.950 ;
        RECT 661.950 631.050 664.050 633.150 ;
        RECT 659.100 628.050 660.900 629.850 ;
        RECT 638.100 625.050 639.900 626.850 ;
        RECT 641.700 621.600 642.900 628.050 ;
        RECT 662.250 623.700 663.450 631.050 ;
        RECT 664.950 629.850 667.050 631.950 ;
        RECT 676.950 631.050 679.050 633.150 ;
        RECT 680.850 630.150 682.050 635.400 ;
        RECT 686.100 630.150 687.900 631.950 ;
        RECT 695.100 630.150 696.900 631.950 ;
        RECT 665.100 628.050 666.900 629.850 ;
        RECT 679.950 628.050 682.050 630.150 ;
        RECT 679.950 624.750 681.150 628.050 ;
        RECT 682.950 626.850 685.050 628.950 ;
        RECT 685.950 628.050 688.050 630.150 ;
        RECT 694.950 628.050 697.050 630.150 ;
        RECT 683.100 625.050 684.900 626.850 ;
        RECT 616.650 615.750 618.450 618.600 ;
        RECT 619.650 615.750 621.450 618.600 ;
        RECT 633.000 615.750 634.800 621.600 ;
        RECT 637.200 619.950 642.900 621.600 ;
        RECT 659.850 622.800 663.450 623.700 ;
        RECT 677.250 623.700 681.000 624.750 ;
        RECT 698.700 624.300 699.900 641.400 ;
        RECT 702.150 635.400 703.950 647.250 ;
        RECT 705.150 635.400 706.950 647.250 ;
        RECT 719.550 635.400 721.350 647.250 ;
        RECT 724.050 635.550 725.850 647.250 ;
        RECT 727.050 636.900 728.850 647.250 ;
        RECT 727.050 635.550 729.450 636.900 ;
        RECT 700.950 629.850 703.050 631.950 ;
        RECT 705.150 630.150 706.350 635.400 ;
        RECT 719.550 634.200 720.750 635.400 ;
        RECT 724.950 634.200 726.750 634.650 ;
        RECT 719.550 633.000 726.750 634.200 ;
        RECT 724.950 632.850 726.750 633.000 ;
        RECT 722.100 630.150 723.900 631.950 ;
        RECT 701.100 628.050 702.900 629.850 ;
        RECT 703.950 628.050 706.350 630.150 ;
        RECT 637.200 615.750 639.000 619.950 ;
        RECT 640.500 615.750 642.300 618.600 ;
        RECT 659.850 615.750 661.650 622.800 ;
        RECT 677.250 621.600 678.450 623.700 ;
        RECT 695.550 623.100 703.050 624.300 ;
        RECT 664.350 615.750 666.150 621.600 ;
        RECT 676.650 615.750 678.450 621.600 ;
        RECT 679.650 620.700 687.450 622.050 ;
        RECT 679.650 615.750 681.450 620.700 ;
        RECT 682.650 615.750 684.450 619.800 ;
        RECT 685.650 615.750 687.450 620.700 ;
        RECT 695.550 615.750 697.350 623.100 ;
        RECT 701.250 622.500 703.050 623.100 ;
        RECT 705.150 621.600 706.350 628.050 ;
        RECT 719.100 627.150 720.900 628.950 ;
        RECT 721.950 628.050 724.050 630.150 ;
        RECT 718.950 625.050 721.050 627.150 ;
        RECT 725.700 624.600 726.600 632.850 ;
        RECT 728.100 628.950 729.450 635.550 ;
        RECT 735.150 635.400 736.950 647.250 ;
        RECT 738.150 641.400 739.950 647.250 ;
        RECT 743.250 641.400 745.050 647.250 ;
        RECT 748.050 641.400 749.850 647.250 ;
        RECT 743.550 640.500 744.750 641.400 ;
        RECT 751.050 640.500 752.850 647.250 ;
        RECT 754.950 641.400 756.750 647.250 ;
        RECT 759.150 641.400 760.950 647.250 ;
        RECT 763.650 644.400 765.450 647.250 ;
        RECT 739.950 638.400 744.750 640.500 ;
        RECT 747.150 638.700 754.050 640.500 ;
        RECT 759.150 639.300 763.050 641.400 ;
        RECT 743.550 637.500 744.750 638.400 ;
        RECT 756.450 637.800 758.250 638.400 ;
        RECT 743.550 636.300 751.050 637.500 ;
        RECT 749.250 635.700 751.050 636.300 ;
        RECT 751.950 636.900 758.250 637.800 ;
        RECT 735.150 634.800 746.250 635.400 ;
        RECT 751.950 634.800 752.850 636.900 ;
        RECT 756.450 636.600 758.250 636.900 ;
        RECT 759.150 636.600 761.850 638.400 ;
        RECT 759.150 635.700 760.050 636.600 ;
        RECT 735.150 634.200 752.850 634.800 ;
        RECT 727.950 626.850 730.050 628.950 ;
        RECT 724.950 623.700 726.750 624.600 ;
        RECT 700.050 615.750 701.850 621.600 ;
        RECT 703.050 620.100 706.350 621.600 ;
        RECT 723.450 622.800 726.750 623.700 ;
        RECT 703.050 615.750 704.850 620.100 ;
        RECT 723.450 618.600 724.350 622.800 ;
        RECT 729.000 621.600 730.050 626.850 ;
        RECT 735.150 621.600 736.050 634.200 ;
        RECT 744.450 633.900 752.850 634.200 ;
        RECT 754.050 634.800 760.050 635.700 ;
        RECT 760.950 634.800 763.050 635.700 ;
        RECT 766.650 635.400 768.450 647.250 ;
        RECT 781.650 646.500 789.450 647.250 ;
        RECT 781.650 635.400 783.450 646.500 ;
        RECT 784.650 635.400 786.450 645.600 ;
        RECT 787.650 636.600 789.450 646.500 ;
        RECT 790.650 637.500 792.450 647.250 ;
        RECT 793.650 636.600 795.450 647.250 ;
        RECT 805.650 641.400 807.450 647.250 ;
        RECT 808.650 641.400 810.450 647.250 ;
        RECT 811.650 641.400 813.450 647.250 ;
        RECT 787.650 635.700 795.450 636.600 ;
        RECT 744.450 633.600 746.250 633.900 ;
        RECT 754.050 630.150 754.950 634.800 ;
        RECT 760.950 633.600 765.150 634.800 ;
        RECT 764.250 631.800 766.050 633.600 ;
        RECT 745.950 629.100 748.050 630.150 ;
        RECT 737.100 627.150 738.900 628.950 ;
        RECT 740.100 628.050 748.050 629.100 ;
        RECT 751.950 628.050 754.950 630.150 ;
        RECT 740.100 627.300 741.900 628.050 ;
        RECT 738.000 626.400 738.900 627.150 ;
        RECT 743.100 626.400 744.900 627.000 ;
        RECT 738.000 625.200 744.900 626.400 ;
        RECT 743.850 624.000 744.900 625.200 ;
        RECT 754.050 624.000 754.950 628.050 ;
        RECT 763.950 627.750 766.050 628.050 ;
        RECT 762.150 625.950 766.050 627.750 ;
        RECT 767.250 625.950 768.450 635.400 ;
        RECT 784.800 634.500 786.600 635.400 ;
        RECT 784.800 633.600 788.850 634.500 ;
        RECT 782.100 630.150 783.900 631.950 ;
        RECT 787.950 630.150 788.850 633.600 ;
        RECT 809.250 633.150 810.450 641.400 ;
        RECT 821.550 635.400 823.350 647.250 ;
        RECT 826.050 635.550 827.850 647.250 ;
        RECT 829.050 636.900 830.850 647.250 ;
        RECT 845.550 641.400 847.350 647.250 ;
        RECT 848.550 641.400 850.350 647.250 ;
        RECT 851.550 641.400 853.350 647.250 ;
        RECT 829.050 635.550 831.450 636.900 ;
        RECT 821.550 634.200 822.750 635.400 ;
        RECT 826.950 634.200 828.750 634.650 ;
        RECT 793.950 630.150 795.750 631.950 ;
        RECT 781.950 628.050 784.050 630.150 ;
        RECT 784.950 626.850 787.050 628.950 ;
        RECT 787.950 628.050 790.050 630.150 ;
        RECT 743.850 623.100 754.950 624.000 ;
        RECT 763.950 623.850 768.450 625.950 ;
        RECT 785.250 625.050 787.050 626.850 ;
        RECT 743.850 622.200 744.900 623.100 ;
        RECT 754.050 622.800 754.950 623.100 ;
        RECT 719.550 615.750 721.350 618.600 ;
        RECT 722.550 615.750 724.350 618.600 ;
        RECT 725.550 615.750 727.350 618.600 ;
        RECT 728.550 615.750 730.350 621.600 ;
        RECT 735.150 615.750 736.950 621.600 ;
        RECT 739.950 619.500 742.050 621.600 ;
        RECT 743.550 620.400 745.350 622.200 ;
        RECT 746.850 621.450 748.650 622.200 ;
        RECT 746.850 620.400 751.800 621.450 ;
        RECT 754.050 621.000 755.850 622.800 ;
        RECT 767.250 621.600 768.450 623.850 ;
        RECT 789.000 621.600 790.050 628.050 ;
        RECT 790.950 626.850 793.050 628.950 ;
        RECT 793.950 628.050 796.050 630.150 ;
        RECT 805.950 629.850 808.050 631.950 ;
        RECT 808.950 631.050 811.050 633.150 ;
        RECT 821.550 633.000 828.750 634.200 ;
        RECT 826.950 632.850 828.750 633.000 ;
        RECT 806.100 628.050 807.900 629.850 ;
        RECT 790.950 625.050 792.750 626.850 ;
        RECT 809.250 623.700 810.450 631.050 ;
        RECT 811.950 629.850 814.050 631.950 ;
        RECT 824.100 630.150 825.900 631.950 ;
        RECT 812.100 628.050 813.900 629.850 ;
        RECT 821.100 627.150 822.900 628.950 ;
        RECT 823.950 628.050 826.050 630.150 ;
        RECT 820.950 625.050 823.050 627.150 ;
        RECT 827.700 624.600 828.600 632.850 ;
        RECT 830.100 628.950 831.450 635.550 ;
        RECT 848.550 633.150 849.750 641.400 ;
        RECT 867.450 635.400 869.250 647.250 ;
        RECT 871.650 635.400 873.450 647.250 ;
        RECT 867.450 634.350 870.000 635.400 ;
        RECT 844.950 629.850 847.050 631.950 ;
        RECT 847.950 631.050 850.050 633.150 ;
        RECT 829.950 626.850 832.050 628.950 ;
        RECT 845.100 628.050 846.900 629.850 ;
        RECT 826.950 623.700 828.750 624.600 ;
        RECT 806.850 622.800 810.450 623.700 ;
        RECT 825.450 622.800 828.750 623.700 ;
        RECT 760.950 620.700 763.050 621.600 ;
        RECT 741.000 618.600 742.050 619.500 ;
        RECT 750.750 618.600 751.800 620.400 ;
        RECT 759.300 619.500 763.050 620.700 ;
        RECT 759.300 618.600 760.350 619.500 ;
        RECT 738.150 615.750 739.950 618.600 ;
        RECT 741.000 617.700 744.750 618.600 ;
        RECT 742.950 615.750 744.750 617.700 ;
        RECT 747.450 615.750 749.250 618.600 ;
        RECT 750.750 615.750 752.550 618.600 ;
        RECT 754.650 615.750 756.450 618.600 ;
        RECT 758.850 615.750 760.650 618.600 ;
        RECT 763.350 615.750 765.150 618.600 ;
        RECT 766.650 615.750 768.450 621.600 ;
        RECT 784.800 615.750 786.600 621.600 ;
        RECT 789.000 615.750 790.800 621.600 ;
        RECT 793.200 615.750 795.000 621.600 ;
        RECT 806.850 615.750 808.650 622.800 ;
        RECT 811.350 615.750 813.150 621.600 ;
        RECT 825.450 618.600 826.350 622.800 ;
        RECT 831.000 621.600 832.050 626.850 ;
        RECT 848.550 623.700 849.750 631.050 ;
        RECT 850.950 629.850 853.050 631.950 ;
        RECT 866.100 630.150 867.900 631.950 ;
        RECT 851.100 628.050 852.900 629.850 ;
        RECT 865.950 628.050 868.050 630.150 ;
        RECT 859.950 625.950 862.050 628.050 ;
        RECT 868.950 627.150 870.000 634.350 ;
        RECT 872.100 630.150 873.900 631.950 ;
        RECT 871.950 628.050 874.050 630.150 ;
        RECT 848.550 622.800 852.150 623.700 ;
        RECT 821.550 615.750 823.350 618.600 ;
        RECT 824.550 615.750 826.350 618.600 ;
        RECT 827.550 615.750 829.350 618.600 ;
        RECT 830.550 615.750 832.350 621.600 ;
        RECT 845.850 615.750 847.650 621.600 ;
        RECT 850.350 615.750 852.150 622.800 ;
        RECT 860.550 621.450 861.450 625.950 ;
        RECT 868.950 625.050 871.050 627.150 ;
        RECT 865.950 621.450 868.050 622.050 ;
        RECT 860.550 620.550 868.050 621.450 ;
        RECT 865.950 619.950 868.050 620.550 ;
        RECT 868.950 618.600 870.000 625.050 ;
        RECT 865.650 615.750 867.450 618.600 ;
        RECT 868.650 615.750 870.450 618.600 ;
        RECT 871.650 615.750 873.450 618.600 ;
        RECT 10.650 608.400 12.450 611.250 ;
        RECT 13.650 608.400 15.450 611.250 ;
        RECT 25.650 608.400 27.450 611.250 ;
        RECT 28.650 608.400 30.450 611.250 ;
        RECT 38.550 608.400 40.350 611.250 ;
        RECT 41.550 608.400 43.350 611.250 ;
        RECT 44.550 608.400 46.350 611.250 ;
        RECT 11.400 600.150 12.600 608.400 ;
        RECT 10.950 598.050 13.050 600.150 ;
        RECT 13.950 599.850 16.050 601.950 ;
        RECT 26.400 600.150 27.600 608.400 ;
        RECT 42.450 604.200 43.350 608.400 ;
        RECT 47.550 605.400 49.350 611.250 ;
        RECT 62.550 606.300 64.350 611.250 ;
        RECT 65.550 607.200 67.350 611.250 ;
        RECT 68.550 606.300 70.350 611.250 ;
        RECT 42.450 603.300 45.750 604.200 ;
        RECT 43.950 602.400 45.750 603.300 ;
        RECT 14.100 598.050 15.900 599.850 ;
        RECT 25.950 598.050 28.050 600.150 ;
        RECT 28.950 599.850 31.050 601.950 ;
        RECT 37.950 599.850 40.050 601.950 ;
        RECT 29.100 598.050 30.900 599.850 ;
        RECT 38.100 598.050 39.900 599.850 ;
        RECT 11.400 585.600 12.600 598.050 ;
        RECT 26.400 585.600 27.600 598.050 ;
        RECT 40.950 596.850 43.050 598.950 ;
        RECT 41.100 595.050 42.900 596.850 ;
        RECT 44.700 594.150 45.600 602.400 ;
        RECT 48.000 600.150 49.050 605.400 ;
        RECT 62.550 604.950 70.350 606.300 ;
        RECT 71.550 605.400 73.350 611.250 ;
        RECT 85.350 605.400 87.150 611.250 ;
        RECT 88.350 605.400 90.150 611.250 ;
        RECT 91.650 608.400 93.450 611.250 ;
        RECT 71.550 603.300 72.750 605.400 ;
        RECT 69.000 602.250 72.750 603.300 ;
        RECT 65.100 600.150 66.900 601.950 ;
        RECT 46.950 598.050 49.050 600.150 ;
        RECT 43.950 594.000 45.750 594.150 ;
        RECT 38.550 592.800 45.750 594.000 ;
        RECT 38.550 591.600 39.750 592.800 ;
        RECT 43.950 592.350 45.750 592.800 ;
        RECT 10.650 579.750 12.450 585.600 ;
        RECT 13.650 579.750 15.450 585.600 ;
        RECT 25.650 579.750 27.450 585.600 ;
        RECT 28.650 579.750 30.450 585.600 ;
        RECT 38.550 579.750 40.350 591.600 ;
        RECT 47.100 591.450 48.450 598.050 ;
        RECT 61.950 596.850 64.050 598.950 ;
        RECT 64.950 598.050 67.050 600.150 ;
        RECT 68.850 598.950 70.050 602.250 ;
        RECT 67.950 596.850 70.050 598.950 ;
        RECT 85.650 598.950 86.850 605.400 ;
        RECT 91.650 604.500 92.850 608.400 ;
        RECT 101.550 605.400 103.350 611.250 ;
        RECT 104.550 605.400 106.350 611.250 ;
        RECT 107.550 605.400 109.350 611.250 ;
        RECT 87.750 603.600 92.850 604.500 ;
        RECT 104.400 604.500 106.200 605.400 ;
        RECT 110.550 604.500 112.350 611.250 ;
        RECT 113.550 605.400 115.350 611.250 ;
        RECT 116.550 605.400 118.350 611.250 ;
        RECT 119.550 605.400 121.350 611.250 ;
        RECT 122.550 605.400 124.350 611.250 ;
        RECT 125.550 605.400 127.350 611.250 ;
        RECT 142.650 605.400 144.450 611.250 ;
        RECT 116.400 604.500 118.200 605.400 ;
        RECT 122.400 604.500 124.200 605.400 ;
        RECT 87.750 602.700 90.000 603.600 ;
        RECT 104.400 603.300 108.450 604.500 ;
        RECT 110.550 603.300 114.300 604.500 ;
        RECT 116.400 603.300 120.300 604.500 ;
        RECT 122.400 604.350 125.100 604.500 ;
        RECT 122.400 603.300 125.250 604.350 ;
        RECT 85.650 596.850 88.050 598.950 ;
        RECT 62.100 595.050 63.900 596.850 ;
        RECT 67.950 591.600 69.150 596.850 ;
        RECT 70.950 593.850 73.050 595.950 ;
        RECT 70.950 592.050 72.750 593.850 ;
        RECT 85.650 591.600 86.850 596.850 ;
        RECT 88.950 594.300 90.000 602.700 ;
        RECT 107.250 602.400 108.450 603.300 ;
        RECT 113.100 602.400 114.300 603.300 ;
        RECT 119.100 602.400 120.300 603.300 ;
        RECT 104.100 600.150 105.900 601.950 ;
        RECT 107.250 600.600 111.300 602.400 ;
        RECT 113.100 600.600 117.300 602.400 ;
        RECT 119.100 600.600 123.300 602.400 ;
        RECT 91.950 596.850 94.050 598.950 ;
        RECT 103.950 598.050 106.050 600.150 ;
        RECT 92.100 595.050 93.900 596.850 ;
        RECT 87.750 593.400 90.000 594.300 ;
        RECT 107.250 593.700 108.450 600.600 ;
        RECT 113.100 593.700 114.300 600.600 ;
        RECT 119.100 593.700 120.300 600.600 ;
        RECT 124.200 600.150 125.250 603.300 ;
        RECT 143.250 603.300 144.450 605.400 ;
        RECT 145.650 606.300 147.450 611.250 ;
        RECT 148.650 607.200 150.450 611.250 ;
        RECT 151.650 606.300 153.450 611.250 ;
        RECT 172.650 608.400 174.450 611.250 ;
        RECT 175.650 608.400 177.450 611.250 ;
        RECT 178.650 608.400 180.450 611.250 ;
        RECT 181.650 608.400 183.750 611.250 ;
        RECT 194.550 608.400 196.350 611.250 ;
        RECT 197.550 608.400 199.350 611.250 ;
        RECT 200.550 608.400 202.350 611.250 ;
        RECT 212.550 608.400 214.350 611.250 ;
        RECT 215.550 608.400 217.350 611.250 ;
        RECT 172.650 607.500 173.700 608.400 ;
        RECT 178.650 607.500 179.700 608.400 ;
        RECT 145.650 604.950 153.450 606.300 ;
        RECT 168.900 606.600 179.700 607.500 ;
        RECT 143.250 602.250 147.000 603.300 ;
        RECT 124.200 598.050 127.050 600.150 ;
        RECT 145.950 598.950 147.150 602.250 ;
        RECT 149.100 600.150 150.900 601.950 ;
        RECT 168.900 600.150 170.100 606.600 ;
        RECT 198.000 601.950 199.050 608.400 ;
        RECT 176.100 600.150 177.900 601.950 ;
        RECT 124.200 593.700 125.250 598.050 ;
        RECT 145.950 596.850 148.050 598.950 ;
        RECT 148.950 598.050 151.050 600.150 ;
        RECT 151.950 596.850 154.050 598.950 ;
        RECT 166.950 598.050 170.100 600.150 ;
        RECT 142.950 593.850 145.050 595.950 ;
        RECT 87.750 592.500 93.450 593.400 ;
        RECT 43.050 579.750 44.850 591.450 ;
        RECT 46.050 590.100 48.450 591.450 ;
        RECT 46.050 579.750 47.850 590.100 ;
        RECT 63.300 579.750 65.100 591.600 ;
        RECT 67.500 579.750 69.300 591.600 ;
        RECT 70.800 579.750 72.600 585.600 ;
        RECT 85.350 579.750 87.150 591.600 ;
        RECT 88.350 579.750 90.150 591.600 ;
        RECT 92.250 585.600 93.450 592.500 ;
        RECT 104.550 592.500 108.450 593.700 ;
        RECT 110.550 592.500 114.300 593.700 ;
        RECT 116.550 592.500 120.300 593.700 ;
        RECT 122.550 592.500 125.250 593.700 ;
        RECT 91.650 579.750 93.450 585.600 ;
        RECT 101.550 579.750 103.350 591.600 ;
        RECT 104.550 579.750 106.350 592.500 ;
        RECT 107.550 579.750 109.350 591.600 ;
        RECT 110.550 579.750 112.350 592.500 ;
        RECT 113.550 579.750 115.350 591.600 ;
        RECT 116.550 579.750 118.350 592.500 ;
        RECT 119.550 579.750 121.350 591.600 ;
        RECT 122.550 579.750 124.350 592.500 ;
        RECT 143.250 592.050 145.050 593.850 ;
        RECT 146.850 591.600 148.050 596.850 ;
        RECT 152.100 595.050 153.900 596.850 ;
        RECT 168.900 592.800 170.100 598.050 ;
        RECT 172.950 596.850 175.050 598.950 ;
        RECT 175.950 598.050 178.050 600.150 ;
        RECT 196.950 599.850 199.050 601.950 ;
        RECT 211.950 599.850 214.050 601.950 ;
        RECT 215.400 600.150 216.600 608.400 ;
        RECT 232.650 605.400 234.450 611.250 ;
        RECT 233.250 603.300 234.450 605.400 ;
        RECT 235.650 606.300 237.450 611.250 ;
        RECT 238.650 607.200 240.450 611.250 ;
        RECT 241.650 606.300 243.450 611.250 ;
        RECT 235.650 604.950 243.450 606.300 ;
        RECT 251.550 605.400 253.350 611.250 ;
        RECT 254.550 605.400 256.350 611.250 ;
        RECT 257.550 605.400 259.350 611.250 ;
        RECT 260.550 605.400 262.350 611.250 ;
        RECT 263.550 605.400 265.350 611.250 ;
        RECT 254.550 604.500 255.750 605.400 ;
        RECT 260.550 604.500 261.750 605.400 ;
        RECT 254.550 603.300 261.750 604.500 ;
        RECT 281.850 604.200 283.650 611.250 ;
        RECT 286.350 605.400 288.150 611.250 ;
        RECT 298.650 605.400 300.450 611.250 ;
        RECT 281.850 603.300 285.450 604.200 ;
        RECT 233.250 602.250 237.000 603.300 ;
        RECT 181.950 596.850 184.050 598.950 ;
        RECT 193.950 596.850 196.050 598.950 ;
        RECT 173.100 595.050 174.900 596.850 ;
        RECT 182.100 595.050 183.900 596.850 ;
        RECT 194.100 595.050 195.900 596.850 ;
        RECT 166.650 591.600 170.100 592.800 ;
        RECT 198.000 592.650 199.050 599.850 ;
        RECT 199.950 596.850 202.050 598.950 ;
        RECT 212.100 598.050 213.900 599.850 ;
        RECT 214.950 598.050 217.050 600.150 ;
        RECT 235.950 598.950 237.150 602.250 ;
        RECT 239.100 600.150 240.900 601.950 ;
        RECT 200.100 595.050 201.900 596.850 ;
        RECT 198.000 591.600 200.550 592.650 ;
        RECT 125.550 579.750 127.350 591.600 ;
        RECT 143.400 579.750 145.200 585.600 ;
        RECT 146.700 579.750 148.500 591.600 ;
        RECT 150.900 579.750 152.700 591.600 ;
        RECT 163.050 580.500 164.850 589.800 ;
        RECT 166.650 589.200 167.850 591.600 ;
        RECT 166.050 581.400 167.850 589.200 ;
        RECT 169.050 589.200 177.450 590.100 ;
        RECT 169.050 580.500 170.850 589.200 ;
        RECT 163.050 579.750 170.850 580.500 ;
        RECT 172.650 580.500 174.450 588.300 ;
        RECT 175.650 581.400 177.450 589.200 ;
        RECT 178.650 589.500 186.450 590.400 ;
        RECT 178.650 580.500 180.450 589.500 ;
        RECT 172.650 579.750 180.450 580.500 ;
        RECT 181.650 579.750 183.450 588.600 ;
        RECT 184.650 579.750 186.450 589.500 ;
        RECT 194.550 579.750 196.350 591.600 ;
        RECT 198.750 579.750 200.550 591.600 ;
        RECT 215.400 585.600 216.600 598.050 ;
        RECT 235.950 596.850 238.050 598.950 ;
        RECT 238.950 598.050 241.050 600.150 ;
        RECT 260.550 598.950 261.750 603.300 ;
        RECT 241.950 596.850 244.050 598.950 ;
        RECT 253.950 596.850 256.050 598.950 ;
        RECT 259.950 596.850 262.050 598.950 ;
        RECT 281.100 597.150 282.900 598.950 ;
        RECT 232.950 593.850 235.050 595.950 ;
        RECT 233.250 592.050 235.050 593.850 ;
        RECT 236.850 591.600 238.050 596.850 ;
        RECT 242.100 595.050 243.900 596.850 ;
        RECT 254.100 595.050 255.900 596.850 ;
        RECT 260.550 593.400 261.750 596.850 ;
        RECT 280.950 595.050 283.050 597.150 ;
        RECT 284.250 595.950 285.450 603.300 ;
        RECT 299.250 603.300 300.450 605.400 ;
        RECT 301.650 606.300 303.450 611.250 ;
        RECT 304.650 607.200 306.450 611.250 ;
        RECT 307.650 606.300 309.450 611.250 ;
        RECT 319.650 608.400 321.450 611.250 ;
        RECT 322.650 608.400 324.450 611.250 ;
        RECT 301.650 604.950 309.450 606.300 ;
        RECT 299.250 602.250 303.000 603.300 ;
        RECT 301.950 598.950 303.150 602.250 ;
        RECT 305.100 600.150 306.900 601.950 ;
        RECT 320.400 600.150 321.600 608.400 ;
        RECT 335.550 606.300 337.350 611.250 ;
        RECT 338.550 607.200 340.350 611.250 ;
        RECT 341.550 606.300 343.350 611.250 ;
        RECT 335.550 604.950 343.350 606.300 ;
        RECT 344.550 605.400 346.350 611.250 ;
        RECT 344.550 603.300 345.750 605.400 ;
        RECT 342.000 602.250 345.750 603.300 ;
        RECT 365.100 603.000 366.900 611.250 ;
        RECT 287.100 597.150 288.900 598.950 ;
        RECT 283.950 593.850 286.050 595.950 ;
        RECT 286.950 595.050 289.050 597.150 ;
        RECT 301.950 596.850 304.050 598.950 ;
        RECT 304.950 598.050 307.050 600.150 ;
        RECT 307.950 596.850 310.050 598.950 ;
        RECT 319.950 598.050 322.050 600.150 ;
        RECT 322.950 599.850 325.050 601.950 ;
        RECT 338.100 600.150 339.900 601.950 ;
        RECT 323.100 598.050 324.900 599.850 ;
        RECT 298.950 593.850 301.050 595.950 ;
        RECT 254.550 592.500 261.750 593.400 ;
        RECT 212.550 579.750 214.350 585.600 ;
        RECT 215.550 579.750 217.350 585.600 ;
        RECT 233.400 579.750 235.200 585.600 ;
        RECT 236.700 579.750 238.500 591.600 ;
        RECT 240.900 579.750 242.700 591.600 ;
        RECT 251.550 579.750 253.350 591.600 ;
        RECT 254.550 579.750 256.350 592.500 ;
        RECT 260.550 591.600 261.750 592.500 ;
        RECT 257.550 579.750 259.350 591.600 ;
        RECT 260.550 579.750 262.350 591.600 ;
        RECT 263.550 579.750 265.350 591.600 ;
        RECT 284.250 585.600 285.450 593.850 ;
        RECT 299.250 592.050 301.050 593.850 ;
        RECT 302.850 591.600 304.050 596.850 ;
        RECT 308.100 595.050 309.900 596.850 ;
        RECT 280.650 579.750 282.450 585.600 ;
        RECT 283.650 579.750 285.450 585.600 ;
        RECT 286.650 579.750 288.450 585.600 ;
        RECT 299.400 579.750 301.200 585.600 ;
        RECT 302.700 579.750 304.500 591.600 ;
        RECT 306.900 579.750 308.700 591.600 ;
        RECT 320.400 585.600 321.600 598.050 ;
        RECT 334.950 596.850 337.050 598.950 ;
        RECT 337.950 598.050 340.050 600.150 ;
        RECT 341.850 598.950 343.050 602.250 ;
        RECT 340.950 596.850 343.050 598.950 ;
        RECT 362.400 601.350 366.900 603.000 ;
        RECT 370.500 602.400 372.300 611.250 ;
        RECT 381.000 605.400 382.800 611.250 ;
        RECT 385.200 607.050 387.000 611.250 ;
        RECT 388.500 608.400 390.300 611.250 ;
        RECT 385.200 605.400 390.900 607.050 ;
        RECT 362.400 597.150 363.600 601.350 ;
        RECT 380.100 600.150 381.900 601.950 ;
        RECT 379.950 598.050 382.050 600.150 ;
        RECT 382.950 599.850 385.050 601.950 ;
        RECT 386.100 600.150 387.900 601.950 ;
        RECT 383.100 598.050 384.900 599.850 ;
        RECT 385.950 598.050 388.050 600.150 ;
        RECT 389.700 598.950 390.900 605.400 ;
        RECT 404.850 604.200 406.650 611.250 ;
        RECT 409.350 605.400 411.150 611.250 ;
        RECT 424.650 605.400 426.450 611.250 ;
        RECT 404.850 603.300 408.450 604.200 ;
        RECT 335.100 595.050 336.900 596.850 ;
        RECT 340.950 591.600 342.150 596.850 ;
        RECT 343.950 593.850 346.050 595.950 ;
        RECT 361.950 595.050 364.050 597.150 ;
        RECT 388.950 596.850 391.050 598.950 ;
        RECT 404.100 597.150 405.900 598.950 ;
        RECT 343.950 592.050 345.750 593.850 ;
        RECT 319.650 579.750 321.450 585.600 ;
        RECT 322.650 579.750 324.450 585.600 ;
        RECT 336.300 579.750 338.100 591.600 ;
        RECT 340.500 579.750 342.300 591.600 ;
        RECT 362.250 586.800 363.300 595.050 ;
        RECT 364.950 593.850 367.050 595.950 ;
        RECT 370.950 593.850 373.050 595.950 ;
        RECT 364.950 592.050 366.750 593.850 ;
        RECT 367.950 590.850 370.050 592.950 ;
        RECT 371.100 592.050 372.900 593.850 ;
        RECT 389.700 591.600 390.900 596.850 ;
        RECT 403.950 595.050 406.050 597.150 ;
        RECT 407.250 595.950 408.450 603.300 ;
        RECT 425.250 603.300 426.450 605.400 ;
        RECT 427.650 606.300 429.450 611.250 ;
        RECT 430.650 607.200 432.450 611.250 ;
        RECT 433.650 606.300 435.450 611.250 ;
        RECT 427.650 604.950 435.450 606.300 ;
        RECT 438.150 605.400 439.950 611.250 ;
        RECT 441.150 608.400 442.950 611.250 ;
        RECT 445.950 609.300 447.750 611.250 ;
        RECT 444.000 608.400 447.750 609.300 ;
        RECT 450.450 608.400 452.250 611.250 ;
        RECT 453.750 608.400 455.550 611.250 ;
        RECT 457.650 608.400 459.450 611.250 ;
        RECT 461.850 608.400 463.650 611.250 ;
        RECT 466.350 608.400 468.150 611.250 ;
        RECT 444.000 607.500 445.050 608.400 ;
        RECT 442.950 605.400 445.050 607.500 ;
        RECT 453.750 606.600 454.800 608.400 ;
        RECT 425.250 602.250 429.000 603.300 ;
        RECT 427.950 598.950 429.150 602.250 ;
        RECT 431.100 600.150 432.900 601.950 ;
        RECT 410.100 597.150 411.900 598.950 ;
        RECT 406.950 593.850 409.050 595.950 ;
        RECT 409.950 595.050 412.050 597.150 ;
        RECT 427.950 596.850 430.050 598.950 ;
        RECT 430.950 598.050 433.050 600.150 ;
        RECT 433.950 596.850 436.050 598.950 ;
        RECT 424.950 593.850 427.050 595.950 ;
        RECT 368.100 589.050 369.900 590.850 ;
        RECT 380.550 590.700 388.350 591.600 ;
        RECT 362.250 585.900 369.300 586.800 ;
        RECT 362.250 585.600 363.450 585.900 ;
        RECT 343.800 579.750 345.600 585.600 ;
        RECT 361.650 579.750 363.450 585.600 ;
        RECT 367.650 585.600 369.300 585.900 ;
        RECT 364.650 579.750 366.450 585.000 ;
        RECT 367.650 579.750 369.450 585.600 ;
        RECT 370.650 579.750 372.450 585.600 ;
        RECT 380.550 579.750 382.350 590.700 ;
        RECT 383.550 579.750 385.350 589.800 ;
        RECT 386.550 579.750 388.350 590.700 ;
        RECT 389.550 579.750 391.350 591.600 ;
        RECT 407.250 585.600 408.450 593.850 ;
        RECT 425.250 592.050 427.050 593.850 ;
        RECT 428.850 591.600 430.050 596.850 ;
        RECT 434.100 595.050 435.900 596.850 ;
        RECT 438.150 592.800 439.050 605.400 ;
        RECT 446.550 604.800 448.350 606.600 ;
        RECT 449.850 605.550 454.800 606.600 ;
        RECT 462.300 607.500 463.350 608.400 ;
        RECT 462.300 606.300 466.050 607.500 ;
        RECT 449.850 604.800 451.650 605.550 ;
        RECT 446.850 603.900 447.900 604.800 ;
        RECT 457.050 604.200 458.850 606.000 ;
        RECT 463.950 605.400 466.050 606.300 ;
        RECT 469.650 605.400 471.450 611.250 ;
        RECT 482.550 608.400 484.350 611.250 ;
        RECT 485.550 608.400 487.350 611.250 ;
        RECT 488.550 608.400 490.350 611.250 ;
        RECT 457.050 603.900 457.950 604.200 ;
        RECT 446.850 603.000 457.950 603.900 ;
        RECT 470.250 603.150 471.450 605.400 ;
        RECT 446.850 601.800 447.900 603.000 ;
        RECT 441.000 600.600 447.900 601.800 ;
        RECT 441.000 599.850 441.900 600.600 ;
        RECT 446.100 600.000 447.900 600.600 ;
        RECT 440.100 598.050 441.900 599.850 ;
        RECT 443.100 598.950 444.900 599.700 ;
        RECT 457.050 598.950 457.950 603.000 ;
        RECT 466.950 601.050 471.450 603.150 ;
        RECT 486.000 601.950 487.050 608.400 ;
        RECT 500.850 605.400 502.650 611.250 ;
        RECT 505.350 604.200 507.150 611.250 ;
        RECT 521.550 608.400 523.350 611.250 ;
        RECT 524.550 608.400 526.350 611.250 ;
        RECT 527.550 608.400 529.350 611.250 ;
        RECT 542.550 608.400 544.350 611.250 ;
        RECT 545.550 608.400 547.350 611.250 ;
        RECT 548.550 608.400 550.350 611.250 ;
        RECT 465.150 599.250 469.050 601.050 ;
        RECT 466.950 598.950 469.050 599.250 ;
        RECT 443.100 597.900 451.050 598.950 ;
        RECT 448.950 596.850 451.050 597.900 ;
        RECT 454.950 596.850 457.950 598.950 ;
        RECT 447.450 593.100 449.250 593.400 ;
        RECT 447.450 592.800 455.850 593.100 ;
        RECT 438.150 592.200 455.850 592.800 ;
        RECT 438.150 591.600 449.250 592.200 ;
        RECT 403.650 579.750 405.450 585.600 ;
        RECT 406.650 579.750 408.450 585.600 ;
        RECT 409.650 579.750 411.450 585.600 ;
        RECT 425.400 579.750 427.200 585.600 ;
        RECT 428.700 579.750 430.500 591.600 ;
        RECT 432.900 579.750 434.700 591.600 ;
        RECT 438.150 579.750 439.950 591.600 ;
        RECT 452.250 590.700 454.050 591.300 ;
        RECT 446.550 589.500 454.050 590.700 ;
        RECT 454.950 590.100 455.850 592.200 ;
        RECT 457.050 592.200 457.950 596.850 ;
        RECT 467.250 593.400 469.050 595.200 ;
        RECT 463.950 592.200 468.150 593.400 ;
        RECT 457.050 591.300 463.050 592.200 ;
        RECT 463.950 591.300 466.050 592.200 ;
        RECT 470.250 591.600 471.450 601.050 ;
        RECT 484.950 599.850 487.050 601.950 ;
        RECT 481.950 596.850 484.050 598.950 ;
        RECT 482.100 595.050 483.900 596.850 ;
        RECT 486.000 592.650 487.050 599.850 ;
        RECT 503.550 603.300 507.150 604.200 ;
        RECT 487.950 596.850 490.050 598.950 ;
        RECT 500.100 597.150 501.900 598.950 ;
        RECT 488.100 595.050 489.900 596.850 ;
        RECT 499.950 595.050 502.050 597.150 ;
        RECT 503.550 595.950 504.750 603.300 ;
        RECT 525.000 601.950 526.050 608.400 ;
        RECT 546.000 601.950 547.050 608.400 ;
        RECT 560.550 603.900 562.350 611.250 ;
        RECT 565.050 605.400 566.850 611.250 ;
        RECT 568.050 606.900 569.850 611.250 ;
        RECT 568.050 605.400 571.350 606.900 ;
        RECT 583.650 605.400 585.450 611.250 ;
        RECT 566.250 603.900 568.050 604.500 ;
        RECT 560.550 602.700 568.050 603.900 ;
        RECT 523.950 599.850 526.050 601.950 ;
        RECT 544.950 599.850 547.050 601.950 ;
        RECT 506.100 597.150 507.900 598.950 ;
        RECT 502.950 593.850 505.050 595.950 ;
        RECT 505.950 595.050 508.050 597.150 ;
        RECT 520.950 596.850 523.050 598.950 ;
        RECT 521.100 595.050 522.900 596.850 ;
        RECT 486.000 591.600 488.550 592.650 ;
        RECT 462.150 590.400 463.050 591.300 ;
        RECT 459.450 590.100 461.250 590.400 ;
        RECT 446.550 588.600 447.750 589.500 ;
        RECT 454.950 589.200 461.250 590.100 ;
        RECT 459.450 588.600 461.250 589.200 ;
        RECT 462.150 588.600 464.850 590.400 ;
        RECT 442.950 586.500 447.750 588.600 ;
        RECT 450.150 586.500 457.050 588.300 ;
        RECT 446.550 585.600 447.750 586.500 ;
        RECT 441.150 579.750 442.950 585.600 ;
        RECT 446.250 579.750 448.050 585.600 ;
        RECT 451.050 579.750 452.850 585.600 ;
        RECT 454.050 579.750 455.850 586.500 ;
        RECT 462.150 585.600 466.050 587.700 ;
        RECT 457.950 579.750 459.750 585.600 ;
        RECT 462.150 579.750 463.950 585.600 ;
        RECT 466.650 579.750 468.450 582.600 ;
        RECT 469.650 579.750 471.450 591.600 ;
        RECT 482.550 579.750 484.350 591.600 ;
        RECT 486.750 579.750 488.550 591.600 ;
        RECT 503.550 585.600 504.750 593.850 ;
        RECT 525.000 592.650 526.050 599.850 ;
        RECT 526.950 596.850 529.050 598.950 ;
        RECT 541.950 596.850 544.050 598.950 ;
        RECT 527.100 595.050 528.900 596.850 ;
        RECT 542.100 595.050 543.900 596.850 ;
        RECT 546.000 592.650 547.050 599.850 ;
        RECT 547.950 596.850 550.050 598.950 ;
        RECT 559.950 596.850 562.050 598.950 ;
        RECT 548.100 595.050 549.900 596.850 ;
        RECT 560.100 595.050 561.900 596.850 ;
        RECT 525.000 591.600 527.550 592.650 ;
        RECT 546.000 591.600 548.550 592.650 ;
        RECT 500.550 579.750 502.350 585.600 ;
        RECT 503.550 579.750 505.350 585.600 ;
        RECT 506.550 579.750 508.350 585.600 ;
        RECT 521.550 579.750 523.350 591.600 ;
        RECT 525.750 579.750 527.550 591.600 ;
        RECT 542.550 579.750 544.350 591.600 ;
        RECT 546.750 579.750 548.550 591.600 ;
        RECT 563.700 585.600 564.900 602.700 ;
        RECT 570.150 598.950 571.350 605.400 ;
        RECT 584.250 603.300 585.450 605.400 ;
        RECT 586.650 606.300 588.450 611.250 ;
        RECT 589.650 607.200 591.450 611.250 ;
        RECT 592.650 606.300 594.450 611.250 ;
        RECT 586.650 604.950 594.450 606.300 ;
        RECT 605.550 606.300 607.350 611.250 ;
        RECT 608.550 607.200 610.350 611.250 ;
        RECT 611.550 606.300 613.350 611.250 ;
        RECT 605.550 604.950 613.350 606.300 ;
        RECT 614.550 605.400 616.350 611.250 ;
        RECT 632.700 608.400 634.500 611.250 ;
        RECT 636.000 607.050 637.800 611.250 ;
        RECT 632.100 605.400 637.800 607.050 ;
        RECT 640.200 605.400 642.000 611.250 ;
        RECT 614.550 603.300 615.750 605.400 ;
        RECT 584.250 602.250 588.000 603.300 ;
        RECT 612.000 602.250 615.750 603.300 ;
        RECT 566.100 597.150 567.900 598.950 ;
        RECT 565.950 595.050 568.050 597.150 ;
        RECT 568.950 596.850 571.350 598.950 ;
        RECT 586.950 598.950 588.150 602.250 ;
        RECT 590.100 600.150 591.900 601.950 ;
        RECT 608.100 600.150 609.900 601.950 ;
        RECT 586.950 596.850 589.050 598.950 ;
        RECT 589.950 598.050 592.050 600.150 ;
        RECT 592.950 596.850 595.050 598.950 ;
        RECT 604.950 596.850 607.050 598.950 ;
        RECT 607.950 598.050 610.050 600.150 ;
        RECT 611.850 598.950 613.050 602.250 ;
        RECT 632.100 598.950 633.300 605.400 ;
        RECT 650.700 602.400 652.500 611.250 ;
        RECT 656.100 603.000 657.900 611.250 ;
        RECT 671.550 608.400 673.350 611.250 ;
        RECT 674.550 608.400 676.350 611.250 ;
        RECT 635.100 600.150 636.900 601.950 ;
        RECT 610.950 596.850 613.050 598.950 ;
        RECT 631.950 596.850 634.050 598.950 ;
        RECT 634.950 598.050 637.050 600.150 ;
        RECT 637.950 599.850 640.050 601.950 ;
        RECT 641.100 600.150 642.900 601.950 ;
        RECT 656.100 601.350 660.600 603.000 ;
        RECT 638.100 598.050 639.900 599.850 ;
        RECT 640.950 598.050 643.050 600.150 ;
        RECT 659.400 597.150 660.600 601.350 ;
        RECT 670.950 599.850 673.050 601.950 ;
        RECT 674.400 600.150 675.600 608.400 ;
        RECT 681.150 605.400 682.950 611.250 ;
        RECT 684.150 608.400 685.950 611.250 ;
        RECT 688.950 609.300 690.750 611.250 ;
        RECT 687.000 608.400 690.750 609.300 ;
        RECT 693.450 608.400 695.250 611.250 ;
        RECT 696.750 608.400 698.550 611.250 ;
        RECT 700.650 608.400 702.450 611.250 ;
        RECT 704.850 608.400 706.650 611.250 ;
        RECT 709.350 608.400 711.150 611.250 ;
        RECT 687.000 607.500 688.050 608.400 ;
        RECT 685.950 605.400 688.050 607.500 ;
        RECT 696.750 606.600 697.800 608.400 ;
        RECT 671.100 598.050 672.900 599.850 ;
        RECT 673.950 598.050 676.050 600.150 ;
        RECT 570.150 591.600 571.350 596.850 ;
        RECT 583.950 593.850 586.050 595.950 ;
        RECT 584.250 592.050 586.050 593.850 ;
        RECT 587.850 591.600 589.050 596.850 ;
        RECT 593.100 595.050 594.900 596.850 ;
        RECT 605.100 595.050 606.900 596.850 ;
        RECT 610.950 591.600 612.150 596.850 ;
        RECT 613.950 593.850 616.050 595.950 ;
        RECT 613.950 592.050 615.750 593.850 ;
        RECT 632.100 591.600 633.300 596.850 ;
        RECT 649.950 593.850 652.050 595.950 ;
        RECT 655.950 593.850 658.050 595.950 ;
        RECT 658.950 595.050 661.050 597.150 ;
        RECT 650.100 592.050 651.900 593.850 ;
        RECT 560.550 579.750 562.350 585.600 ;
        RECT 563.550 579.750 565.350 585.600 ;
        RECT 567.150 579.750 568.950 591.600 ;
        RECT 570.150 579.750 571.950 591.600 ;
        RECT 584.400 579.750 586.200 585.600 ;
        RECT 587.700 579.750 589.500 591.600 ;
        RECT 591.900 579.750 593.700 591.600 ;
        RECT 606.300 579.750 608.100 591.600 ;
        RECT 610.500 579.750 612.300 591.600 ;
        RECT 613.800 579.750 615.600 585.600 ;
        RECT 631.650 579.750 633.450 591.600 ;
        RECT 634.650 590.700 642.450 591.600 ;
        RECT 652.950 590.850 655.050 592.950 ;
        RECT 656.250 592.050 658.050 593.850 ;
        RECT 634.650 579.750 636.450 590.700 ;
        RECT 637.650 579.750 639.450 589.800 ;
        RECT 640.650 579.750 642.450 590.700 ;
        RECT 653.100 589.050 654.900 590.850 ;
        RECT 659.700 586.800 660.750 595.050 ;
        RECT 653.700 585.900 660.750 586.800 ;
        RECT 653.700 585.600 655.350 585.900 ;
        RECT 650.550 579.750 652.350 585.600 ;
        RECT 653.550 579.750 655.350 585.600 ;
        RECT 659.550 585.600 660.750 585.900 ;
        RECT 674.400 585.600 675.600 598.050 ;
        RECT 681.150 592.800 682.050 605.400 ;
        RECT 689.550 604.800 691.350 606.600 ;
        RECT 692.850 605.550 697.800 606.600 ;
        RECT 705.300 607.500 706.350 608.400 ;
        RECT 705.300 606.300 709.050 607.500 ;
        RECT 692.850 604.800 694.650 605.550 ;
        RECT 689.850 603.900 690.900 604.800 ;
        RECT 700.050 604.200 701.850 606.000 ;
        RECT 706.950 605.400 709.050 606.300 ;
        RECT 712.650 605.400 714.450 611.250 ;
        RECT 725.550 608.400 727.350 611.250 ;
        RECT 728.550 608.400 730.350 611.250 ;
        RECT 740.550 608.400 742.350 611.250 ;
        RECT 743.550 608.400 745.350 611.250 ;
        RECT 746.550 608.400 748.350 611.250 ;
        RECT 758.550 608.400 760.350 611.250 ;
        RECT 761.550 608.400 763.350 611.250 ;
        RECT 700.050 603.900 700.950 604.200 ;
        RECT 689.850 603.000 700.950 603.900 ;
        RECT 713.250 603.150 714.450 605.400 ;
        RECT 689.850 601.800 690.900 603.000 ;
        RECT 684.000 600.600 690.900 601.800 ;
        RECT 684.000 599.850 684.900 600.600 ;
        RECT 689.100 600.000 690.900 600.600 ;
        RECT 683.100 598.050 684.900 599.850 ;
        RECT 686.100 598.950 687.900 599.700 ;
        RECT 700.050 598.950 700.950 603.000 ;
        RECT 709.950 601.050 714.450 603.150 ;
        RECT 708.150 599.250 712.050 601.050 ;
        RECT 709.950 598.950 712.050 599.250 ;
        RECT 686.100 597.900 694.050 598.950 ;
        RECT 691.950 596.850 694.050 597.900 ;
        RECT 697.950 596.850 700.950 598.950 ;
        RECT 690.450 593.100 692.250 593.400 ;
        RECT 690.450 592.800 698.850 593.100 ;
        RECT 681.150 592.200 698.850 592.800 ;
        RECT 681.150 591.600 692.250 592.200 ;
        RECT 656.550 579.750 658.350 585.000 ;
        RECT 659.550 579.750 661.350 585.600 ;
        RECT 671.550 579.750 673.350 585.600 ;
        RECT 674.550 579.750 676.350 585.600 ;
        RECT 681.150 579.750 682.950 591.600 ;
        RECT 695.250 590.700 697.050 591.300 ;
        RECT 689.550 589.500 697.050 590.700 ;
        RECT 697.950 590.100 698.850 592.200 ;
        RECT 700.050 592.200 700.950 596.850 ;
        RECT 710.250 593.400 712.050 595.200 ;
        RECT 706.950 592.200 711.150 593.400 ;
        RECT 700.050 591.300 706.050 592.200 ;
        RECT 706.950 591.300 709.050 592.200 ;
        RECT 713.250 591.600 714.450 601.050 ;
        RECT 724.950 599.850 727.050 601.950 ;
        RECT 728.400 600.150 729.600 608.400 ;
        RECT 744.000 601.950 745.050 608.400 ;
        RECT 725.100 598.050 726.900 599.850 ;
        RECT 727.950 598.050 730.050 600.150 ;
        RECT 742.950 599.850 745.050 601.950 ;
        RECT 757.950 599.850 760.050 601.950 ;
        RECT 761.400 600.150 762.600 608.400 ;
        RECT 776.850 604.200 778.650 611.250 ;
        RECT 781.350 605.400 783.150 611.250 ;
        RECT 794.850 604.200 796.650 611.250 ;
        RECT 799.350 605.400 801.150 611.250 ;
        RECT 803.550 605.400 805.350 611.250 ;
        RECT 806.850 608.400 808.650 611.250 ;
        RECT 811.350 608.400 813.150 611.250 ;
        RECT 815.550 608.400 817.350 611.250 ;
        RECT 819.450 608.400 821.250 611.250 ;
        RECT 822.750 608.400 824.550 611.250 ;
        RECT 827.250 609.300 829.050 611.250 ;
        RECT 827.250 608.400 831.000 609.300 ;
        RECT 832.050 608.400 833.850 611.250 ;
        RECT 811.650 607.500 812.700 608.400 ;
        RECT 808.950 606.300 812.700 607.500 ;
        RECT 820.200 606.600 821.250 608.400 ;
        RECT 829.950 607.500 831.000 608.400 ;
        RECT 808.950 605.400 811.050 606.300 ;
        RECT 776.850 603.300 780.450 604.200 ;
        RECT 794.850 603.300 798.450 604.200 ;
        RECT 705.150 590.400 706.050 591.300 ;
        RECT 702.450 590.100 704.250 590.400 ;
        RECT 689.550 588.600 690.750 589.500 ;
        RECT 697.950 589.200 704.250 590.100 ;
        RECT 702.450 588.600 704.250 589.200 ;
        RECT 705.150 588.600 707.850 590.400 ;
        RECT 685.950 586.500 690.750 588.600 ;
        RECT 693.150 586.500 700.050 588.300 ;
        RECT 689.550 585.600 690.750 586.500 ;
        RECT 684.150 579.750 685.950 585.600 ;
        RECT 689.250 579.750 691.050 585.600 ;
        RECT 694.050 579.750 695.850 585.600 ;
        RECT 697.050 579.750 698.850 586.500 ;
        RECT 705.150 585.600 709.050 587.700 ;
        RECT 700.950 579.750 702.750 585.600 ;
        RECT 705.150 579.750 706.950 585.600 ;
        RECT 709.650 579.750 711.450 582.600 ;
        RECT 712.650 579.750 714.450 591.600 ;
        RECT 728.400 585.600 729.600 598.050 ;
        RECT 739.950 596.850 742.050 598.950 ;
        RECT 740.100 595.050 741.900 596.850 ;
        RECT 744.000 592.650 745.050 599.850 ;
        RECT 745.950 596.850 748.050 598.950 ;
        RECT 758.100 598.050 759.900 599.850 ;
        RECT 760.950 598.050 763.050 600.150 ;
        RECT 746.100 595.050 747.900 596.850 ;
        RECT 744.000 591.600 746.550 592.650 ;
        RECT 725.550 579.750 727.350 585.600 ;
        RECT 728.550 579.750 730.350 585.600 ;
        RECT 740.550 579.750 742.350 591.600 ;
        RECT 744.750 579.750 746.550 591.600 ;
        RECT 761.400 585.600 762.600 598.050 ;
        RECT 776.100 597.150 777.900 598.950 ;
        RECT 775.950 595.050 778.050 597.150 ;
        RECT 779.250 595.950 780.450 603.300 ;
        RECT 782.100 597.150 783.900 598.950 ;
        RECT 794.100 597.150 795.900 598.950 ;
        RECT 778.950 593.850 781.050 595.950 ;
        RECT 781.950 595.050 784.050 597.150 ;
        RECT 793.950 595.050 796.050 597.150 ;
        RECT 797.250 595.950 798.450 603.300 ;
        RECT 803.550 603.150 804.750 605.400 ;
        RECT 816.150 604.200 817.950 606.000 ;
        RECT 820.200 605.550 825.150 606.600 ;
        RECT 823.350 604.800 825.150 605.550 ;
        RECT 826.650 604.800 828.450 606.600 ;
        RECT 829.950 605.400 832.050 607.500 ;
        RECT 835.050 605.400 836.850 611.250 ;
        RECT 847.650 605.400 849.450 611.250 ;
        RECT 817.050 603.900 817.950 604.200 ;
        RECT 827.100 603.900 828.150 604.800 ;
        RECT 803.550 601.050 808.050 603.150 ;
        RECT 817.050 603.000 828.150 603.900 ;
        RECT 800.100 597.150 801.900 598.950 ;
        RECT 796.950 593.850 799.050 595.950 ;
        RECT 799.950 595.050 802.050 597.150 ;
        RECT 779.250 585.600 780.450 593.850 ;
        RECT 797.250 585.600 798.450 593.850 ;
        RECT 803.550 591.600 804.750 601.050 ;
        RECT 805.950 599.250 809.850 601.050 ;
        RECT 805.950 598.950 808.050 599.250 ;
        RECT 817.050 598.950 817.950 603.000 ;
        RECT 827.100 601.800 828.150 603.000 ;
        RECT 827.100 600.600 834.000 601.800 ;
        RECT 827.100 600.000 828.900 600.600 ;
        RECT 833.100 599.850 834.000 600.600 ;
        RECT 830.100 598.950 831.900 599.700 ;
        RECT 817.050 596.850 820.050 598.950 ;
        RECT 823.950 597.900 831.900 598.950 ;
        RECT 833.100 598.050 834.900 599.850 ;
        RECT 823.950 596.850 826.050 597.900 ;
        RECT 805.950 593.400 807.750 595.200 ;
        RECT 806.850 592.200 811.050 593.400 ;
        RECT 817.050 592.200 817.950 596.850 ;
        RECT 825.750 593.100 827.550 593.400 ;
        RECT 758.550 579.750 760.350 585.600 ;
        RECT 761.550 579.750 763.350 585.600 ;
        RECT 775.650 579.750 777.450 585.600 ;
        RECT 778.650 579.750 780.450 585.600 ;
        RECT 781.650 579.750 783.450 585.600 ;
        RECT 793.650 579.750 795.450 585.600 ;
        RECT 796.650 579.750 798.450 585.600 ;
        RECT 799.650 579.750 801.450 585.600 ;
        RECT 803.550 579.750 805.350 591.600 ;
        RECT 808.950 591.300 811.050 592.200 ;
        RECT 811.950 591.300 817.950 592.200 ;
        RECT 819.150 592.800 827.550 593.100 ;
        RECT 835.950 592.800 836.850 605.400 ;
        RECT 848.250 603.300 849.450 605.400 ;
        RECT 850.650 606.300 852.450 611.250 ;
        RECT 853.650 607.200 855.450 611.250 ;
        RECT 856.650 606.300 858.450 611.250 ;
        RECT 850.650 604.950 858.450 606.300 ;
        RECT 866.550 606.300 868.350 611.250 ;
        RECT 869.550 607.200 871.350 611.250 ;
        RECT 872.550 606.300 874.350 611.250 ;
        RECT 866.550 604.950 874.350 606.300 ;
        RECT 875.550 605.400 877.350 611.250 ;
        RECT 856.950 603.450 859.050 604.050 ;
        RECT 848.250 602.250 852.000 603.300 ;
        RECT 856.950 602.550 864.450 603.450 ;
        RECT 875.550 603.300 876.750 605.400 ;
        RECT 850.950 598.950 852.150 602.250 ;
        RECT 856.950 601.950 859.050 602.550 ;
        RECT 854.100 600.150 855.900 601.950 ;
        RECT 850.950 596.850 853.050 598.950 ;
        RECT 853.950 598.050 856.050 600.150 ;
        RECT 856.950 596.850 859.050 598.950 ;
        RECT 847.950 593.850 850.050 595.950 ;
        RECT 819.150 592.200 836.850 592.800 ;
        RECT 811.950 590.400 812.850 591.300 ;
        RECT 810.150 588.600 812.850 590.400 ;
        RECT 813.750 590.100 815.550 590.400 ;
        RECT 819.150 590.100 820.050 592.200 ;
        RECT 825.750 591.600 836.850 592.200 ;
        RECT 848.250 592.050 850.050 593.850 ;
        RECT 851.850 591.600 853.050 596.850 ;
        RECT 857.100 595.050 858.900 596.850 ;
        RECT 863.550 595.050 864.450 602.550 ;
        RECT 873.000 602.250 876.750 603.300 ;
        RECT 869.100 600.150 870.900 601.950 ;
        RECT 865.950 596.850 868.050 598.950 ;
        RECT 868.950 598.050 871.050 600.150 ;
        RECT 872.850 598.950 874.050 602.250 ;
        RECT 871.950 596.850 874.050 598.950 ;
        RECT 866.100 595.050 867.900 596.850 ;
        RECT 862.950 592.950 865.050 595.050 ;
        RECT 871.950 591.600 873.150 596.850 ;
        RECT 874.950 593.850 877.050 595.950 ;
        RECT 874.950 592.050 876.750 593.850 ;
        RECT 813.750 589.200 820.050 590.100 ;
        RECT 820.950 590.700 822.750 591.300 ;
        RECT 820.950 589.500 828.450 590.700 ;
        RECT 813.750 588.600 815.550 589.200 ;
        RECT 827.250 588.600 828.450 589.500 ;
        RECT 808.950 585.600 812.850 587.700 ;
        RECT 817.950 586.500 824.850 588.300 ;
        RECT 827.250 586.500 832.050 588.600 ;
        RECT 806.550 579.750 808.350 582.600 ;
        RECT 811.050 579.750 812.850 585.600 ;
        RECT 815.250 579.750 817.050 585.600 ;
        RECT 819.150 579.750 820.950 586.500 ;
        RECT 827.250 585.600 828.450 586.500 ;
        RECT 822.150 579.750 823.950 585.600 ;
        RECT 826.950 579.750 828.750 585.600 ;
        RECT 832.050 579.750 833.850 585.600 ;
        RECT 835.050 579.750 836.850 591.600 ;
        RECT 848.400 579.750 850.200 585.600 ;
        RECT 851.700 579.750 853.500 591.600 ;
        RECT 855.900 579.750 857.700 591.600 ;
        RECT 867.300 579.750 869.100 591.600 ;
        RECT 871.500 579.750 873.300 591.600 ;
        RECT 874.800 579.750 876.600 585.600 ;
        RECT 11.550 563.400 13.350 575.250 ;
        RECT 16.050 563.550 17.850 575.250 ;
        RECT 19.050 564.900 20.850 575.250 ;
        RECT 34.650 569.400 36.450 575.250 ;
        RECT 37.650 570.000 39.450 575.250 ;
        RECT 35.250 569.100 36.450 569.400 ;
        RECT 40.650 569.400 42.450 575.250 ;
        RECT 43.650 569.400 45.450 575.250 ;
        RECT 53.550 569.400 55.350 575.250 ;
        RECT 56.550 569.400 58.350 575.250 ;
        RECT 59.550 569.400 61.350 575.250 ;
        RECT 74.400 569.400 76.200 575.250 ;
        RECT 40.650 569.100 42.300 569.400 ;
        RECT 35.250 568.200 42.300 569.100 ;
        RECT 19.050 563.550 21.450 564.900 ;
        RECT 11.550 562.200 12.750 563.400 ;
        RECT 16.950 562.200 18.750 562.650 ;
        RECT 11.550 561.000 18.750 562.200 ;
        RECT 16.950 560.850 18.750 561.000 ;
        RECT 14.100 558.150 15.900 559.950 ;
        RECT 11.100 555.150 12.900 556.950 ;
        RECT 13.950 556.050 16.050 558.150 ;
        RECT 10.950 553.050 13.050 555.150 ;
        RECT 17.700 552.600 18.600 560.850 ;
        RECT 20.100 556.950 21.450 563.550 ;
        RECT 35.250 559.950 36.300 568.200 ;
        RECT 41.100 564.150 42.900 565.950 ;
        RECT 37.950 561.150 39.750 562.950 ;
        RECT 40.950 562.050 43.050 564.150 ;
        RECT 44.100 561.150 45.900 562.950 ;
        RECT 56.550 561.150 57.750 569.400 ;
        RECT 77.700 563.400 79.500 575.250 ;
        RECT 81.900 563.400 83.700 575.250 ;
        RECT 95.550 563.400 97.350 575.250 ;
        RECT 99.750 563.400 101.550 575.250 ;
        RECT 113.550 563.400 115.350 575.250 ;
        RECT 117.750 563.400 119.550 575.250 ;
        RECT 136.650 569.400 138.450 575.250 ;
        RECT 139.650 569.400 141.450 575.250 ;
        RECT 142.650 569.400 144.450 575.250 ;
        RECT 74.250 561.150 76.050 562.950 ;
        RECT 34.950 557.850 37.050 559.950 ;
        RECT 37.950 559.050 40.050 561.150 ;
        RECT 43.950 559.050 46.050 561.150 ;
        RECT 52.950 557.850 55.050 559.950 ;
        RECT 55.950 559.050 58.050 561.150 ;
        RECT 19.950 554.850 22.050 556.950 ;
        RECT 16.950 551.700 18.750 552.600 ;
        RECT 15.450 550.800 18.750 551.700 ;
        RECT 15.450 546.600 16.350 550.800 ;
        RECT 21.000 549.600 22.050 554.850 ;
        RECT 35.400 553.650 36.600 557.850 ;
        RECT 53.100 556.050 54.900 557.850 ;
        RECT 35.400 552.000 39.900 553.650 ;
        RECT 11.550 543.750 13.350 546.600 ;
        RECT 14.550 543.750 16.350 546.600 ;
        RECT 17.550 543.750 19.350 546.600 ;
        RECT 20.550 543.750 22.350 549.600 ;
        RECT 38.100 543.750 39.900 552.000 ;
        RECT 43.500 543.750 45.300 552.600 ;
        RECT 56.550 551.700 57.750 559.050 ;
        RECT 58.950 557.850 61.050 559.950 ;
        RECT 73.950 559.050 76.050 561.150 ;
        RECT 77.850 558.150 79.050 563.400 ;
        RECT 99.000 562.350 101.550 563.400 ;
        RECT 117.000 562.350 119.550 563.400 ;
        RECT 83.100 558.150 84.900 559.950 ;
        RECT 95.100 558.150 96.900 559.950 ;
        RECT 59.100 556.050 60.900 557.850 ;
        RECT 76.950 556.050 79.050 558.150 ;
        RECT 76.950 552.750 78.150 556.050 ;
        RECT 79.950 554.850 82.050 556.950 ;
        RECT 82.950 556.050 85.050 558.150 ;
        RECT 94.950 556.050 97.050 558.150 ;
        RECT 99.000 555.150 100.050 562.350 ;
        RECT 101.100 558.150 102.900 559.950 ;
        RECT 113.100 558.150 114.900 559.950 ;
        RECT 100.950 556.050 103.050 558.150 ;
        RECT 112.950 556.050 115.050 558.150 ;
        RECT 117.000 555.150 118.050 562.350 ;
        RECT 140.250 561.150 141.450 569.400 ;
        RECT 154.350 563.400 156.150 575.250 ;
        RECT 157.350 563.400 159.150 575.250 ;
        RECT 160.650 569.400 162.450 575.250 ;
        RECT 119.100 558.150 120.900 559.950 ;
        RECT 118.950 556.050 121.050 558.150 ;
        RECT 136.950 557.850 139.050 559.950 ;
        RECT 139.950 559.050 142.050 561.150 ;
        RECT 137.100 556.050 138.900 557.850 ;
        RECT 80.100 553.050 81.900 554.850 ;
        RECT 97.950 553.050 100.050 555.150 ;
        RECT 115.950 553.050 118.050 555.150 ;
        RECT 74.250 551.700 78.000 552.750 ;
        RECT 56.550 550.800 60.150 551.700 ;
        RECT 53.850 543.750 55.650 549.600 ;
        RECT 58.350 543.750 60.150 550.800 ;
        RECT 74.250 549.600 75.450 551.700 ;
        RECT 73.650 543.750 75.450 549.600 ;
        RECT 76.650 548.700 84.450 550.050 ;
        RECT 76.650 543.750 78.450 548.700 ;
        RECT 79.650 543.750 81.450 547.800 ;
        RECT 82.650 543.750 84.450 548.700 ;
        RECT 99.000 546.600 100.050 553.050 ;
        RECT 117.000 546.600 118.050 553.050 ;
        RECT 140.250 551.700 141.450 559.050 ;
        RECT 142.950 557.850 145.050 559.950 ;
        RECT 154.650 558.150 155.850 563.400 ;
        RECT 161.250 562.500 162.450 569.400 ;
        RECT 156.750 561.600 162.450 562.500 ;
        RECT 164.550 563.400 166.350 575.250 ;
        RECT 167.550 572.400 169.350 575.250 ;
        RECT 172.050 569.400 173.850 575.250 ;
        RECT 176.250 569.400 178.050 575.250 ;
        RECT 169.950 567.300 173.850 569.400 ;
        RECT 180.150 568.500 181.950 575.250 ;
        RECT 183.150 569.400 184.950 575.250 ;
        RECT 187.950 569.400 189.750 575.250 ;
        RECT 193.050 569.400 194.850 575.250 ;
        RECT 188.250 568.500 189.450 569.400 ;
        RECT 178.950 566.700 185.850 568.500 ;
        RECT 188.250 566.400 193.050 568.500 ;
        RECT 171.150 564.600 173.850 566.400 ;
        RECT 174.750 565.800 176.550 566.400 ;
        RECT 174.750 564.900 181.050 565.800 ;
        RECT 188.250 565.500 189.450 566.400 ;
        RECT 174.750 564.600 176.550 564.900 ;
        RECT 172.950 563.700 173.850 564.600 ;
        RECT 156.750 560.700 159.000 561.600 ;
        RECT 143.100 556.050 144.900 557.850 ;
        RECT 154.650 556.050 157.050 558.150 ;
        RECT 137.850 550.800 141.450 551.700 ;
        RECT 95.550 543.750 97.350 546.600 ;
        RECT 98.550 543.750 100.350 546.600 ;
        RECT 101.550 543.750 103.350 546.600 ;
        RECT 113.550 543.750 115.350 546.600 ;
        RECT 116.550 543.750 118.350 546.600 ;
        RECT 119.550 543.750 121.350 546.600 ;
        RECT 137.850 543.750 139.650 550.800 ;
        RECT 154.650 549.600 155.850 556.050 ;
        RECT 157.950 552.300 159.000 560.700 ;
        RECT 161.100 558.150 162.900 559.950 ;
        RECT 160.950 556.050 163.050 558.150 ;
        RECT 156.750 551.400 159.000 552.300 ;
        RECT 164.550 553.950 165.750 563.400 ;
        RECT 169.950 562.800 172.050 563.700 ;
        RECT 172.950 562.800 178.950 563.700 ;
        RECT 167.850 561.600 172.050 562.800 ;
        RECT 166.950 559.800 168.750 561.600 ;
        RECT 178.050 558.150 178.950 562.800 ;
        RECT 180.150 562.800 181.050 564.900 ;
        RECT 181.950 564.300 189.450 565.500 ;
        RECT 181.950 563.700 183.750 564.300 ;
        RECT 196.050 563.400 197.850 575.250 ;
        RECT 208.650 569.400 210.450 575.250 ;
        RECT 211.650 569.400 213.450 575.250 ;
        RECT 214.650 569.400 216.450 575.250 ;
        RECT 227.400 569.400 229.200 575.250 ;
        RECT 186.750 562.800 197.850 563.400 ;
        RECT 180.150 562.200 197.850 562.800 ;
        RECT 180.150 561.900 188.550 562.200 ;
        RECT 186.750 561.600 188.550 561.900 ;
        RECT 178.050 556.050 181.050 558.150 ;
        RECT 184.950 557.100 187.050 558.150 ;
        RECT 184.950 556.050 192.900 557.100 ;
        RECT 166.950 555.750 169.050 556.050 ;
        RECT 166.950 553.950 170.850 555.750 ;
        RECT 164.550 551.850 169.050 553.950 ;
        RECT 178.050 552.000 178.950 556.050 ;
        RECT 191.100 555.300 192.900 556.050 ;
        RECT 194.100 555.150 195.900 556.950 ;
        RECT 188.100 554.400 189.900 555.000 ;
        RECT 194.100 554.400 195.000 555.150 ;
        RECT 188.100 553.200 195.000 554.400 ;
        RECT 188.100 552.000 189.150 553.200 ;
        RECT 156.750 550.500 161.850 551.400 ;
        RECT 142.350 543.750 144.150 549.600 ;
        RECT 154.350 543.750 156.150 549.600 ;
        RECT 157.350 543.750 159.150 549.600 ;
        RECT 160.650 546.600 161.850 550.500 ;
        RECT 164.550 549.600 165.750 551.850 ;
        RECT 178.050 551.100 189.150 552.000 ;
        RECT 178.050 550.800 178.950 551.100 ;
        RECT 160.650 543.750 162.450 546.600 ;
        RECT 164.550 543.750 166.350 549.600 ;
        RECT 169.950 548.700 172.050 549.600 ;
        RECT 177.150 549.000 178.950 550.800 ;
        RECT 188.100 550.200 189.150 551.100 ;
        RECT 184.350 549.450 186.150 550.200 ;
        RECT 169.950 547.500 173.700 548.700 ;
        RECT 172.650 546.600 173.700 547.500 ;
        RECT 181.200 548.400 186.150 549.450 ;
        RECT 187.650 548.400 189.450 550.200 ;
        RECT 196.950 549.600 197.850 562.200 ;
        RECT 212.250 561.150 213.450 569.400 ;
        RECT 230.700 563.400 232.500 575.250 ;
        RECT 234.900 563.400 236.700 575.250 ;
        RECT 245.550 564.300 247.350 575.250 ;
        RECT 248.550 565.200 250.350 575.250 ;
        RECT 251.550 564.300 253.350 575.250 ;
        RECT 245.550 563.400 253.350 564.300 ;
        RECT 254.550 563.400 256.350 575.250 ;
        RECT 266.550 569.400 268.350 575.250 ;
        RECT 269.550 569.400 271.350 575.250 ;
        RECT 272.550 570.000 274.350 575.250 ;
        RECT 269.700 569.100 271.350 569.400 ;
        RECT 275.550 569.400 277.350 575.250 ;
        RECT 287.550 569.400 289.350 575.250 ;
        RECT 290.550 569.400 292.350 575.250 ;
        RECT 293.550 570.000 295.350 575.250 ;
        RECT 275.550 569.100 276.750 569.400 ;
        RECT 269.700 568.200 276.750 569.100 ;
        RECT 290.700 569.100 292.350 569.400 ;
        RECT 296.550 569.400 298.350 575.250 ;
        RECT 308.550 569.400 310.350 575.250 ;
        RECT 311.550 569.400 313.350 575.250 ;
        RECT 314.550 569.400 316.350 575.250 ;
        RECT 332.400 569.400 334.200 575.250 ;
        RECT 296.550 569.100 297.750 569.400 ;
        RECT 290.700 568.200 297.750 569.100 ;
        RECT 269.100 564.150 270.900 565.950 ;
        RECT 227.250 561.150 229.050 562.950 ;
        RECT 208.950 557.850 211.050 559.950 ;
        RECT 211.950 559.050 214.050 561.150 ;
        RECT 209.100 556.050 210.900 557.850 ;
        RECT 212.250 551.700 213.450 559.050 ;
        RECT 214.950 557.850 217.050 559.950 ;
        RECT 226.950 559.050 229.050 561.150 ;
        RECT 230.850 558.150 232.050 563.400 ;
        RECT 236.100 558.150 237.900 559.950 ;
        RECT 254.700 558.150 255.900 563.400 ;
        RECT 266.100 561.150 267.900 562.950 ;
        RECT 268.950 562.050 271.050 564.150 ;
        RECT 272.250 561.150 274.050 562.950 ;
        RECT 265.950 559.050 268.050 561.150 ;
        RECT 271.950 559.050 274.050 561.150 ;
        RECT 275.700 559.950 276.750 568.200 ;
        RECT 290.100 564.150 291.900 565.950 ;
        RECT 287.100 561.150 288.900 562.950 ;
        RECT 289.950 562.050 292.050 564.150 ;
        RECT 293.250 561.150 295.050 562.950 ;
        RECT 215.100 556.050 216.900 557.850 ;
        RECT 229.950 556.050 232.050 558.150 ;
        RECT 229.950 552.750 231.150 556.050 ;
        RECT 232.950 554.850 235.050 556.950 ;
        RECT 235.950 556.050 238.050 558.150 ;
        RECT 244.950 554.850 247.050 556.950 ;
        RECT 248.100 555.150 249.900 556.950 ;
        RECT 233.100 553.050 234.900 554.850 ;
        RECT 245.100 553.050 246.900 554.850 ;
        RECT 247.950 553.050 250.050 555.150 ;
        RECT 250.950 554.850 253.050 556.950 ;
        RECT 253.950 556.050 256.050 558.150 ;
        RECT 274.950 557.850 277.050 559.950 ;
        RECT 286.950 559.050 289.050 561.150 ;
        RECT 292.950 559.050 295.050 561.150 ;
        RECT 296.700 559.950 297.750 568.200 ;
        RECT 311.550 561.150 312.750 569.400 ;
        RECT 335.700 563.400 337.500 575.250 ;
        RECT 339.900 563.400 341.700 575.250 ;
        RECT 352.650 569.400 354.450 575.250 ;
        RECT 355.650 569.400 357.450 575.250 ;
        RECT 370.650 569.400 372.450 575.250 ;
        RECT 373.650 570.000 375.450 575.250 ;
        RECT 332.250 561.150 334.050 562.950 ;
        RECT 295.950 557.850 298.050 559.950 ;
        RECT 307.950 557.850 310.050 559.950 ;
        RECT 310.950 559.050 313.050 561.150 ;
        RECT 251.100 553.050 252.900 554.850 ;
        RECT 181.200 546.600 182.250 548.400 ;
        RECT 190.950 547.500 193.050 549.600 ;
        RECT 190.950 546.600 192.000 547.500 ;
        RECT 167.850 543.750 169.650 546.600 ;
        RECT 172.350 543.750 174.150 546.600 ;
        RECT 176.550 543.750 178.350 546.600 ;
        RECT 180.450 543.750 182.250 546.600 ;
        RECT 183.750 543.750 185.550 546.600 ;
        RECT 188.250 545.700 192.000 546.600 ;
        RECT 188.250 543.750 190.050 545.700 ;
        RECT 193.050 543.750 194.850 546.600 ;
        RECT 196.050 543.750 197.850 549.600 ;
        RECT 209.850 550.800 213.450 551.700 ;
        RECT 227.250 551.700 231.000 552.750 ;
        RECT 209.850 543.750 211.650 550.800 ;
        RECT 227.250 549.600 228.450 551.700 ;
        RECT 214.350 543.750 216.150 549.600 ;
        RECT 226.650 543.750 228.450 549.600 ;
        RECT 229.650 548.700 237.450 550.050 ;
        RECT 254.700 549.600 255.900 556.050 ;
        RECT 275.400 553.650 276.600 557.850 ;
        RECT 296.400 553.650 297.600 557.850 ;
        RECT 308.100 556.050 309.900 557.850 ;
        RECT 229.650 543.750 231.450 548.700 ;
        RECT 232.650 543.750 234.450 547.800 ;
        RECT 235.650 543.750 237.450 548.700 ;
        RECT 246.000 543.750 247.800 549.600 ;
        RECT 250.200 547.950 255.900 549.600 ;
        RECT 250.200 543.750 252.000 547.950 ;
        RECT 253.500 543.750 255.300 546.600 ;
        RECT 266.700 543.750 268.500 552.600 ;
        RECT 272.100 552.000 276.600 553.650 ;
        RECT 272.100 543.750 273.900 552.000 ;
        RECT 287.700 543.750 289.500 552.600 ;
        RECT 293.100 552.000 297.600 553.650 ;
        RECT 293.100 543.750 294.900 552.000 ;
        RECT 311.550 551.700 312.750 559.050 ;
        RECT 313.950 557.850 316.050 559.950 ;
        RECT 331.950 559.050 334.050 561.150 ;
        RECT 335.850 558.150 337.050 563.400 ;
        RECT 341.100 558.150 342.900 559.950 ;
        RECT 314.100 556.050 315.900 557.850 ;
        RECT 334.950 556.050 337.050 558.150 ;
        RECT 334.950 552.750 336.150 556.050 ;
        RECT 337.950 554.850 340.050 556.950 ;
        RECT 340.950 556.050 343.050 558.150 ;
        RECT 353.400 556.950 354.600 569.400 ;
        RECT 371.250 569.100 372.450 569.400 ;
        RECT 376.650 569.400 378.450 575.250 ;
        RECT 379.650 569.400 381.450 575.250 ;
        RECT 391.650 569.400 393.450 575.250 ;
        RECT 394.650 570.000 396.450 575.250 ;
        RECT 376.650 569.100 378.300 569.400 ;
        RECT 371.250 568.200 378.300 569.100 ;
        RECT 392.250 569.100 393.450 569.400 ;
        RECT 397.650 569.400 399.450 575.250 ;
        RECT 400.650 569.400 402.450 575.250 ;
        RECT 410.550 569.400 412.350 575.250 ;
        RECT 413.550 569.400 415.350 575.250 ;
        RECT 416.550 569.400 418.350 575.250 ;
        RECT 428.550 569.400 430.350 575.250 ;
        RECT 431.550 569.400 433.350 575.250 ;
        RECT 434.550 569.400 436.350 575.250 ;
        RECT 397.650 569.100 399.300 569.400 ;
        RECT 392.250 568.200 399.300 569.100 ;
        RECT 371.250 559.950 372.300 568.200 ;
        RECT 377.100 564.150 378.900 565.950 ;
        RECT 373.950 561.150 375.750 562.950 ;
        RECT 376.950 562.050 379.050 564.150 ;
        RECT 380.100 561.150 381.900 562.950 ;
        RECT 370.950 557.850 373.050 559.950 ;
        RECT 373.950 559.050 376.050 561.150 ;
        RECT 379.950 559.050 382.050 561.150 ;
        RECT 392.250 559.950 393.300 568.200 ;
        RECT 398.100 564.150 399.900 565.950 ;
        RECT 394.950 561.150 396.750 562.950 ;
        RECT 397.950 562.050 400.050 564.150 ;
        RECT 401.100 561.150 402.900 562.950 ;
        RECT 413.550 561.150 414.750 569.400 ;
        RECT 431.550 561.150 432.750 569.400 ;
        RECT 451.350 563.400 453.150 575.250 ;
        RECT 454.350 563.400 456.150 575.250 ;
        RECT 457.650 569.400 459.450 575.250 ;
        RECT 391.950 557.850 394.050 559.950 ;
        RECT 394.950 559.050 397.050 561.150 ;
        RECT 400.950 559.050 403.050 561.150 ;
        RECT 409.950 557.850 412.050 559.950 ;
        RECT 412.950 559.050 415.050 561.150 ;
        RECT 352.950 554.850 355.050 556.950 ;
        RECT 356.100 555.150 357.900 556.950 ;
        RECT 338.100 553.050 339.900 554.850 ;
        RECT 332.250 551.700 336.000 552.750 ;
        RECT 343.950 552.450 346.050 553.050 ;
        RECT 349.950 552.450 352.050 553.050 ;
        RECT 311.550 550.800 315.150 551.700 ;
        RECT 308.850 543.750 310.650 549.600 ;
        RECT 313.350 543.750 315.150 550.800 ;
        RECT 332.250 549.600 333.450 551.700 ;
        RECT 343.950 551.550 352.050 552.450 ;
        RECT 343.950 550.950 346.050 551.550 ;
        RECT 349.950 550.950 352.050 551.550 ;
        RECT 331.650 543.750 333.450 549.600 ;
        RECT 334.650 548.700 342.450 550.050 ;
        RECT 334.650 543.750 336.450 548.700 ;
        RECT 337.650 543.750 339.450 547.800 ;
        RECT 340.650 543.750 342.450 548.700 ;
        RECT 353.400 546.600 354.600 554.850 ;
        RECT 355.950 553.050 358.050 555.150 ;
        RECT 371.400 553.650 372.600 557.850 ;
        RECT 392.400 553.650 393.600 557.850 ;
        RECT 410.100 556.050 411.900 557.850 ;
        RECT 400.950 555.450 403.050 556.050 ;
        RECT 406.950 555.450 409.050 556.050 ;
        RECT 400.950 554.550 409.050 555.450 ;
        RECT 400.950 553.950 403.050 554.550 ;
        RECT 406.950 553.950 409.050 554.550 ;
        RECT 371.400 552.000 375.900 553.650 ;
        RECT 352.650 543.750 354.450 546.600 ;
        RECT 355.650 543.750 357.450 546.600 ;
        RECT 374.100 543.750 375.900 552.000 ;
        RECT 379.500 543.750 381.300 552.600 ;
        RECT 392.400 552.000 396.900 553.650 ;
        RECT 395.100 543.750 396.900 552.000 ;
        RECT 400.500 543.750 402.300 552.600 ;
        RECT 413.550 551.700 414.750 559.050 ;
        RECT 415.950 557.850 418.050 559.950 ;
        RECT 427.950 557.850 430.050 559.950 ;
        RECT 430.950 559.050 433.050 561.150 ;
        RECT 416.100 556.050 417.900 557.850 ;
        RECT 428.100 556.050 429.900 557.850 ;
        RECT 431.550 551.700 432.750 559.050 ;
        RECT 433.950 557.850 436.050 559.950 ;
        RECT 451.650 558.150 452.850 563.400 ;
        RECT 458.250 562.500 459.450 569.400 ;
        RECT 453.750 561.600 459.450 562.500 ;
        RECT 467.550 569.400 469.350 575.250 ;
        RECT 467.550 562.500 468.750 569.400 ;
        RECT 470.850 563.400 472.650 575.250 ;
        RECT 473.850 563.400 475.650 575.250 ;
        RECT 485.550 569.400 487.350 575.250 ;
        RECT 467.550 561.600 473.250 562.500 ;
        RECT 453.750 560.700 456.000 561.600 ;
        RECT 434.100 556.050 435.900 557.850 ;
        RECT 451.650 556.050 454.050 558.150 ;
        RECT 413.550 550.800 417.150 551.700 ;
        RECT 431.550 550.800 435.150 551.700 ;
        RECT 410.850 543.750 412.650 549.600 ;
        RECT 415.350 543.750 417.150 550.800 ;
        RECT 428.850 543.750 430.650 549.600 ;
        RECT 433.350 543.750 435.150 550.800 ;
        RECT 451.650 549.600 452.850 556.050 ;
        RECT 454.950 552.300 456.000 560.700 ;
        RECT 471.000 560.700 473.250 561.600 ;
        RECT 458.100 558.150 459.900 559.950 ;
        RECT 467.100 558.150 468.900 559.950 ;
        RECT 457.950 556.050 460.050 558.150 ;
        RECT 466.950 556.050 469.050 558.150 ;
        RECT 453.750 551.400 456.000 552.300 ;
        RECT 471.000 552.300 472.050 560.700 ;
        RECT 474.150 558.150 475.350 563.400 ;
        RECT 485.550 562.500 486.750 569.400 ;
        RECT 488.850 563.400 490.650 575.250 ;
        RECT 491.850 563.400 493.650 575.250 ;
        RECT 503.550 569.400 505.350 575.250 ;
        RECT 485.550 561.600 491.250 562.500 ;
        RECT 489.000 560.700 491.250 561.600 ;
        RECT 485.100 558.150 486.900 559.950 ;
        RECT 472.950 556.050 475.350 558.150 ;
        RECT 484.950 556.050 487.050 558.150 ;
        RECT 471.000 551.400 473.250 552.300 ;
        RECT 453.750 550.500 458.850 551.400 ;
        RECT 451.350 543.750 453.150 549.600 ;
        RECT 454.350 543.750 456.150 549.600 ;
        RECT 457.650 546.600 458.850 550.500 ;
        RECT 468.150 550.500 473.250 551.400 ;
        RECT 468.150 546.600 469.350 550.500 ;
        RECT 474.150 549.600 475.350 556.050 ;
        RECT 489.000 552.300 490.050 560.700 ;
        RECT 492.150 558.150 493.350 563.400 ;
        RECT 503.550 562.500 504.750 569.400 ;
        RECT 506.850 563.400 508.650 575.250 ;
        RECT 509.850 563.400 511.650 575.250 ;
        RECT 525.300 563.400 527.100 575.250 ;
        RECT 529.500 563.400 531.300 575.250 ;
        RECT 532.800 569.400 534.600 575.250 ;
        RECT 547.650 563.400 549.450 575.250 ;
        RECT 550.650 564.300 552.450 575.250 ;
        RECT 553.650 565.200 555.450 575.250 ;
        RECT 556.650 564.300 558.450 575.250 ;
        RECT 566.550 569.400 568.350 575.250 ;
        RECT 569.550 569.400 571.350 575.250 ;
        RECT 572.550 570.000 574.350 575.250 ;
        RECT 569.700 569.100 571.350 569.400 ;
        RECT 575.550 569.400 577.350 575.250 ;
        RECT 575.550 569.100 576.750 569.400 ;
        RECT 569.700 568.200 576.750 569.100 ;
        RECT 550.650 563.400 558.450 564.300 ;
        RECT 569.100 564.150 570.900 565.950 ;
        RECT 503.550 561.600 509.250 562.500 ;
        RECT 507.000 560.700 509.250 561.600 ;
        RECT 503.100 558.150 504.900 559.950 ;
        RECT 490.950 556.050 493.350 558.150 ;
        RECT 502.950 556.050 505.050 558.150 ;
        RECT 489.000 551.400 491.250 552.300 ;
        RECT 486.150 550.500 491.250 551.400 ;
        RECT 457.650 543.750 459.450 546.600 ;
        RECT 467.550 543.750 469.350 546.600 ;
        RECT 470.850 543.750 472.650 549.600 ;
        RECT 473.850 543.750 475.650 549.600 ;
        RECT 486.150 546.600 487.350 550.500 ;
        RECT 492.150 549.600 493.350 556.050 ;
        RECT 507.000 552.300 508.050 560.700 ;
        RECT 510.150 558.150 511.350 563.400 ;
        RECT 524.100 558.150 525.900 559.950 ;
        RECT 529.950 558.150 531.150 563.400 ;
        RECT 532.950 561.150 534.750 562.950 ;
        RECT 532.950 559.050 535.050 561.150 ;
        RECT 548.100 558.150 549.300 563.400 ;
        RECT 566.100 561.150 567.900 562.950 ;
        RECT 568.950 562.050 571.050 564.150 ;
        RECT 572.250 561.150 574.050 562.950 ;
        RECT 565.950 559.050 568.050 561.150 ;
        RECT 571.950 559.050 574.050 561.150 ;
        RECT 575.700 559.950 576.750 568.200 ;
        RECT 587.550 563.400 589.350 575.250 ;
        RECT 592.050 563.550 593.850 575.250 ;
        RECT 595.050 564.900 596.850 575.250 ;
        RECT 595.050 563.550 597.450 564.900 ;
        RECT 587.550 562.200 588.750 563.400 ;
        RECT 592.950 562.200 594.750 562.650 ;
        RECT 587.550 561.000 594.750 562.200 ;
        RECT 592.950 560.850 594.750 561.000 ;
        RECT 508.950 556.050 511.350 558.150 ;
        RECT 523.950 556.050 526.050 558.150 ;
        RECT 507.000 551.400 509.250 552.300 ;
        RECT 504.150 550.500 509.250 551.400 ;
        RECT 485.550 543.750 487.350 546.600 ;
        RECT 488.850 543.750 490.650 549.600 ;
        RECT 491.850 543.750 493.650 549.600 ;
        RECT 504.150 546.600 505.350 550.500 ;
        RECT 510.150 549.600 511.350 556.050 ;
        RECT 526.950 554.850 529.050 556.950 ;
        RECT 529.950 556.050 532.050 558.150 ;
        RECT 547.950 556.050 550.050 558.150 ;
        RECT 574.950 557.850 577.050 559.950 ;
        RECT 590.100 558.150 591.900 559.950 ;
        RECT 527.100 553.050 528.900 554.850 ;
        RECT 530.850 552.750 532.050 556.050 ;
        RECT 531.000 551.700 534.750 552.750 ;
        RECT 503.550 543.750 505.350 546.600 ;
        RECT 506.850 543.750 508.650 549.600 ;
        RECT 509.850 543.750 511.650 549.600 ;
        RECT 524.550 548.700 532.350 550.050 ;
        RECT 524.550 543.750 526.350 548.700 ;
        RECT 527.550 543.750 529.350 547.800 ;
        RECT 530.550 543.750 532.350 548.700 ;
        RECT 533.550 549.600 534.750 551.700 ;
        RECT 548.100 549.600 549.300 556.050 ;
        RECT 550.950 554.850 553.050 556.950 ;
        RECT 554.100 555.150 555.900 556.950 ;
        RECT 551.100 553.050 552.900 554.850 ;
        RECT 553.950 553.050 556.050 555.150 ;
        RECT 556.950 554.850 559.050 556.950 ;
        RECT 557.100 553.050 558.900 554.850 ;
        RECT 575.400 553.650 576.600 557.850 ;
        RECT 587.100 555.150 588.900 556.950 ;
        RECT 589.950 556.050 592.050 558.150 ;
        RECT 533.550 543.750 535.350 549.600 ;
        RECT 548.100 547.950 553.800 549.600 ;
        RECT 548.700 543.750 550.500 546.600 ;
        RECT 552.000 543.750 553.800 547.950 ;
        RECT 556.200 543.750 558.000 549.600 ;
        RECT 566.700 543.750 568.500 552.600 ;
        RECT 572.100 552.000 576.600 553.650 ;
        RECT 586.950 553.050 589.050 555.150 ;
        RECT 593.700 552.600 594.600 560.850 ;
        RECT 596.100 556.950 597.450 563.550 ;
        RECT 609.300 563.400 611.100 575.250 ;
        RECT 613.500 563.400 615.300 575.250 ;
        RECT 616.800 569.400 618.600 575.250 ;
        RECT 632.550 569.400 634.350 575.250 ;
        RECT 635.550 569.400 637.350 575.250 ;
        RECT 638.550 570.000 640.350 575.250 ;
        RECT 635.700 569.100 637.350 569.400 ;
        RECT 641.550 569.400 643.350 575.250 ;
        RECT 641.550 569.100 642.750 569.400 ;
        RECT 635.700 568.200 642.750 569.100 ;
        RECT 635.100 564.150 636.900 565.950 ;
        RECT 608.100 558.150 609.900 559.950 ;
        RECT 613.950 558.150 615.150 563.400 ;
        RECT 616.950 561.150 618.750 562.950 ;
        RECT 632.100 561.150 633.900 562.950 ;
        RECT 634.950 562.050 637.050 564.150 ;
        RECT 638.250 561.150 640.050 562.950 ;
        RECT 616.950 559.050 619.050 561.150 ;
        RECT 631.950 559.050 634.050 561.150 ;
        RECT 637.950 559.050 640.050 561.150 ;
        RECT 641.700 559.950 642.750 568.200 ;
        RECT 653.550 564.300 655.350 575.250 ;
        RECT 656.550 565.200 658.350 575.250 ;
        RECT 659.550 564.300 661.350 575.250 ;
        RECT 653.550 563.400 661.350 564.300 ;
        RECT 662.550 563.400 664.350 575.250 ;
        RECT 668.550 563.400 670.350 575.250 ;
        RECT 671.550 572.400 673.350 575.250 ;
        RECT 676.050 569.400 677.850 575.250 ;
        RECT 680.250 569.400 682.050 575.250 ;
        RECT 673.950 567.300 677.850 569.400 ;
        RECT 684.150 568.500 685.950 575.250 ;
        RECT 687.150 569.400 688.950 575.250 ;
        RECT 691.950 569.400 693.750 575.250 ;
        RECT 697.050 569.400 698.850 575.250 ;
        RECT 692.250 568.500 693.450 569.400 ;
        RECT 682.950 566.700 689.850 568.500 ;
        RECT 692.250 566.400 697.050 568.500 ;
        RECT 675.150 564.600 677.850 566.400 ;
        RECT 678.750 565.800 680.550 566.400 ;
        RECT 678.750 564.900 685.050 565.800 ;
        RECT 692.250 565.500 693.450 566.400 ;
        RECT 678.750 564.600 680.550 564.900 ;
        RECT 676.950 563.700 677.850 564.600 ;
        RECT 595.950 554.850 598.050 556.950 ;
        RECT 607.950 556.050 610.050 558.150 ;
        RECT 610.950 554.850 613.050 556.950 ;
        RECT 613.950 556.050 616.050 558.150 ;
        RECT 640.950 557.850 643.050 559.950 ;
        RECT 662.700 558.150 663.900 563.400 ;
        RECT 572.100 543.750 573.900 552.000 ;
        RECT 592.950 551.700 594.750 552.600 ;
        RECT 591.450 550.800 594.750 551.700 ;
        RECT 591.450 546.600 592.350 550.800 ;
        RECT 597.000 549.600 598.050 554.850 ;
        RECT 611.100 553.050 612.900 554.850 ;
        RECT 614.850 552.750 616.050 556.050 ;
        RECT 641.400 553.650 642.600 557.850 ;
        RECT 652.950 554.850 655.050 556.950 ;
        RECT 656.100 555.150 657.900 556.950 ;
        RECT 615.000 551.700 618.750 552.750 ;
        RECT 587.550 543.750 589.350 546.600 ;
        RECT 590.550 543.750 592.350 546.600 ;
        RECT 593.550 543.750 595.350 546.600 ;
        RECT 596.550 543.750 598.350 549.600 ;
        RECT 608.550 548.700 616.350 550.050 ;
        RECT 608.550 543.750 610.350 548.700 ;
        RECT 611.550 543.750 613.350 547.800 ;
        RECT 614.550 543.750 616.350 548.700 ;
        RECT 617.550 549.600 618.750 551.700 ;
        RECT 617.550 543.750 619.350 549.600 ;
        RECT 632.700 543.750 634.500 552.600 ;
        RECT 638.100 552.000 642.600 553.650 ;
        RECT 653.100 553.050 654.900 554.850 ;
        RECT 655.950 553.050 658.050 555.150 ;
        RECT 658.950 554.850 661.050 556.950 ;
        RECT 661.950 556.050 664.050 558.150 ;
        RECT 659.100 553.050 660.900 554.850 ;
        RECT 638.100 543.750 639.900 552.000 ;
        RECT 662.700 549.600 663.900 556.050 ;
        RECT 654.000 543.750 655.800 549.600 ;
        RECT 658.200 547.950 663.900 549.600 ;
        RECT 668.550 553.950 669.750 563.400 ;
        RECT 673.950 562.800 676.050 563.700 ;
        RECT 676.950 562.800 682.950 563.700 ;
        RECT 671.850 561.600 676.050 562.800 ;
        RECT 670.950 559.800 672.750 561.600 ;
        RECT 682.050 558.150 682.950 562.800 ;
        RECT 684.150 562.800 685.050 564.900 ;
        RECT 685.950 564.300 693.450 565.500 ;
        RECT 685.950 563.700 687.750 564.300 ;
        RECT 700.050 563.400 701.850 575.250 ;
        RECT 712.350 563.400 714.150 575.250 ;
        RECT 715.350 563.400 717.150 575.250 ;
        RECT 718.650 569.400 720.450 575.250 ;
        RECT 731.400 569.400 733.200 575.250 ;
        RECT 690.750 562.800 701.850 563.400 ;
        RECT 684.150 562.200 701.850 562.800 ;
        RECT 684.150 561.900 692.550 562.200 ;
        RECT 690.750 561.600 692.550 561.900 ;
        RECT 682.050 556.050 685.050 558.150 ;
        RECT 688.950 557.100 691.050 558.150 ;
        RECT 688.950 556.050 696.900 557.100 ;
        RECT 670.950 555.750 673.050 556.050 ;
        RECT 670.950 553.950 674.850 555.750 ;
        RECT 668.550 551.850 673.050 553.950 ;
        RECT 682.050 552.000 682.950 556.050 ;
        RECT 695.100 555.300 696.900 556.050 ;
        RECT 698.100 555.150 699.900 556.950 ;
        RECT 692.100 554.400 693.900 555.000 ;
        RECT 698.100 554.400 699.000 555.150 ;
        RECT 692.100 553.200 699.000 554.400 ;
        RECT 692.100 552.000 693.150 553.200 ;
        RECT 668.550 549.600 669.750 551.850 ;
        RECT 682.050 551.100 693.150 552.000 ;
        RECT 682.050 550.800 682.950 551.100 ;
        RECT 658.200 543.750 660.000 547.950 ;
        RECT 661.500 543.750 663.300 546.600 ;
        RECT 668.550 543.750 670.350 549.600 ;
        RECT 673.950 548.700 676.050 549.600 ;
        RECT 681.150 549.000 682.950 550.800 ;
        RECT 692.100 550.200 693.150 551.100 ;
        RECT 688.350 549.450 690.150 550.200 ;
        RECT 673.950 547.500 677.700 548.700 ;
        RECT 676.650 546.600 677.700 547.500 ;
        RECT 685.200 548.400 690.150 549.450 ;
        RECT 691.650 548.400 693.450 550.200 ;
        RECT 700.950 549.600 701.850 562.200 ;
        RECT 712.650 558.150 713.850 563.400 ;
        RECT 719.250 562.500 720.450 569.400 ;
        RECT 734.700 563.400 736.500 575.250 ;
        RECT 738.900 563.400 740.700 575.250 ;
        RECT 752.550 569.400 754.350 575.250 ;
        RECT 755.550 569.400 757.350 575.250 ;
        RECT 714.750 561.600 720.450 562.500 ;
        RECT 714.750 560.700 717.000 561.600 ;
        RECT 731.250 561.150 733.050 562.950 ;
        RECT 712.650 556.050 715.050 558.150 ;
        RECT 712.650 549.600 713.850 556.050 ;
        RECT 715.950 552.300 717.000 560.700 ;
        RECT 719.100 558.150 720.900 559.950 ;
        RECT 730.950 559.050 733.050 561.150 ;
        RECT 734.850 558.150 736.050 563.400 ;
        RECT 740.100 558.150 741.900 559.950 ;
        RECT 718.950 556.050 721.050 558.150 ;
        RECT 733.950 556.050 736.050 558.150 ;
        RECT 733.950 552.750 735.150 556.050 ;
        RECT 736.950 554.850 739.050 556.950 ;
        RECT 739.950 556.050 742.050 558.150 ;
        RECT 755.400 556.950 756.600 569.400 ;
        RECT 768.300 563.400 770.100 575.250 ;
        RECT 772.500 563.400 774.300 575.250 ;
        RECT 775.800 569.400 777.600 575.250 ;
        RECT 788.550 569.400 790.350 575.250 ;
        RECT 791.550 569.400 793.350 575.250 ;
        RECT 806.550 569.400 808.350 575.250 ;
        RECT 809.550 569.400 811.350 575.250 ;
        RECT 812.550 570.000 814.350 575.250 ;
        RECT 767.100 558.150 768.900 559.950 ;
        RECT 772.950 558.150 774.150 563.400 ;
        RECT 778.950 562.950 781.050 565.050 ;
        RECT 775.950 561.150 777.750 562.950 ;
        RECT 775.950 559.050 778.050 561.150 ;
        RECT 752.100 555.150 753.900 556.950 ;
        RECT 737.100 553.050 738.900 554.850 ;
        RECT 751.950 553.050 754.050 555.150 ;
        RECT 754.950 554.850 757.050 556.950 ;
        RECT 766.950 556.050 769.050 558.150 ;
        RECT 769.950 554.850 772.050 556.950 ;
        RECT 772.950 556.050 775.050 558.150 ;
        RECT 714.750 551.400 717.000 552.300 ;
        RECT 731.250 551.700 735.000 552.750 ;
        RECT 714.750 550.500 719.850 551.400 ;
        RECT 685.200 546.600 686.250 548.400 ;
        RECT 694.950 547.500 697.050 549.600 ;
        RECT 694.950 546.600 696.000 547.500 ;
        RECT 671.850 543.750 673.650 546.600 ;
        RECT 676.350 543.750 678.150 546.600 ;
        RECT 680.550 543.750 682.350 546.600 ;
        RECT 684.450 543.750 686.250 546.600 ;
        RECT 687.750 543.750 689.550 546.600 ;
        RECT 692.250 545.700 696.000 546.600 ;
        RECT 692.250 543.750 694.050 545.700 ;
        RECT 697.050 543.750 698.850 546.600 ;
        RECT 700.050 543.750 701.850 549.600 ;
        RECT 712.350 543.750 714.150 549.600 ;
        RECT 715.350 543.750 717.150 549.600 ;
        RECT 718.650 546.600 719.850 550.500 ;
        RECT 731.250 549.600 732.450 551.700 ;
        RECT 718.650 543.750 720.450 546.600 ;
        RECT 730.650 543.750 732.450 549.600 ;
        RECT 733.650 548.700 741.450 550.050 ;
        RECT 733.650 543.750 735.450 548.700 ;
        RECT 736.650 543.750 738.450 547.800 ;
        RECT 739.650 543.750 741.450 548.700 ;
        RECT 755.400 546.600 756.600 554.850 ;
        RECT 770.100 553.050 771.900 554.850 ;
        RECT 773.850 552.750 775.050 556.050 ;
        RECT 775.950 555.450 778.050 556.050 ;
        RECT 779.550 555.450 780.450 562.950 ;
        RECT 791.400 556.950 792.600 569.400 ;
        RECT 809.700 569.100 811.350 569.400 ;
        RECT 815.550 569.400 817.350 575.250 ;
        RECT 830.550 569.400 832.350 575.250 ;
        RECT 833.550 569.400 835.350 575.250 ;
        RECT 845.550 569.400 847.350 575.250 ;
        RECT 848.550 569.400 850.350 575.250 ;
        RECT 851.550 569.400 853.350 575.250 ;
        RECT 866.550 569.400 868.350 575.250 ;
        RECT 869.550 569.400 871.350 575.250 ;
        RECT 872.550 569.400 874.350 575.250 ;
        RECT 815.550 569.100 816.750 569.400 ;
        RECT 809.700 568.200 816.750 569.100 ;
        RECT 809.100 564.150 810.900 565.950 ;
        RECT 806.100 561.150 807.900 562.950 ;
        RECT 808.950 562.050 811.050 564.150 ;
        RECT 812.250 561.150 814.050 562.950 ;
        RECT 805.950 559.050 808.050 561.150 ;
        RECT 811.950 559.050 814.050 561.150 ;
        RECT 815.700 559.950 816.750 568.200 ;
        RECT 814.950 557.850 817.050 559.950 ;
        RECT 775.950 554.550 780.450 555.450 ;
        RECT 788.100 555.150 789.900 556.950 ;
        RECT 775.950 553.950 778.050 554.550 ;
        RECT 787.950 553.050 790.050 555.150 ;
        RECT 790.950 554.850 793.050 556.950 ;
        RECT 774.000 551.700 777.750 552.750 ;
        RECT 767.550 548.700 775.350 550.050 ;
        RECT 752.550 543.750 754.350 546.600 ;
        RECT 755.550 543.750 757.350 546.600 ;
        RECT 767.550 543.750 769.350 548.700 ;
        RECT 770.550 543.750 772.350 547.800 ;
        RECT 773.550 543.750 775.350 548.700 ;
        RECT 776.550 549.600 777.750 551.700 ;
        RECT 776.550 543.750 778.350 549.600 ;
        RECT 791.400 546.600 792.600 554.850 ;
        RECT 815.400 553.650 816.600 557.850 ;
        RECT 833.400 556.950 834.600 569.400 ;
        RECT 848.550 561.150 849.750 569.400 ;
        RECT 869.550 561.150 870.750 569.400 ;
        RECT 844.950 557.850 847.050 559.950 ;
        RECT 847.950 559.050 850.050 561.150 ;
        RECT 830.100 555.150 831.900 556.950 ;
        RECT 788.550 543.750 790.350 546.600 ;
        RECT 791.550 543.750 793.350 546.600 ;
        RECT 806.700 543.750 808.500 552.600 ;
        RECT 812.100 552.000 816.600 553.650 ;
        RECT 829.950 553.050 832.050 555.150 ;
        RECT 832.950 554.850 835.050 556.950 ;
        RECT 845.100 556.050 846.900 557.850 ;
        RECT 812.100 543.750 813.900 552.000 ;
        RECT 833.400 546.600 834.600 554.850 ;
        RECT 848.550 551.700 849.750 559.050 ;
        RECT 850.950 557.850 853.050 559.950 ;
        RECT 865.950 557.850 868.050 559.950 ;
        RECT 868.950 559.050 871.050 561.150 ;
        RECT 851.100 556.050 852.900 557.850 ;
        RECT 866.100 556.050 867.900 557.850 ;
        RECT 869.550 551.700 870.750 559.050 ;
        RECT 871.950 557.850 874.050 559.950 ;
        RECT 872.100 556.050 873.900 557.850 ;
        RECT 848.550 550.800 852.150 551.700 ;
        RECT 869.550 550.800 873.150 551.700 ;
        RECT 830.550 543.750 832.350 546.600 ;
        RECT 833.550 543.750 835.350 546.600 ;
        RECT 845.850 543.750 847.650 549.600 ;
        RECT 850.350 543.750 852.150 550.800 ;
        RECT 866.850 543.750 868.650 549.600 ;
        RECT 871.350 543.750 873.150 550.800 ;
        RECT 3.150 533.400 4.950 539.250 ;
        RECT 6.150 536.400 7.950 539.250 ;
        RECT 10.950 537.300 12.750 539.250 ;
        RECT 9.000 536.400 12.750 537.300 ;
        RECT 15.450 536.400 17.250 539.250 ;
        RECT 18.750 536.400 20.550 539.250 ;
        RECT 22.650 536.400 24.450 539.250 ;
        RECT 26.850 536.400 28.650 539.250 ;
        RECT 31.350 536.400 33.150 539.250 ;
        RECT 9.000 535.500 10.050 536.400 ;
        RECT 7.950 533.400 10.050 535.500 ;
        RECT 18.750 534.600 19.800 536.400 ;
        RECT 3.150 520.800 4.050 533.400 ;
        RECT 11.550 532.800 13.350 534.600 ;
        RECT 14.850 533.550 19.800 534.600 ;
        RECT 27.300 535.500 28.350 536.400 ;
        RECT 27.300 534.300 31.050 535.500 ;
        RECT 14.850 532.800 16.650 533.550 ;
        RECT 11.850 531.900 12.900 532.800 ;
        RECT 22.050 532.200 23.850 534.000 ;
        RECT 28.950 533.400 31.050 534.300 ;
        RECT 34.650 533.400 36.450 539.250 ;
        RECT 22.050 531.900 22.950 532.200 ;
        RECT 11.850 531.000 22.950 531.900 ;
        RECT 35.250 531.150 36.450 533.400 ;
        RECT 47.550 534.300 49.350 539.250 ;
        RECT 50.550 535.200 52.350 539.250 ;
        RECT 53.550 534.300 55.350 539.250 ;
        RECT 47.550 532.950 55.350 534.300 ;
        RECT 56.550 533.400 58.350 539.250 ;
        RECT 56.550 531.300 57.750 533.400 ;
        RECT 71.850 532.200 73.650 539.250 ;
        RECT 76.350 533.400 78.150 539.250 ;
        RECT 88.650 536.400 90.450 539.250 ;
        RECT 91.650 536.400 93.450 539.250 ;
        RECT 94.650 536.400 96.450 539.250 ;
        RECT 71.850 531.300 75.450 532.200 ;
        RECT 11.850 529.800 12.900 531.000 ;
        RECT 6.000 528.600 12.900 529.800 ;
        RECT 6.000 527.850 6.900 528.600 ;
        RECT 11.100 528.000 12.900 528.600 ;
        RECT 5.100 526.050 6.900 527.850 ;
        RECT 8.100 526.950 9.900 527.700 ;
        RECT 22.050 526.950 22.950 531.000 ;
        RECT 31.950 529.050 36.450 531.150 ;
        RECT 54.000 530.250 57.750 531.300 ;
        RECT 30.150 527.250 34.050 529.050 ;
        RECT 31.950 526.950 34.050 527.250 ;
        RECT 8.100 525.900 16.050 526.950 ;
        RECT 13.950 524.850 16.050 525.900 ;
        RECT 19.950 524.850 22.950 526.950 ;
        RECT 12.450 521.100 14.250 521.400 ;
        RECT 12.450 520.800 20.850 521.100 ;
        RECT 3.150 520.200 20.850 520.800 ;
        RECT 3.150 519.600 14.250 520.200 ;
        RECT 3.150 507.750 4.950 519.600 ;
        RECT 17.250 518.700 19.050 519.300 ;
        RECT 11.550 517.500 19.050 518.700 ;
        RECT 19.950 518.100 20.850 520.200 ;
        RECT 22.050 520.200 22.950 524.850 ;
        RECT 32.250 521.400 34.050 523.200 ;
        RECT 28.950 520.200 33.150 521.400 ;
        RECT 22.050 519.300 28.050 520.200 ;
        RECT 28.950 519.300 31.050 520.200 ;
        RECT 35.250 519.600 36.450 529.050 ;
        RECT 50.100 528.150 51.900 529.950 ;
        RECT 46.950 524.850 49.050 526.950 ;
        RECT 49.950 526.050 52.050 528.150 ;
        RECT 53.850 526.950 55.050 530.250 ;
        RECT 52.950 524.850 55.050 526.950 ;
        RECT 71.100 525.150 72.900 526.950 ;
        RECT 47.100 523.050 48.900 524.850 ;
        RECT 52.950 519.600 54.150 524.850 ;
        RECT 55.950 521.850 58.050 523.950 ;
        RECT 70.950 523.050 73.050 525.150 ;
        RECT 74.250 523.950 75.450 531.300 ;
        RECT 91.950 529.950 93.000 536.400 ;
        RECT 106.650 533.400 108.450 539.250 ;
        RECT 107.250 531.300 108.450 533.400 ;
        RECT 109.650 534.300 111.450 539.250 ;
        RECT 112.650 535.200 114.450 539.250 ;
        RECT 115.650 534.300 117.450 539.250 ;
        RECT 125.550 536.400 127.350 539.250 ;
        RECT 128.550 536.400 130.350 539.250 ;
        RECT 131.550 536.400 133.350 539.250 ;
        RECT 109.650 532.950 117.450 534.300 ;
        RECT 107.250 530.250 111.000 531.300 ;
        RECT 91.950 527.850 94.050 529.950 ;
        RECT 77.100 525.150 78.900 526.950 ;
        RECT 73.950 521.850 76.050 523.950 ;
        RECT 76.950 523.050 79.050 525.150 ;
        RECT 88.950 524.850 91.050 526.950 ;
        RECT 89.100 523.050 90.900 524.850 ;
        RECT 55.950 520.050 57.750 521.850 ;
        RECT 27.150 518.400 28.050 519.300 ;
        RECT 24.450 518.100 26.250 518.400 ;
        RECT 11.550 516.600 12.750 517.500 ;
        RECT 19.950 517.200 26.250 518.100 ;
        RECT 24.450 516.600 26.250 517.200 ;
        RECT 27.150 516.600 29.850 518.400 ;
        RECT 7.950 514.500 12.750 516.600 ;
        RECT 15.150 514.500 22.050 516.300 ;
        RECT 11.550 513.600 12.750 514.500 ;
        RECT 6.150 507.750 7.950 513.600 ;
        RECT 11.250 507.750 13.050 513.600 ;
        RECT 16.050 507.750 17.850 513.600 ;
        RECT 19.050 507.750 20.850 514.500 ;
        RECT 27.150 513.600 31.050 515.700 ;
        RECT 22.950 507.750 24.750 513.600 ;
        RECT 27.150 507.750 28.950 513.600 ;
        RECT 31.650 507.750 33.450 510.600 ;
        RECT 34.650 507.750 36.450 519.600 ;
        RECT 48.300 507.750 50.100 519.600 ;
        RECT 52.500 507.750 54.300 519.600 ;
        RECT 74.250 513.600 75.450 521.850 ;
        RECT 91.950 520.650 93.000 527.850 ;
        RECT 109.950 526.950 111.150 530.250 ;
        RECT 129.000 529.950 130.050 536.400 ;
        RECT 148.650 533.400 150.450 539.250 ;
        RECT 149.250 531.300 150.450 533.400 ;
        RECT 151.650 534.300 153.450 539.250 ;
        RECT 154.650 535.200 156.450 539.250 ;
        RECT 157.650 534.300 159.450 539.250 ;
        RECT 167.550 536.400 169.350 539.250 ;
        RECT 170.550 536.400 172.350 539.250 ;
        RECT 151.650 532.950 159.450 534.300 ;
        RECT 149.250 530.250 153.000 531.300 ;
        RECT 113.100 528.150 114.900 529.950 ;
        RECT 94.950 524.850 97.050 526.950 ;
        RECT 109.950 524.850 112.050 526.950 ;
        RECT 112.950 526.050 115.050 528.150 ;
        RECT 127.950 527.850 130.050 529.950 ;
        RECT 115.950 524.850 118.050 526.950 ;
        RECT 124.950 524.850 127.050 526.950 ;
        RECT 95.100 523.050 96.900 524.850 ;
        RECT 106.950 521.850 109.050 523.950 ;
        RECT 90.450 519.600 93.000 520.650 ;
        RECT 107.250 520.050 109.050 521.850 ;
        RECT 110.850 519.600 112.050 524.850 ;
        RECT 116.100 523.050 117.900 524.850 ;
        RECT 125.100 523.050 126.900 524.850 ;
        RECT 129.000 520.650 130.050 527.850 ;
        RECT 151.950 526.950 153.150 530.250 ;
        RECT 155.100 528.150 156.900 529.950 ;
        RECT 130.950 524.850 133.050 526.950 ;
        RECT 151.950 524.850 154.050 526.950 ;
        RECT 154.950 526.050 157.050 528.150 ;
        RECT 166.950 527.850 169.050 529.950 ;
        RECT 170.400 528.150 171.600 536.400 ;
        RECT 182.550 534.300 184.350 539.250 ;
        RECT 185.550 535.200 187.350 539.250 ;
        RECT 188.550 534.300 190.350 539.250 ;
        RECT 182.550 532.950 190.350 534.300 ;
        RECT 191.550 533.400 193.350 539.250 ;
        RECT 191.550 531.300 192.750 533.400 ;
        RECT 206.850 532.200 208.650 539.250 ;
        RECT 211.350 533.400 213.150 539.250 ;
        RECT 216.150 533.400 217.950 539.250 ;
        RECT 219.150 536.400 220.950 539.250 ;
        RECT 223.950 537.300 225.750 539.250 ;
        RECT 222.000 536.400 225.750 537.300 ;
        RECT 228.450 536.400 230.250 539.250 ;
        RECT 231.750 536.400 233.550 539.250 ;
        RECT 235.650 536.400 237.450 539.250 ;
        RECT 239.850 536.400 241.650 539.250 ;
        RECT 244.350 536.400 246.150 539.250 ;
        RECT 222.000 535.500 223.050 536.400 ;
        RECT 220.950 533.400 223.050 535.500 ;
        RECT 231.750 534.600 232.800 536.400 ;
        RECT 206.850 531.300 210.450 532.200 ;
        RECT 189.000 530.250 192.750 531.300 ;
        RECT 185.100 528.150 186.900 529.950 ;
        RECT 157.950 524.850 160.050 526.950 ;
        RECT 167.100 526.050 168.900 527.850 ;
        RECT 169.950 526.050 172.050 528.150 ;
        RECT 131.100 523.050 132.900 524.850 ;
        RECT 148.950 521.850 151.050 523.950 ;
        RECT 129.000 519.600 131.550 520.650 ;
        RECT 149.250 520.050 151.050 521.850 ;
        RECT 152.850 519.600 154.050 524.850 ;
        RECT 158.100 523.050 159.900 524.850 ;
        RECT 55.800 507.750 57.600 513.600 ;
        RECT 70.650 507.750 72.450 513.600 ;
        RECT 73.650 507.750 75.450 513.600 ;
        RECT 76.650 507.750 78.450 513.600 ;
        RECT 90.450 507.750 92.250 519.600 ;
        RECT 94.650 507.750 96.450 519.600 ;
        RECT 107.400 507.750 109.200 513.600 ;
        RECT 110.700 507.750 112.500 519.600 ;
        RECT 114.900 507.750 116.700 519.600 ;
        RECT 125.550 507.750 127.350 519.600 ;
        RECT 129.750 507.750 131.550 519.600 ;
        RECT 149.400 507.750 151.200 513.600 ;
        RECT 152.700 507.750 154.500 519.600 ;
        RECT 156.900 507.750 158.700 519.600 ;
        RECT 170.400 513.600 171.600 526.050 ;
        RECT 181.950 524.850 184.050 526.950 ;
        RECT 184.950 526.050 187.050 528.150 ;
        RECT 188.850 526.950 190.050 530.250 ;
        RECT 187.950 524.850 190.050 526.950 ;
        RECT 206.100 525.150 207.900 526.950 ;
        RECT 182.100 523.050 183.900 524.850 ;
        RECT 187.950 519.600 189.150 524.850 ;
        RECT 190.950 521.850 193.050 523.950 ;
        RECT 205.950 523.050 208.050 525.150 ;
        RECT 209.250 523.950 210.450 531.300 ;
        RECT 212.100 525.150 213.900 526.950 ;
        RECT 208.950 521.850 211.050 523.950 ;
        RECT 211.950 523.050 214.050 525.150 ;
        RECT 190.950 520.050 192.750 521.850 ;
        RECT 167.550 507.750 169.350 513.600 ;
        RECT 170.550 507.750 172.350 513.600 ;
        RECT 183.300 507.750 185.100 519.600 ;
        RECT 187.500 507.750 189.300 519.600 ;
        RECT 209.250 513.600 210.450 521.850 ;
        RECT 216.150 520.800 217.050 533.400 ;
        RECT 224.550 532.800 226.350 534.600 ;
        RECT 227.850 533.550 232.800 534.600 ;
        RECT 240.300 535.500 241.350 536.400 ;
        RECT 240.300 534.300 244.050 535.500 ;
        RECT 227.850 532.800 229.650 533.550 ;
        RECT 224.850 531.900 225.900 532.800 ;
        RECT 235.050 532.200 236.850 534.000 ;
        RECT 241.950 533.400 244.050 534.300 ;
        RECT 247.650 533.400 249.450 539.250 ;
        RECT 259.650 536.400 261.450 539.250 ;
        RECT 262.650 536.400 264.450 539.250 ;
        RECT 235.050 531.900 235.950 532.200 ;
        RECT 224.850 531.000 235.950 531.900 ;
        RECT 248.250 531.150 249.450 533.400 ;
        RECT 224.850 529.800 225.900 531.000 ;
        RECT 219.000 528.600 225.900 529.800 ;
        RECT 219.000 527.850 219.900 528.600 ;
        RECT 224.100 528.000 225.900 528.600 ;
        RECT 218.100 526.050 219.900 527.850 ;
        RECT 221.100 526.950 222.900 527.700 ;
        RECT 235.050 526.950 235.950 531.000 ;
        RECT 244.950 529.050 249.450 531.150 ;
        RECT 243.150 527.250 247.050 529.050 ;
        RECT 244.950 526.950 247.050 527.250 ;
        RECT 221.100 525.900 229.050 526.950 ;
        RECT 226.950 524.850 229.050 525.900 ;
        RECT 232.950 524.850 235.950 526.950 ;
        RECT 225.450 521.100 227.250 521.400 ;
        RECT 225.450 520.800 233.850 521.100 ;
        RECT 216.150 520.200 233.850 520.800 ;
        RECT 216.150 519.600 227.250 520.200 ;
        RECT 190.800 507.750 192.600 513.600 ;
        RECT 205.650 507.750 207.450 513.600 ;
        RECT 208.650 507.750 210.450 513.600 ;
        RECT 211.650 507.750 213.450 513.600 ;
        RECT 216.150 507.750 217.950 519.600 ;
        RECT 230.250 518.700 232.050 519.300 ;
        RECT 224.550 517.500 232.050 518.700 ;
        RECT 232.950 518.100 233.850 520.200 ;
        RECT 235.050 520.200 235.950 524.850 ;
        RECT 245.250 521.400 247.050 523.200 ;
        RECT 241.950 520.200 246.150 521.400 ;
        RECT 235.050 519.300 241.050 520.200 ;
        RECT 241.950 519.300 244.050 520.200 ;
        RECT 248.250 519.600 249.450 529.050 ;
        RECT 260.400 528.150 261.600 536.400 ;
        RECT 272.550 534.300 274.350 539.250 ;
        RECT 275.550 535.200 277.350 539.250 ;
        RECT 278.550 534.300 280.350 539.250 ;
        RECT 272.550 532.950 280.350 534.300 ;
        RECT 281.550 533.400 283.350 539.250 ;
        RECT 296.550 536.400 298.350 539.250 ;
        RECT 299.550 536.400 301.350 539.250 ;
        RECT 281.550 531.300 282.750 533.400 ;
        RECT 279.000 530.250 282.750 531.300 ;
        RECT 259.950 526.050 262.050 528.150 ;
        RECT 262.950 527.850 265.050 529.950 ;
        RECT 275.100 528.150 276.900 529.950 ;
        RECT 263.100 526.050 264.900 527.850 ;
        RECT 240.150 518.400 241.050 519.300 ;
        RECT 237.450 518.100 239.250 518.400 ;
        RECT 224.550 516.600 225.750 517.500 ;
        RECT 232.950 517.200 239.250 518.100 ;
        RECT 237.450 516.600 239.250 517.200 ;
        RECT 240.150 516.600 242.850 518.400 ;
        RECT 220.950 514.500 225.750 516.600 ;
        RECT 228.150 514.500 235.050 516.300 ;
        RECT 224.550 513.600 225.750 514.500 ;
        RECT 219.150 507.750 220.950 513.600 ;
        RECT 224.250 507.750 226.050 513.600 ;
        RECT 229.050 507.750 230.850 513.600 ;
        RECT 232.050 507.750 233.850 514.500 ;
        RECT 240.150 513.600 244.050 515.700 ;
        RECT 235.950 507.750 237.750 513.600 ;
        RECT 240.150 507.750 241.950 513.600 ;
        RECT 244.650 507.750 246.450 510.600 ;
        RECT 247.650 507.750 249.450 519.600 ;
        RECT 260.400 513.600 261.600 526.050 ;
        RECT 271.950 524.850 274.050 526.950 ;
        RECT 274.950 526.050 277.050 528.150 ;
        RECT 278.850 526.950 280.050 530.250 ;
        RECT 295.950 527.850 298.050 529.950 ;
        RECT 299.400 528.150 300.600 536.400 ;
        RECT 314.850 532.200 316.650 539.250 ;
        RECT 319.350 533.400 321.150 539.250 ;
        RECT 332.550 536.400 334.350 539.250 ;
        RECT 335.550 536.400 337.350 539.250 ;
        RECT 314.850 531.300 318.450 532.200 ;
        RECT 277.950 524.850 280.050 526.950 ;
        RECT 296.100 526.050 297.900 527.850 ;
        RECT 298.950 526.050 301.050 528.150 ;
        RECT 272.100 523.050 273.900 524.850 ;
        RECT 277.950 519.600 279.150 524.850 ;
        RECT 280.950 521.850 283.050 523.950 ;
        RECT 280.950 520.050 282.750 521.850 ;
        RECT 259.650 507.750 261.450 513.600 ;
        RECT 262.650 507.750 264.450 513.600 ;
        RECT 273.300 507.750 275.100 519.600 ;
        RECT 277.500 507.750 279.300 519.600 ;
        RECT 299.400 513.600 300.600 526.050 ;
        RECT 314.100 525.150 315.900 526.950 ;
        RECT 313.950 523.050 316.050 525.150 ;
        RECT 317.250 523.950 318.450 531.300 ;
        RECT 331.950 527.850 334.050 529.950 ;
        RECT 335.400 528.150 336.600 536.400 ;
        RECT 347.850 533.400 349.650 539.250 ;
        RECT 352.350 532.200 354.150 539.250 ;
        RECT 370.650 536.400 372.450 539.250 ;
        RECT 373.650 536.400 375.450 539.250 ;
        RECT 350.550 531.300 354.150 532.200 ;
        RECT 320.100 525.150 321.900 526.950 ;
        RECT 332.100 526.050 333.900 527.850 ;
        RECT 334.950 526.050 337.050 528.150 ;
        RECT 316.950 521.850 319.050 523.950 ;
        RECT 319.950 523.050 322.050 525.150 ;
        RECT 317.250 513.600 318.450 521.850 ;
        RECT 335.400 513.600 336.600 526.050 ;
        RECT 347.100 525.150 348.900 526.950 ;
        RECT 346.950 523.050 349.050 525.150 ;
        RECT 350.550 523.950 351.750 531.300 ;
        RECT 371.400 528.150 372.600 536.400 ;
        RECT 386.550 534.300 388.350 539.250 ;
        RECT 389.550 535.200 391.350 539.250 ;
        RECT 392.550 534.300 394.350 539.250 ;
        RECT 386.550 532.950 394.350 534.300 ;
        RECT 395.550 533.400 397.350 539.250 ;
        RECT 410.550 534.300 412.350 539.250 ;
        RECT 413.550 535.200 415.350 539.250 ;
        RECT 416.550 534.300 418.350 539.250 ;
        RECT 395.550 531.300 396.750 533.400 ;
        RECT 410.550 532.950 418.350 534.300 ;
        RECT 419.550 533.400 421.350 539.250 ;
        RECT 426.150 533.400 427.950 539.250 ;
        RECT 429.150 536.400 430.950 539.250 ;
        RECT 433.950 537.300 435.750 539.250 ;
        RECT 432.000 536.400 435.750 537.300 ;
        RECT 438.450 536.400 440.250 539.250 ;
        RECT 441.750 536.400 443.550 539.250 ;
        RECT 445.650 536.400 447.450 539.250 ;
        RECT 449.850 536.400 451.650 539.250 ;
        RECT 454.350 536.400 456.150 539.250 ;
        RECT 432.000 535.500 433.050 536.400 ;
        RECT 430.950 533.400 433.050 535.500 ;
        RECT 441.750 534.600 442.800 536.400 ;
        RECT 419.550 531.300 420.750 533.400 ;
        RECT 393.000 530.250 396.750 531.300 ;
        RECT 417.000 530.250 420.750 531.300 ;
        RECT 353.100 525.150 354.900 526.950 ;
        RECT 370.950 526.050 373.050 528.150 ;
        RECT 373.950 527.850 376.050 529.950 ;
        RECT 389.100 528.150 390.900 529.950 ;
        RECT 374.100 526.050 375.900 527.850 ;
        RECT 349.950 521.850 352.050 523.950 ;
        RECT 352.950 523.050 355.050 525.150 ;
        RECT 350.550 513.600 351.750 521.850 ;
        RECT 371.400 513.600 372.600 526.050 ;
        RECT 385.950 524.850 388.050 526.950 ;
        RECT 388.950 526.050 391.050 528.150 ;
        RECT 392.850 526.950 394.050 530.250 ;
        RECT 413.100 528.150 414.900 529.950 ;
        RECT 391.950 524.850 394.050 526.950 ;
        RECT 409.950 524.850 412.050 526.950 ;
        RECT 412.950 526.050 415.050 528.150 ;
        RECT 416.850 526.950 418.050 530.250 ;
        RECT 415.950 524.850 418.050 526.950 ;
        RECT 386.100 523.050 387.900 524.850 ;
        RECT 391.950 519.600 393.150 524.850 ;
        RECT 394.950 521.850 397.050 523.950 ;
        RECT 410.100 523.050 411.900 524.850 ;
        RECT 394.950 520.050 396.750 521.850 ;
        RECT 415.950 519.600 417.150 524.850 ;
        RECT 418.950 521.850 421.050 523.950 ;
        RECT 418.950 520.050 420.750 521.850 ;
        RECT 426.150 520.800 427.050 533.400 ;
        RECT 434.550 532.800 436.350 534.600 ;
        RECT 437.850 533.550 442.800 534.600 ;
        RECT 450.300 535.500 451.350 536.400 ;
        RECT 450.300 534.300 454.050 535.500 ;
        RECT 437.850 532.800 439.650 533.550 ;
        RECT 434.850 531.900 435.900 532.800 ;
        RECT 445.050 532.200 446.850 534.000 ;
        RECT 451.950 533.400 454.050 534.300 ;
        RECT 457.650 533.400 459.450 539.250 ;
        RECT 445.050 531.900 445.950 532.200 ;
        RECT 434.850 531.000 445.950 531.900 ;
        RECT 458.250 531.150 459.450 533.400 ;
        RECT 434.850 529.800 435.900 531.000 ;
        RECT 429.000 528.600 435.900 529.800 ;
        RECT 429.000 527.850 429.900 528.600 ;
        RECT 434.100 528.000 435.900 528.600 ;
        RECT 428.100 526.050 429.900 527.850 ;
        RECT 431.100 526.950 432.900 527.700 ;
        RECT 445.050 526.950 445.950 531.000 ;
        RECT 454.950 529.050 459.450 531.150 ;
        RECT 453.150 527.250 457.050 529.050 ;
        RECT 454.950 526.950 457.050 527.250 ;
        RECT 431.100 525.900 439.050 526.950 ;
        RECT 436.950 524.850 439.050 525.900 ;
        RECT 442.950 524.850 445.950 526.950 ;
        RECT 435.450 521.100 437.250 521.400 ;
        RECT 435.450 520.800 443.850 521.100 ;
        RECT 426.150 520.200 443.850 520.800 ;
        RECT 426.150 519.600 437.250 520.200 ;
        RECT 280.800 507.750 282.600 513.600 ;
        RECT 296.550 507.750 298.350 513.600 ;
        RECT 299.550 507.750 301.350 513.600 ;
        RECT 313.650 507.750 315.450 513.600 ;
        RECT 316.650 507.750 318.450 513.600 ;
        RECT 319.650 507.750 321.450 513.600 ;
        RECT 332.550 507.750 334.350 513.600 ;
        RECT 335.550 507.750 337.350 513.600 ;
        RECT 347.550 507.750 349.350 513.600 ;
        RECT 350.550 507.750 352.350 513.600 ;
        RECT 353.550 507.750 355.350 513.600 ;
        RECT 370.650 507.750 372.450 513.600 ;
        RECT 373.650 507.750 375.450 513.600 ;
        RECT 387.300 507.750 389.100 519.600 ;
        RECT 391.500 507.750 393.300 519.600 ;
        RECT 394.800 507.750 396.600 513.600 ;
        RECT 411.300 507.750 413.100 519.600 ;
        RECT 415.500 507.750 417.300 519.600 ;
        RECT 418.800 507.750 420.600 513.600 ;
        RECT 426.150 507.750 427.950 519.600 ;
        RECT 440.250 518.700 442.050 519.300 ;
        RECT 434.550 517.500 442.050 518.700 ;
        RECT 442.950 518.100 443.850 520.200 ;
        RECT 445.050 520.200 445.950 524.850 ;
        RECT 455.250 521.400 457.050 523.200 ;
        RECT 451.950 520.200 456.150 521.400 ;
        RECT 445.050 519.300 451.050 520.200 ;
        RECT 451.950 519.300 454.050 520.200 ;
        RECT 458.250 519.600 459.450 529.050 ;
        RECT 450.150 518.400 451.050 519.300 ;
        RECT 447.450 518.100 449.250 518.400 ;
        RECT 434.550 516.600 435.750 517.500 ;
        RECT 442.950 517.200 449.250 518.100 ;
        RECT 447.450 516.600 449.250 517.200 ;
        RECT 450.150 516.600 452.850 518.400 ;
        RECT 430.950 514.500 435.750 516.600 ;
        RECT 438.150 514.500 445.050 516.300 ;
        RECT 434.550 513.600 435.750 514.500 ;
        RECT 429.150 507.750 430.950 513.600 ;
        RECT 434.250 507.750 436.050 513.600 ;
        RECT 439.050 507.750 440.850 513.600 ;
        RECT 442.050 507.750 443.850 514.500 ;
        RECT 450.150 513.600 454.050 515.700 ;
        RECT 445.950 507.750 447.750 513.600 ;
        RECT 450.150 507.750 451.950 513.600 ;
        RECT 454.650 507.750 456.450 510.600 ;
        RECT 457.650 507.750 459.450 519.600 ;
        RECT 462.150 533.400 463.950 539.250 ;
        RECT 465.150 536.400 466.950 539.250 ;
        RECT 469.950 537.300 471.750 539.250 ;
        RECT 468.000 536.400 471.750 537.300 ;
        RECT 474.450 536.400 476.250 539.250 ;
        RECT 477.750 536.400 479.550 539.250 ;
        RECT 481.650 536.400 483.450 539.250 ;
        RECT 485.850 536.400 487.650 539.250 ;
        RECT 490.350 536.400 492.150 539.250 ;
        RECT 468.000 535.500 469.050 536.400 ;
        RECT 466.950 533.400 469.050 535.500 ;
        RECT 477.750 534.600 478.800 536.400 ;
        RECT 462.150 520.800 463.050 533.400 ;
        RECT 470.550 532.800 472.350 534.600 ;
        RECT 473.850 533.550 478.800 534.600 ;
        RECT 486.300 535.500 487.350 536.400 ;
        RECT 486.300 534.300 490.050 535.500 ;
        RECT 473.850 532.800 475.650 533.550 ;
        RECT 470.850 531.900 471.900 532.800 ;
        RECT 481.050 532.200 482.850 534.000 ;
        RECT 487.950 533.400 490.050 534.300 ;
        RECT 493.650 533.400 495.450 539.250 ;
        RECT 506.700 536.400 508.500 539.250 ;
        RECT 510.000 535.050 511.800 539.250 ;
        RECT 481.050 531.900 481.950 532.200 ;
        RECT 470.850 531.000 481.950 531.900 ;
        RECT 494.250 531.150 495.450 533.400 ;
        RECT 470.850 529.800 471.900 531.000 ;
        RECT 465.000 528.600 471.900 529.800 ;
        RECT 465.000 527.850 465.900 528.600 ;
        RECT 470.100 528.000 471.900 528.600 ;
        RECT 464.100 526.050 465.900 527.850 ;
        RECT 467.100 526.950 468.900 527.700 ;
        RECT 481.050 526.950 481.950 531.000 ;
        RECT 490.950 529.050 495.450 531.150 ;
        RECT 489.150 527.250 493.050 529.050 ;
        RECT 490.950 526.950 493.050 527.250 ;
        RECT 467.100 525.900 475.050 526.950 ;
        RECT 472.950 524.850 475.050 525.900 ;
        RECT 478.950 524.850 481.950 526.950 ;
        RECT 471.450 521.100 473.250 521.400 ;
        RECT 471.450 520.800 479.850 521.100 ;
        RECT 462.150 520.200 479.850 520.800 ;
        RECT 462.150 519.600 473.250 520.200 ;
        RECT 462.150 507.750 463.950 519.600 ;
        RECT 476.250 518.700 478.050 519.300 ;
        RECT 470.550 517.500 478.050 518.700 ;
        RECT 478.950 518.100 479.850 520.200 ;
        RECT 481.050 520.200 481.950 524.850 ;
        RECT 491.250 521.400 493.050 523.200 ;
        RECT 487.950 520.200 492.150 521.400 ;
        RECT 481.050 519.300 487.050 520.200 ;
        RECT 487.950 519.300 490.050 520.200 ;
        RECT 494.250 519.600 495.450 529.050 ;
        RECT 506.100 533.400 511.800 535.050 ;
        RECT 514.200 533.400 516.000 539.250 ;
        RECT 506.100 526.950 507.300 533.400 ;
        RECT 524.550 531.900 526.350 539.250 ;
        RECT 529.050 533.400 530.850 539.250 ;
        RECT 532.050 534.900 533.850 539.250 ;
        RECT 532.050 533.400 535.350 534.900 ;
        RECT 550.650 533.400 552.450 539.250 ;
        RECT 530.250 531.900 532.050 532.500 ;
        RECT 524.550 530.700 532.050 531.900 ;
        RECT 509.100 528.150 510.900 529.950 ;
        RECT 505.950 524.850 508.050 526.950 ;
        RECT 508.950 526.050 511.050 528.150 ;
        RECT 511.950 527.850 514.050 529.950 ;
        RECT 515.100 528.150 516.900 529.950 ;
        RECT 512.100 526.050 513.900 527.850 ;
        RECT 514.950 526.050 517.050 528.150 ;
        RECT 523.950 524.850 526.050 526.950 ;
        RECT 506.100 519.600 507.300 524.850 ;
        RECT 524.100 523.050 525.900 524.850 ;
        RECT 486.150 518.400 487.050 519.300 ;
        RECT 483.450 518.100 485.250 518.400 ;
        RECT 470.550 516.600 471.750 517.500 ;
        RECT 478.950 517.200 485.250 518.100 ;
        RECT 483.450 516.600 485.250 517.200 ;
        RECT 486.150 516.600 488.850 518.400 ;
        RECT 466.950 514.500 471.750 516.600 ;
        RECT 474.150 514.500 481.050 516.300 ;
        RECT 470.550 513.600 471.750 514.500 ;
        RECT 465.150 507.750 466.950 513.600 ;
        RECT 470.250 507.750 472.050 513.600 ;
        RECT 475.050 507.750 476.850 513.600 ;
        RECT 478.050 507.750 479.850 514.500 ;
        RECT 486.150 513.600 490.050 515.700 ;
        RECT 481.950 507.750 483.750 513.600 ;
        RECT 486.150 507.750 487.950 513.600 ;
        RECT 490.650 507.750 492.450 510.600 ;
        RECT 493.650 507.750 495.450 519.600 ;
        RECT 505.650 507.750 507.450 519.600 ;
        RECT 508.650 518.700 516.450 519.600 ;
        RECT 508.650 507.750 510.450 518.700 ;
        RECT 511.650 507.750 513.450 517.800 ;
        RECT 514.650 507.750 516.450 518.700 ;
        RECT 527.700 513.600 528.900 530.700 ;
        RECT 534.150 526.950 535.350 533.400 ;
        RECT 551.250 531.300 552.450 533.400 ;
        RECT 553.650 534.300 555.450 539.250 ;
        RECT 556.650 535.200 558.450 539.250 ;
        RECT 559.650 534.300 561.450 539.250 ;
        RECT 571.650 536.400 573.450 539.250 ;
        RECT 574.650 536.400 576.450 539.250 ;
        RECT 553.650 532.950 561.450 534.300 ;
        RECT 551.250 530.250 555.000 531.300 ;
        RECT 530.100 525.150 531.900 526.950 ;
        RECT 529.950 523.050 532.050 525.150 ;
        RECT 532.950 524.850 535.350 526.950 ;
        RECT 553.950 526.950 555.150 530.250 ;
        RECT 557.100 528.150 558.900 529.950 ;
        RECT 572.400 528.150 573.600 536.400 ;
        RECT 587.700 530.400 589.500 539.250 ;
        RECT 593.100 531.000 594.900 539.250 ;
        RECT 611.550 536.400 613.350 539.250 ;
        RECT 614.550 536.400 616.350 539.250 ;
        RECT 617.550 536.400 619.350 539.250 ;
        RECT 553.950 524.850 556.050 526.950 ;
        RECT 556.950 526.050 559.050 528.150 ;
        RECT 559.950 524.850 562.050 526.950 ;
        RECT 571.950 526.050 574.050 528.150 ;
        RECT 574.950 527.850 577.050 529.950 ;
        RECT 593.100 529.350 597.600 531.000 ;
        RECT 615.000 529.950 616.050 536.400 ;
        RECT 632.550 534.300 634.350 539.250 ;
        RECT 635.550 535.200 637.350 539.250 ;
        RECT 638.550 534.300 640.350 539.250 ;
        RECT 632.550 532.950 640.350 534.300 ;
        RECT 641.550 533.400 643.350 539.250 ;
        RECT 653.550 534.300 655.350 539.250 ;
        RECT 656.550 535.200 658.350 539.250 ;
        RECT 659.550 534.300 661.350 539.250 ;
        RECT 641.550 531.300 642.750 533.400 ;
        RECT 653.550 532.950 661.350 534.300 ;
        RECT 662.550 533.400 664.350 539.250 ;
        RECT 674.850 533.400 676.650 539.250 ;
        RECT 662.550 531.300 663.750 533.400 ;
        RECT 679.350 532.200 681.150 539.250 ;
        RECT 639.000 530.250 642.750 531.300 ;
        RECT 660.000 530.250 663.750 531.300 ;
        RECT 677.550 531.300 681.150 532.200 ;
        RECT 687.150 533.400 688.950 539.250 ;
        RECT 690.150 536.400 691.950 539.250 ;
        RECT 694.950 537.300 696.750 539.250 ;
        RECT 693.000 536.400 696.750 537.300 ;
        RECT 699.450 536.400 701.250 539.250 ;
        RECT 702.750 536.400 704.550 539.250 ;
        RECT 706.650 536.400 708.450 539.250 ;
        RECT 710.850 536.400 712.650 539.250 ;
        RECT 715.350 536.400 717.150 539.250 ;
        RECT 693.000 535.500 694.050 536.400 ;
        RECT 691.950 533.400 694.050 535.500 ;
        RECT 702.750 534.600 703.800 536.400 ;
        RECT 575.100 526.050 576.900 527.850 ;
        RECT 534.150 519.600 535.350 524.850 ;
        RECT 550.950 521.850 553.050 523.950 ;
        RECT 551.250 520.050 553.050 521.850 ;
        RECT 554.850 519.600 556.050 524.850 ;
        RECT 560.100 523.050 561.900 524.850 ;
        RECT 524.550 507.750 526.350 513.600 ;
        RECT 527.550 507.750 529.350 513.600 ;
        RECT 531.150 507.750 532.950 519.600 ;
        RECT 534.150 507.750 535.950 519.600 ;
        RECT 551.400 507.750 553.200 513.600 ;
        RECT 554.700 507.750 556.500 519.600 ;
        RECT 558.900 507.750 560.700 519.600 ;
        RECT 572.400 513.600 573.600 526.050 ;
        RECT 596.400 525.150 597.600 529.350 ;
        RECT 613.950 527.850 616.050 529.950 ;
        RECT 635.100 528.150 636.900 529.950 ;
        RECT 586.950 521.850 589.050 523.950 ;
        RECT 592.950 521.850 595.050 523.950 ;
        RECT 595.950 523.050 598.050 525.150 ;
        RECT 610.950 524.850 613.050 526.950 ;
        RECT 611.100 523.050 612.900 524.850 ;
        RECT 587.100 520.050 588.900 521.850 ;
        RECT 589.950 518.850 592.050 520.950 ;
        RECT 593.250 520.050 595.050 521.850 ;
        RECT 590.100 517.050 591.900 518.850 ;
        RECT 596.700 514.800 597.750 523.050 ;
        RECT 615.000 520.650 616.050 527.850 ;
        RECT 616.950 524.850 619.050 526.950 ;
        RECT 631.950 524.850 634.050 526.950 ;
        RECT 634.950 526.050 637.050 528.150 ;
        RECT 638.850 526.950 640.050 530.250 ;
        RECT 656.100 528.150 657.900 529.950 ;
        RECT 637.950 524.850 640.050 526.950 ;
        RECT 652.950 524.850 655.050 526.950 ;
        RECT 655.950 526.050 658.050 528.150 ;
        RECT 659.850 526.950 661.050 530.250 ;
        RECT 658.950 524.850 661.050 526.950 ;
        RECT 674.100 525.150 675.900 526.950 ;
        RECT 617.100 523.050 618.900 524.850 ;
        RECT 632.100 523.050 633.900 524.850 ;
        RECT 615.000 519.600 617.550 520.650 ;
        RECT 637.950 519.600 639.150 524.850 ;
        RECT 640.950 521.850 643.050 523.950 ;
        RECT 653.100 523.050 654.900 524.850 ;
        RECT 640.950 520.050 642.750 521.850 ;
        RECT 658.950 519.600 660.150 524.850 ;
        RECT 661.950 521.850 664.050 523.950 ;
        RECT 673.950 523.050 676.050 525.150 ;
        RECT 677.550 523.950 678.750 531.300 ;
        RECT 680.100 525.150 681.900 526.950 ;
        RECT 676.950 521.850 679.050 523.950 ;
        RECT 679.950 523.050 682.050 525.150 ;
        RECT 661.950 520.050 663.750 521.850 ;
        RECT 590.700 513.900 597.750 514.800 ;
        RECT 590.700 513.600 592.350 513.900 ;
        RECT 571.650 507.750 573.450 513.600 ;
        RECT 574.650 507.750 576.450 513.600 ;
        RECT 587.550 507.750 589.350 513.600 ;
        RECT 590.550 507.750 592.350 513.600 ;
        RECT 596.550 513.600 597.750 513.900 ;
        RECT 593.550 507.750 595.350 513.000 ;
        RECT 596.550 507.750 598.350 513.600 ;
        RECT 611.550 507.750 613.350 519.600 ;
        RECT 615.750 507.750 617.550 519.600 ;
        RECT 633.300 507.750 635.100 519.600 ;
        RECT 637.500 507.750 639.300 519.600 ;
        RECT 640.800 507.750 642.600 513.600 ;
        RECT 654.300 507.750 656.100 519.600 ;
        RECT 658.500 507.750 660.300 519.600 ;
        RECT 677.550 513.600 678.750 521.850 ;
        RECT 687.150 520.800 688.050 533.400 ;
        RECT 695.550 532.800 697.350 534.600 ;
        RECT 698.850 533.550 703.800 534.600 ;
        RECT 711.300 535.500 712.350 536.400 ;
        RECT 711.300 534.300 715.050 535.500 ;
        RECT 698.850 532.800 700.650 533.550 ;
        RECT 695.850 531.900 696.900 532.800 ;
        RECT 706.050 532.200 707.850 534.000 ;
        RECT 712.950 533.400 715.050 534.300 ;
        RECT 718.650 533.400 720.450 539.250 ;
        RECT 728.550 536.400 730.350 539.250 ;
        RECT 731.550 536.400 733.350 539.250 ;
        RECT 706.050 531.900 706.950 532.200 ;
        RECT 695.850 531.000 706.950 531.900 ;
        RECT 719.250 531.150 720.450 533.400 ;
        RECT 695.850 529.800 696.900 531.000 ;
        RECT 690.000 528.600 696.900 529.800 ;
        RECT 690.000 527.850 690.900 528.600 ;
        RECT 695.100 528.000 696.900 528.600 ;
        RECT 689.100 526.050 690.900 527.850 ;
        RECT 692.100 526.950 693.900 527.700 ;
        RECT 706.050 526.950 706.950 531.000 ;
        RECT 715.950 529.050 720.450 531.150 ;
        RECT 714.150 527.250 718.050 529.050 ;
        RECT 715.950 526.950 718.050 527.250 ;
        RECT 692.100 525.900 700.050 526.950 ;
        RECT 697.950 524.850 700.050 525.900 ;
        RECT 703.950 524.850 706.950 526.950 ;
        RECT 696.450 521.100 698.250 521.400 ;
        RECT 696.450 520.800 704.850 521.100 ;
        RECT 687.150 520.200 704.850 520.800 ;
        RECT 687.150 519.600 698.250 520.200 ;
        RECT 661.800 507.750 663.600 513.600 ;
        RECT 674.550 507.750 676.350 513.600 ;
        RECT 677.550 507.750 679.350 513.600 ;
        RECT 680.550 507.750 682.350 513.600 ;
        RECT 687.150 507.750 688.950 519.600 ;
        RECT 701.250 518.700 703.050 519.300 ;
        RECT 695.550 517.500 703.050 518.700 ;
        RECT 703.950 518.100 704.850 520.200 ;
        RECT 706.050 520.200 706.950 524.850 ;
        RECT 716.250 521.400 718.050 523.200 ;
        RECT 712.950 520.200 717.150 521.400 ;
        RECT 706.050 519.300 712.050 520.200 ;
        RECT 712.950 519.300 715.050 520.200 ;
        RECT 719.250 519.600 720.450 529.050 ;
        RECT 727.950 527.850 730.050 529.950 ;
        RECT 731.400 528.150 732.600 536.400 ;
        RECT 746.850 532.200 748.650 539.250 ;
        RECT 751.350 533.400 753.150 539.250 ;
        RECT 761.550 536.400 763.350 539.250 ;
        RECT 764.550 536.400 766.350 539.250 ;
        RECT 767.550 536.400 769.350 539.250 ;
        RECT 746.850 531.300 750.450 532.200 ;
        RECT 728.100 526.050 729.900 527.850 ;
        RECT 730.950 526.050 733.050 528.150 ;
        RECT 711.150 518.400 712.050 519.300 ;
        RECT 708.450 518.100 710.250 518.400 ;
        RECT 695.550 516.600 696.750 517.500 ;
        RECT 703.950 517.200 710.250 518.100 ;
        RECT 708.450 516.600 710.250 517.200 ;
        RECT 711.150 516.600 713.850 518.400 ;
        RECT 691.950 514.500 696.750 516.600 ;
        RECT 699.150 514.500 706.050 516.300 ;
        RECT 695.550 513.600 696.750 514.500 ;
        RECT 690.150 507.750 691.950 513.600 ;
        RECT 695.250 507.750 697.050 513.600 ;
        RECT 700.050 507.750 701.850 513.600 ;
        RECT 703.050 507.750 704.850 514.500 ;
        RECT 711.150 513.600 715.050 515.700 ;
        RECT 706.950 507.750 708.750 513.600 ;
        RECT 711.150 507.750 712.950 513.600 ;
        RECT 715.650 507.750 717.450 510.600 ;
        RECT 718.650 507.750 720.450 519.600 ;
        RECT 731.400 513.600 732.600 526.050 ;
        RECT 746.100 525.150 747.900 526.950 ;
        RECT 745.950 523.050 748.050 525.150 ;
        RECT 749.250 523.950 750.450 531.300 ;
        RECT 765.000 529.950 766.050 536.400 ;
        RECT 784.650 533.400 786.450 539.250 ;
        RECT 787.650 533.400 789.450 539.250 ;
        RECT 763.950 527.850 766.050 529.950 ;
        RECT 752.100 525.150 753.900 526.950 ;
        RECT 748.950 521.850 751.050 523.950 ;
        RECT 751.950 523.050 754.050 525.150 ;
        RECT 760.950 524.850 763.050 526.950 ;
        RECT 761.100 523.050 762.900 524.850 ;
        RECT 749.250 513.600 750.450 521.850 ;
        RECT 765.000 520.650 766.050 527.850 ;
        RECT 785.400 526.950 786.600 533.400 ;
        RECT 800.850 532.200 802.650 539.250 ;
        RECT 805.350 533.400 807.150 539.250 ;
        RECT 820.650 533.400 822.450 539.250 ;
        RECT 800.850 531.300 804.450 532.200 ;
        RECT 788.100 528.150 789.900 529.950 ;
        RECT 766.950 524.850 769.050 526.950 ;
        RECT 784.950 524.850 787.050 526.950 ;
        RECT 787.950 526.050 790.050 528.150 ;
        RECT 800.100 525.150 801.900 526.950 ;
        RECT 767.100 523.050 768.900 524.850 ;
        RECT 765.000 519.600 767.550 520.650 ;
        RECT 785.400 519.600 786.600 524.850 ;
        RECT 799.950 523.050 802.050 525.150 ;
        RECT 803.250 523.950 804.450 531.300 ;
        RECT 821.250 531.300 822.450 533.400 ;
        RECT 823.650 534.300 825.450 539.250 ;
        RECT 826.650 535.200 828.450 539.250 ;
        RECT 829.650 534.300 831.450 539.250 ;
        RECT 823.650 532.950 831.450 534.300 ;
        RECT 834.150 533.400 835.950 539.250 ;
        RECT 837.150 536.400 838.950 539.250 ;
        RECT 841.950 537.300 843.750 539.250 ;
        RECT 840.000 536.400 843.750 537.300 ;
        RECT 846.450 536.400 848.250 539.250 ;
        RECT 849.750 536.400 851.550 539.250 ;
        RECT 853.650 536.400 855.450 539.250 ;
        RECT 857.850 536.400 859.650 539.250 ;
        RECT 862.350 536.400 864.150 539.250 ;
        RECT 840.000 535.500 841.050 536.400 ;
        RECT 838.950 533.400 841.050 535.500 ;
        RECT 849.750 534.600 850.800 536.400 ;
        RECT 821.250 530.250 825.000 531.300 ;
        RECT 811.950 528.450 814.050 529.050 ;
        RECT 820.950 528.450 823.050 529.050 ;
        RECT 811.950 527.550 823.050 528.450 ;
        RECT 811.950 526.950 814.050 527.550 ;
        RECT 820.950 526.950 823.050 527.550 ;
        RECT 823.950 526.950 825.150 530.250 ;
        RECT 827.100 528.150 828.900 529.950 ;
        RECT 806.100 525.150 807.900 526.950 ;
        RECT 802.950 521.850 805.050 523.950 ;
        RECT 805.950 523.050 808.050 525.150 ;
        RECT 823.950 524.850 826.050 526.950 ;
        RECT 826.950 526.050 829.050 528.150 ;
        RECT 829.950 524.850 832.050 526.950 ;
        RECT 820.950 521.850 823.050 523.950 ;
        RECT 728.550 507.750 730.350 513.600 ;
        RECT 731.550 507.750 733.350 513.600 ;
        RECT 745.650 507.750 747.450 513.600 ;
        RECT 748.650 507.750 750.450 513.600 ;
        RECT 751.650 507.750 753.450 513.600 ;
        RECT 761.550 507.750 763.350 519.600 ;
        RECT 765.750 507.750 767.550 519.600 ;
        RECT 784.650 507.750 786.450 519.600 ;
        RECT 787.650 507.750 789.450 519.600 ;
        RECT 803.250 513.600 804.450 521.850 ;
        RECT 821.250 520.050 823.050 521.850 ;
        RECT 824.850 519.600 826.050 524.850 ;
        RECT 830.100 523.050 831.900 524.850 ;
        RECT 834.150 520.800 835.050 533.400 ;
        RECT 842.550 532.800 844.350 534.600 ;
        RECT 845.850 533.550 850.800 534.600 ;
        RECT 858.300 535.500 859.350 536.400 ;
        RECT 858.300 534.300 862.050 535.500 ;
        RECT 845.850 532.800 847.650 533.550 ;
        RECT 842.850 531.900 843.900 532.800 ;
        RECT 853.050 532.200 854.850 534.000 ;
        RECT 859.950 533.400 862.050 534.300 ;
        RECT 865.650 533.400 867.450 539.250 ;
        RECT 878.550 536.400 880.350 539.250 ;
        RECT 881.550 536.400 883.350 539.250 ;
        RECT 853.050 531.900 853.950 532.200 ;
        RECT 842.850 531.000 853.950 531.900 ;
        RECT 866.250 531.150 867.450 533.400 ;
        RECT 842.850 529.800 843.900 531.000 ;
        RECT 837.000 528.600 843.900 529.800 ;
        RECT 837.000 527.850 837.900 528.600 ;
        RECT 842.100 528.000 843.900 528.600 ;
        RECT 836.100 526.050 837.900 527.850 ;
        RECT 839.100 526.950 840.900 527.700 ;
        RECT 853.050 526.950 853.950 531.000 ;
        RECT 862.950 529.050 867.450 531.150 ;
        RECT 861.150 527.250 865.050 529.050 ;
        RECT 862.950 526.950 865.050 527.250 ;
        RECT 839.100 525.900 847.050 526.950 ;
        RECT 844.950 524.850 847.050 525.900 ;
        RECT 850.950 524.850 853.950 526.950 ;
        RECT 843.450 521.100 845.250 521.400 ;
        RECT 843.450 520.800 851.850 521.100 ;
        RECT 834.150 520.200 851.850 520.800 ;
        RECT 834.150 519.600 845.250 520.200 ;
        RECT 799.650 507.750 801.450 513.600 ;
        RECT 802.650 507.750 804.450 513.600 ;
        RECT 805.650 507.750 807.450 513.600 ;
        RECT 821.400 507.750 823.200 513.600 ;
        RECT 824.700 507.750 826.500 519.600 ;
        RECT 828.900 507.750 830.700 519.600 ;
        RECT 834.150 507.750 835.950 519.600 ;
        RECT 848.250 518.700 850.050 519.300 ;
        RECT 842.550 517.500 850.050 518.700 ;
        RECT 850.950 518.100 851.850 520.200 ;
        RECT 853.050 520.200 853.950 524.850 ;
        RECT 863.250 521.400 865.050 523.200 ;
        RECT 859.950 520.200 864.150 521.400 ;
        RECT 853.050 519.300 859.050 520.200 ;
        RECT 859.950 519.300 862.050 520.200 ;
        RECT 866.250 519.600 867.450 529.050 ;
        RECT 877.950 527.850 880.050 529.950 ;
        RECT 881.400 528.150 882.600 536.400 ;
        RECT 878.100 526.050 879.900 527.850 ;
        RECT 880.950 526.050 883.050 528.150 ;
        RECT 858.150 518.400 859.050 519.300 ;
        RECT 855.450 518.100 857.250 518.400 ;
        RECT 842.550 516.600 843.750 517.500 ;
        RECT 850.950 517.200 857.250 518.100 ;
        RECT 855.450 516.600 857.250 517.200 ;
        RECT 858.150 516.600 860.850 518.400 ;
        RECT 838.950 514.500 843.750 516.600 ;
        RECT 846.150 514.500 853.050 516.300 ;
        RECT 842.550 513.600 843.750 514.500 ;
        RECT 837.150 507.750 838.950 513.600 ;
        RECT 842.250 507.750 844.050 513.600 ;
        RECT 847.050 507.750 848.850 513.600 ;
        RECT 850.050 507.750 851.850 514.500 ;
        RECT 858.150 513.600 862.050 515.700 ;
        RECT 853.950 507.750 855.750 513.600 ;
        RECT 858.150 507.750 859.950 513.600 ;
        RECT 862.650 507.750 864.450 510.600 ;
        RECT 865.650 507.750 867.450 519.600 ;
        RECT 881.400 513.600 882.600 526.050 ;
        RECT 878.550 507.750 880.350 513.600 ;
        RECT 881.550 507.750 883.350 513.600 ;
        RECT 12.450 491.400 14.250 503.250 ;
        RECT 16.650 491.400 18.450 503.250 ;
        RECT 21.150 491.400 22.950 503.250 ;
        RECT 24.150 497.400 25.950 503.250 ;
        RECT 29.250 497.400 31.050 503.250 ;
        RECT 34.050 497.400 35.850 503.250 ;
        RECT 29.550 496.500 30.750 497.400 ;
        RECT 37.050 496.500 38.850 503.250 ;
        RECT 40.950 497.400 42.750 503.250 ;
        RECT 45.150 497.400 46.950 503.250 ;
        RECT 49.650 500.400 51.450 503.250 ;
        RECT 25.950 494.400 30.750 496.500 ;
        RECT 33.150 494.700 40.050 496.500 ;
        RECT 45.150 495.300 49.050 497.400 ;
        RECT 29.550 493.500 30.750 494.400 ;
        RECT 42.450 493.800 44.250 494.400 ;
        RECT 29.550 492.300 37.050 493.500 ;
        RECT 35.250 491.700 37.050 492.300 ;
        RECT 37.950 492.900 44.250 493.800 ;
        RECT 12.450 490.350 15.000 491.400 ;
        RECT 11.100 486.150 12.900 487.950 ;
        RECT 10.950 484.050 13.050 486.150 ;
        RECT 13.950 483.150 15.000 490.350 ;
        RECT 21.150 490.800 32.250 491.400 ;
        RECT 37.950 490.800 38.850 492.900 ;
        RECT 42.450 492.600 44.250 492.900 ;
        RECT 45.150 492.600 47.850 494.400 ;
        RECT 45.150 491.700 46.050 492.600 ;
        RECT 21.150 490.200 38.850 490.800 ;
        RECT 17.100 486.150 18.900 487.950 ;
        RECT 16.950 484.050 19.050 486.150 ;
        RECT 13.950 481.050 16.050 483.150 ;
        RECT 13.950 474.600 15.000 481.050 ;
        RECT 21.150 477.600 22.050 490.200 ;
        RECT 30.450 489.900 38.850 490.200 ;
        RECT 40.050 490.800 46.050 491.700 ;
        RECT 46.950 490.800 49.050 491.700 ;
        RECT 52.650 491.400 54.450 503.250 ;
        RECT 68.400 497.400 70.200 503.250 ;
        RECT 71.700 491.400 73.500 503.250 ;
        RECT 75.900 491.400 77.700 503.250 ;
        RECT 88.650 497.400 90.450 503.250 ;
        RECT 91.650 497.400 93.450 503.250 ;
        RECT 30.450 489.600 32.250 489.900 ;
        RECT 40.050 486.150 40.950 490.800 ;
        RECT 46.950 489.600 51.150 490.800 ;
        RECT 50.250 487.800 52.050 489.600 ;
        RECT 31.950 485.100 34.050 486.150 ;
        RECT 23.100 483.150 24.900 484.950 ;
        RECT 26.100 484.050 34.050 485.100 ;
        RECT 37.950 484.050 40.950 486.150 ;
        RECT 26.100 483.300 27.900 484.050 ;
        RECT 24.000 482.400 24.900 483.150 ;
        RECT 29.100 482.400 30.900 483.000 ;
        RECT 24.000 481.200 30.900 482.400 ;
        RECT 29.850 480.000 30.900 481.200 ;
        RECT 40.050 480.000 40.950 484.050 ;
        RECT 49.950 483.750 52.050 484.050 ;
        RECT 48.150 481.950 52.050 483.750 ;
        RECT 53.250 481.950 54.450 491.400 ;
        RECT 68.250 489.150 70.050 490.950 ;
        RECT 67.950 487.050 70.050 489.150 ;
        RECT 71.850 486.150 73.050 491.400 ;
        RECT 77.100 486.150 78.900 487.950 ;
        RECT 29.850 479.100 40.950 480.000 ;
        RECT 49.950 479.850 54.450 481.950 ;
        RECT 70.950 484.050 73.050 486.150 ;
        RECT 70.950 480.750 72.150 484.050 ;
        RECT 73.950 482.850 76.050 484.950 ;
        RECT 76.950 484.050 79.050 486.150 ;
        RECT 89.400 484.950 90.600 497.400 ;
        RECT 105.450 491.400 107.250 503.250 ;
        RECT 109.650 491.400 111.450 503.250 ;
        RECT 120.300 491.400 122.100 503.250 ;
        RECT 124.500 491.400 126.300 503.250 ;
        RECT 127.800 497.400 129.600 503.250 ;
        RECT 145.650 497.400 147.450 503.250 ;
        RECT 148.650 497.400 150.450 503.250 ;
        RECT 151.650 497.400 153.450 503.250 ;
        RECT 164.400 497.400 166.200 503.250 ;
        RECT 105.450 490.350 108.000 491.400 ;
        RECT 104.100 486.150 105.900 487.950 ;
        RECT 88.950 482.850 91.050 484.950 ;
        RECT 92.100 483.150 93.900 484.950 ;
        RECT 103.950 484.050 106.050 486.150 ;
        RECT 106.950 483.150 108.000 490.350 ;
        RECT 110.100 486.150 111.900 487.950 ;
        RECT 119.100 486.150 120.900 487.950 ;
        RECT 124.950 486.150 126.150 491.400 ;
        RECT 127.950 489.150 129.750 490.950 ;
        RECT 149.250 489.150 150.450 497.400 ;
        RECT 167.700 491.400 169.500 503.250 ;
        RECT 171.900 491.400 173.700 503.250 ;
        RECT 176.550 491.400 178.350 503.250 ;
        RECT 179.550 500.400 181.350 503.250 ;
        RECT 184.050 497.400 185.850 503.250 ;
        RECT 188.250 497.400 190.050 503.250 ;
        RECT 181.950 495.300 185.850 497.400 ;
        RECT 192.150 496.500 193.950 503.250 ;
        RECT 195.150 497.400 196.950 503.250 ;
        RECT 199.950 497.400 201.750 503.250 ;
        RECT 205.050 497.400 206.850 503.250 ;
        RECT 200.250 496.500 201.450 497.400 ;
        RECT 190.950 494.700 197.850 496.500 ;
        RECT 200.250 494.400 205.050 496.500 ;
        RECT 183.150 492.600 185.850 494.400 ;
        RECT 186.750 493.800 188.550 494.400 ;
        RECT 186.750 492.900 193.050 493.800 ;
        RECT 200.250 493.500 201.450 494.400 ;
        RECT 186.750 492.600 188.550 492.900 ;
        RECT 184.950 491.700 185.850 492.600 ;
        RECT 164.250 489.150 166.050 490.950 ;
        RECT 127.950 487.050 130.050 489.150 ;
        RECT 109.950 484.050 112.050 486.150 ;
        RECT 118.950 484.050 121.050 486.150 ;
        RECT 74.100 481.050 75.900 482.850 ;
        RECT 29.850 478.200 30.900 479.100 ;
        RECT 40.050 478.800 40.950 479.100 ;
        RECT 10.650 471.750 12.450 474.600 ;
        RECT 13.650 471.750 15.450 474.600 ;
        RECT 16.650 471.750 18.450 474.600 ;
        RECT 21.150 471.750 22.950 477.600 ;
        RECT 25.950 475.500 28.050 477.600 ;
        RECT 29.550 476.400 31.350 478.200 ;
        RECT 32.850 477.450 34.650 478.200 ;
        RECT 32.850 476.400 37.800 477.450 ;
        RECT 40.050 477.000 41.850 478.800 ;
        RECT 53.250 477.600 54.450 479.850 ;
        RECT 68.250 479.700 72.000 480.750 ;
        RECT 68.250 477.600 69.450 479.700 ;
        RECT 46.950 476.700 49.050 477.600 ;
        RECT 27.000 474.600 28.050 475.500 ;
        RECT 36.750 474.600 37.800 476.400 ;
        RECT 45.300 475.500 49.050 476.700 ;
        RECT 45.300 474.600 46.350 475.500 ;
        RECT 24.150 471.750 25.950 474.600 ;
        RECT 27.000 473.700 30.750 474.600 ;
        RECT 28.950 471.750 30.750 473.700 ;
        RECT 33.450 471.750 35.250 474.600 ;
        RECT 36.750 471.750 38.550 474.600 ;
        RECT 40.650 471.750 42.450 474.600 ;
        RECT 44.850 471.750 46.650 474.600 ;
        RECT 49.350 471.750 51.150 474.600 ;
        RECT 52.650 471.750 54.450 477.600 ;
        RECT 67.650 471.750 69.450 477.600 ;
        RECT 70.650 476.700 78.450 478.050 ;
        RECT 70.650 471.750 72.450 476.700 ;
        RECT 73.650 471.750 75.450 475.800 ;
        RECT 76.650 471.750 78.450 476.700 ;
        RECT 89.400 474.600 90.600 482.850 ;
        RECT 91.950 481.050 94.050 483.150 ;
        RECT 106.950 481.050 109.050 483.150 ;
        RECT 121.950 482.850 124.050 484.950 ;
        RECT 124.950 484.050 127.050 486.150 ;
        RECT 145.950 485.850 148.050 487.950 ;
        RECT 148.950 487.050 151.050 489.150 ;
        RECT 146.100 484.050 147.900 485.850 ;
        RECT 122.100 481.050 123.900 482.850 ;
        RECT 94.950 480.450 97.050 481.050 ;
        RECT 103.950 480.450 106.050 481.050 ;
        RECT 94.950 479.550 106.050 480.450 ;
        RECT 94.950 478.950 97.050 479.550 ;
        RECT 103.950 478.950 106.050 479.550 ;
        RECT 106.950 474.600 108.000 481.050 ;
        RECT 125.850 480.750 127.050 484.050 ;
        RECT 126.000 479.700 129.750 480.750 ;
        RECT 149.250 479.700 150.450 487.050 ;
        RECT 151.950 485.850 154.050 487.950 ;
        RECT 163.950 487.050 166.050 489.150 ;
        RECT 167.850 486.150 169.050 491.400 ;
        RECT 173.100 486.150 174.900 487.950 ;
        RECT 152.100 484.050 153.900 485.850 ;
        RECT 166.950 484.050 169.050 486.150 ;
        RECT 166.950 480.750 168.150 484.050 ;
        RECT 169.950 482.850 172.050 484.950 ;
        RECT 172.950 484.050 175.050 486.150 ;
        RECT 170.100 481.050 171.900 482.850 ;
        RECT 176.550 481.950 177.750 491.400 ;
        RECT 181.950 490.800 184.050 491.700 ;
        RECT 184.950 490.800 190.950 491.700 ;
        RECT 179.850 489.600 184.050 490.800 ;
        RECT 178.950 487.800 180.750 489.600 ;
        RECT 190.050 486.150 190.950 490.800 ;
        RECT 192.150 490.800 193.050 492.900 ;
        RECT 193.950 492.300 201.450 493.500 ;
        RECT 193.950 491.700 195.750 492.300 ;
        RECT 208.050 491.400 209.850 503.250 ;
        RECT 221.550 497.400 223.350 503.250 ;
        RECT 224.550 497.400 226.350 503.250 ;
        RECT 227.550 497.400 229.350 503.250 ;
        RECT 198.750 490.800 209.850 491.400 ;
        RECT 192.150 490.200 209.850 490.800 ;
        RECT 192.150 489.900 200.550 490.200 ;
        RECT 198.750 489.600 200.550 489.900 ;
        RECT 190.050 484.050 193.050 486.150 ;
        RECT 196.950 485.100 199.050 486.150 ;
        RECT 196.950 484.050 204.900 485.100 ;
        RECT 178.950 483.750 181.050 484.050 ;
        RECT 178.950 481.950 182.850 483.750 ;
        RECT 119.550 476.700 127.350 478.050 ;
        RECT 88.650 471.750 90.450 474.600 ;
        RECT 91.650 471.750 93.450 474.600 ;
        RECT 103.650 471.750 105.450 474.600 ;
        RECT 106.650 471.750 108.450 474.600 ;
        RECT 109.650 471.750 111.450 474.600 ;
        RECT 119.550 471.750 121.350 476.700 ;
        RECT 122.550 471.750 124.350 475.800 ;
        RECT 125.550 471.750 127.350 476.700 ;
        RECT 128.550 477.600 129.750 479.700 ;
        RECT 146.850 478.800 150.450 479.700 ;
        RECT 164.250 479.700 168.000 480.750 ;
        RECT 176.550 479.850 181.050 481.950 ;
        RECT 190.050 480.000 190.950 484.050 ;
        RECT 203.100 483.300 204.900 484.050 ;
        RECT 206.100 483.150 207.900 484.950 ;
        RECT 200.100 482.400 201.900 483.000 ;
        RECT 206.100 482.400 207.000 483.150 ;
        RECT 200.100 481.200 207.000 482.400 ;
        RECT 200.100 480.000 201.150 481.200 ;
        RECT 128.550 471.750 130.350 477.600 ;
        RECT 146.850 471.750 148.650 478.800 ;
        RECT 164.250 477.600 165.450 479.700 ;
        RECT 151.350 471.750 153.150 477.600 ;
        RECT 163.650 471.750 165.450 477.600 ;
        RECT 166.650 476.700 174.450 478.050 ;
        RECT 166.650 471.750 168.450 476.700 ;
        RECT 169.650 471.750 171.450 475.800 ;
        RECT 172.650 471.750 174.450 476.700 ;
        RECT 176.550 477.600 177.750 479.850 ;
        RECT 190.050 479.100 201.150 480.000 ;
        RECT 190.050 478.800 190.950 479.100 ;
        RECT 176.550 471.750 178.350 477.600 ;
        RECT 181.950 476.700 184.050 477.600 ;
        RECT 189.150 477.000 190.950 478.800 ;
        RECT 200.100 478.200 201.150 479.100 ;
        RECT 196.350 477.450 198.150 478.200 ;
        RECT 181.950 475.500 185.700 476.700 ;
        RECT 184.650 474.600 185.700 475.500 ;
        RECT 193.200 476.400 198.150 477.450 ;
        RECT 199.650 476.400 201.450 478.200 ;
        RECT 208.950 477.600 209.850 490.200 ;
        RECT 224.550 489.150 225.750 497.400 ;
        RECT 241.350 491.400 243.150 503.250 ;
        RECT 244.350 491.400 246.150 503.250 ;
        RECT 247.650 497.400 249.450 503.250 ;
        RECT 260.400 497.400 262.200 503.250 ;
        RECT 220.950 485.850 223.050 487.950 ;
        RECT 223.950 487.050 226.050 489.150 ;
        RECT 221.100 484.050 222.900 485.850 ;
        RECT 224.550 479.700 225.750 487.050 ;
        RECT 226.950 485.850 229.050 487.950 ;
        RECT 241.650 486.150 242.850 491.400 ;
        RECT 248.250 490.500 249.450 497.400 ;
        RECT 263.700 491.400 265.500 503.250 ;
        RECT 267.900 491.400 269.700 503.250 ;
        RECT 279.300 491.400 281.100 503.250 ;
        RECT 283.500 491.400 285.300 503.250 ;
        RECT 286.800 497.400 288.600 503.250 ;
        RECT 299.550 497.400 301.350 503.250 ;
        RECT 302.550 497.400 304.350 503.250 ;
        RECT 305.550 497.400 307.350 503.250 ;
        RECT 243.750 489.600 249.450 490.500 ;
        RECT 243.750 488.700 246.000 489.600 ;
        RECT 260.250 489.150 262.050 490.950 ;
        RECT 227.100 484.050 228.900 485.850 ;
        RECT 241.650 484.050 244.050 486.150 ;
        RECT 224.550 478.800 228.150 479.700 ;
        RECT 193.200 474.600 194.250 476.400 ;
        RECT 202.950 475.500 205.050 477.600 ;
        RECT 202.950 474.600 204.000 475.500 ;
        RECT 179.850 471.750 181.650 474.600 ;
        RECT 184.350 471.750 186.150 474.600 ;
        RECT 188.550 471.750 190.350 474.600 ;
        RECT 192.450 471.750 194.250 474.600 ;
        RECT 195.750 471.750 197.550 474.600 ;
        RECT 200.250 473.700 204.000 474.600 ;
        RECT 200.250 471.750 202.050 473.700 ;
        RECT 205.050 471.750 206.850 474.600 ;
        RECT 208.050 471.750 209.850 477.600 ;
        RECT 221.850 471.750 223.650 477.600 ;
        RECT 226.350 471.750 228.150 478.800 ;
        RECT 241.650 477.600 242.850 484.050 ;
        RECT 244.950 480.300 246.000 488.700 ;
        RECT 248.100 486.150 249.900 487.950 ;
        RECT 259.950 487.050 262.050 489.150 ;
        RECT 263.850 486.150 265.050 491.400 ;
        RECT 269.100 486.150 270.900 487.950 ;
        RECT 278.100 486.150 279.900 487.950 ;
        RECT 283.950 486.150 285.150 491.400 ;
        RECT 286.950 489.150 288.750 490.950 ;
        RECT 302.550 489.150 303.750 497.400 ;
        RECT 319.650 491.400 321.450 503.250 ;
        RECT 322.650 491.400 324.450 503.250 ;
        RECT 334.650 497.400 336.450 503.250 ;
        RECT 337.650 497.400 339.450 503.250 ;
        RECT 340.650 497.400 342.450 503.250 ;
        RECT 353.400 497.400 355.200 503.250 ;
        RECT 286.950 487.050 289.050 489.150 ;
        RECT 247.950 484.050 250.050 486.150 ;
        RECT 262.950 484.050 265.050 486.150 ;
        RECT 262.950 480.750 264.150 484.050 ;
        RECT 265.950 482.850 268.050 484.950 ;
        RECT 268.950 484.050 271.050 486.150 ;
        RECT 277.950 484.050 280.050 486.150 ;
        RECT 280.950 482.850 283.050 484.950 ;
        RECT 283.950 484.050 286.050 486.150 ;
        RECT 298.950 485.850 301.050 487.950 ;
        RECT 301.950 487.050 304.050 489.150 ;
        RECT 299.100 484.050 300.900 485.850 ;
        RECT 266.100 481.050 267.900 482.850 ;
        RECT 281.100 481.050 282.900 482.850 ;
        RECT 284.850 480.750 286.050 484.050 ;
        RECT 243.750 479.400 246.000 480.300 ;
        RECT 260.250 479.700 264.000 480.750 ;
        RECT 285.000 479.700 288.750 480.750 ;
        RECT 243.750 478.500 248.850 479.400 ;
        RECT 241.350 471.750 243.150 477.600 ;
        RECT 244.350 471.750 246.150 477.600 ;
        RECT 247.650 474.600 248.850 478.500 ;
        RECT 260.250 477.600 261.450 479.700 ;
        RECT 247.650 471.750 249.450 474.600 ;
        RECT 259.650 471.750 261.450 477.600 ;
        RECT 262.650 476.700 270.450 478.050 ;
        RECT 262.650 471.750 264.450 476.700 ;
        RECT 265.650 471.750 267.450 475.800 ;
        RECT 268.650 471.750 270.450 476.700 ;
        RECT 278.550 476.700 286.350 478.050 ;
        RECT 278.550 471.750 280.350 476.700 ;
        RECT 281.550 471.750 283.350 475.800 ;
        RECT 284.550 471.750 286.350 476.700 ;
        RECT 287.550 477.600 288.750 479.700 ;
        RECT 302.550 479.700 303.750 487.050 ;
        RECT 304.950 485.850 307.050 487.950 ;
        RECT 320.400 486.150 321.600 491.400 ;
        RECT 338.250 489.150 339.450 497.400 ;
        RECT 356.700 491.400 358.500 503.250 ;
        RECT 360.900 491.400 362.700 503.250 ;
        RECT 373.650 497.400 375.450 503.250 ;
        RECT 376.650 497.400 378.450 503.250 ;
        RECT 379.650 497.400 381.450 503.250 ;
        RECT 391.650 497.400 393.450 503.250 ;
        RECT 394.650 497.400 396.450 503.250 ;
        RECT 397.650 497.400 399.450 503.250 ;
        RECT 409.650 497.400 411.450 503.250 ;
        RECT 412.650 497.400 414.450 503.250 ;
        RECT 415.650 497.400 417.450 503.250 ;
        RECT 431.400 497.400 433.200 503.250 ;
        RECT 353.250 489.150 355.050 490.950 ;
        RECT 305.100 484.050 306.900 485.850 ;
        RECT 319.950 484.050 322.050 486.150 ;
        RECT 334.950 485.850 337.050 487.950 ;
        RECT 337.950 487.050 340.050 489.150 ;
        RECT 302.550 478.800 306.150 479.700 ;
        RECT 287.550 471.750 289.350 477.600 ;
        RECT 299.850 471.750 301.650 477.600 ;
        RECT 304.350 471.750 306.150 478.800 ;
        RECT 320.400 477.600 321.600 484.050 ;
        RECT 322.950 482.850 325.050 484.950 ;
        RECT 335.100 484.050 336.900 485.850 ;
        RECT 323.100 481.050 324.900 482.850 ;
        RECT 338.250 479.700 339.450 487.050 ;
        RECT 340.950 485.850 343.050 487.950 ;
        RECT 352.950 487.050 355.050 489.150 ;
        RECT 356.850 486.150 358.050 491.400 ;
        RECT 377.250 489.150 378.450 497.400 ;
        RECT 395.250 489.150 396.450 497.400 ;
        RECT 413.250 489.150 414.450 497.400 ;
        RECT 434.700 491.400 436.500 503.250 ;
        RECT 438.900 491.400 440.700 503.250 ;
        RECT 451.650 497.400 453.450 503.250 ;
        RECT 454.650 497.400 456.450 503.250 ;
        RECT 431.250 489.150 433.050 490.950 ;
        RECT 362.100 486.150 363.900 487.950 ;
        RECT 341.100 484.050 342.900 485.850 ;
        RECT 355.950 484.050 358.050 486.150 ;
        RECT 355.950 480.750 357.150 484.050 ;
        RECT 358.950 482.850 361.050 484.950 ;
        RECT 361.950 484.050 364.050 486.150 ;
        RECT 373.950 485.850 376.050 487.950 ;
        RECT 376.950 487.050 379.050 489.150 ;
        RECT 374.100 484.050 375.900 485.850 ;
        RECT 359.100 481.050 360.900 482.850 ;
        RECT 335.850 478.800 339.450 479.700 ;
        RECT 353.250 479.700 357.000 480.750 ;
        RECT 377.250 479.700 378.450 487.050 ;
        RECT 379.950 485.850 382.050 487.950 ;
        RECT 391.950 485.850 394.050 487.950 ;
        RECT 394.950 487.050 397.050 489.150 ;
        RECT 380.100 484.050 381.900 485.850 ;
        RECT 392.100 484.050 393.900 485.850 ;
        RECT 395.250 479.700 396.450 487.050 ;
        RECT 397.950 485.850 400.050 487.950 ;
        RECT 409.950 485.850 412.050 487.950 ;
        RECT 412.950 487.050 415.050 489.150 ;
        RECT 398.100 484.050 399.900 485.850 ;
        RECT 410.100 484.050 411.900 485.850 ;
        RECT 413.250 479.700 414.450 487.050 ;
        RECT 415.950 485.850 418.050 487.950 ;
        RECT 430.950 487.050 433.050 489.150 ;
        RECT 434.850 486.150 436.050 491.400 ;
        RECT 440.100 486.150 441.900 487.950 ;
        RECT 416.100 484.050 417.900 485.850 ;
        RECT 433.950 484.050 436.050 486.150 ;
        RECT 433.950 480.750 435.150 484.050 ;
        RECT 436.950 482.850 439.050 484.950 ;
        RECT 439.950 484.050 442.050 486.150 ;
        RECT 452.400 484.950 453.600 497.400 ;
        RECT 466.650 491.400 468.450 503.250 ;
        RECT 469.650 492.300 471.450 503.250 ;
        RECT 472.650 493.200 474.450 503.250 ;
        RECT 475.650 492.300 477.450 503.250 ;
        RECT 491.400 497.400 493.200 503.250 ;
        RECT 469.650 491.400 477.450 492.300 ;
        RECT 494.700 491.400 496.500 503.250 ;
        RECT 498.900 491.400 500.700 503.250 ;
        RECT 512.400 497.400 514.200 503.250 ;
        RECT 515.700 491.400 517.500 503.250 ;
        RECT 519.900 491.400 521.700 503.250 ;
        RECT 531.300 491.400 533.100 503.250 ;
        RECT 535.500 491.400 537.300 503.250 ;
        RECT 538.800 497.400 540.600 503.250 ;
        RECT 557.400 497.400 559.200 503.250 ;
        RECT 560.700 491.400 562.500 503.250 ;
        RECT 564.900 491.400 566.700 503.250 ;
        RECT 579.450 491.400 581.250 503.250 ;
        RECT 583.650 491.400 585.450 503.250 ;
        RECT 597.450 491.400 599.250 503.250 ;
        RECT 601.650 491.400 603.450 503.250 ;
        RECT 611.550 497.400 613.350 503.250 ;
        RECT 614.550 497.400 616.350 503.250 ;
        RECT 467.100 486.150 468.300 491.400 ;
        RECT 491.250 489.150 493.050 490.950 ;
        RECT 490.950 487.050 493.050 489.150 ;
        RECT 494.850 486.150 496.050 491.400 ;
        RECT 512.250 489.150 514.050 490.950 ;
        RECT 500.100 486.150 501.900 487.950 ;
        RECT 511.950 487.050 514.050 489.150 ;
        RECT 515.850 486.150 517.050 491.400 ;
        RECT 521.100 486.150 522.900 487.950 ;
        RECT 530.100 486.150 531.900 487.950 ;
        RECT 535.950 486.150 537.150 491.400 ;
        RECT 538.950 489.150 540.750 490.950 ;
        RECT 557.250 489.150 559.050 490.950 ;
        RECT 538.950 487.050 541.050 489.150 ;
        RECT 556.950 487.050 559.050 489.150 ;
        RECT 560.850 486.150 562.050 491.400 ;
        RECT 579.450 490.350 582.000 491.400 ;
        RECT 597.450 490.350 600.000 491.400 ;
        RECT 566.100 486.150 567.900 487.950 ;
        RECT 578.100 486.150 579.900 487.950 ;
        RECT 451.950 482.850 454.050 484.950 ;
        RECT 455.100 483.150 456.900 484.950 ;
        RECT 466.950 484.050 469.050 486.150 ;
        RECT 437.100 481.050 438.900 482.850 ;
        RECT 319.650 471.750 321.450 477.600 ;
        RECT 322.650 471.750 324.450 477.600 ;
        RECT 335.850 471.750 337.650 478.800 ;
        RECT 353.250 477.600 354.450 479.700 ;
        RECT 374.850 478.800 378.450 479.700 ;
        RECT 392.850 478.800 396.450 479.700 ;
        RECT 410.850 478.800 414.450 479.700 ;
        RECT 431.250 479.700 435.000 480.750 ;
        RECT 340.350 471.750 342.150 477.600 ;
        RECT 352.650 471.750 354.450 477.600 ;
        RECT 355.650 476.700 363.450 478.050 ;
        RECT 355.650 471.750 357.450 476.700 ;
        RECT 358.650 471.750 360.450 475.800 ;
        RECT 361.650 471.750 363.450 476.700 ;
        RECT 374.850 471.750 376.650 478.800 ;
        RECT 379.350 471.750 381.150 477.600 ;
        RECT 392.850 471.750 394.650 478.800 ;
        RECT 397.350 471.750 399.150 477.600 ;
        RECT 410.850 471.750 412.650 478.800 ;
        RECT 431.250 477.600 432.450 479.700 ;
        RECT 415.350 471.750 417.150 477.600 ;
        RECT 430.650 471.750 432.450 477.600 ;
        RECT 433.650 476.700 441.450 478.050 ;
        RECT 433.650 471.750 435.450 476.700 ;
        RECT 436.650 471.750 438.450 475.800 ;
        RECT 439.650 471.750 441.450 476.700 ;
        RECT 452.400 474.600 453.600 482.850 ;
        RECT 454.950 481.050 457.050 483.150 ;
        RECT 467.100 477.600 468.300 484.050 ;
        RECT 469.950 482.850 472.050 484.950 ;
        RECT 473.100 483.150 474.900 484.950 ;
        RECT 470.100 481.050 471.900 482.850 ;
        RECT 472.950 481.050 475.050 483.150 ;
        RECT 475.950 482.850 478.050 484.950 ;
        RECT 493.950 484.050 496.050 486.150 ;
        RECT 476.100 481.050 477.900 482.850 ;
        RECT 493.950 480.750 495.150 484.050 ;
        RECT 496.950 482.850 499.050 484.950 ;
        RECT 499.950 484.050 502.050 486.150 ;
        RECT 514.950 484.050 517.050 486.150 ;
        RECT 497.100 481.050 498.900 482.850 ;
        RECT 514.950 480.750 516.150 484.050 ;
        RECT 517.950 482.850 520.050 484.950 ;
        RECT 520.950 484.050 523.050 486.150 ;
        RECT 529.950 484.050 532.050 486.150 ;
        RECT 532.950 482.850 535.050 484.950 ;
        RECT 535.950 484.050 538.050 486.150 ;
        RECT 518.100 481.050 519.900 482.850 ;
        RECT 533.100 481.050 534.900 482.850 ;
        RECT 536.850 480.750 538.050 484.050 ;
        RECT 559.950 484.050 562.050 486.150 ;
        RECT 559.950 480.750 561.150 484.050 ;
        RECT 562.950 482.850 565.050 484.950 ;
        RECT 565.950 484.050 568.050 486.150 ;
        RECT 577.950 484.050 580.050 486.150 ;
        RECT 580.950 483.150 582.000 490.350 ;
        RECT 584.100 486.150 585.900 487.950 ;
        RECT 596.100 486.150 597.900 487.950 ;
        RECT 583.950 484.050 586.050 486.150 ;
        RECT 595.950 484.050 598.050 486.150 ;
        RECT 598.950 483.150 600.000 490.350 ;
        RECT 602.100 486.150 603.900 487.950 ;
        RECT 601.950 484.050 604.050 486.150 ;
        RECT 614.400 484.950 615.600 497.400 ;
        RECT 620.550 491.400 622.350 503.250 ;
        RECT 623.550 500.400 625.350 503.250 ;
        RECT 628.050 497.400 629.850 503.250 ;
        RECT 632.250 497.400 634.050 503.250 ;
        RECT 625.950 495.300 629.850 497.400 ;
        RECT 636.150 496.500 637.950 503.250 ;
        RECT 639.150 497.400 640.950 503.250 ;
        RECT 643.950 497.400 645.750 503.250 ;
        RECT 649.050 497.400 650.850 503.250 ;
        RECT 644.250 496.500 645.450 497.400 ;
        RECT 634.950 494.700 641.850 496.500 ;
        RECT 644.250 494.400 649.050 496.500 ;
        RECT 627.150 492.600 629.850 494.400 ;
        RECT 630.750 493.800 632.550 494.400 ;
        RECT 630.750 492.900 637.050 493.800 ;
        RECT 644.250 493.500 645.450 494.400 ;
        RECT 630.750 492.600 632.550 492.900 ;
        RECT 628.950 491.700 629.850 492.600 ;
        RECT 611.100 483.150 612.900 484.950 ;
        RECT 563.100 481.050 564.900 482.850 ;
        RECT 580.950 481.050 583.050 483.150 ;
        RECT 598.950 481.050 601.050 483.150 ;
        RECT 610.950 481.050 613.050 483.150 ;
        RECT 613.950 482.850 616.050 484.950 ;
        RECT 491.250 479.700 495.000 480.750 ;
        RECT 512.250 479.700 516.000 480.750 ;
        RECT 537.000 479.700 540.750 480.750 ;
        RECT 491.250 477.600 492.450 479.700 ;
        RECT 467.100 475.950 472.800 477.600 ;
        RECT 451.650 471.750 453.450 474.600 ;
        RECT 454.650 471.750 456.450 474.600 ;
        RECT 467.700 471.750 469.500 474.600 ;
        RECT 471.000 471.750 472.800 475.950 ;
        RECT 475.200 471.750 477.000 477.600 ;
        RECT 490.650 471.750 492.450 477.600 ;
        RECT 493.650 476.700 501.450 478.050 ;
        RECT 512.250 477.600 513.450 479.700 ;
        RECT 493.650 471.750 495.450 476.700 ;
        RECT 496.650 471.750 498.450 475.800 ;
        RECT 499.650 471.750 501.450 476.700 ;
        RECT 511.650 471.750 513.450 477.600 ;
        RECT 514.650 476.700 522.450 478.050 ;
        RECT 514.650 471.750 516.450 476.700 ;
        RECT 517.650 471.750 519.450 475.800 ;
        RECT 520.650 471.750 522.450 476.700 ;
        RECT 530.550 476.700 538.350 478.050 ;
        RECT 530.550 471.750 532.350 476.700 ;
        RECT 533.550 471.750 535.350 475.800 ;
        RECT 536.550 471.750 538.350 476.700 ;
        RECT 539.550 477.600 540.750 479.700 ;
        RECT 557.250 479.700 561.000 480.750 ;
        RECT 557.250 477.600 558.450 479.700 ;
        RECT 539.550 471.750 541.350 477.600 ;
        RECT 556.650 471.750 558.450 477.600 ;
        RECT 559.650 476.700 567.450 478.050 ;
        RECT 559.650 471.750 561.450 476.700 ;
        RECT 562.650 471.750 564.450 475.800 ;
        RECT 565.650 471.750 567.450 476.700 ;
        RECT 580.950 474.600 582.000 481.050 ;
        RECT 598.950 474.600 600.000 481.050 ;
        RECT 614.400 474.600 615.600 482.850 ;
        RECT 620.550 481.950 621.750 491.400 ;
        RECT 625.950 490.800 628.050 491.700 ;
        RECT 628.950 490.800 634.950 491.700 ;
        RECT 623.850 489.600 628.050 490.800 ;
        RECT 622.950 487.800 624.750 489.600 ;
        RECT 634.050 486.150 634.950 490.800 ;
        RECT 636.150 490.800 637.050 492.900 ;
        RECT 637.950 492.300 645.450 493.500 ;
        RECT 637.950 491.700 639.750 492.300 ;
        RECT 652.050 491.400 653.850 503.250 ;
        RECT 667.650 491.400 669.450 503.250 ;
        RECT 670.650 492.300 672.450 503.250 ;
        RECT 673.650 493.200 675.450 503.250 ;
        RECT 676.650 492.300 678.450 503.250 ;
        RECT 688.650 497.400 690.450 503.250 ;
        RECT 691.650 497.400 693.450 503.250 ;
        RECT 670.650 491.400 678.450 492.300 ;
        RECT 642.750 490.800 653.850 491.400 ;
        RECT 636.150 490.200 653.850 490.800 ;
        RECT 636.150 489.900 644.550 490.200 ;
        RECT 642.750 489.600 644.550 489.900 ;
        RECT 634.050 484.050 637.050 486.150 ;
        RECT 640.950 485.100 643.050 486.150 ;
        RECT 640.950 484.050 648.900 485.100 ;
        RECT 622.950 483.750 625.050 484.050 ;
        RECT 622.950 481.950 626.850 483.750 ;
        RECT 620.550 479.850 625.050 481.950 ;
        RECT 634.050 480.000 634.950 484.050 ;
        RECT 647.100 483.300 648.900 484.050 ;
        RECT 650.100 483.150 651.900 484.950 ;
        RECT 644.100 482.400 645.900 483.000 ;
        RECT 650.100 482.400 651.000 483.150 ;
        RECT 644.100 481.200 651.000 482.400 ;
        RECT 644.100 480.000 645.150 481.200 ;
        RECT 620.550 477.600 621.750 479.850 ;
        RECT 634.050 479.100 645.150 480.000 ;
        RECT 634.050 478.800 634.950 479.100 ;
        RECT 577.650 471.750 579.450 474.600 ;
        RECT 580.650 471.750 582.450 474.600 ;
        RECT 583.650 471.750 585.450 474.600 ;
        RECT 595.650 471.750 597.450 474.600 ;
        RECT 598.650 471.750 600.450 474.600 ;
        RECT 601.650 471.750 603.450 474.600 ;
        RECT 611.550 471.750 613.350 474.600 ;
        RECT 614.550 471.750 616.350 474.600 ;
        RECT 620.550 471.750 622.350 477.600 ;
        RECT 625.950 476.700 628.050 477.600 ;
        RECT 633.150 477.000 634.950 478.800 ;
        RECT 644.100 478.200 645.150 479.100 ;
        RECT 640.350 477.450 642.150 478.200 ;
        RECT 625.950 475.500 629.700 476.700 ;
        RECT 628.650 474.600 629.700 475.500 ;
        RECT 637.200 476.400 642.150 477.450 ;
        RECT 643.650 476.400 645.450 478.200 ;
        RECT 652.950 477.600 653.850 490.200 ;
        RECT 668.100 486.150 669.300 491.400 ;
        RECT 667.950 484.050 670.050 486.150 ;
        RECT 689.400 484.950 690.600 497.400 ;
        RECT 702.300 491.400 704.100 503.250 ;
        RECT 706.500 491.400 708.300 503.250 ;
        RECT 709.800 497.400 711.600 503.250 ;
        RECT 725.550 497.400 727.350 503.250 ;
        RECT 728.550 497.400 730.350 503.250 ;
        RECT 746.400 497.400 748.200 503.250 ;
        RECT 701.100 486.150 702.900 487.950 ;
        RECT 706.950 486.150 708.150 491.400 ;
        RECT 709.950 489.150 711.750 490.950 ;
        RECT 709.950 487.050 712.050 489.150 ;
        RECT 637.200 474.600 638.250 476.400 ;
        RECT 646.950 475.500 649.050 477.600 ;
        RECT 646.950 474.600 648.000 475.500 ;
        RECT 623.850 471.750 625.650 474.600 ;
        RECT 628.350 471.750 630.150 474.600 ;
        RECT 632.550 471.750 634.350 474.600 ;
        RECT 636.450 471.750 638.250 474.600 ;
        RECT 639.750 471.750 641.550 474.600 ;
        RECT 644.250 473.700 648.000 474.600 ;
        RECT 644.250 471.750 646.050 473.700 ;
        RECT 649.050 471.750 650.850 474.600 ;
        RECT 652.050 471.750 653.850 477.600 ;
        RECT 668.100 477.600 669.300 484.050 ;
        RECT 670.950 482.850 673.050 484.950 ;
        RECT 674.100 483.150 675.900 484.950 ;
        RECT 671.100 481.050 672.900 482.850 ;
        RECT 673.950 481.050 676.050 483.150 ;
        RECT 676.950 482.850 679.050 484.950 ;
        RECT 688.950 482.850 691.050 484.950 ;
        RECT 692.100 483.150 693.900 484.950 ;
        RECT 700.950 484.050 703.050 486.150 ;
        RECT 677.100 481.050 678.900 482.850 ;
        RECT 668.100 475.950 673.800 477.600 ;
        RECT 668.700 471.750 670.500 474.600 ;
        RECT 672.000 471.750 673.800 475.950 ;
        RECT 676.200 471.750 678.000 477.600 ;
        RECT 689.400 474.600 690.600 482.850 ;
        RECT 691.950 481.050 694.050 483.150 ;
        RECT 703.950 482.850 706.050 484.950 ;
        RECT 706.950 484.050 709.050 486.150 ;
        RECT 728.400 484.950 729.600 497.400 ;
        RECT 749.700 491.400 751.500 503.250 ;
        RECT 753.900 491.400 755.700 503.250 ;
        RECT 765.300 491.400 767.100 503.250 ;
        RECT 769.500 491.400 771.300 503.250 ;
        RECT 772.800 497.400 774.600 503.250 ;
        RECT 786.300 491.400 788.100 503.250 ;
        RECT 790.500 491.400 792.300 503.250 ;
        RECT 793.800 497.400 795.600 503.250 ;
        RECT 801.150 491.400 802.950 503.250 ;
        RECT 804.150 497.400 805.950 503.250 ;
        RECT 809.250 497.400 811.050 503.250 ;
        RECT 814.050 497.400 815.850 503.250 ;
        RECT 809.550 496.500 810.750 497.400 ;
        RECT 817.050 496.500 818.850 503.250 ;
        RECT 820.950 497.400 822.750 503.250 ;
        RECT 825.150 497.400 826.950 503.250 ;
        RECT 829.650 500.400 831.450 503.250 ;
        RECT 805.950 494.400 810.750 496.500 ;
        RECT 813.150 494.700 820.050 496.500 ;
        RECT 825.150 495.300 829.050 497.400 ;
        RECT 809.550 493.500 810.750 494.400 ;
        RECT 822.450 493.800 824.250 494.400 ;
        RECT 809.550 492.300 817.050 493.500 ;
        RECT 815.250 491.700 817.050 492.300 ;
        RECT 817.950 492.900 824.250 493.800 ;
        RECT 746.250 489.150 748.050 490.950 ;
        RECT 745.950 487.050 748.050 489.150 ;
        RECT 749.850 486.150 751.050 491.400 ;
        RECT 755.100 486.150 756.900 487.950 ;
        RECT 764.100 486.150 765.900 487.950 ;
        RECT 769.950 486.150 771.150 491.400 ;
        RECT 772.950 489.150 774.750 490.950 ;
        RECT 772.950 487.050 775.050 489.150 ;
        RECT 785.100 486.150 786.900 487.950 ;
        RECT 790.950 486.150 792.150 491.400 ;
        RECT 793.950 489.150 795.750 490.950 ;
        RECT 801.150 490.800 812.250 491.400 ;
        RECT 817.950 490.800 818.850 492.900 ;
        RECT 822.450 492.600 824.250 492.900 ;
        RECT 825.150 492.600 827.850 494.400 ;
        RECT 825.150 491.700 826.050 492.600 ;
        RECT 801.150 490.200 818.850 490.800 ;
        RECT 793.950 487.050 796.050 489.150 ;
        RECT 704.100 481.050 705.900 482.850 ;
        RECT 707.850 480.750 709.050 484.050 ;
        RECT 725.100 483.150 726.900 484.950 ;
        RECT 724.950 481.050 727.050 483.150 ;
        RECT 727.950 482.850 730.050 484.950 ;
        RECT 748.950 484.050 751.050 486.150 ;
        RECT 708.000 479.700 711.750 480.750 ;
        RECT 701.550 476.700 709.350 478.050 ;
        RECT 688.650 471.750 690.450 474.600 ;
        RECT 691.650 471.750 693.450 474.600 ;
        RECT 701.550 471.750 703.350 476.700 ;
        RECT 704.550 471.750 706.350 475.800 ;
        RECT 707.550 471.750 709.350 476.700 ;
        RECT 710.550 477.600 711.750 479.700 ;
        RECT 710.550 471.750 712.350 477.600 ;
        RECT 728.400 474.600 729.600 482.850 ;
        RECT 748.950 480.750 750.150 484.050 ;
        RECT 751.950 482.850 754.050 484.950 ;
        RECT 754.950 484.050 757.050 486.150 ;
        RECT 763.950 484.050 766.050 486.150 ;
        RECT 766.950 482.850 769.050 484.950 ;
        RECT 769.950 484.050 772.050 486.150 ;
        RECT 784.950 484.050 787.050 486.150 ;
        RECT 752.100 481.050 753.900 482.850 ;
        RECT 767.100 481.050 768.900 482.850 ;
        RECT 770.850 480.750 772.050 484.050 ;
        RECT 787.950 482.850 790.050 484.950 ;
        RECT 790.950 484.050 793.050 486.150 ;
        RECT 788.100 481.050 789.900 482.850 ;
        RECT 791.850 480.750 793.050 484.050 ;
        RECT 746.250 479.700 750.000 480.750 ;
        RECT 771.000 479.700 774.750 480.750 ;
        RECT 792.000 479.700 795.750 480.750 ;
        RECT 746.250 477.600 747.450 479.700 ;
        RECT 725.550 471.750 727.350 474.600 ;
        RECT 728.550 471.750 730.350 474.600 ;
        RECT 745.650 471.750 747.450 477.600 ;
        RECT 748.650 476.700 756.450 478.050 ;
        RECT 748.650 471.750 750.450 476.700 ;
        RECT 751.650 471.750 753.450 475.800 ;
        RECT 754.650 471.750 756.450 476.700 ;
        RECT 764.550 476.700 772.350 478.050 ;
        RECT 764.550 471.750 766.350 476.700 ;
        RECT 767.550 471.750 769.350 475.800 ;
        RECT 770.550 471.750 772.350 476.700 ;
        RECT 773.550 477.600 774.750 479.700 ;
        RECT 773.550 471.750 775.350 477.600 ;
        RECT 785.550 476.700 793.350 478.050 ;
        RECT 785.550 471.750 787.350 476.700 ;
        RECT 788.550 471.750 790.350 475.800 ;
        RECT 791.550 471.750 793.350 476.700 ;
        RECT 794.550 477.600 795.750 479.700 ;
        RECT 801.150 477.600 802.050 490.200 ;
        RECT 810.450 489.900 818.850 490.200 ;
        RECT 820.050 490.800 826.050 491.700 ;
        RECT 826.950 490.800 829.050 491.700 ;
        RECT 832.650 491.400 834.450 503.250 ;
        RECT 845.550 497.400 847.350 503.250 ;
        RECT 848.550 497.400 850.350 503.250 ;
        RECT 851.550 497.400 853.350 503.250 ;
        RECT 863.550 497.400 865.350 503.250 ;
        RECT 866.550 497.400 868.350 503.250 ;
        RECT 869.550 497.400 871.350 503.250 ;
        RECT 810.450 489.600 812.250 489.900 ;
        RECT 820.050 486.150 820.950 490.800 ;
        RECT 826.950 489.600 831.150 490.800 ;
        RECT 830.250 487.800 832.050 489.600 ;
        RECT 811.950 485.100 814.050 486.150 ;
        RECT 803.100 483.150 804.900 484.950 ;
        RECT 806.100 484.050 814.050 485.100 ;
        RECT 817.950 484.050 820.950 486.150 ;
        RECT 806.100 483.300 807.900 484.050 ;
        RECT 804.000 482.400 804.900 483.150 ;
        RECT 809.100 482.400 810.900 483.000 ;
        RECT 804.000 481.200 810.900 482.400 ;
        RECT 809.850 480.000 810.900 481.200 ;
        RECT 820.050 480.000 820.950 484.050 ;
        RECT 829.950 483.750 832.050 484.050 ;
        RECT 828.150 481.950 832.050 483.750 ;
        RECT 833.250 481.950 834.450 491.400 ;
        RECT 848.550 489.150 849.750 497.400 ;
        RECT 866.550 489.150 867.750 497.400 ;
        RECT 844.950 485.850 847.050 487.950 ;
        RECT 847.950 487.050 850.050 489.150 ;
        RECT 845.100 484.050 846.900 485.850 ;
        RECT 809.850 479.100 820.950 480.000 ;
        RECT 829.950 479.850 834.450 481.950 ;
        RECT 809.850 478.200 810.900 479.100 ;
        RECT 820.050 478.800 820.950 479.100 ;
        RECT 794.550 471.750 796.350 477.600 ;
        RECT 801.150 471.750 802.950 477.600 ;
        RECT 805.950 475.500 808.050 477.600 ;
        RECT 809.550 476.400 811.350 478.200 ;
        RECT 812.850 477.450 814.650 478.200 ;
        RECT 812.850 476.400 817.800 477.450 ;
        RECT 820.050 477.000 821.850 478.800 ;
        RECT 833.250 477.600 834.450 479.850 ;
        RECT 848.550 479.700 849.750 487.050 ;
        RECT 850.950 485.850 853.050 487.950 ;
        RECT 862.950 485.850 865.050 487.950 ;
        RECT 865.950 487.050 868.050 489.150 ;
        RECT 851.100 484.050 852.900 485.850 ;
        RECT 863.100 484.050 864.900 485.850 ;
        RECT 866.550 479.700 867.750 487.050 ;
        RECT 868.950 485.850 871.050 487.950 ;
        RECT 869.100 484.050 870.900 485.850 ;
        RECT 848.550 478.800 852.150 479.700 ;
        RECT 866.550 478.800 870.150 479.700 ;
        RECT 826.950 476.700 829.050 477.600 ;
        RECT 807.000 474.600 808.050 475.500 ;
        RECT 816.750 474.600 817.800 476.400 ;
        RECT 825.300 475.500 829.050 476.700 ;
        RECT 825.300 474.600 826.350 475.500 ;
        RECT 804.150 471.750 805.950 474.600 ;
        RECT 807.000 473.700 810.750 474.600 ;
        RECT 808.950 471.750 810.750 473.700 ;
        RECT 813.450 471.750 815.250 474.600 ;
        RECT 816.750 471.750 818.550 474.600 ;
        RECT 820.650 471.750 822.450 474.600 ;
        RECT 824.850 471.750 826.650 474.600 ;
        RECT 829.350 471.750 831.150 474.600 ;
        RECT 832.650 471.750 834.450 477.600 ;
        RECT 845.850 471.750 847.650 477.600 ;
        RECT 850.350 471.750 852.150 478.800 ;
        RECT 863.850 471.750 865.650 477.600 ;
        RECT 868.350 471.750 870.150 478.800 ;
        RECT 8.550 462.300 10.350 467.250 ;
        RECT 11.550 463.200 13.350 467.250 ;
        RECT 14.550 462.300 16.350 467.250 ;
        RECT 8.550 460.950 16.350 462.300 ;
        RECT 17.550 461.400 19.350 467.250 ;
        RECT 17.550 459.300 18.750 461.400 ;
        RECT 15.000 458.250 18.750 459.300 ;
        RECT 32.550 459.900 34.350 467.250 ;
        RECT 37.050 461.400 38.850 467.250 ;
        RECT 40.050 462.900 41.850 467.250 ;
        RECT 55.650 464.400 57.450 467.250 ;
        RECT 58.650 464.400 60.450 467.250 ;
        RECT 40.050 461.400 43.350 462.900 ;
        RECT 38.250 459.900 40.050 460.500 ;
        RECT 32.550 458.700 40.050 459.900 ;
        RECT 11.100 456.150 12.900 457.950 ;
        RECT 7.950 452.850 10.050 454.950 ;
        RECT 10.950 454.050 13.050 456.150 ;
        RECT 14.850 454.950 16.050 458.250 ;
        RECT 13.950 452.850 16.050 454.950 ;
        RECT 31.950 452.850 34.050 454.950 ;
        RECT 8.100 451.050 9.900 452.850 ;
        RECT 13.950 447.600 15.150 452.850 ;
        RECT 16.950 449.850 19.050 451.950 ;
        RECT 32.100 451.050 33.900 452.850 ;
        RECT 16.950 448.050 18.750 449.850 ;
        RECT 9.300 435.750 11.100 447.600 ;
        RECT 13.500 435.750 15.300 447.600 ;
        RECT 35.700 441.600 36.900 458.700 ;
        RECT 42.150 454.950 43.350 461.400 ;
        RECT 56.400 456.150 57.600 464.400 ;
        RECT 62.550 461.400 64.350 467.250 ;
        RECT 65.850 464.400 67.650 467.250 ;
        RECT 70.350 464.400 72.150 467.250 ;
        RECT 74.550 464.400 76.350 467.250 ;
        RECT 78.450 464.400 80.250 467.250 ;
        RECT 81.750 464.400 83.550 467.250 ;
        RECT 86.250 465.300 88.050 467.250 ;
        RECT 86.250 464.400 90.000 465.300 ;
        RECT 91.050 464.400 92.850 467.250 ;
        RECT 70.650 463.500 71.700 464.400 ;
        RECT 67.950 462.300 71.700 463.500 ;
        RECT 79.200 462.600 80.250 464.400 ;
        RECT 88.950 463.500 90.000 464.400 ;
        RECT 67.950 461.400 70.050 462.300 ;
        RECT 62.550 459.150 63.750 461.400 ;
        RECT 75.150 460.200 76.950 462.000 ;
        RECT 79.200 461.550 84.150 462.600 ;
        RECT 82.350 460.800 84.150 461.550 ;
        RECT 85.650 460.800 87.450 462.600 ;
        RECT 88.950 461.400 91.050 463.500 ;
        RECT 94.050 461.400 95.850 467.250 ;
        RECT 76.050 459.900 76.950 460.200 ;
        RECT 86.100 459.900 87.150 460.800 ;
        RECT 38.100 453.150 39.900 454.950 ;
        RECT 37.950 451.050 40.050 453.150 ;
        RECT 40.950 452.850 43.350 454.950 ;
        RECT 55.950 454.050 58.050 456.150 ;
        RECT 58.950 455.850 61.050 457.950 ;
        RECT 62.550 457.050 67.050 459.150 ;
        RECT 76.050 459.000 87.150 459.900 ;
        RECT 59.100 454.050 60.900 455.850 ;
        RECT 42.150 447.600 43.350 452.850 ;
        RECT 16.800 435.750 18.600 441.600 ;
        RECT 32.550 435.750 34.350 441.600 ;
        RECT 35.550 435.750 37.350 441.600 ;
        RECT 39.150 435.750 40.950 447.600 ;
        RECT 42.150 435.750 43.950 447.600 ;
        RECT 56.400 441.600 57.600 454.050 ;
        RECT 62.550 447.600 63.750 457.050 ;
        RECT 64.950 455.250 68.850 457.050 ;
        RECT 64.950 454.950 67.050 455.250 ;
        RECT 76.050 454.950 76.950 459.000 ;
        RECT 86.100 457.800 87.150 459.000 ;
        RECT 86.100 456.600 93.000 457.800 ;
        RECT 86.100 456.000 87.900 456.600 ;
        RECT 92.100 455.850 93.000 456.600 ;
        RECT 89.100 454.950 90.900 455.700 ;
        RECT 76.050 452.850 79.050 454.950 ;
        RECT 82.950 453.900 90.900 454.950 ;
        RECT 92.100 454.050 93.900 455.850 ;
        RECT 82.950 452.850 85.050 453.900 ;
        RECT 64.950 449.400 66.750 451.200 ;
        RECT 65.850 448.200 70.050 449.400 ;
        RECT 76.050 448.200 76.950 452.850 ;
        RECT 84.750 449.100 86.550 449.400 ;
        RECT 55.650 435.750 57.450 441.600 ;
        RECT 58.650 435.750 60.450 441.600 ;
        RECT 62.550 435.750 64.350 447.600 ;
        RECT 67.950 447.300 70.050 448.200 ;
        RECT 70.950 447.300 76.950 448.200 ;
        RECT 78.150 448.800 86.550 449.100 ;
        RECT 94.950 448.800 95.850 461.400 ;
        RECT 107.550 462.300 109.350 467.250 ;
        RECT 110.550 463.200 112.350 467.250 ;
        RECT 113.550 462.300 115.350 467.250 ;
        RECT 107.550 460.950 115.350 462.300 ;
        RECT 116.550 461.400 118.350 467.250 ;
        RECT 128.850 461.400 130.650 467.250 ;
        RECT 116.550 459.300 117.750 461.400 ;
        RECT 133.350 460.200 135.150 467.250 ;
        RECT 151.350 461.400 153.150 467.250 ;
        RECT 154.350 461.400 156.150 467.250 ;
        RECT 157.650 464.400 159.450 467.250 ;
        RECT 114.000 458.250 117.750 459.300 ;
        RECT 131.550 459.300 135.150 460.200 ;
        RECT 110.100 456.150 111.900 457.950 ;
        RECT 106.950 452.850 109.050 454.950 ;
        RECT 109.950 454.050 112.050 456.150 ;
        RECT 113.850 454.950 115.050 458.250 ;
        RECT 112.950 452.850 115.050 454.950 ;
        RECT 128.100 453.150 129.900 454.950 ;
        RECT 107.100 451.050 108.900 452.850 ;
        RECT 78.150 448.200 95.850 448.800 ;
        RECT 70.950 446.400 71.850 447.300 ;
        RECT 69.150 444.600 71.850 446.400 ;
        RECT 72.750 446.100 74.550 446.400 ;
        RECT 78.150 446.100 79.050 448.200 ;
        RECT 84.750 447.600 95.850 448.200 ;
        RECT 112.950 447.600 114.150 452.850 ;
        RECT 115.950 449.850 118.050 451.950 ;
        RECT 127.950 451.050 130.050 453.150 ;
        RECT 131.550 451.950 132.750 459.300 ;
        RECT 151.650 454.950 152.850 461.400 ;
        RECT 157.650 460.500 158.850 464.400 ;
        RECT 153.750 459.600 158.850 460.500 ;
        RECT 169.650 460.200 171.450 467.250 ;
        RECT 174.150 461.700 175.950 466.200 ;
        RECT 178.650 463.200 180.450 467.250 ;
        RECT 181.650 463.200 183.450 466.200 ;
        RECT 191.550 464.400 193.350 467.250 ;
        RECT 194.550 464.400 196.350 467.250 ;
        RECT 173.850 460.800 175.950 461.700 ;
        RECT 153.750 458.700 156.000 459.600 ;
        RECT 134.100 453.150 135.900 454.950 ;
        RECT 130.950 449.850 133.050 451.950 ;
        RECT 133.950 451.050 136.050 453.150 ;
        RECT 151.650 452.850 154.050 454.950 ;
        RECT 115.950 448.050 117.750 449.850 ;
        RECT 72.750 445.200 79.050 446.100 ;
        RECT 79.950 446.700 81.750 447.300 ;
        RECT 79.950 445.500 87.450 446.700 ;
        RECT 72.750 444.600 74.550 445.200 ;
        RECT 86.250 444.600 87.450 445.500 ;
        RECT 67.950 441.600 71.850 443.700 ;
        RECT 76.950 442.500 83.850 444.300 ;
        RECT 86.250 442.500 91.050 444.600 ;
        RECT 65.550 435.750 67.350 438.600 ;
        RECT 70.050 435.750 71.850 441.600 ;
        RECT 74.250 435.750 76.050 441.600 ;
        RECT 78.150 435.750 79.950 442.500 ;
        RECT 86.250 441.600 87.450 442.500 ;
        RECT 81.150 435.750 82.950 441.600 ;
        RECT 85.950 435.750 87.750 441.600 ;
        RECT 91.050 435.750 92.850 441.600 ;
        RECT 94.050 435.750 95.850 447.600 ;
        RECT 108.300 435.750 110.100 447.600 ;
        RECT 112.500 435.750 114.300 447.600 ;
        RECT 131.550 441.600 132.750 449.850 ;
        RECT 151.650 447.600 152.850 452.850 ;
        RECT 154.950 450.300 156.000 458.700 ;
        RECT 173.850 456.150 174.750 460.800 ;
        RECT 181.650 459.900 182.700 463.200 ;
        RECT 176.400 459.000 182.700 459.900 ;
        RECT 157.950 452.850 160.050 454.950 ;
        RECT 169.950 452.850 172.050 454.950 ;
        RECT 172.950 454.050 175.050 456.150 ;
        RECT 158.100 451.050 159.900 452.850 ;
        RECT 170.100 451.050 171.900 452.850 ;
        RECT 153.750 449.400 156.000 450.300 ;
        RECT 153.750 448.500 159.450 449.400 ;
        RECT 115.800 435.750 117.600 441.600 ;
        RECT 128.550 435.750 130.350 441.600 ;
        RECT 131.550 435.750 133.350 441.600 ;
        RECT 134.550 435.750 136.350 441.600 ;
        RECT 151.350 435.750 153.150 447.600 ;
        RECT 154.350 435.750 156.150 447.600 ;
        RECT 158.250 441.600 159.450 448.500 ;
        RECT 157.650 435.750 159.450 441.600 ;
        RECT 169.650 435.750 171.450 447.600 ;
        RECT 173.850 447.000 174.750 454.050 ;
        RECT 176.400 453.300 177.750 459.000 ;
        RECT 181.950 456.150 183.750 457.950 ;
        RECT 175.950 451.500 177.750 453.300 ;
        RECT 176.400 448.800 177.750 451.500 ;
        RECT 178.950 452.850 181.050 454.950 ;
        RECT 181.950 454.050 184.050 456.150 ;
        RECT 190.950 455.850 193.050 457.950 ;
        RECT 194.400 456.150 195.600 464.400 ;
        RECT 209.550 462.300 211.350 467.250 ;
        RECT 212.550 463.200 214.350 467.250 ;
        RECT 215.550 462.300 217.350 467.250 ;
        RECT 209.550 460.950 217.350 462.300 ;
        RECT 218.550 461.400 220.350 467.250 ;
        RECT 230.850 461.400 232.650 467.250 ;
        RECT 218.550 459.300 219.750 461.400 ;
        RECT 235.350 460.200 237.150 467.250 ;
        RECT 253.650 460.200 255.450 467.250 ;
        RECT 258.150 461.700 259.950 466.200 ;
        RECT 262.650 463.200 264.450 467.250 ;
        RECT 265.650 463.200 267.450 466.200 ;
        RECT 275.550 464.400 277.350 467.250 ;
        RECT 257.850 460.800 259.950 461.700 ;
        RECT 216.000 458.250 219.750 459.300 ;
        RECT 233.550 459.300 237.150 460.200 ;
        RECT 212.100 456.150 213.900 457.950 ;
        RECT 191.100 454.050 192.900 455.850 ;
        RECT 193.950 454.050 196.050 456.150 ;
        RECT 178.950 451.050 180.750 452.850 ;
        RECT 176.400 447.900 182.550 448.800 ;
        RECT 173.850 446.100 175.950 447.000 ;
        RECT 174.150 436.800 175.950 446.100 ;
        RECT 181.650 442.800 182.550 447.900 ;
        RECT 178.650 435.750 180.450 442.800 ;
        RECT 181.650 436.800 183.450 442.800 ;
        RECT 194.400 441.600 195.600 454.050 ;
        RECT 208.950 452.850 211.050 454.950 ;
        RECT 211.950 454.050 214.050 456.150 ;
        RECT 215.850 454.950 217.050 458.250 ;
        RECT 214.950 452.850 217.050 454.950 ;
        RECT 230.100 453.150 231.900 454.950 ;
        RECT 209.100 451.050 210.900 452.850 ;
        RECT 214.950 447.600 216.150 452.850 ;
        RECT 217.950 449.850 220.050 451.950 ;
        RECT 229.950 451.050 232.050 453.150 ;
        RECT 233.550 451.950 234.750 459.300 ;
        RECT 257.850 456.150 258.750 460.800 ;
        RECT 265.650 459.900 266.700 463.200 ;
        RECT 260.400 459.000 266.700 459.900 ;
        RECT 276.150 460.500 277.350 464.400 ;
        RECT 278.850 461.400 280.650 467.250 ;
        RECT 281.850 461.400 283.650 467.250 ;
        RECT 276.150 459.600 281.250 460.500 ;
        RECT 236.100 453.150 237.900 454.950 ;
        RECT 232.950 449.850 235.050 451.950 ;
        RECT 235.950 451.050 238.050 453.150 ;
        RECT 253.950 452.850 256.050 454.950 ;
        RECT 256.950 454.050 259.050 456.150 ;
        RECT 254.100 451.050 255.900 452.850 ;
        RECT 217.950 448.050 219.750 449.850 ;
        RECT 191.550 435.750 193.350 441.600 ;
        RECT 194.550 435.750 196.350 441.600 ;
        RECT 210.300 435.750 212.100 447.600 ;
        RECT 214.500 435.750 216.300 447.600 ;
        RECT 233.550 441.600 234.750 449.850 ;
        RECT 217.800 435.750 219.600 441.600 ;
        RECT 230.550 435.750 232.350 441.600 ;
        RECT 233.550 435.750 235.350 441.600 ;
        RECT 236.550 435.750 238.350 441.600 ;
        RECT 253.650 435.750 255.450 447.600 ;
        RECT 257.850 447.000 258.750 454.050 ;
        RECT 260.400 453.300 261.750 459.000 ;
        RECT 279.000 458.700 281.250 459.600 ;
        RECT 265.950 456.150 267.750 457.950 ;
        RECT 259.950 451.500 261.750 453.300 ;
        RECT 260.400 448.800 261.750 451.500 ;
        RECT 262.950 452.850 265.050 454.950 ;
        RECT 265.950 454.050 268.050 456.150 ;
        RECT 274.950 452.850 277.050 454.950 ;
        RECT 262.950 451.050 264.750 452.850 ;
        RECT 275.100 451.050 276.900 452.850 ;
        RECT 279.000 450.300 280.050 458.700 ;
        RECT 282.150 454.950 283.350 461.400 ;
        RECT 299.850 460.200 301.650 467.250 ;
        RECT 304.350 461.400 306.150 467.250 ;
        RECT 319.650 460.200 321.450 467.250 ;
        RECT 324.150 461.700 325.950 466.200 ;
        RECT 328.650 463.200 330.450 467.250 ;
        RECT 331.650 463.200 333.450 466.200 ;
        RECT 323.850 460.800 325.950 461.700 ;
        RECT 299.850 459.300 303.450 460.200 ;
        RECT 280.950 452.850 283.350 454.950 ;
        RECT 299.100 453.150 300.900 454.950 ;
        RECT 279.000 449.400 281.250 450.300 ;
        RECT 260.400 447.900 266.550 448.800 ;
        RECT 257.850 446.100 259.950 447.000 ;
        RECT 258.150 436.800 259.950 446.100 ;
        RECT 265.650 442.800 266.550 447.900 ;
        RECT 275.550 448.500 281.250 449.400 ;
        RECT 262.650 435.750 264.450 442.800 ;
        RECT 265.650 436.800 267.450 442.800 ;
        RECT 275.550 441.600 276.750 448.500 ;
        RECT 282.150 447.600 283.350 452.850 ;
        RECT 298.950 451.050 301.050 453.150 ;
        RECT 302.250 451.950 303.450 459.300 ;
        RECT 323.850 456.150 324.750 460.800 ;
        RECT 331.650 459.900 332.700 463.200 ;
        RECT 341.550 462.300 343.350 467.250 ;
        RECT 344.550 463.200 346.350 467.250 ;
        RECT 347.550 462.300 349.350 467.250 ;
        RECT 341.550 460.950 349.350 462.300 ;
        RECT 350.550 461.400 352.350 467.250 ;
        RECT 356.550 461.400 358.350 467.250 ;
        RECT 359.850 464.400 361.650 467.250 ;
        RECT 364.350 464.400 366.150 467.250 ;
        RECT 368.550 464.400 370.350 467.250 ;
        RECT 372.450 464.400 374.250 467.250 ;
        RECT 375.750 464.400 377.550 467.250 ;
        RECT 380.250 465.300 382.050 467.250 ;
        RECT 380.250 464.400 384.000 465.300 ;
        RECT 385.050 464.400 386.850 467.250 ;
        RECT 364.650 463.500 365.700 464.400 ;
        RECT 361.950 462.300 365.700 463.500 ;
        RECT 373.200 462.600 374.250 464.400 ;
        RECT 382.950 463.500 384.000 464.400 ;
        RECT 361.950 461.400 364.050 462.300 ;
        RECT 326.400 459.000 332.700 459.900 ;
        RECT 350.550 459.300 351.750 461.400 ;
        RECT 305.100 453.150 306.900 454.950 ;
        RECT 301.950 449.850 304.050 451.950 ;
        RECT 304.950 451.050 307.050 453.150 ;
        RECT 319.950 452.850 322.050 454.950 ;
        RECT 322.950 454.050 325.050 456.150 ;
        RECT 320.100 451.050 321.900 452.850 ;
        RECT 275.550 435.750 277.350 441.600 ;
        RECT 278.850 435.750 280.650 447.600 ;
        RECT 281.850 435.750 283.650 447.600 ;
        RECT 302.250 441.600 303.450 449.850 ;
        RECT 298.650 435.750 300.450 441.600 ;
        RECT 301.650 435.750 303.450 441.600 ;
        RECT 304.650 435.750 306.450 441.600 ;
        RECT 319.650 435.750 321.450 447.600 ;
        RECT 323.850 447.000 324.750 454.050 ;
        RECT 326.400 453.300 327.750 459.000 ;
        RECT 348.000 458.250 351.750 459.300 ;
        RECT 356.550 459.150 357.750 461.400 ;
        RECT 369.150 460.200 370.950 462.000 ;
        RECT 373.200 461.550 378.150 462.600 ;
        RECT 376.350 460.800 378.150 461.550 ;
        RECT 379.650 460.800 381.450 462.600 ;
        RECT 382.950 461.400 385.050 463.500 ;
        RECT 388.050 461.400 389.850 467.250 ;
        RECT 370.050 459.900 370.950 460.200 ;
        RECT 380.100 459.900 381.150 460.800 ;
        RECT 331.950 456.150 333.750 457.950 ;
        RECT 344.100 456.150 345.900 457.950 ;
        RECT 325.950 451.500 327.750 453.300 ;
        RECT 326.400 448.800 327.750 451.500 ;
        RECT 328.950 452.850 331.050 454.950 ;
        RECT 331.950 454.050 334.050 456.150 ;
        RECT 340.950 452.850 343.050 454.950 ;
        RECT 343.950 454.050 346.050 456.150 ;
        RECT 347.850 454.950 349.050 458.250 ;
        RECT 346.950 452.850 349.050 454.950 ;
        RECT 356.550 457.050 361.050 459.150 ;
        RECT 370.050 459.000 381.150 459.900 ;
        RECT 328.950 451.050 330.750 452.850 ;
        RECT 341.100 451.050 342.900 452.850 ;
        RECT 326.400 447.900 332.550 448.800 ;
        RECT 323.850 446.100 325.950 447.000 ;
        RECT 324.150 436.800 325.950 446.100 ;
        RECT 331.650 442.800 332.550 447.900 ;
        RECT 346.950 447.600 348.150 452.850 ;
        RECT 349.950 449.850 352.050 451.950 ;
        RECT 349.950 448.050 351.750 449.850 ;
        RECT 356.550 447.600 357.750 457.050 ;
        RECT 358.950 455.250 362.850 457.050 ;
        RECT 358.950 454.950 361.050 455.250 ;
        RECT 370.050 454.950 370.950 459.000 ;
        RECT 380.100 457.800 381.150 459.000 ;
        RECT 380.100 456.600 387.000 457.800 ;
        RECT 380.100 456.000 381.900 456.600 ;
        RECT 386.100 455.850 387.000 456.600 ;
        RECT 383.100 454.950 384.900 455.700 ;
        RECT 370.050 452.850 373.050 454.950 ;
        RECT 376.950 453.900 384.900 454.950 ;
        RECT 386.100 454.050 387.900 455.850 ;
        RECT 376.950 452.850 379.050 453.900 ;
        RECT 358.950 449.400 360.750 451.200 ;
        RECT 359.850 448.200 364.050 449.400 ;
        RECT 370.050 448.200 370.950 452.850 ;
        RECT 378.750 449.100 380.550 449.400 ;
        RECT 328.650 435.750 330.450 442.800 ;
        RECT 331.650 436.800 333.450 442.800 ;
        RECT 342.300 435.750 344.100 447.600 ;
        RECT 346.500 435.750 348.300 447.600 ;
        RECT 349.800 435.750 351.600 441.600 ;
        RECT 356.550 435.750 358.350 447.600 ;
        RECT 361.950 447.300 364.050 448.200 ;
        RECT 364.950 447.300 370.950 448.200 ;
        RECT 372.150 448.800 380.550 449.100 ;
        RECT 388.950 448.800 389.850 461.400 ;
        RECT 401.700 458.400 403.500 467.250 ;
        RECT 407.100 459.000 408.900 467.250 ;
        RECT 422.850 461.400 424.650 467.250 ;
        RECT 427.350 460.200 429.150 467.250 ;
        RECT 425.550 459.300 429.150 460.200 ;
        RECT 443.850 460.200 445.650 467.250 ;
        RECT 448.350 461.400 450.150 467.250 ;
        RECT 463.650 461.400 465.450 467.250 ;
        RECT 443.850 459.300 447.450 460.200 ;
        RECT 407.100 457.350 411.600 459.000 ;
        RECT 410.400 453.150 411.600 457.350 ;
        RECT 422.100 453.150 423.900 454.950 ;
        RECT 400.950 449.850 403.050 451.950 ;
        RECT 406.950 449.850 409.050 451.950 ;
        RECT 409.950 451.050 412.050 453.150 ;
        RECT 421.950 451.050 424.050 453.150 ;
        RECT 425.550 451.950 426.750 459.300 ;
        RECT 428.100 453.150 429.900 454.950 ;
        RECT 443.100 453.150 444.900 454.950 ;
        RECT 372.150 448.200 389.850 448.800 ;
        RECT 364.950 446.400 365.850 447.300 ;
        RECT 363.150 444.600 365.850 446.400 ;
        RECT 366.750 446.100 368.550 446.400 ;
        RECT 372.150 446.100 373.050 448.200 ;
        RECT 378.750 447.600 389.850 448.200 ;
        RECT 401.100 448.050 402.900 449.850 ;
        RECT 366.750 445.200 373.050 446.100 ;
        RECT 373.950 446.700 375.750 447.300 ;
        RECT 373.950 445.500 381.450 446.700 ;
        RECT 366.750 444.600 368.550 445.200 ;
        RECT 380.250 444.600 381.450 445.500 ;
        RECT 361.950 441.600 365.850 443.700 ;
        RECT 370.950 442.500 377.850 444.300 ;
        RECT 380.250 442.500 385.050 444.600 ;
        RECT 359.550 435.750 361.350 438.600 ;
        RECT 364.050 435.750 365.850 441.600 ;
        RECT 368.250 435.750 370.050 441.600 ;
        RECT 372.150 435.750 373.950 442.500 ;
        RECT 380.250 441.600 381.450 442.500 ;
        RECT 375.150 435.750 376.950 441.600 ;
        RECT 379.950 435.750 381.750 441.600 ;
        RECT 385.050 435.750 386.850 441.600 ;
        RECT 388.050 435.750 389.850 447.600 ;
        RECT 403.950 446.850 406.050 448.950 ;
        RECT 407.250 448.050 409.050 449.850 ;
        RECT 404.100 445.050 405.900 446.850 ;
        RECT 410.700 442.800 411.750 451.050 ;
        RECT 424.950 449.850 427.050 451.950 ;
        RECT 427.950 451.050 430.050 453.150 ;
        RECT 442.950 451.050 445.050 453.150 ;
        RECT 446.250 451.950 447.450 459.300 ;
        RECT 464.250 459.300 465.450 461.400 ;
        RECT 466.650 462.300 468.450 467.250 ;
        RECT 469.650 463.200 471.450 467.250 ;
        RECT 472.650 462.300 474.450 467.250 ;
        RECT 466.650 460.950 474.450 462.300 ;
        RECT 464.250 458.250 468.000 459.300 ;
        RECT 482.700 458.400 484.500 467.250 ;
        RECT 488.100 459.000 489.900 467.250 ;
        RECT 506.850 461.400 508.650 467.250 ;
        RECT 511.350 460.200 513.150 467.250 ;
        RECT 529.650 464.400 531.450 467.250 ;
        RECT 532.650 464.400 534.450 467.250 ;
        RECT 509.550 459.300 513.150 460.200 ;
        RECT 466.950 454.950 468.150 458.250 ;
        RECT 470.100 456.150 471.900 457.950 ;
        RECT 488.100 457.350 492.600 459.000 ;
        RECT 475.950 456.450 478.050 457.050 ;
        RECT 484.950 456.450 487.050 457.050 ;
        RECT 449.100 453.150 450.900 454.950 ;
        RECT 445.950 449.850 448.050 451.950 ;
        RECT 448.950 451.050 451.050 453.150 ;
        RECT 466.950 452.850 469.050 454.950 ;
        RECT 469.950 454.050 472.050 456.150 ;
        RECT 475.950 455.550 487.050 456.450 ;
        RECT 475.950 454.950 478.050 455.550 ;
        RECT 484.950 454.950 487.050 455.550 ;
        RECT 472.950 452.850 475.050 454.950 ;
        RECT 491.400 453.150 492.600 457.350 ;
        RECT 506.100 453.150 507.900 454.950 ;
        RECT 463.950 449.850 466.050 451.950 ;
        RECT 404.700 441.900 411.750 442.800 ;
        RECT 404.700 441.600 406.350 441.900 ;
        RECT 401.550 435.750 403.350 441.600 ;
        RECT 404.550 435.750 406.350 441.600 ;
        RECT 410.550 441.600 411.750 441.900 ;
        RECT 425.550 441.600 426.750 449.850 ;
        RECT 446.250 441.600 447.450 449.850 ;
        RECT 464.250 448.050 466.050 449.850 ;
        RECT 467.850 447.600 469.050 452.850 ;
        RECT 473.100 451.050 474.900 452.850 ;
        RECT 481.950 449.850 484.050 451.950 ;
        RECT 487.950 449.850 490.050 451.950 ;
        RECT 490.950 451.050 493.050 453.150 ;
        RECT 505.950 451.050 508.050 453.150 ;
        RECT 509.550 451.950 510.750 459.300 ;
        RECT 530.400 456.150 531.600 464.400 ;
        RECT 544.650 461.400 546.450 467.250 ;
        RECT 545.250 459.300 546.450 461.400 ;
        RECT 547.650 462.300 549.450 467.250 ;
        RECT 550.650 463.200 552.450 467.250 ;
        RECT 553.650 462.300 555.450 467.250 ;
        RECT 547.650 460.950 555.450 462.300 ;
        RECT 545.250 458.250 549.000 459.300 ;
        RECT 566.700 458.400 568.500 467.250 ;
        RECT 572.100 459.000 573.900 467.250 ;
        RECT 590.850 460.200 592.650 467.250 ;
        RECT 595.350 461.400 597.150 467.250 ;
        RECT 610.650 461.400 612.450 467.250 ;
        RECT 590.850 459.300 594.450 460.200 ;
        RECT 512.100 453.150 513.900 454.950 ;
        RECT 529.950 454.050 532.050 456.150 ;
        RECT 532.950 455.850 535.050 457.950 ;
        RECT 533.100 454.050 534.900 455.850 ;
        RECT 547.950 454.950 549.150 458.250 ;
        RECT 551.100 456.150 552.900 457.950 ;
        RECT 572.100 457.350 576.600 459.000 ;
        RECT 482.100 448.050 483.900 449.850 ;
        RECT 407.550 435.750 409.350 441.000 ;
        RECT 410.550 435.750 412.350 441.600 ;
        RECT 422.550 435.750 424.350 441.600 ;
        RECT 425.550 435.750 427.350 441.600 ;
        RECT 428.550 435.750 430.350 441.600 ;
        RECT 442.650 435.750 444.450 441.600 ;
        RECT 445.650 435.750 447.450 441.600 ;
        RECT 448.650 435.750 450.450 441.600 ;
        RECT 464.400 435.750 466.200 441.600 ;
        RECT 467.700 435.750 469.500 447.600 ;
        RECT 471.900 435.750 473.700 447.600 ;
        RECT 484.950 446.850 487.050 448.950 ;
        RECT 488.250 448.050 490.050 449.850 ;
        RECT 485.100 445.050 486.900 446.850 ;
        RECT 491.700 442.800 492.750 451.050 ;
        RECT 508.950 449.850 511.050 451.950 ;
        RECT 511.950 451.050 514.050 453.150 ;
        RECT 485.700 441.900 492.750 442.800 ;
        RECT 485.700 441.600 487.350 441.900 ;
        RECT 482.550 435.750 484.350 441.600 ;
        RECT 485.550 435.750 487.350 441.600 ;
        RECT 491.550 441.600 492.750 441.900 ;
        RECT 509.550 441.600 510.750 449.850 ;
        RECT 530.400 441.600 531.600 454.050 ;
        RECT 547.950 452.850 550.050 454.950 ;
        RECT 550.950 454.050 553.050 456.150 ;
        RECT 553.950 452.850 556.050 454.950 ;
        RECT 575.400 453.150 576.600 457.350 ;
        RECT 590.100 453.150 591.900 454.950 ;
        RECT 544.950 449.850 547.050 451.950 ;
        RECT 545.250 448.050 547.050 449.850 ;
        RECT 548.850 447.600 550.050 452.850 ;
        RECT 554.100 451.050 555.900 452.850 ;
        RECT 565.950 449.850 568.050 451.950 ;
        RECT 571.950 449.850 574.050 451.950 ;
        RECT 574.950 451.050 577.050 453.150 ;
        RECT 589.950 451.050 592.050 453.150 ;
        RECT 593.250 451.950 594.450 459.300 ;
        RECT 611.250 459.300 612.450 461.400 ;
        RECT 613.650 462.300 615.450 467.250 ;
        RECT 616.650 463.200 618.450 467.250 ;
        RECT 619.650 462.300 621.450 467.250 ;
        RECT 613.650 460.950 621.450 462.300 ;
        RECT 635.850 460.200 637.650 467.250 ;
        RECT 640.350 461.400 642.150 467.250 ;
        RECT 652.650 461.400 654.450 467.250 ;
        RECT 635.850 459.300 639.450 460.200 ;
        RECT 611.250 458.250 615.000 459.300 ;
        RECT 613.950 454.950 615.150 458.250 ;
        RECT 617.100 456.150 618.900 457.950 ;
        RECT 596.100 453.150 597.900 454.950 ;
        RECT 566.100 448.050 567.900 449.850 ;
        RECT 488.550 435.750 490.350 441.000 ;
        RECT 491.550 435.750 493.350 441.600 ;
        RECT 506.550 435.750 508.350 441.600 ;
        RECT 509.550 435.750 511.350 441.600 ;
        RECT 512.550 435.750 514.350 441.600 ;
        RECT 529.650 435.750 531.450 441.600 ;
        RECT 532.650 435.750 534.450 441.600 ;
        RECT 545.400 435.750 547.200 441.600 ;
        RECT 548.700 435.750 550.500 447.600 ;
        RECT 552.900 435.750 554.700 447.600 ;
        RECT 568.950 446.850 571.050 448.950 ;
        RECT 572.250 448.050 574.050 449.850 ;
        RECT 569.100 445.050 570.900 446.850 ;
        RECT 575.700 442.800 576.750 451.050 ;
        RECT 592.950 449.850 595.050 451.950 ;
        RECT 595.950 451.050 598.050 453.150 ;
        RECT 613.950 452.850 616.050 454.950 ;
        RECT 616.950 454.050 619.050 456.150 ;
        RECT 619.950 452.850 622.050 454.950 ;
        RECT 635.100 453.150 636.900 454.950 ;
        RECT 610.950 449.850 613.050 451.950 ;
        RECT 569.700 441.900 576.750 442.800 ;
        RECT 569.700 441.600 571.350 441.900 ;
        RECT 566.550 435.750 568.350 441.600 ;
        RECT 569.550 435.750 571.350 441.600 ;
        RECT 575.550 441.600 576.750 441.900 ;
        RECT 593.250 441.600 594.450 449.850 ;
        RECT 611.250 448.050 613.050 449.850 ;
        RECT 614.850 447.600 616.050 452.850 ;
        RECT 620.100 451.050 621.900 452.850 ;
        RECT 634.950 451.050 637.050 453.150 ;
        RECT 638.250 451.950 639.450 459.300 ;
        RECT 653.250 459.300 654.450 461.400 ;
        RECT 655.650 462.300 657.450 467.250 ;
        RECT 658.650 463.200 660.450 467.250 ;
        RECT 661.650 462.300 663.450 467.250 ;
        RECT 655.650 460.950 663.450 462.300 ;
        RECT 674.550 462.300 676.350 467.250 ;
        RECT 677.550 463.200 679.350 467.250 ;
        RECT 680.550 462.300 682.350 467.250 ;
        RECT 674.550 460.950 682.350 462.300 ;
        RECT 683.550 461.400 685.350 467.250 ;
        RECT 661.950 459.450 664.050 460.050 ;
        RECT 670.950 459.450 673.050 460.050 ;
        RECT 653.250 458.250 657.000 459.300 ;
        RECT 661.950 458.550 673.050 459.450 ;
        RECT 683.550 459.300 684.750 461.400 ;
        RECT 655.950 454.950 657.150 458.250 ;
        RECT 661.950 457.950 664.050 458.550 ;
        RECT 670.950 457.950 673.050 458.550 ;
        RECT 681.000 458.250 684.750 459.300 ;
        RECT 695.700 458.400 697.500 467.250 ;
        RECT 701.100 459.000 702.900 467.250 ;
        RECT 718.650 461.400 720.450 467.250 ;
        RECT 719.250 459.300 720.450 461.400 ;
        RECT 721.650 462.300 723.450 467.250 ;
        RECT 724.650 463.200 726.450 467.250 ;
        RECT 727.650 462.300 729.450 467.250 ;
        RECT 740.550 464.400 742.350 467.250 ;
        RECT 743.550 464.400 745.350 467.250 ;
        RECT 746.550 464.400 748.350 467.250 ;
        RECT 761.550 464.400 763.350 467.250 ;
        RECT 721.650 460.950 729.450 462.300 ;
        RECT 659.100 456.150 660.900 457.950 ;
        RECT 677.100 456.150 678.900 457.950 ;
        RECT 641.100 453.150 642.900 454.950 ;
        RECT 637.950 449.850 640.050 451.950 ;
        RECT 640.950 451.050 643.050 453.150 ;
        RECT 655.950 452.850 658.050 454.950 ;
        RECT 658.950 454.050 661.050 456.150 ;
        RECT 661.950 452.850 664.050 454.950 ;
        RECT 673.950 452.850 676.050 454.950 ;
        RECT 676.950 454.050 679.050 456.150 ;
        RECT 680.850 454.950 682.050 458.250 ;
        RECT 701.100 457.350 705.600 459.000 ;
        RECT 719.250 458.250 723.000 459.300 ;
        RECT 679.950 452.850 682.050 454.950 ;
        RECT 704.400 453.150 705.600 457.350 ;
        RECT 721.950 454.950 723.150 458.250 ;
        RECT 744.000 457.950 745.050 464.400 ;
        RECT 762.150 460.500 763.350 464.400 ;
        RECT 764.850 461.400 766.650 467.250 ;
        RECT 767.850 461.400 769.650 467.250 ;
        RECT 782.550 464.400 784.350 467.250 ;
        RECT 762.150 459.600 767.250 460.500 ;
        RECT 725.100 456.150 726.900 457.950 ;
        RECT 652.950 449.850 655.050 451.950 ;
        RECT 572.550 435.750 574.350 441.000 ;
        RECT 575.550 435.750 577.350 441.600 ;
        RECT 589.650 435.750 591.450 441.600 ;
        RECT 592.650 435.750 594.450 441.600 ;
        RECT 595.650 435.750 597.450 441.600 ;
        RECT 611.400 435.750 613.200 441.600 ;
        RECT 614.700 435.750 616.500 447.600 ;
        RECT 618.900 435.750 620.700 447.600 ;
        RECT 638.250 441.600 639.450 449.850 ;
        RECT 653.250 448.050 655.050 449.850 ;
        RECT 656.850 447.600 658.050 452.850 ;
        RECT 662.100 451.050 663.900 452.850 ;
        RECT 674.100 451.050 675.900 452.850 ;
        RECT 679.950 447.600 681.150 452.850 ;
        RECT 682.950 449.850 685.050 451.950 ;
        RECT 694.950 449.850 697.050 451.950 ;
        RECT 700.950 449.850 703.050 451.950 ;
        RECT 703.950 451.050 706.050 453.150 ;
        RECT 721.950 452.850 724.050 454.950 ;
        RECT 724.950 454.050 727.050 456.150 ;
        RECT 742.950 455.850 745.050 457.950 ;
        RECT 727.950 452.850 730.050 454.950 ;
        RECT 739.950 452.850 742.050 454.950 ;
        RECT 682.950 448.050 684.750 449.850 ;
        RECT 695.100 448.050 696.900 449.850 ;
        RECT 634.650 435.750 636.450 441.600 ;
        RECT 637.650 435.750 639.450 441.600 ;
        RECT 640.650 435.750 642.450 441.600 ;
        RECT 653.400 435.750 655.200 441.600 ;
        RECT 656.700 435.750 658.500 447.600 ;
        RECT 660.900 435.750 662.700 447.600 ;
        RECT 675.300 435.750 677.100 447.600 ;
        RECT 679.500 435.750 681.300 447.600 ;
        RECT 697.950 446.850 700.050 448.950 ;
        RECT 701.250 448.050 703.050 449.850 ;
        RECT 698.100 445.050 699.900 446.850 ;
        RECT 704.700 442.800 705.750 451.050 ;
        RECT 718.950 449.850 721.050 451.950 ;
        RECT 719.250 448.050 721.050 449.850 ;
        RECT 722.850 447.600 724.050 452.850 ;
        RECT 728.100 451.050 729.900 452.850 ;
        RECT 740.100 451.050 741.900 452.850 ;
        RECT 744.000 448.650 745.050 455.850 ;
        RECT 765.000 458.700 767.250 459.600 ;
        RECT 745.950 452.850 748.050 454.950 ;
        RECT 760.950 452.850 763.050 454.950 ;
        RECT 746.100 451.050 747.900 452.850 ;
        RECT 761.100 451.050 762.900 452.850 ;
        RECT 765.000 450.300 766.050 458.700 ;
        RECT 768.150 454.950 769.350 461.400 ;
        RECT 783.150 460.500 784.350 464.400 ;
        RECT 785.850 461.400 787.650 467.250 ;
        RECT 788.850 461.400 790.650 467.250 ;
        RECT 800.550 464.400 802.350 467.250 ;
        RECT 803.550 464.400 805.350 467.250 ;
        RECT 806.550 464.400 808.350 467.250 ;
        RECT 820.650 464.400 822.450 467.250 ;
        RECT 823.650 464.400 825.450 467.250 ;
        RECT 833.550 464.400 835.350 467.250 ;
        RECT 836.550 464.400 838.350 467.250 ;
        RECT 839.550 464.400 841.350 467.250 ;
        RECT 783.150 459.600 788.250 460.500 ;
        RECT 786.000 458.700 788.250 459.600 ;
        RECT 766.950 452.850 769.350 454.950 ;
        RECT 781.950 452.850 784.050 454.950 ;
        RECT 765.000 449.400 767.250 450.300 ;
        RECT 744.000 447.600 746.550 448.650 ;
        RECT 698.700 441.900 705.750 442.800 ;
        RECT 698.700 441.600 700.350 441.900 ;
        RECT 682.800 435.750 684.600 441.600 ;
        RECT 695.550 435.750 697.350 441.600 ;
        RECT 698.550 435.750 700.350 441.600 ;
        RECT 704.550 441.600 705.750 441.900 ;
        RECT 701.550 435.750 703.350 441.000 ;
        RECT 704.550 435.750 706.350 441.600 ;
        RECT 719.400 435.750 721.200 441.600 ;
        RECT 722.700 435.750 724.500 447.600 ;
        RECT 726.900 435.750 728.700 447.600 ;
        RECT 740.550 435.750 742.350 447.600 ;
        RECT 744.750 435.750 746.550 447.600 ;
        RECT 761.550 448.500 767.250 449.400 ;
        RECT 761.550 441.600 762.750 448.500 ;
        RECT 768.150 447.600 769.350 452.850 ;
        RECT 782.100 451.050 783.900 452.850 ;
        RECT 786.000 450.300 787.050 458.700 ;
        RECT 789.150 454.950 790.350 461.400 ;
        RECT 804.000 457.950 805.050 464.400 ;
        RECT 802.950 455.850 805.050 457.950 ;
        RECT 821.400 456.150 822.600 464.400 ;
        RECT 837.450 460.200 838.350 464.400 ;
        RECT 842.550 461.400 844.350 467.250 ;
        RECT 848.550 461.400 850.350 467.250 ;
        RECT 851.850 464.400 853.650 467.250 ;
        RECT 856.350 464.400 858.150 467.250 ;
        RECT 860.550 464.400 862.350 467.250 ;
        RECT 864.450 464.400 866.250 467.250 ;
        RECT 867.750 464.400 869.550 467.250 ;
        RECT 872.250 465.300 874.050 467.250 ;
        RECT 872.250 464.400 876.000 465.300 ;
        RECT 877.050 464.400 878.850 467.250 ;
        RECT 856.650 463.500 857.700 464.400 ;
        RECT 853.950 462.300 857.700 463.500 ;
        RECT 865.200 462.600 866.250 464.400 ;
        RECT 874.950 463.500 876.000 464.400 ;
        RECT 853.950 461.400 856.050 462.300 ;
        RECT 837.450 459.300 840.750 460.200 ;
        RECT 838.950 458.400 840.750 459.300 ;
        RECT 787.950 452.850 790.350 454.950 ;
        RECT 799.950 452.850 802.050 454.950 ;
        RECT 786.000 449.400 788.250 450.300 ;
        RECT 782.550 448.500 788.250 449.400 ;
        RECT 761.550 435.750 763.350 441.600 ;
        RECT 764.850 435.750 766.650 447.600 ;
        RECT 767.850 435.750 769.650 447.600 ;
        RECT 782.550 441.600 783.750 448.500 ;
        RECT 789.150 447.600 790.350 452.850 ;
        RECT 800.100 451.050 801.900 452.850 ;
        RECT 804.000 448.650 805.050 455.850 ;
        RECT 805.950 452.850 808.050 454.950 ;
        RECT 820.950 454.050 823.050 456.150 ;
        RECT 823.950 455.850 826.050 457.950 ;
        RECT 832.950 455.850 835.050 457.950 ;
        RECT 824.100 454.050 825.900 455.850 ;
        RECT 833.100 454.050 834.900 455.850 ;
        RECT 806.100 451.050 807.900 452.850 ;
        RECT 804.000 447.600 806.550 448.650 ;
        RECT 782.550 435.750 784.350 441.600 ;
        RECT 785.850 435.750 787.650 447.600 ;
        RECT 788.850 435.750 790.650 447.600 ;
        RECT 800.550 435.750 802.350 447.600 ;
        RECT 804.750 435.750 806.550 447.600 ;
        RECT 821.400 441.600 822.600 454.050 ;
        RECT 835.950 452.850 838.050 454.950 ;
        RECT 836.100 451.050 837.900 452.850 ;
        RECT 839.700 450.150 840.600 458.400 ;
        RECT 843.000 456.150 844.050 461.400 ;
        RECT 841.950 454.050 844.050 456.150 ;
        RECT 848.550 459.150 849.750 461.400 ;
        RECT 861.150 460.200 862.950 462.000 ;
        RECT 865.200 461.550 870.150 462.600 ;
        RECT 868.350 460.800 870.150 461.550 ;
        RECT 871.650 460.800 873.450 462.600 ;
        RECT 874.950 461.400 877.050 463.500 ;
        RECT 880.050 461.400 881.850 467.250 ;
        RECT 862.050 459.900 862.950 460.200 ;
        RECT 872.100 459.900 873.150 460.800 ;
        RECT 848.550 457.050 853.050 459.150 ;
        RECT 862.050 459.000 873.150 459.900 ;
        RECT 838.950 450.000 840.750 450.150 ;
        RECT 833.550 448.800 840.750 450.000 ;
        RECT 833.550 447.600 834.750 448.800 ;
        RECT 838.950 448.350 840.750 448.800 ;
        RECT 820.650 435.750 822.450 441.600 ;
        RECT 823.650 435.750 825.450 441.600 ;
        RECT 833.550 435.750 835.350 447.600 ;
        RECT 842.100 447.450 843.450 454.050 ;
        RECT 838.050 435.750 839.850 447.450 ;
        RECT 841.050 446.100 843.450 447.450 ;
        RECT 848.550 447.600 849.750 457.050 ;
        RECT 850.950 455.250 854.850 457.050 ;
        RECT 850.950 454.950 853.050 455.250 ;
        RECT 862.050 454.950 862.950 459.000 ;
        RECT 872.100 457.800 873.150 459.000 ;
        RECT 872.100 456.600 879.000 457.800 ;
        RECT 872.100 456.000 873.900 456.600 ;
        RECT 878.100 455.850 879.000 456.600 ;
        RECT 875.100 454.950 876.900 455.700 ;
        RECT 862.050 452.850 865.050 454.950 ;
        RECT 868.950 453.900 876.900 454.950 ;
        RECT 878.100 454.050 879.900 455.850 ;
        RECT 868.950 452.850 871.050 453.900 ;
        RECT 850.950 449.400 852.750 451.200 ;
        RECT 851.850 448.200 856.050 449.400 ;
        RECT 862.050 448.200 862.950 452.850 ;
        RECT 870.750 449.100 872.550 449.400 ;
        RECT 841.050 435.750 842.850 446.100 ;
        RECT 848.550 435.750 850.350 447.600 ;
        RECT 853.950 447.300 856.050 448.200 ;
        RECT 856.950 447.300 862.950 448.200 ;
        RECT 864.150 448.800 872.550 449.100 ;
        RECT 880.950 448.800 881.850 461.400 ;
        RECT 864.150 448.200 881.850 448.800 ;
        RECT 856.950 446.400 857.850 447.300 ;
        RECT 855.150 444.600 857.850 446.400 ;
        RECT 858.750 446.100 860.550 446.400 ;
        RECT 864.150 446.100 865.050 448.200 ;
        RECT 870.750 447.600 881.850 448.200 ;
        RECT 858.750 445.200 865.050 446.100 ;
        RECT 865.950 446.700 867.750 447.300 ;
        RECT 865.950 445.500 873.450 446.700 ;
        RECT 858.750 444.600 860.550 445.200 ;
        RECT 872.250 444.600 873.450 445.500 ;
        RECT 853.950 441.600 857.850 443.700 ;
        RECT 862.950 442.500 869.850 444.300 ;
        RECT 872.250 442.500 877.050 444.600 ;
        RECT 851.550 435.750 853.350 438.600 ;
        RECT 856.050 435.750 857.850 441.600 ;
        RECT 860.250 435.750 862.050 441.600 ;
        RECT 864.150 435.750 865.950 442.500 ;
        RECT 872.250 441.600 873.450 442.500 ;
        RECT 867.150 435.750 868.950 441.600 ;
        RECT 871.950 435.750 873.750 441.600 ;
        RECT 877.050 435.750 878.850 441.600 ;
        RECT 880.050 435.750 881.850 447.600 ;
        RECT 11.400 425.400 13.200 431.250 ;
        RECT 14.700 419.400 16.500 431.250 ;
        RECT 18.900 419.400 20.700 431.250 ;
        RECT 24.150 419.400 25.950 431.250 ;
        RECT 27.150 425.400 28.950 431.250 ;
        RECT 32.250 425.400 34.050 431.250 ;
        RECT 37.050 425.400 38.850 431.250 ;
        RECT 32.550 424.500 33.750 425.400 ;
        RECT 40.050 424.500 41.850 431.250 ;
        RECT 43.950 425.400 45.750 431.250 ;
        RECT 48.150 425.400 49.950 431.250 ;
        RECT 52.650 428.400 54.450 431.250 ;
        RECT 28.950 422.400 33.750 424.500 ;
        RECT 36.150 422.700 43.050 424.500 ;
        RECT 48.150 423.300 52.050 425.400 ;
        RECT 32.550 421.500 33.750 422.400 ;
        RECT 45.450 421.800 47.250 422.400 ;
        RECT 32.550 420.300 40.050 421.500 ;
        RECT 38.250 419.700 40.050 420.300 ;
        RECT 40.950 420.900 47.250 421.800 ;
        RECT 11.250 417.150 13.050 418.950 ;
        RECT 10.950 415.050 13.050 417.150 ;
        RECT 14.850 414.150 16.050 419.400 ;
        RECT 24.150 418.800 35.250 419.400 ;
        RECT 40.950 418.800 41.850 420.900 ;
        RECT 45.450 420.600 47.250 420.900 ;
        RECT 48.150 420.600 50.850 422.400 ;
        RECT 48.150 419.700 49.050 420.600 ;
        RECT 24.150 418.200 41.850 418.800 ;
        RECT 20.100 414.150 21.900 415.950 ;
        RECT 13.950 412.050 16.050 414.150 ;
        RECT 13.950 408.750 15.150 412.050 ;
        RECT 16.950 410.850 19.050 412.950 ;
        RECT 19.950 412.050 22.050 414.150 ;
        RECT 17.100 409.050 18.900 410.850 ;
        RECT 11.250 407.700 15.000 408.750 ;
        RECT 11.250 405.600 12.450 407.700 ;
        RECT 10.650 399.750 12.450 405.600 ;
        RECT 13.650 404.700 21.450 406.050 ;
        RECT 13.650 399.750 15.450 404.700 ;
        RECT 16.650 399.750 18.450 403.800 ;
        RECT 19.650 399.750 21.450 404.700 ;
        RECT 24.150 405.600 25.050 418.200 ;
        RECT 33.450 417.900 41.850 418.200 ;
        RECT 43.050 418.800 49.050 419.700 ;
        RECT 49.950 418.800 52.050 419.700 ;
        RECT 55.650 419.400 57.450 431.250 ;
        RECT 69.300 419.400 71.100 431.250 ;
        RECT 73.500 419.400 75.300 431.250 ;
        RECT 76.800 425.400 78.600 431.250 ;
        RECT 89.550 425.400 91.350 431.250 ;
        RECT 92.550 425.400 94.350 431.250 ;
        RECT 95.550 425.400 97.350 431.250 ;
        RECT 110.400 425.400 112.200 431.250 ;
        RECT 33.450 417.600 35.250 417.900 ;
        RECT 43.050 414.150 43.950 418.800 ;
        RECT 49.950 417.600 54.150 418.800 ;
        RECT 53.250 415.800 55.050 417.600 ;
        RECT 34.950 413.100 37.050 414.150 ;
        RECT 26.100 411.150 27.900 412.950 ;
        RECT 29.100 412.050 37.050 413.100 ;
        RECT 40.950 412.050 43.950 414.150 ;
        RECT 29.100 411.300 30.900 412.050 ;
        RECT 27.000 410.400 27.900 411.150 ;
        RECT 32.100 410.400 33.900 411.000 ;
        RECT 27.000 409.200 33.900 410.400 ;
        RECT 32.850 408.000 33.900 409.200 ;
        RECT 43.050 408.000 43.950 412.050 ;
        RECT 52.950 411.750 55.050 412.050 ;
        RECT 51.150 409.950 55.050 411.750 ;
        RECT 56.250 409.950 57.450 419.400 ;
        RECT 68.100 414.150 69.900 415.950 ;
        RECT 73.950 414.150 75.150 419.400 ;
        RECT 76.950 417.150 78.750 418.950 ;
        RECT 92.550 417.150 93.750 425.400 ;
        RECT 113.700 419.400 115.500 431.250 ;
        RECT 117.900 419.400 119.700 431.250 ;
        RECT 130.650 425.400 132.450 431.250 ;
        RECT 133.650 425.400 135.450 431.250 ;
        RECT 110.250 417.150 112.050 418.950 ;
        RECT 76.950 415.050 79.050 417.150 ;
        RECT 67.950 412.050 70.050 414.150 ;
        RECT 70.950 410.850 73.050 412.950 ;
        RECT 73.950 412.050 76.050 414.150 ;
        RECT 88.950 413.850 91.050 415.950 ;
        RECT 91.950 415.050 94.050 417.150 ;
        RECT 89.100 412.050 90.900 413.850 ;
        RECT 32.850 407.100 43.950 408.000 ;
        RECT 52.950 407.850 57.450 409.950 ;
        RECT 71.100 409.050 72.900 410.850 ;
        RECT 74.850 408.750 76.050 412.050 ;
        RECT 32.850 406.200 33.900 407.100 ;
        RECT 43.050 406.800 43.950 407.100 ;
        RECT 24.150 399.750 25.950 405.600 ;
        RECT 28.950 403.500 31.050 405.600 ;
        RECT 32.550 404.400 34.350 406.200 ;
        RECT 35.850 405.450 37.650 406.200 ;
        RECT 35.850 404.400 40.800 405.450 ;
        RECT 43.050 405.000 44.850 406.800 ;
        RECT 56.250 405.600 57.450 407.850 ;
        RECT 75.000 407.700 78.750 408.750 ;
        RECT 49.950 404.700 52.050 405.600 ;
        RECT 30.000 402.600 31.050 403.500 ;
        RECT 39.750 402.600 40.800 404.400 ;
        RECT 48.300 403.500 52.050 404.700 ;
        RECT 48.300 402.600 49.350 403.500 ;
        RECT 27.150 399.750 28.950 402.600 ;
        RECT 30.000 401.700 33.750 402.600 ;
        RECT 31.950 399.750 33.750 401.700 ;
        RECT 36.450 399.750 38.250 402.600 ;
        RECT 39.750 399.750 41.550 402.600 ;
        RECT 43.650 399.750 45.450 402.600 ;
        RECT 47.850 399.750 49.650 402.600 ;
        RECT 52.350 399.750 54.150 402.600 ;
        RECT 55.650 399.750 57.450 405.600 ;
        RECT 68.550 404.700 76.350 406.050 ;
        RECT 68.550 399.750 70.350 404.700 ;
        RECT 71.550 399.750 73.350 403.800 ;
        RECT 74.550 399.750 76.350 404.700 ;
        RECT 77.550 405.600 78.750 407.700 ;
        RECT 92.550 407.700 93.750 415.050 ;
        RECT 94.950 413.850 97.050 415.950 ;
        RECT 109.950 415.050 112.050 417.150 ;
        RECT 113.850 414.150 115.050 419.400 ;
        RECT 119.100 414.150 120.900 415.950 ;
        RECT 95.100 412.050 96.900 413.850 ;
        RECT 112.950 412.050 115.050 414.150 ;
        RECT 112.950 408.750 114.150 412.050 ;
        RECT 115.950 410.850 118.050 412.950 ;
        RECT 118.950 412.050 121.050 414.150 ;
        RECT 131.400 412.950 132.600 425.400 ;
        RECT 145.350 419.400 147.150 431.250 ;
        RECT 148.350 419.400 150.150 431.250 ;
        RECT 151.650 425.400 153.450 431.250 ;
        RECT 166.650 425.400 168.450 431.250 ;
        RECT 169.650 425.400 171.450 431.250 ;
        RECT 172.650 425.400 174.450 431.250 ;
        RECT 185.400 425.400 187.200 431.250 ;
        RECT 145.650 414.150 146.850 419.400 ;
        RECT 152.250 418.500 153.450 425.400 ;
        RECT 147.750 417.600 153.450 418.500 ;
        RECT 147.750 416.700 150.000 417.600 ;
        RECT 170.250 417.150 171.450 425.400 ;
        RECT 188.700 419.400 190.500 431.250 ;
        RECT 192.900 419.400 194.700 431.250 ;
        RECT 205.650 425.400 207.450 431.250 ;
        RECT 208.650 425.400 210.450 431.250 ;
        RECT 211.650 425.400 213.450 431.250 ;
        RECT 226.650 425.400 228.450 431.250 ;
        RECT 229.650 425.400 231.450 431.250 ;
        RECT 232.650 425.400 234.450 431.250 ;
        RECT 248.400 425.400 250.200 431.250 ;
        RECT 185.250 417.150 187.050 418.950 ;
        RECT 130.950 410.850 133.050 412.950 ;
        RECT 134.100 411.150 135.900 412.950 ;
        RECT 145.650 412.050 148.050 414.150 ;
        RECT 116.100 409.050 117.900 410.850 ;
        RECT 110.250 407.700 114.000 408.750 ;
        RECT 92.550 406.800 96.150 407.700 ;
        RECT 77.550 399.750 79.350 405.600 ;
        RECT 89.850 399.750 91.650 405.600 ;
        RECT 94.350 399.750 96.150 406.800 ;
        RECT 110.250 405.600 111.450 407.700 ;
        RECT 109.650 399.750 111.450 405.600 ;
        RECT 112.650 404.700 120.450 406.050 ;
        RECT 112.650 399.750 114.450 404.700 ;
        RECT 115.650 399.750 117.450 403.800 ;
        RECT 118.650 399.750 120.450 404.700 ;
        RECT 131.400 402.600 132.600 410.850 ;
        RECT 133.950 409.050 136.050 411.150 ;
        RECT 145.650 405.600 146.850 412.050 ;
        RECT 148.950 408.300 150.000 416.700 ;
        RECT 152.100 414.150 153.900 415.950 ;
        RECT 151.950 412.050 154.050 414.150 ;
        RECT 166.950 413.850 169.050 415.950 ;
        RECT 169.950 415.050 172.050 417.150 ;
        RECT 167.100 412.050 168.900 413.850 ;
        RECT 147.750 407.400 150.000 408.300 ;
        RECT 170.250 407.700 171.450 415.050 ;
        RECT 172.950 413.850 175.050 415.950 ;
        RECT 184.950 415.050 187.050 417.150 ;
        RECT 188.850 414.150 190.050 419.400 ;
        RECT 209.250 417.150 210.450 425.400 ;
        RECT 230.250 417.150 231.450 425.400 ;
        RECT 251.700 419.400 253.500 431.250 ;
        RECT 255.900 419.400 257.700 431.250 ;
        RECT 266.550 425.400 268.350 431.250 ;
        RECT 269.550 425.400 271.350 431.250 ;
        RECT 272.550 426.000 274.350 431.250 ;
        RECT 269.700 425.100 271.350 425.400 ;
        RECT 275.550 425.400 277.350 431.250 ;
        RECT 289.650 425.400 291.450 431.250 ;
        RECT 292.650 426.000 294.450 431.250 ;
        RECT 275.550 425.100 276.750 425.400 ;
        RECT 269.700 424.200 276.750 425.100 ;
        RECT 269.100 420.150 270.900 421.950 ;
        RECT 248.250 417.150 250.050 418.950 ;
        RECT 194.100 414.150 195.900 415.950 ;
        RECT 173.100 412.050 174.900 413.850 ;
        RECT 187.950 412.050 190.050 414.150 ;
        RECT 187.950 408.750 189.150 412.050 ;
        RECT 190.950 410.850 193.050 412.950 ;
        RECT 193.950 412.050 196.050 414.150 ;
        RECT 205.950 413.850 208.050 415.950 ;
        RECT 208.950 415.050 211.050 417.150 ;
        RECT 206.100 412.050 207.900 413.850 ;
        RECT 191.100 409.050 192.900 410.850 ;
        RECT 147.750 406.500 152.850 407.400 ;
        RECT 130.650 399.750 132.450 402.600 ;
        RECT 133.650 399.750 135.450 402.600 ;
        RECT 145.350 399.750 147.150 405.600 ;
        RECT 148.350 399.750 150.150 405.600 ;
        RECT 151.650 402.600 152.850 406.500 ;
        RECT 167.850 406.800 171.450 407.700 ;
        RECT 185.250 407.700 189.000 408.750 ;
        RECT 209.250 407.700 210.450 415.050 ;
        RECT 211.950 413.850 214.050 415.950 ;
        RECT 226.950 413.850 229.050 415.950 ;
        RECT 229.950 415.050 232.050 417.150 ;
        RECT 212.100 412.050 213.900 413.850 ;
        RECT 227.100 412.050 228.900 413.850 ;
        RECT 230.250 407.700 231.450 415.050 ;
        RECT 232.950 413.850 235.050 415.950 ;
        RECT 247.950 415.050 250.050 417.150 ;
        RECT 251.850 414.150 253.050 419.400 ;
        RECT 266.100 417.150 267.900 418.950 ;
        RECT 268.950 418.050 271.050 420.150 ;
        RECT 272.250 417.150 274.050 418.950 ;
        RECT 257.100 414.150 258.900 415.950 ;
        RECT 265.950 415.050 268.050 417.150 ;
        RECT 271.950 415.050 274.050 417.150 ;
        RECT 275.700 415.950 276.750 424.200 ;
        RECT 290.250 425.100 291.450 425.400 ;
        RECT 295.650 425.400 297.450 431.250 ;
        RECT 298.650 425.400 300.450 431.250 ;
        RECT 295.650 425.100 297.300 425.400 ;
        RECT 290.250 424.200 297.300 425.100 ;
        RECT 277.950 417.450 280.050 418.050 ;
        RECT 286.950 417.450 289.050 418.050 ;
        RECT 277.950 416.550 289.050 417.450 ;
        RECT 277.950 415.950 280.050 416.550 ;
        RECT 286.950 415.950 289.050 416.550 ;
        RECT 290.250 415.950 291.300 424.200 ;
        RECT 296.100 420.150 297.900 421.950 ;
        RECT 311.550 420.600 313.350 431.250 ;
        RECT 314.550 421.500 316.350 431.250 ;
        RECT 317.550 430.500 325.350 431.250 ;
        RECT 317.550 420.600 319.350 430.500 ;
        RECT 292.950 417.150 294.750 418.950 ;
        RECT 295.950 418.050 298.050 420.150 ;
        RECT 311.550 419.700 319.350 420.600 ;
        RECT 320.550 419.400 322.350 429.600 ;
        RECT 323.550 419.400 325.350 430.500 ;
        RECT 337.650 425.400 339.450 431.250 ;
        RECT 340.650 426.000 342.450 431.250 ;
        RECT 338.250 425.100 339.450 425.400 ;
        RECT 343.650 425.400 345.450 431.250 ;
        RECT 346.650 425.400 348.450 431.250 ;
        RECT 359.550 425.400 361.350 431.250 ;
        RECT 362.550 425.400 364.350 431.250 ;
        RECT 365.550 425.400 367.350 431.250 ;
        RECT 377.550 425.400 379.350 431.250 ;
        RECT 380.550 425.400 382.350 431.250 ;
        RECT 383.550 426.000 385.350 431.250 ;
        RECT 343.650 425.100 345.300 425.400 ;
        RECT 338.250 424.200 345.300 425.100 ;
        RECT 299.100 417.150 300.900 418.950 ;
        RECT 320.400 418.500 322.200 419.400 ;
        RECT 318.150 417.600 322.200 418.500 ;
        RECT 233.100 412.050 234.900 413.850 ;
        RECT 250.950 412.050 253.050 414.150 ;
        RECT 250.950 408.750 252.150 412.050 ;
        RECT 253.950 410.850 256.050 412.950 ;
        RECT 256.950 412.050 259.050 414.150 ;
        RECT 274.950 413.850 277.050 415.950 ;
        RECT 289.950 413.850 292.050 415.950 ;
        RECT 292.950 415.050 295.050 417.150 ;
        RECT 298.950 415.050 301.050 417.150 ;
        RECT 311.250 414.150 313.050 415.950 ;
        RECT 318.150 414.150 319.050 417.600 ;
        RECT 338.250 415.950 339.300 424.200 ;
        RECT 344.100 420.150 345.900 421.950 ;
        RECT 340.950 417.150 342.750 418.950 ;
        RECT 343.950 418.050 346.050 420.150 ;
        RECT 347.100 417.150 348.900 418.950 ;
        RECT 362.550 417.150 363.750 425.400 ;
        RECT 380.700 425.100 382.350 425.400 ;
        RECT 386.550 425.400 388.350 431.250 ;
        RECT 398.550 425.400 400.350 431.250 ;
        RECT 401.550 425.400 403.350 431.250 ;
        RECT 404.550 425.400 406.350 431.250 ;
        RECT 416.550 425.400 418.350 431.250 ;
        RECT 419.550 425.400 421.350 431.250 ;
        RECT 422.550 425.400 424.350 431.250 ;
        RECT 386.550 425.100 387.750 425.400 ;
        RECT 380.700 424.200 387.750 425.100 ;
        RECT 380.100 420.150 381.900 421.950 ;
        RECT 377.100 417.150 378.900 418.950 ;
        RECT 379.950 418.050 382.050 420.150 ;
        RECT 383.250 417.150 385.050 418.950 ;
        RECT 323.100 414.150 324.900 415.950 ;
        RECT 254.100 409.050 255.900 410.850 ;
        RECT 275.400 409.650 276.600 413.850 ;
        RECT 151.650 399.750 153.450 402.600 ;
        RECT 167.850 399.750 169.650 406.800 ;
        RECT 185.250 405.600 186.450 407.700 ;
        RECT 206.850 406.800 210.450 407.700 ;
        RECT 227.850 406.800 231.450 407.700 ;
        RECT 248.250 407.700 252.000 408.750 ;
        RECT 172.350 399.750 174.150 405.600 ;
        RECT 184.650 399.750 186.450 405.600 ;
        RECT 187.650 404.700 195.450 406.050 ;
        RECT 187.650 399.750 189.450 404.700 ;
        RECT 190.650 399.750 192.450 403.800 ;
        RECT 193.650 399.750 195.450 404.700 ;
        RECT 206.850 399.750 208.650 406.800 ;
        RECT 211.350 399.750 213.150 405.600 ;
        RECT 227.850 399.750 229.650 406.800 ;
        RECT 248.250 405.600 249.450 407.700 ;
        RECT 232.350 399.750 234.150 405.600 ;
        RECT 247.650 399.750 249.450 405.600 ;
        RECT 250.650 404.700 258.450 406.050 ;
        RECT 250.650 399.750 252.450 404.700 ;
        RECT 253.650 399.750 255.450 403.800 ;
        RECT 256.650 399.750 258.450 404.700 ;
        RECT 266.700 399.750 268.500 408.600 ;
        RECT 272.100 408.000 276.600 409.650 ;
        RECT 290.400 409.650 291.600 413.850 ;
        RECT 310.950 412.050 313.050 414.150 ;
        RECT 313.950 410.850 316.050 412.950 ;
        RECT 290.400 408.000 294.900 409.650 ;
        RECT 314.250 409.050 316.050 410.850 ;
        RECT 316.950 412.050 319.050 414.150 ;
        RECT 272.100 399.750 273.900 408.000 ;
        RECT 293.100 399.750 294.900 408.000 ;
        RECT 298.500 399.750 300.300 408.600 ;
        RECT 316.950 405.600 318.000 412.050 ;
        RECT 319.950 410.850 322.050 412.950 ;
        RECT 322.950 412.050 325.050 414.150 ;
        RECT 337.950 413.850 340.050 415.950 ;
        RECT 340.950 415.050 343.050 417.150 ;
        RECT 346.950 415.050 349.050 417.150 ;
        RECT 358.950 413.850 361.050 415.950 ;
        RECT 361.950 415.050 364.050 417.150 ;
        RECT 319.950 409.050 321.750 410.850 ;
        RECT 338.400 409.650 339.600 413.850 ;
        RECT 359.100 412.050 360.900 413.850 ;
        RECT 338.400 408.000 342.900 409.650 ;
        RECT 312.000 399.750 313.800 405.600 ;
        RECT 316.200 399.750 318.000 405.600 ;
        RECT 320.400 399.750 322.200 405.600 ;
        RECT 341.100 399.750 342.900 408.000 ;
        RECT 346.500 399.750 348.300 408.600 ;
        RECT 362.550 407.700 363.750 415.050 ;
        RECT 364.950 413.850 367.050 415.950 ;
        RECT 376.950 415.050 379.050 417.150 ;
        RECT 382.950 415.050 385.050 417.150 ;
        RECT 386.700 415.950 387.750 424.200 ;
        RECT 401.550 417.150 402.750 425.400 ;
        RECT 419.550 417.150 420.750 425.400 ;
        RECT 437.550 424.200 439.350 430.200 ;
        RECT 440.550 424.200 442.350 431.250 ;
        RECT 438.450 419.100 439.350 424.200 ;
        RECT 445.050 420.900 446.850 430.200 ;
        RECT 445.050 420.000 447.150 420.900 ;
        RECT 438.450 418.200 444.600 419.100 ;
        RECT 385.950 413.850 388.050 415.950 ;
        RECT 397.950 413.850 400.050 415.950 ;
        RECT 400.950 415.050 403.050 417.150 ;
        RECT 365.100 412.050 366.900 413.850 ;
        RECT 386.400 409.650 387.600 413.850 ;
        RECT 398.100 412.050 399.900 413.850 ;
        RECT 362.550 406.800 366.150 407.700 ;
        RECT 359.850 399.750 361.650 405.600 ;
        RECT 364.350 399.750 366.150 406.800 ;
        RECT 377.700 399.750 379.500 408.600 ;
        RECT 383.100 408.000 387.600 409.650 ;
        RECT 383.100 399.750 384.900 408.000 ;
        RECT 401.550 407.700 402.750 415.050 ;
        RECT 403.950 413.850 406.050 415.950 ;
        RECT 415.950 413.850 418.050 415.950 ;
        RECT 418.950 415.050 421.050 417.150 ;
        RECT 404.100 412.050 405.900 413.850 ;
        RECT 416.100 412.050 417.900 413.850 ;
        RECT 419.550 407.700 420.750 415.050 ;
        RECT 421.950 413.850 424.050 415.950 ;
        RECT 440.250 414.150 442.050 415.950 ;
        RECT 422.100 412.050 423.900 413.850 ;
        RECT 436.950 410.850 439.050 412.950 ;
        RECT 439.950 412.050 442.050 414.150 ;
        RECT 443.250 415.500 444.600 418.200 ;
        RECT 443.250 413.700 445.050 415.500 ;
        RECT 437.250 409.050 439.050 410.850 ;
        RECT 443.250 408.000 444.600 413.700 ;
        RECT 446.250 412.950 447.150 420.000 ;
        RECT 449.550 419.400 451.350 431.250 ;
        RECT 461.550 424.200 463.350 430.200 ;
        RECT 464.550 424.200 466.350 431.250 ;
        RECT 462.450 419.100 463.350 424.200 ;
        RECT 469.050 420.900 470.850 430.200 ;
        RECT 469.050 420.000 471.150 420.900 ;
        RECT 462.450 418.200 468.600 419.100 ;
        RECT 449.100 414.150 450.900 415.950 ;
        RECT 464.250 414.150 466.050 415.950 ;
        RECT 445.950 410.850 448.050 412.950 ;
        RECT 448.950 412.050 451.050 414.150 ;
        RECT 460.950 410.850 463.050 412.950 ;
        RECT 463.950 412.050 466.050 414.150 ;
        RECT 467.250 415.500 468.600 418.200 ;
        RECT 467.250 413.700 469.050 415.500 ;
        RECT 401.550 406.800 405.150 407.700 ;
        RECT 419.550 406.800 423.150 407.700 ;
        RECT 398.850 399.750 400.650 405.600 ;
        RECT 403.350 399.750 405.150 406.800 ;
        RECT 416.850 399.750 418.650 405.600 ;
        RECT 421.350 399.750 423.150 406.800 ;
        RECT 438.300 407.100 444.600 408.000 ;
        RECT 438.300 403.800 439.350 407.100 ;
        RECT 446.250 406.200 447.150 410.850 ;
        RECT 461.250 409.050 463.050 410.850 ;
        RECT 467.250 408.000 468.600 413.700 ;
        RECT 470.250 412.950 471.150 420.000 ;
        RECT 473.550 419.400 475.350 431.250 ;
        RECT 487.350 419.400 489.150 431.250 ;
        RECT 490.350 419.400 492.150 431.250 ;
        RECT 493.650 425.400 495.450 431.250 ;
        RECT 505.650 425.400 507.450 431.250 ;
        RECT 508.650 425.400 510.450 431.250 ;
        RECT 521.400 425.400 523.200 431.250 ;
        RECT 473.100 414.150 474.900 415.950 ;
        RECT 487.650 414.150 488.850 419.400 ;
        RECT 494.250 418.500 495.450 425.400 ;
        RECT 489.750 417.600 495.450 418.500 ;
        RECT 489.750 416.700 492.000 417.600 ;
        RECT 469.950 410.850 472.050 412.950 ;
        RECT 472.950 412.050 475.050 414.150 ;
        RECT 487.650 412.050 490.050 414.150 ;
        RECT 462.300 407.100 468.600 408.000 ;
        RECT 445.050 405.300 447.150 406.200 ;
        RECT 437.550 400.800 439.350 403.800 ;
        RECT 440.550 399.750 442.350 403.800 ;
        RECT 445.050 400.800 446.850 405.300 ;
        RECT 449.550 399.750 451.350 406.800 ;
        RECT 462.300 403.800 463.350 407.100 ;
        RECT 470.250 406.200 471.150 410.850 ;
        RECT 469.050 405.300 471.150 406.200 ;
        RECT 461.550 400.800 463.350 403.800 ;
        RECT 464.550 399.750 466.350 403.800 ;
        RECT 469.050 400.800 470.850 405.300 ;
        RECT 473.550 399.750 475.350 406.800 ;
        RECT 487.650 405.600 488.850 412.050 ;
        RECT 490.950 408.300 492.000 416.700 ;
        RECT 494.100 414.150 495.900 415.950 ;
        RECT 493.950 412.050 496.050 414.150 ;
        RECT 506.400 412.950 507.600 425.400 ;
        RECT 524.700 419.400 526.500 431.250 ;
        RECT 528.900 419.400 530.700 431.250 ;
        RECT 539.550 425.400 541.350 431.250 ;
        RECT 542.550 425.400 544.350 431.250 ;
        RECT 545.550 425.400 547.350 431.250 ;
        RECT 560.400 425.400 562.200 431.250 ;
        RECT 521.250 417.150 523.050 418.950 ;
        RECT 520.950 415.050 523.050 417.150 ;
        RECT 524.850 414.150 526.050 419.400 ;
        RECT 542.550 417.150 543.750 425.400 ;
        RECT 563.700 419.400 565.500 431.250 ;
        RECT 567.900 419.400 569.700 431.250 ;
        RECT 584.400 425.400 586.200 431.250 ;
        RECT 587.700 419.400 589.500 431.250 ;
        RECT 591.900 419.400 593.700 431.250 ;
        RECT 608.400 425.400 610.200 431.250 ;
        RECT 611.700 419.400 613.500 431.250 ;
        RECT 615.900 419.400 617.700 431.250 ;
        RECT 626.550 425.400 628.350 431.250 ;
        RECT 629.550 425.400 631.350 431.250 ;
        RECT 632.550 425.400 634.350 431.250 ;
        RECT 644.550 425.400 646.350 431.250 ;
        RECT 647.550 425.400 649.350 431.250 ;
        RECT 560.250 417.150 562.050 418.950 ;
        RECT 530.100 414.150 531.900 415.950 ;
        RECT 505.950 410.850 508.050 412.950 ;
        RECT 509.100 411.150 510.900 412.950 ;
        RECT 523.950 412.050 526.050 414.150 ;
        RECT 489.750 407.400 492.000 408.300 ;
        RECT 489.750 406.500 494.850 407.400 ;
        RECT 487.350 399.750 489.150 405.600 ;
        RECT 490.350 399.750 492.150 405.600 ;
        RECT 493.650 402.600 494.850 406.500 ;
        RECT 506.400 402.600 507.600 410.850 ;
        RECT 508.950 409.050 511.050 411.150 ;
        RECT 523.950 408.750 525.150 412.050 ;
        RECT 526.950 410.850 529.050 412.950 ;
        RECT 529.950 412.050 532.050 414.150 ;
        RECT 538.950 413.850 541.050 415.950 ;
        RECT 541.950 415.050 544.050 417.150 ;
        RECT 539.100 412.050 540.900 413.850 ;
        RECT 527.100 409.050 528.900 410.850 ;
        RECT 521.250 407.700 525.000 408.750 ;
        RECT 542.550 407.700 543.750 415.050 ;
        RECT 544.950 413.850 547.050 415.950 ;
        RECT 559.950 415.050 562.050 417.150 ;
        RECT 563.850 414.150 565.050 419.400 ;
        RECT 584.250 417.150 586.050 418.950 ;
        RECT 569.100 414.150 570.900 415.950 ;
        RECT 583.950 415.050 586.050 417.150 ;
        RECT 587.850 414.150 589.050 419.400 ;
        RECT 608.250 417.150 610.050 418.950 ;
        RECT 593.100 414.150 594.900 415.950 ;
        RECT 607.950 415.050 610.050 417.150 ;
        RECT 611.850 414.150 613.050 419.400 ;
        RECT 629.550 417.150 630.750 425.400 ;
        RECT 617.100 414.150 618.900 415.950 ;
        RECT 545.100 412.050 546.900 413.850 ;
        RECT 562.950 412.050 565.050 414.150 ;
        RECT 562.950 408.750 564.150 412.050 ;
        RECT 565.950 410.850 568.050 412.950 ;
        RECT 568.950 412.050 571.050 414.150 ;
        RECT 586.950 412.050 589.050 414.150 ;
        RECT 566.100 409.050 567.900 410.850 ;
        RECT 586.950 408.750 588.150 412.050 ;
        RECT 589.950 410.850 592.050 412.950 ;
        RECT 592.950 412.050 595.050 414.150 ;
        RECT 610.950 412.050 613.050 414.150 ;
        RECT 590.100 409.050 591.900 410.850 ;
        RECT 610.950 408.750 612.150 412.050 ;
        RECT 613.950 410.850 616.050 412.950 ;
        RECT 616.950 412.050 619.050 414.150 ;
        RECT 625.950 413.850 628.050 415.950 ;
        RECT 628.950 415.050 631.050 417.150 ;
        RECT 626.100 412.050 627.900 413.850 ;
        RECT 614.100 409.050 615.900 410.850 ;
        RECT 560.250 407.700 564.000 408.750 ;
        RECT 584.250 407.700 588.000 408.750 ;
        RECT 608.250 407.700 612.000 408.750 ;
        RECT 629.550 407.700 630.750 415.050 ;
        RECT 631.950 413.850 634.050 415.950 ;
        RECT 632.100 412.050 633.900 413.850 ;
        RECT 647.400 412.950 648.600 425.400 ;
        RECT 660.300 419.400 662.100 431.250 ;
        RECT 664.500 419.400 666.300 431.250 ;
        RECT 667.800 425.400 669.600 431.250 ;
        RECT 682.650 425.400 684.450 431.250 ;
        RECT 685.650 425.400 687.450 431.250 ;
        RECT 688.650 425.400 690.450 431.250 ;
        RECT 700.650 425.400 702.450 431.250 ;
        RECT 703.650 425.400 705.450 431.250 ;
        RECT 706.650 425.400 708.450 431.250 ;
        RECT 659.100 414.150 660.900 415.950 ;
        RECT 664.950 414.150 666.150 419.400 ;
        RECT 667.950 417.150 669.750 418.950 ;
        RECT 686.250 417.150 687.450 425.400 ;
        RECT 704.250 417.150 705.450 425.400 ;
        RECT 717.300 419.400 719.100 431.250 ;
        RECT 721.500 419.400 723.300 431.250 ;
        RECT 724.800 425.400 726.600 431.250 ;
        RECT 731.550 419.400 733.350 431.250 ;
        RECT 734.550 428.400 736.350 431.250 ;
        RECT 739.050 425.400 740.850 431.250 ;
        RECT 743.250 425.400 745.050 431.250 ;
        RECT 736.950 423.300 740.850 425.400 ;
        RECT 747.150 424.500 748.950 431.250 ;
        RECT 750.150 425.400 751.950 431.250 ;
        RECT 754.950 425.400 756.750 431.250 ;
        RECT 760.050 425.400 761.850 431.250 ;
        RECT 755.250 424.500 756.450 425.400 ;
        RECT 745.950 422.700 752.850 424.500 ;
        RECT 755.250 422.400 760.050 424.500 ;
        RECT 738.150 420.600 740.850 422.400 ;
        RECT 741.750 421.800 743.550 422.400 ;
        RECT 741.750 420.900 748.050 421.800 ;
        RECT 755.250 421.500 756.450 422.400 ;
        RECT 741.750 420.600 743.550 420.900 ;
        RECT 739.950 419.700 740.850 420.600 ;
        RECT 667.950 415.050 670.050 417.150 ;
        RECT 644.100 411.150 645.900 412.950 ;
        RECT 643.950 409.050 646.050 411.150 ;
        RECT 646.950 410.850 649.050 412.950 ;
        RECT 658.950 412.050 661.050 414.150 ;
        RECT 661.950 410.850 664.050 412.950 ;
        RECT 664.950 412.050 667.050 414.150 ;
        RECT 682.950 413.850 685.050 415.950 ;
        RECT 685.950 415.050 688.050 417.150 ;
        RECT 683.100 412.050 684.900 413.850 ;
        RECT 521.250 405.600 522.450 407.700 ;
        RECT 542.550 406.800 546.150 407.700 ;
        RECT 493.650 399.750 495.450 402.600 ;
        RECT 505.650 399.750 507.450 402.600 ;
        RECT 508.650 399.750 510.450 402.600 ;
        RECT 520.650 399.750 522.450 405.600 ;
        RECT 523.650 404.700 531.450 406.050 ;
        RECT 523.650 399.750 525.450 404.700 ;
        RECT 526.650 399.750 528.450 403.800 ;
        RECT 529.650 399.750 531.450 404.700 ;
        RECT 539.850 399.750 541.650 405.600 ;
        RECT 544.350 399.750 546.150 406.800 ;
        RECT 560.250 405.600 561.450 407.700 ;
        RECT 559.650 399.750 561.450 405.600 ;
        RECT 562.650 404.700 570.450 406.050 ;
        RECT 584.250 405.600 585.450 407.700 ;
        RECT 562.650 399.750 564.450 404.700 ;
        RECT 565.650 399.750 567.450 403.800 ;
        RECT 568.650 399.750 570.450 404.700 ;
        RECT 583.650 399.750 585.450 405.600 ;
        RECT 586.650 404.700 594.450 406.050 ;
        RECT 608.250 405.600 609.450 407.700 ;
        RECT 629.550 406.800 633.150 407.700 ;
        RECT 586.650 399.750 588.450 404.700 ;
        RECT 589.650 399.750 591.450 403.800 ;
        RECT 592.650 399.750 594.450 404.700 ;
        RECT 607.650 399.750 609.450 405.600 ;
        RECT 610.650 404.700 618.450 406.050 ;
        RECT 610.650 399.750 612.450 404.700 ;
        RECT 613.650 399.750 615.450 403.800 ;
        RECT 616.650 399.750 618.450 404.700 ;
        RECT 626.850 399.750 628.650 405.600 ;
        RECT 631.350 399.750 633.150 406.800 ;
        RECT 647.400 402.600 648.600 410.850 ;
        RECT 662.100 409.050 663.900 410.850 ;
        RECT 665.850 408.750 667.050 412.050 ;
        RECT 666.000 407.700 669.750 408.750 ;
        RECT 686.250 407.700 687.450 415.050 ;
        RECT 688.950 413.850 691.050 415.950 ;
        RECT 700.950 413.850 703.050 415.950 ;
        RECT 703.950 415.050 706.050 417.150 ;
        RECT 689.100 412.050 690.900 413.850 ;
        RECT 701.100 412.050 702.900 413.850 ;
        RECT 704.250 407.700 705.450 415.050 ;
        RECT 706.950 413.850 709.050 415.950 ;
        RECT 716.100 414.150 717.900 415.950 ;
        RECT 721.950 414.150 723.150 419.400 ;
        RECT 724.950 417.150 726.750 418.950 ;
        RECT 724.950 415.050 727.050 417.150 ;
        RECT 707.100 412.050 708.900 413.850 ;
        RECT 715.950 412.050 718.050 414.150 ;
        RECT 718.950 410.850 721.050 412.950 ;
        RECT 721.950 412.050 724.050 414.150 ;
        RECT 719.100 409.050 720.900 410.850 ;
        RECT 722.850 408.750 724.050 412.050 ;
        RECT 731.550 409.950 732.750 419.400 ;
        RECT 736.950 418.800 739.050 419.700 ;
        RECT 739.950 418.800 745.950 419.700 ;
        RECT 734.850 417.600 739.050 418.800 ;
        RECT 733.950 415.800 735.750 417.600 ;
        RECT 745.050 414.150 745.950 418.800 ;
        RECT 747.150 418.800 748.050 420.900 ;
        RECT 748.950 420.300 756.450 421.500 ;
        RECT 748.950 419.700 750.750 420.300 ;
        RECT 763.050 419.400 764.850 431.250 ;
        RECT 753.750 418.800 764.850 419.400 ;
        RECT 747.150 418.200 764.850 418.800 ;
        RECT 747.150 417.900 755.550 418.200 ;
        RECT 753.750 417.600 755.550 417.900 ;
        RECT 745.050 412.050 748.050 414.150 ;
        RECT 751.950 413.100 754.050 414.150 ;
        RECT 751.950 412.050 759.900 413.100 ;
        RECT 733.950 411.750 736.050 412.050 ;
        RECT 733.950 409.950 737.850 411.750 ;
        RECT 723.000 407.700 726.750 408.750 ;
        RECT 659.550 404.700 667.350 406.050 ;
        RECT 644.550 399.750 646.350 402.600 ;
        RECT 647.550 399.750 649.350 402.600 ;
        RECT 659.550 399.750 661.350 404.700 ;
        RECT 662.550 399.750 664.350 403.800 ;
        RECT 665.550 399.750 667.350 404.700 ;
        RECT 668.550 405.600 669.750 407.700 ;
        RECT 683.850 406.800 687.450 407.700 ;
        RECT 701.850 406.800 705.450 407.700 ;
        RECT 668.550 399.750 670.350 405.600 ;
        RECT 683.850 399.750 685.650 406.800 ;
        RECT 688.350 399.750 690.150 405.600 ;
        RECT 701.850 399.750 703.650 406.800 ;
        RECT 706.350 399.750 708.150 405.600 ;
        RECT 716.550 404.700 724.350 406.050 ;
        RECT 716.550 399.750 718.350 404.700 ;
        RECT 719.550 399.750 721.350 403.800 ;
        RECT 722.550 399.750 724.350 404.700 ;
        RECT 725.550 405.600 726.750 407.700 ;
        RECT 731.550 407.850 736.050 409.950 ;
        RECT 745.050 408.000 745.950 412.050 ;
        RECT 758.100 411.300 759.900 412.050 ;
        RECT 761.100 411.150 762.900 412.950 ;
        RECT 755.100 410.400 756.900 411.000 ;
        RECT 761.100 410.400 762.000 411.150 ;
        RECT 755.100 409.200 762.000 410.400 ;
        RECT 755.100 408.000 756.150 409.200 ;
        RECT 731.550 405.600 732.750 407.850 ;
        RECT 745.050 407.100 756.150 408.000 ;
        RECT 745.050 406.800 745.950 407.100 ;
        RECT 725.550 399.750 727.350 405.600 ;
        RECT 731.550 399.750 733.350 405.600 ;
        RECT 736.950 404.700 739.050 405.600 ;
        RECT 744.150 405.000 745.950 406.800 ;
        RECT 755.100 406.200 756.150 407.100 ;
        RECT 751.350 405.450 753.150 406.200 ;
        RECT 736.950 403.500 740.700 404.700 ;
        RECT 739.650 402.600 740.700 403.500 ;
        RECT 748.200 404.400 753.150 405.450 ;
        RECT 754.650 404.400 756.450 406.200 ;
        RECT 763.950 405.600 764.850 418.200 ;
        RECT 773.550 425.400 775.350 431.250 ;
        RECT 773.550 418.500 774.750 425.400 ;
        RECT 776.850 419.400 778.650 431.250 ;
        RECT 779.850 419.400 781.650 431.250 ;
        RECT 791.550 425.400 793.350 431.250 ;
        RECT 773.550 417.600 779.250 418.500 ;
        RECT 777.000 416.700 779.250 417.600 ;
        RECT 773.100 414.150 774.900 415.950 ;
        RECT 772.950 412.050 775.050 414.150 ;
        RECT 777.000 408.300 778.050 416.700 ;
        RECT 780.150 414.150 781.350 419.400 ;
        RECT 791.550 418.500 792.750 425.400 ;
        RECT 794.850 419.400 796.650 431.250 ;
        RECT 797.850 419.400 799.650 431.250 ;
        RECT 811.350 419.400 813.150 431.250 ;
        RECT 814.350 419.400 816.150 431.250 ;
        RECT 817.650 425.400 819.450 431.250 ;
        RECT 791.550 417.600 797.250 418.500 ;
        RECT 795.000 416.700 797.250 417.600 ;
        RECT 791.100 414.150 792.900 415.950 ;
        RECT 778.950 412.050 781.350 414.150 ;
        RECT 790.950 412.050 793.050 414.150 ;
        RECT 777.000 407.400 779.250 408.300 ;
        RECT 748.200 402.600 749.250 404.400 ;
        RECT 757.950 403.500 760.050 405.600 ;
        RECT 757.950 402.600 759.000 403.500 ;
        RECT 734.850 399.750 736.650 402.600 ;
        RECT 739.350 399.750 741.150 402.600 ;
        RECT 743.550 399.750 745.350 402.600 ;
        RECT 747.450 399.750 749.250 402.600 ;
        RECT 750.750 399.750 752.550 402.600 ;
        RECT 755.250 401.700 759.000 402.600 ;
        RECT 755.250 399.750 757.050 401.700 ;
        RECT 760.050 399.750 761.850 402.600 ;
        RECT 763.050 399.750 764.850 405.600 ;
        RECT 774.150 406.500 779.250 407.400 ;
        RECT 774.150 402.600 775.350 406.500 ;
        RECT 780.150 405.600 781.350 412.050 ;
        RECT 795.000 408.300 796.050 416.700 ;
        RECT 798.150 414.150 799.350 419.400 ;
        RECT 796.950 412.050 799.350 414.150 ;
        RECT 795.000 407.400 797.250 408.300 ;
        RECT 792.150 406.500 797.250 407.400 ;
        RECT 773.550 399.750 775.350 402.600 ;
        RECT 776.850 399.750 778.650 405.600 ;
        RECT 779.850 399.750 781.650 405.600 ;
        RECT 792.150 402.600 793.350 406.500 ;
        RECT 798.150 405.600 799.350 412.050 ;
        RECT 811.650 414.150 812.850 419.400 ;
        RECT 818.250 418.500 819.450 425.400 ;
        RECT 813.750 417.600 819.450 418.500 ;
        RECT 822.150 419.400 823.950 431.250 ;
        RECT 825.150 425.400 826.950 431.250 ;
        RECT 830.250 425.400 832.050 431.250 ;
        RECT 835.050 425.400 836.850 431.250 ;
        RECT 830.550 424.500 831.750 425.400 ;
        RECT 838.050 424.500 839.850 431.250 ;
        RECT 841.950 425.400 843.750 431.250 ;
        RECT 846.150 425.400 847.950 431.250 ;
        RECT 850.650 428.400 852.450 431.250 ;
        RECT 826.950 422.400 831.750 424.500 ;
        RECT 834.150 422.700 841.050 424.500 ;
        RECT 846.150 423.300 850.050 425.400 ;
        RECT 830.550 421.500 831.750 422.400 ;
        RECT 843.450 421.800 845.250 422.400 ;
        RECT 830.550 420.300 838.050 421.500 ;
        RECT 836.250 419.700 838.050 420.300 ;
        RECT 838.950 420.900 845.250 421.800 ;
        RECT 822.150 418.800 833.250 419.400 ;
        RECT 838.950 418.800 839.850 420.900 ;
        RECT 843.450 420.600 845.250 420.900 ;
        RECT 846.150 420.600 848.850 422.400 ;
        RECT 846.150 419.700 847.050 420.600 ;
        RECT 822.150 418.200 839.850 418.800 ;
        RECT 813.750 416.700 816.000 417.600 ;
        RECT 811.650 412.050 814.050 414.150 ;
        RECT 811.650 405.600 812.850 412.050 ;
        RECT 814.950 408.300 816.000 416.700 ;
        RECT 818.100 414.150 819.900 415.950 ;
        RECT 817.950 412.050 820.050 414.150 ;
        RECT 813.750 407.400 816.000 408.300 ;
        RECT 813.750 406.500 818.850 407.400 ;
        RECT 791.550 399.750 793.350 402.600 ;
        RECT 794.850 399.750 796.650 405.600 ;
        RECT 797.850 399.750 799.650 405.600 ;
        RECT 811.350 399.750 813.150 405.600 ;
        RECT 814.350 399.750 816.150 405.600 ;
        RECT 817.650 402.600 818.850 406.500 ;
        RECT 822.150 405.600 823.050 418.200 ;
        RECT 831.450 417.900 839.850 418.200 ;
        RECT 841.050 418.800 847.050 419.700 ;
        RECT 847.950 418.800 850.050 419.700 ;
        RECT 853.650 419.400 855.450 431.250 ;
        RECT 863.550 419.400 865.350 431.250 ;
        RECT 867.750 419.400 869.550 431.250 ;
        RECT 831.450 417.600 833.250 417.900 ;
        RECT 841.050 414.150 841.950 418.800 ;
        RECT 847.950 417.600 852.150 418.800 ;
        RECT 851.250 415.800 853.050 417.600 ;
        RECT 832.950 413.100 835.050 414.150 ;
        RECT 824.100 411.150 825.900 412.950 ;
        RECT 827.100 412.050 835.050 413.100 ;
        RECT 838.950 412.050 841.950 414.150 ;
        RECT 827.100 411.300 828.900 412.050 ;
        RECT 825.000 410.400 825.900 411.150 ;
        RECT 830.100 410.400 831.900 411.000 ;
        RECT 825.000 409.200 831.900 410.400 ;
        RECT 830.850 408.000 831.900 409.200 ;
        RECT 841.050 408.000 841.950 412.050 ;
        RECT 850.950 411.750 853.050 412.050 ;
        RECT 849.150 409.950 853.050 411.750 ;
        RECT 854.250 409.950 855.450 419.400 ;
        RECT 867.000 418.350 869.550 419.400 ;
        RECT 863.100 414.150 864.900 415.950 ;
        RECT 862.950 412.050 865.050 414.150 ;
        RECT 867.000 411.150 868.050 418.350 ;
        RECT 869.100 414.150 870.900 415.950 ;
        RECT 868.950 412.050 871.050 414.150 ;
        RECT 830.850 407.100 841.950 408.000 ;
        RECT 850.950 407.850 855.450 409.950 ;
        RECT 865.950 409.050 868.050 411.150 ;
        RECT 830.850 406.200 831.900 407.100 ;
        RECT 841.050 406.800 841.950 407.100 ;
        RECT 817.650 399.750 819.450 402.600 ;
        RECT 822.150 399.750 823.950 405.600 ;
        RECT 826.950 403.500 829.050 405.600 ;
        RECT 830.550 404.400 832.350 406.200 ;
        RECT 833.850 405.450 835.650 406.200 ;
        RECT 833.850 404.400 838.800 405.450 ;
        RECT 841.050 405.000 842.850 406.800 ;
        RECT 854.250 405.600 855.450 407.850 ;
        RECT 847.950 404.700 850.050 405.600 ;
        RECT 828.000 402.600 829.050 403.500 ;
        RECT 837.750 402.600 838.800 404.400 ;
        RECT 846.300 403.500 850.050 404.700 ;
        RECT 846.300 402.600 847.350 403.500 ;
        RECT 825.150 399.750 826.950 402.600 ;
        RECT 828.000 401.700 831.750 402.600 ;
        RECT 829.950 399.750 831.750 401.700 ;
        RECT 834.450 399.750 836.250 402.600 ;
        RECT 837.750 399.750 839.550 402.600 ;
        RECT 841.650 399.750 843.450 402.600 ;
        RECT 845.850 399.750 847.650 402.600 ;
        RECT 850.350 399.750 852.150 402.600 ;
        RECT 853.650 399.750 855.450 405.600 ;
        RECT 867.000 402.600 868.050 409.050 ;
        RECT 863.550 399.750 865.350 402.600 ;
        RECT 866.550 399.750 868.350 402.600 ;
        RECT 869.550 399.750 871.350 402.600 ;
        RECT 11.850 388.200 13.650 395.250 ;
        RECT 16.350 389.400 18.150 395.250 ;
        RECT 31.650 392.400 33.450 395.250 ;
        RECT 34.650 392.400 36.450 395.250 ;
        RECT 11.850 387.300 15.450 388.200 ;
        RECT 11.100 381.150 12.900 382.950 ;
        RECT 10.950 379.050 13.050 381.150 ;
        RECT 14.250 379.950 15.450 387.300 ;
        RECT 32.400 384.150 33.600 392.400 ;
        RECT 47.850 388.200 49.650 395.250 ;
        RECT 52.350 389.400 54.150 395.250 ;
        RECT 67.650 389.400 69.450 395.250 ;
        RECT 47.850 387.300 51.450 388.200 ;
        RECT 17.100 381.150 18.900 382.950 ;
        RECT 31.950 382.050 34.050 384.150 ;
        RECT 34.950 383.850 37.050 385.950 ;
        RECT 35.100 382.050 36.900 383.850 ;
        RECT 13.950 377.850 16.050 379.950 ;
        RECT 16.950 379.050 19.050 381.150 ;
        RECT 14.250 369.600 15.450 377.850 ;
        RECT 32.400 369.600 33.600 382.050 ;
        RECT 47.100 381.150 48.900 382.950 ;
        RECT 46.950 379.050 49.050 381.150 ;
        RECT 50.250 379.950 51.450 387.300 ;
        RECT 68.250 387.300 69.450 389.400 ;
        RECT 70.650 390.300 72.450 395.250 ;
        RECT 73.650 391.200 75.450 395.250 ;
        RECT 76.650 390.300 78.450 395.250 ;
        RECT 70.650 388.950 78.450 390.300 ;
        RECT 88.650 388.200 90.450 395.250 ;
        RECT 93.150 389.700 94.950 394.200 ;
        RECT 97.650 391.200 99.450 395.250 ;
        RECT 100.650 391.200 102.450 394.200 ;
        RECT 92.850 388.800 94.950 389.700 ;
        RECT 68.250 386.250 72.000 387.300 ;
        RECT 70.950 382.950 72.150 386.250 ;
        RECT 74.100 384.150 75.900 385.950 ;
        RECT 92.850 384.150 93.750 388.800 ;
        RECT 100.650 387.900 101.700 391.200 ;
        RECT 115.650 389.400 117.450 395.250 ;
        RECT 95.400 387.000 101.700 387.900 ;
        RECT 116.250 387.300 117.450 389.400 ;
        RECT 118.650 390.300 120.450 395.250 ;
        RECT 121.650 391.200 123.450 395.250 ;
        RECT 124.650 390.300 126.450 395.250 ;
        RECT 134.550 391.200 136.350 394.200 ;
        RECT 137.550 391.200 139.350 395.250 ;
        RECT 118.650 388.950 126.450 390.300 ;
        RECT 135.300 387.900 136.350 391.200 ;
        RECT 142.050 389.700 143.850 394.200 ;
        RECT 142.050 388.800 144.150 389.700 ;
        RECT 53.100 381.150 54.900 382.950 ;
        RECT 49.950 377.850 52.050 379.950 ;
        RECT 52.950 379.050 55.050 381.150 ;
        RECT 70.950 380.850 73.050 382.950 ;
        RECT 73.950 382.050 76.050 384.150 ;
        RECT 76.950 380.850 79.050 382.950 ;
        RECT 88.950 380.850 91.050 382.950 ;
        RECT 91.950 382.050 94.050 384.150 ;
        RECT 67.950 377.850 70.050 379.950 ;
        RECT 50.250 369.600 51.450 377.850 ;
        RECT 68.250 376.050 70.050 377.850 ;
        RECT 71.850 375.600 73.050 380.850 ;
        RECT 77.100 379.050 78.900 380.850 ;
        RECT 89.100 379.050 90.900 380.850 ;
        RECT 10.650 363.750 12.450 369.600 ;
        RECT 13.650 363.750 15.450 369.600 ;
        RECT 16.650 363.750 18.450 369.600 ;
        RECT 31.650 363.750 33.450 369.600 ;
        RECT 34.650 363.750 36.450 369.600 ;
        RECT 46.650 363.750 48.450 369.600 ;
        RECT 49.650 363.750 51.450 369.600 ;
        RECT 52.650 363.750 54.450 369.600 ;
        RECT 68.400 363.750 70.200 369.600 ;
        RECT 71.700 363.750 73.500 375.600 ;
        RECT 75.900 363.750 77.700 375.600 ;
        RECT 88.650 363.750 90.450 375.600 ;
        RECT 92.850 375.000 93.750 382.050 ;
        RECT 95.400 381.300 96.750 387.000 ;
        RECT 116.250 386.250 120.000 387.300 ;
        RECT 135.300 387.000 141.600 387.900 ;
        RECT 100.950 384.150 102.750 385.950 ;
        RECT 94.950 379.500 96.750 381.300 ;
        RECT 95.400 376.800 96.750 379.500 ;
        RECT 97.950 380.850 100.050 382.950 ;
        RECT 100.950 382.050 103.050 384.150 ;
        RECT 118.950 382.950 120.150 386.250 ;
        RECT 122.100 384.150 123.900 385.950 ;
        RECT 134.250 384.150 136.050 385.950 ;
        RECT 118.950 380.850 121.050 382.950 ;
        RECT 121.950 382.050 124.050 384.150 ;
        RECT 124.950 380.850 127.050 382.950 ;
        RECT 133.950 382.050 136.050 384.150 ;
        RECT 136.950 380.850 139.050 382.950 ;
        RECT 97.950 379.050 99.750 380.850 ;
        RECT 115.950 377.850 118.050 379.950 ;
        RECT 95.400 375.900 101.550 376.800 ;
        RECT 116.250 376.050 118.050 377.850 ;
        RECT 92.850 374.100 94.950 375.000 ;
        RECT 93.150 364.800 94.950 374.100 ;
        RECT 100.650 370.800 101.550 375.900 ;
        RECT 119.850 375.600 121.050 380.850 ;
        RECT 125.100 379.050 126.900 380.850 ;
        RECT 137.250 379.050 139.050 380.850 ;
        RECT 140.250 381.300 141.600 387.000 ;
        RECT 143.250 384.150 144.150 388.800 ;
        RECT 146.550 388.200 148.350 395.250 ;
        RECT 161.550 389.400 163.350 395.250 ;
        RECT 164.550 389.400 166.350 395.250 ;
        RECT 167.550 389.400 169.350 395.250 ;
        RECT 170.550 389.400 172.350 395.250 ;
        RECT 173.550 389.400 175.350 395.250 ;
        RECT 185.550 390.300 187.350 395.250 ;
        RECT 188.550 391.200 190.350 395.250 ;
        RECT 191.550 390.300 193.350 395.250 ;
        RECT 164.550 388.500 165.750 389.400 ;
        RECT 170.550 388.500 171.750 389.400 ;
        RECT 185.550 388.950 193.350 390.300 ;
        RECT 194.550 389.400 196.350 395.250 ;
        RECT 206.850 389.400 208.650 395.250 ;
        RECT 164.550 387.300 171.750 388.500 ;
        RECT 194.550 387.300 195.750 389.400 ;
        RECT 211.350 388.200 213.150 395.250 ;
        RECT 227.550 391.200 229.350 394.200 ;
        RECT 230.550 391.200 232.350 395.250 ;
        RECT 142.950 382.050 145.050 384.150 ;
        RECT 170.550 382.950 171.750 387.300 ;
        RECT 192.000 386.250 195.750 387.300 ;
        RECT 209.550 387.300 213.150 388.200 ;
        RECT 228.300 387.900 229.350 391.200 ;
        RECT 235.050 389.700 236.850 394.200 ;
        RECT 235.050 388.800 237.150 389.700 ;
        RECT 188.100 384.150 189.900 385.950 ;
        RECT 140.250 379.500 142.050 381.300 ;
        RECT 140.250 376.800 141.600 379.500 ;
        RECT 135.450 375.900 141.600 376.800 ;
        RECT 97.650 363.750 99.450 370.800 ;
        RECT 100.650 364.800 102.450 370.800 ;
        RECT 116.400 363.750 118.200 369.600 ;
        RECT 119.700 363.750 121.500 375.600 ;
        RECT 123.900 363.750 125.700 375.600 ;
        RECT 135.450 370.800 136.350 375.900 ;
        RECT 143.250 375.000 144.150 382.050 ;
        RECT 145.950 380.850 148.050 382.950 ;
        RECT 163.950 380.850 166.050 382.950 ;
        RECT 169.950 380.850 172.050 382.950 ;
        RECT 184.950 380.850 187.050 382.950 ;
        RECT 187.950 382.050 190.050 384.150 ;
        RECT 191.850 382.950 193.050 386.250 ;
        RECT 190.950 380.850 193.050 382.950 ;
        RECT 206.100 381.150 207.900 382.950 ;
        RECT 146.100 379.050 147.900 380.850 ;
        RECT 164.100 379.050 165.900 380.850 ;
        RECT 170.550 377.400 171.750 380.850 ;
        RECT 185.100 379.050 186.900 380.850 ;
        RECT 164.550 376.500 171.750 377.400 ;
        RECT 142.050 374.100 144.150 375.000 ;
        RECT 134.550 364.800 136.350 370.800 ;
        RECT 137.550 363.750 139.350 370.800 ;
        RECT 142.050 364.800 143.850 374.100 ;
        RECT 146.550 363.750 148.350 375.600 ;
        RECT 161.550 363.750 163.350 375.600 ;
        RECT 164.550 363.750 166.350 376.500 ;
        RECT 170.550 375.600 171.750 376.500 ;
        RECT 190.950 375.600 192.150 380.850 ;
        RECT 193.950 377.850 196.050 379.950 ;
        RECT 205.950 379.050 208.050 381.150 ;
        RECT 209.550 379.950 210.750 387.300 ;
        RECT 228.300 387.000 234.600 387.900 ;
        RECT 227.250 384.150 229.050 385.950 ;
        RECT 212.100 381.150 213.900 382.950 ;
        RECT 226.950 382.050 229.050 384.150 ;
        RECT 208.950 377.850 211.050 379.950 ;
        RECT 211.950 379.050 214.050 381.150 ;
        RECT 229.950 380.850 232.050 382.950 ;
        RECT 230.250 379.050 232.050 380.850 ;
        RECT 233.250 381.300 234.600 387.000 ;
        RECT 236.250 384.150 237.150 388.800 ;
        RECT 239.550 388.200 241.350 395.250 ;
        RECT 251.850 389.400 253.650 395.250 ;
        RECT 256.350 388.200 258.150 395.250 ;
        RECT 269.550 391.200 271.350 394.200 ;
        RECT 272.550 391.200 274.350 395.250 ;
        RECT 254.550 387.300 258.150 388.200 ;
        RECT 270.300 387.900 271.350 391.200 ;
        RECT 277.050 389.700 278.850 394.200 ;
        RECT 277.050 388.800 279.150 389.700 ;
        RECT 235.950 382.050 238.050 384.150 ;
        RECT 233.250 379.500 235.050 381.300 ;
        RECT 193.950 376.050 195.750 377.850 ;
        RECT 167.550 363.750 169.350 375.600 ;
        RECT 170.550 363.750 172.350 375.600 ;
        RECT 173.550 363.750 175.350 375.600 ;
        RECT 186.300 363.750 188.100 375.600 ;
        RECT 190.500 363.750 192.300 375.600 ;
        RECT 209.550 369.600 210.750 377.850 ;
        RECT 233.250 376.800 234.600 379.500 ;
        RECT 228.450 375.900 234.600 376.800 ;
        RECT 228.450 370.800 229.350 375.900 ;
        RECT 236.250 375.000 237.150 382.050 ;
        RECT 238.950 380.850 241.050 382.950 ;
        RECT 251.100 381.150 252.900 382.950 ;
        RECT 239.100 379.050 240.900 380.850 ;
        RECT 250.950 379.050 253.050 381.150 ;
        RECT 254.550 379.950 255.750 387.300 ;
        RECT 270.300 387.000 276.600 387.900 ;
        RECT 269.250 384.150 271.050 385.950 ;
        RECT 257.100 381.150 258.900 382.950 ;
        RECT 268.950 382.050 271.050 384.150 ;
        RECT 253.950 377.850 256.050 379.950 ;
        RECT 256.950 379.050 259.050 381.150 ;
        RECT 271.950 380.850 274.050 382.950 ;
        RECT 272.250 379.050 274.050 380.850 ;
        RECT 275.250 381.300 276.600 387.000 ;
        RECT 278.250 384.150 279.150 388.800 ;
        RECT 281.550 388.200 283.350 395.250 ;
        RECT 296.850 389.400 298.650 395.250 ;
        RECT 301.350 388.200 303.150 395.250 ;
        RECT 299.550 387.300 303.150 388.200 ;
        RECT 277.950 382.050 280.050 384.150 ;
        RECT 275.250 379.500 277.050 381.300 ;
        RECT 235.050 374.100 237.150 375.000 ;
        RECT 193.800 363.750 195.600 369.600 ;
        RECT 206.550 363.750 208.350 369.600 ;
        RECT 209.550 363.750 211.350 369.600 ;
        RECT 212.550 363.750 214.350 369.600 ;
        RECT 227.550 364.800 229.350 370.800 ;
        RECT 230.550 363.750 232.350 370.800 ;
        RECT 235.050 364.800 236.850 374.100 ;
        RECT 239.550 363.750 241.350 375.600 ;
        RECT 254.550 369.600 255.750 377.850 ;
        RECT 275.250 376.800 276.600 379.500 ;
        RECT 270.450 375.900 276.600 376.800 ;
        RECT 270.450 370.800 271.350 375.900 ;
        RECT 278.250 375.000 279.150 382.050 ;
        RECT 280.950 380.850 283.050 382.950 ;
        RECT 296.100 381.150 297.900 382.950 ;
        RECT 281.100 379.050 282.900 380.850 ;
        RECT 295.950 379.050 298.050 381.150 ;
        RECT 299.550 379.950 300.750 387.300 ;
        RECT 320.100 387.000 321.900 395.250 ;
        RECT 317.400 385.350 321.900 387.000 ;
        RECT 325.500 386.400 327.300 395.250 ;
        RECT 341.850 388.200 343.650 395.250 ;
        RECT 346.350 389.400 348.150 395.250 ;
        RECT 358.650 388.200 360.450 395.250 ;
        RECT 363.150 389.700 364.950 394.200 ;
        RECT 367.650 391.200 369.450 395.250 ;
        RECT 370.650 391.200 372.450 394.200 ;
        RECT 380.550 391.200 382.350 394.200 ;
        RECT 383.550 391.200 385.350 395.250 ;
        RECT 362.850 388.800 364.950 389.700 ;
        RECT 341.850 387.300 345.450 388.200 ;
        RECT 302.100 381.150 303.900 382.950 ;
        RECT 317.400 381.150 318.600 385.350 ;
        RECT 341.100 381.150 342.900 382.950 ;
        RECT 298.950 377.850 301.050 379.950 ;
        RECT 301.950 379.050 304.050 381.150 ;
        RECT 316.950 379.050 319.050 381.150 ;
        RECT 277.050 374.100 279.150 375.000 ;
        RECT 251.550 363.750 253.350 369.600 ;
        RECT 254.550 363.750 256.350 369.600 ;
        RECT 257.550 363.750 259.350 369.600 ;
        RECT 269.550 364.800 271.350 370.800 ;
        RECT 272.550 363.750 274.350 370.800 ;
        RECT 277.050 364.800 278.850 374.100 ;
        RECT 281.550 363.750 283.350 375.600 ;
        RECT 299.550 369.600 300.750 377.850 ;
        RECT 317.250 370.800 318.300 379.050 ;
        RECT 319.950 377.850 322.050 379.950 ;
        RECT 325.950 377.850 328.050 379.950 ;
        RECT 340.950 379.050 343.050 381.150 ;
        RECT 344.250 379.950 345.450 387.300 ;
        RECT 362.850 384.150 363.750 388.800 ;
        RECT 370.650 387.900 371.700 391.200 ;
        RECT 365.400 387.000 371.700 387.900 ;
        RECT 381.300 387.900 382.350 391.200 ;
        RECT 388.050 389.700 389.850 394.200 ;
        RECT 388.050 388.800 390.150 389.700 ;
        RECT 381.300 387.000 387.600 387.900 ;
        RECT 347.100 381.150 348.900 382.950 ;
        RECT 343.950 377.850 346.050 379.950 ;
        RECT 346.950 379.050 349.050 381.150 ;
        RECT 358.950 380.850 361.050 382.950 ;
        RECT 361.950 382.050 364.050 384.150 ;
        RECT 359.100 379.050 360.900 380.850 ;
        RECT 319.950 376.050 321.750 377.850 ;
        RECT 322.950 374.850 325.050 376.950 ;
        RECT 326.100 376.050 327.900 377.850 ;
        RECT 323.100 373.050 324.900 374.850 ;
        RECT 317.250 369.900 324.300 370.800 ;
        RECT 317.250 369.600 318.450 369.900 ;
        RECT 296.550 363.750 298.350 369.600 ;
        RECT 299.550 363.750 301.350 369.600 ;
        RECT 302.550 363.750 304.350 369.600 ;
        RECT 316.650 363.750 318.450 369.600 ;
        RECT 322.650 369.600 324.300 369.900 ;
        RECT 344.250 369.600 345.450 377.850 ;
        RECT 319.650 363.750 321.450 369.000 ;
        RECT 322.650 363.750 324.450 369.600 ;
        RECT 325.650 363.750 327.450 369.600 ;
        RECT 340.650 363.750 342.450 369.600 ;
        RECT 343.650 363.750 345.450 369.600 ;
        RECT 346.650 363.750 348.450 369.600 ;
        RECT 358.650 363.750 360.450 375.600 ;
        RECT 362.850 375.000 363.750 382.050 ;
        RECT 365.400 381.300 366.750 387.000 ;
        RECT 370.950 384.150 372.750 385.950 ;
        RECT 380.250 384.150 382.050 385.950 ;
        RECT 364.950 379.500 366.750 381.300 ;
        RECT 365.400 376.800 366.750 379.500 ;
        RECT 367.950 380.850 370.050 382.950 ;
        RECT 370.950 382.050 373.050 384.150 ;
        RECT 379.950 382.050 382.050 384.150 ;
        RECT 382.950 380.850 385.050 382.950 ;
        RECT 367.950 379.050 369.750 380.850 ;
        RECT 383.250 379.050 385.050 380.850 ;
        RECT 386.250 381.300 387.600 387.000 ;
        RECT 389.250 384.150 390.150 388.800 ;
        RECT 392.550 388.200 394.350 395.250 ;
        RECT 407.550 392.400 409.350 395.250 ;
        RECT 408.150 388.500 409.350 392.400 ;
        RECT 410.850 389.400 412.650 395.250 ;
        RECT 413.850 389.400 415.650 395.250 ;
        RECT 425.550 391.200 427.350 394.200 ;
        RECT 428.550 391.200 430.350 395.250 ;
        RECT 408.150 387.600 413.250 388.500 ;
        RECT 411.000 386.700 413.250 387.600 ;
        RECT 388.950 382.050 391.050 384.150 ;
        RECT 386.250 379.500 388.050 381.300 ;
        RECT 386.250 376.800 387.600 379.500 ;
        RECT 365.400 375.900 371.550 376.800 ;
        RECT 362.850 374.100 364.950 375.000 ;
        RECT 363.150 364.800 364.950 374.100 ;
        RECT 370.650 370.800 371.550 375.900 ;
        RECT 381.450 375.900 387.600 376.800 ;
        RECT 381.450 370.800 382.350 375.900 ;
        RECT 389.250 375.000 390.150 382.050 ;
        RECT 391.950 380.850 394.050 382.950 ;
        RECT 406.950 380.850 409.050 382.950 ;
        RECT 392.100 379.050 393.900 380.850 ;
        RECT 407.100 379.050 408.900 380.850 ;
        RECT 411.000 378.300 412.050 386.700 ;
        RECT 414.150 382.950 415.350 389.400 ;
        RECT 426.300 387.900 427.350 391.200 ;
        RECT 433.050 389.700 434.850 394.200 ;
        RECT 433.050 388.800 435.150 389.700 ;
        RECT 426.300 387.000 432.600 387.900 ;
        RECT 425.250 384.150 427.050 385.950 ;
        RECT 412.950 380.850 415.350 382.950 ;
        RECT 424.950 382.050 427.050 384.150 ;
        RECT 427.950 380.850 430.050 382.950 ;
        RECT 411.000 377.400 413.250 378.300 ;
        RECT 407.550 376.500 413.250 377.400 ;
        RECT 388.050 374.100 390.150 375.000 ;
        RECT 367.650 363.750 369.450 370.800 ;
        RECT 370.650 364.800 372.450 370.800 ;
        RECT 380.550 364.800 382.350 370.800 ;
        RECT 383.550 363.750 385.350 370.800 ;
        RECT 388.050 364.800 389.850 374.100 ;
        RECT 392.550 363.750 394.350 375.600 ;
        RECT 407.550 369.600 408.750 376.500 ;
        RECT 414.150 375.600 415.350 380.850 ;
        RECT 428.250 379.050 430.050 380.850 ;
        RECT 431.250 381.300 432.600 387.000 ;
        RECT 434.250 384.150 435.150 388.800 ;
        RECT 437.550 388.200 439.350 395.250 ;
        RECT 451.650 388.200 453.450 395.250 ;
        RECT 456.150 389.700 457.950 394.200 ;
        RECT 460.650 391.200 462.450 395.250 ;
        RECT 463.650 391.200 465.450 394.200 ;
        RECT 476.550 391.200 478.350 394.200 ;
        RECT 479.550 391.200 481.350 395.250 ;
        RECT 455.850 388.800 457.950 389.700 ;
        RECT 455.850 384.150 456.750 388.800 ;
        RECT 463.650 387.900 464.700 391.200 ;
        RECT 458.400 387.000 464.700 387.900 ;
        RECT 477.300 387.900 478.350 391.200 ;
        RECT 484.050 389.700 485.850 394.200 ;
        RECT 484.050 388.800 486.150 389.700 ;
        RECT 477.300 387.000 483.600 387.900 ;
        RECT 433.950 382.050 436.050 384.150 ;
        RECT 431.250 379.500 433.050 381.300 ;
        RECT 431.250 376.800 432.600 379.500 ;
        RECT 426.450 375.900 432.600 376.800 ;
        RECT 407.550 363.750 409.350 369.600 ;
        RECT 410.850 363.750 412.650 375.600 ;
        RECT 413.850 363.750 415.650 375.600 ;
        RECT 426.450 370.800 427.350 375.900 ;
        RECT 434.250 375.000 435.150 382.050 ;
        RECT 436.950 380.850 439.050 382.950 ;
        RECT 451.950 380.850 454.050 382.950 ;
        RECT 454.950 382.050 457.050 384.150 ;
        RECT 437.100 379.050 438.900 380.850 ;
        RECT 452.100 379.050 453.900 380.850 ;
        RECT 433.050 374.100 435.150 375.000 ;
        RECT 425.550 364.800 427.350 370.800 ;
        RECT 428.550 363.750 430.350 370.800 ;
        RECT 433.050 364.800 434.850 374.100 ;
        RECT 437.550 363.750 439.350 375.600 ;
        RECT 451.650 363.750 453.450 375.600 ;
        RECT 455.850 375.000 456.750 382.050 ;
        RECT 458.400 381.300 459.750 387.000 ;
        RECT 463.950 384.150 465.750 385.950 ;
        RECT 476.250 384.150 478.050 385.950 ;
        RECT 457.950 379.500 459.750 381.300 ;
        RECT 458.400 376.800 459.750 379.500 ;
        RECT 460.950 380.850 463.050 382.950 ;
        RECT 463.950 382.050 466.050 384.150 ;
        RECT 475.950 382.050 478.050 384.150 ;
        RECT 478.950 380.850 481.050 382.950 ;
        RECT 460.950 379.050 462.750 380.850 ;
        RECT 479.250 379.050 481.050 380.850 ;
        RECT 482.250 381.300 483.600 387.000 ;
        RECT 485.250 384.150 486.150 388.800 ;
        RECT 488.550 388.200 490.350 395.250 ;
        RECT 503.550 392.400 505.350 395.250 ;
        RECT 504.150 388.500 505.350 392.400 ;
        RECT 506.850 389.400 508.650 395.250 ;
        RECT 509.850 389.400 511.650 395.250 ;
        RECT 524.850 389.400 526.650 395.250 ;
        RECT 504.150 387.600 509.250 388.500 ;
        RECT 507.000 386.700 509.250 387.600 ;
        RECT 484.950 382.050 487.050 384.150 ;
        RECT 482.250 379.500 484.050 381.300 ;
        RECT 482.250 376.800 483.600 379.500 ;
        RECT 458.400 375.900 464.550 376.800 ;
        RECT 455.850 374.100 457.950 375.000 ;
        RECT 456.150 364.800 457.950 374.100 ;
        RECT 463.650 370.800 464.550 375.900 ;
        RECT 477.450 375.900 483.600 376.800 ;
        RECT 477.450 370.800 478.350 375.900 ;
        RECT 485.250 375.000 486.150 382.050 ;
        RECT 487.950 380.850 490.050 382.950 ;
        RECT 502.950 380.850 505.050 382.950 ;
        RECT 488.100 379.050 489.900 380.850 ;
        RECT 503.100 379.050 504.900 380.850 ;
        RECT 507.000 378.300 508.050 386.700 ;
        RECT 510.150 382.950 511.350 389.400 ;
        RECT 529.350 388.200 531.150 395.250 ;
        RECT 547.650 388.200 549.450 395.250 ;
        RECT 552.150 389.700 553.950 394.200 ;
        RECT 556.650 391.200 558.450 395.250 ;
        RECT 559.650 391.200 561.450 394.200 ;
        RECT 551.850 388.800 553.950 389.700 ;
        RECT 527.550 387.300 531.150 388.200 ;
        RECT 508.950 380.850 511.350 382.950 ;
        RECT 524.100 381.150 525.900 382.950 ;
        RECT 507.000 377.400 509.250 378.300 ;
        RECT 503.550 376.500 509.250 377.400 ;
        RECT 484.050 374.100 486.150 375.000 ;
        RECT 460.650 363.750 462.450 370.800 ;
        RECT 463.650 364.800 465.450 370.800 ;
        RECT 476.550 364.800 478.350 370.800 ;
        RECT 479.550 363.750 481.350 370.800 ;
        RECT 484.050 364.800 485.850 374.100 ;
        RECT 488.550 363.750 490.350 375.600 ;
        RECT 503.550 369.600 504.750 376.500 ;
        RECT 510.150 375.600 511.350 380.850 ;
        RECT 523.950 379.050 526.050 381.150 ;
        RECT 527.550 379.950 528.750 387.300 ;
        RECT 551.850 384.150 552.750 388.800 ;
        RECT 559.650 387.900 560.700 391.200 ;
        RECT 574.650 388.200 576.450 395.250 ;
        RECT 579.150 389.700 580.950 394.200 ;
        RECT 583.650 391.200 585.450 395.250 ;
        RECT 586.650 391.200 588.450 394.200 ;
        RECT 578.850 388.800 580.950 389.700 ;
        RECT 554.400 387.000 560.700 387.900 ;
        RECT 530.100 381.150 531.900 382.950 ;
        RECT 526.950 377.850 529.050 379.950 ;
        RECT 529.950 379.050 532.050 381.150 ;
        RECT 547.950 380.850 550.050 382.950 ;
        RECT 550.950 382.050 553.050 384.150 ;
        RECT 548.100 379.050 549.900 380.850 ;
        RECT 503.550 363.750 505.350 369.600 ;
        RECT 506.850 363.750 508.650 375.600 ;
        RECT 509.850 363.750 511.650 375.600 ;
        RECT 527.550 369.600 528.750 377.850 ;
        RECT 524.550 363.750 526.350 369.600 ;
        RECT 527.550 363.750 529.350 369.600 ;
        RECT 530.550 363.750 532.350 369.600 ;
        RECT 547.650 363.750 549.450 375.600 ;
        RECT 551.850 375.000 552.750 382.050 ;
        RECT 554.400 381.300 555.750 387.000 ;
        RECT 559.950 384.150 561.750 385.950 ;
        RECT 578.850 384.150 579.750 388.800 ;
        RECT 586.650 387.900 587.700 391.200 ;
        RECT 581.400 387.000 587.700 387.900 ;
        RECT 599.850 388.200 601.650 395.250 ;
        RECT 604.350 389.400 606.150 395.250 ;
        RECT 616.650 392.400 618.450 395.250 ;
        RECT 619.650 392.400 621.450 395.250 ;
        RECT 622.650 392.400 624.450 395.250 ;
        RECT 637.650 392.400 639.450 395.250 ;
        RECT 640.650 392.400 642.450 395.250 ;
        RECT 599.850 387.300 603.450 388.200 ;
        RECT 553.950 379.500 555.750 381.300 ;
        RECT 554.400 376.800 555.750 379.500 ;
        RECT 556.950 380.850 559.050 382.950 ;
        RECT 559.950 382.050 562.050 384.150 ;
        RECT 574.950 380.850 577.050 382.950 ;
        RECT 577.950 382.050 580.050 384.150 ;
        RECT 556.950 379.050 558.750 380.850 ;
        RECT 575.100 379.050 576.900 380.850 ;
        RECT 554.400 375.900 560.550 376.800 ;
        RECT 551.850 374.100 553.950 375.000 ;
        RECT 552.150 364.800 553.950 374.100 ;
        RECT 559.650 370.800 560.550 375.900 ;
        RECT 556.650 363.750 558.450 370.800 ;
        RECT 559.650 364.800 561.450 370.800 ;
        RECT 574.650 363.750 576.450 375.600 ;
        RECT 578.850 375.000 579.750 382.050 ;
        RECT 581.400 381.300 582.750 387.000 ;
        RECT 586.950 384.150 588.750 385.950 ;
        RECT 580.950 379.500 582.750 381.300 ;
        RECT 581.400 376.800 582.750 379.500 ;
        RECT 583.950 380.850 586.050 382.950 ;
        RECT 586.950 382.050 589.050 384.150 ;
        RECT 599.100 381.150 600.900 382.950 ;
        RECT 583.950 379.050 585.750 380.850 ;
        RECT 598.950 379.050 601.050 381.150 ;
        RECT 602.250 379.950 603.450 387.300 ;
        RECT 619.950 385.950 621.000 392.400 ;
        RECT 619.950 383.850 622.050 385.950 ;
        RECT 638.400 384.150 639.600 392.400 ;
        RECT 656.850 388.200 658.650 395.250 ;
        RECT 661.350 389.400 663.150 395.250 ;
        RECT 673.650 389.400 675.450 395.250 ;
        RECT 656.850 387.300 660.450 388.200 ;
        RECT 605.100 381.150 606.900 382.950 ;
        RECT 601.950 377.850 604.050 379.950 ;
        RECT 604.950 379.050 607.050 381.150 ;
        RECT 616.950 380.850 619.050 382.950 ;
        RECT 617.100 379.050 618.900 380.850 ;
        RECT 581.400 375.900 587.550 376.800 ;
        RECT 578.850 374.100 580.950 375.000 ;
        RECT 579.150 364.800 580.950 374.100 ;
        RECT 586.650 370.800 587.550 375.900 ;
        RECT 583.650 363.750 585.450 370.800 ;
        RECT 586.650 364.800 588.450 370.800 ;
        RECT 602.250 369.600 603.450 377.850 ;
        RECT 619.950 376.650 621.000 383.850 ;
        RECT 622.950 380.850 625.050 382.950 ;
        RECT 637.950 382.050 640.050 384.150 ;
        RECT 640.950 383.850 643.050 385.950 ;
        RECT 641.100 382.050 642.900 383.850 ;
        RECT 623.100 379.050 624.900 380.850 ;
        RECT 618.450 375.600 621.000 376.650 ;
        RECT 598.650 363.750 600.450 369.600 ;
        RECT 601.650 363.750 603.450 369.600 ;
        RECT 604.650 363.750 606.450 369.600 ;
        RECT 618.450 363.750 620.250 375.600 ;
        RECT 622.650 363.750 624.450 375.600 ;
        RECT 638.400 369.600 639.600 382.050 ;
        RECT 656.100 381.150 657.900 382.950 ;
        RECT 655.950 379.050 658.050 381.150 ;
        RECT 659.250 379.950 660.450 387.300 ;
        RECT 674.250 387.300 675.450 389.400 ;
        RECT 676.650 390.300 678.450 395.250 ;
        RECT 679.650 391.200 681.450 395.250 ;
        RECT 682.650 390.300 684.450 395.250 ;
        RECT 676.650 388.950 684.450 390.300 ;
        RECT 686.550 389.400 688.350 395.250 ;
        RECT 689.850 392.400 691.650 395.250 ;
        RECT 694.350 392.400 696.150 395.250 ;
        RECT 698.550 392.400 700.350 395.250 ;
        RECT 702.450 392.400 704.250 395.250 ;
        RECT 705.750 392.400 707.550 395.250 ;
        RECT 710.250 393.300 712.050 395.250 ;
        RECT 710.250 392.400 714.000 393.300 ;
        RECT 715.050 392.400 716.850 395.250 ;
        RECT 694.650 391.500 695.700 392.400 ;
        RECT 691.950 390.300 695.700 391.500 ;
        RECT 703.200 390.600 704.250 392.400 ;
        RECT 712.950 391.500 714.000 392.400 ;
        RECT 691.950 389.400 694.050 390.300 ;
        RECT 674.250 386.250 678.000 387.300 ;
        RECT 686.550 387.150 687.750 389.400 ;
        RECT 699.150 388.200 700.950 390.000 ;
        RECT 703.200 389.550 708.150 390.600 ;
        RECT 706.350 388.800 708.150 389.550 ;
        RECT 709.650 388.800 711.450 390.600 ;
        RECT 712.950 389.400 715.050 391.500 ;
        RECT 718.050 389.400 719.850 395.250 ;
        RECT 730.350 389.400 732.150 395.250 ;
        RECT 733.350 389.400 735.150 395.250 ;
        RECT 736.650 392.400 738.450 395.250 ;
        RECT 700.050 387.900 700.950 388.200 ;
        RECT 710.100 387.900 711.150 388.800 ;
        RECT 676.950 382.950 678.150 386.250 ;
        RECT 680.100 384.150 681.900 385.950 ;
        RECT 686.550 385.050 691.050 387.150 ;
        RECT 700.050 387.000 711.150 387.900 ;
        RECT 662.100 381.150 663.900 382.950 ;
        RECT 658.950 377.850 661.050 379.950 ;
        RECT 661.950 379.050 664.050 381.150 ;
        RECT 676.950 380.850 679.050 382.950 ;
        RECT 679.950 382.050 682.050 384.150 ;
        RECT 682.950 380.850 685.050 382.950 ;
        RECT 673.950 377.850 676.050 379.950 ;
        RECT 659.250 369.600 660.450 377.850 ;
        RECT 674.250 376.050 676.050 377.850 ;
        RECT 677.850 375.600 679.050 380.850 ;
        RECT 683.100 379.050 684.900 380.850 ;
        RECT 686.550 375.600 687.750 385.050 ;
        RECT 688.950 383.250 692.850 385.050 ;
        RECT 688.950 382.950 691.050 383.250 ;
        RECT 700.050 382.950 700.950 387.000 ;
        RECT 710.100 385.800 711.150 387.000 ;
        RECT 710.100 384.600 717.000 385.800 ;
        RECT 710.100 384.000 711.900 384.600 ;
        RECT 716.100 383.850 717.000 384.600 ;
        RECT 713.100 382.950 714.900 383.700 ;
        RECT 700.050 380.850 703.050 382.950 ;
        RECT 706.950 381.900 714.900 382.950 ;
        RECT 716.100 382.050 717.900 383.850 ;
        RECT 706.950 380.850 709.050 381.900 ;
        RECT 688.950 377.400 690.750 379.200 ;
        RECT 689.850 376.200 694.050 377.400 ;
        RECT 700.050 376.200 700.950 380.850 ;
        RECT 708.750 377.100 710.550 377.400 ;
        RECT 637.650 363.750 639.450 369.600 ;
        RECT 640.650 363.750 642.450 369.600 ;
        RECT 655.650 363.750 657.450 369.600 ;
        RECT 658.650 363.750 660.450 369.600 ;
        RECT 661.650 363.750 663.450 369.600 ;
        RECT 674.400 363.750 676.200 369.600 ;
        RECT 677.700 363.750 679.500 375.600 ;
        RECT 681.900 363.750 683.700 375.600 ;
        RECT 686.550 363.750 688.350 375.600 ;
        RECT 691.950 375.300 694.050 376.200 ;
        RECT 694.950 375.300 700.950 376.200 ;
        RECT 702.150 376.800 710.550 377.100 ;
        RECT 718.950 376.800 719.850 389.400 ;
        RECT 702.150 376.200 719.850 376.800 ;
        RECT 694.950 374.400 695.850 375.300 ;
        RECT 693.150 372.600 695.850 374.400 ;
        RECT 696.750 374.100 698.550 374.400 ;
        RECT 702.150 374.100 703.050 376.200 ;
        RECT 708.750 375.600 719.850 376.200 ;
        RECT 730.650 382.950 731.850 389.400 ;
        RECT 736.650 388.500 737.850 392.400 ;
        RECT 732.750 387.600 737.850 388.500 ;
        RECT 740.550 389.400 742.350 395.250 ;
        RECT 743.850 392.400 745.650 395.250 ;
        RECT 748.350 392.400 750.150 395.250 ;
        RECT 752.550 392.400 754.350 395.250 ;
        RECT 756.450 392.400 758.250 395.250 ;
        RECT 759.750 392.400 761.550 395.250 ;
        RECT 764.250 393.300 766.050 395.250 ;
        RECT 764.250 392.400 768.000 393.300 ;
        RECT 769.050 392.400 770.850 395.250 ;
        RECT 748.650 391.500 749.700 392.400 ;
        RECT 745.950 390.300 749.700 391.500 ;
        RECT 757.200 390.600 758.250 392.400 ;
        RECT 766.950 391.500 768.000 392.400 ;
        RECT 745.950 389.400 748.050 390.300 ;
        RECT 732.750 386.700 735.000 387.600 ;
        RECT 730.650 380.850 733.050 382.950 ;
        RECT 730.650 375.600 731.850 380.850 ;
        RECT 733.950 378.300 735.000 386.700 ;
        RECT 740.550 387.150 741.750 389.400 ;
        RECT 753.150 388.200 754.950 390.000 ;
        RECT 757.200 389.550 762.150 390.600 ;
        RECT 760.350 388.800 762.150 389.550 ;
        RECT 763.650 388.800 765.450 390.600 ;
        RECT 766.950 389.400 769.050 391.500 ;
        RECT 772.050 389.400 773.850 395.250 ;
        RECT 754.050 387.900 754.950 388.200 ;
        RECT 764.100 387.900 765.150 388.800 ;
        RECT 740.550 385.050 745.050 387.150 ;
        RECT 754.050 387.000 765.150 387.900 ;
        RECT 736.950 380.850 739.050 382.950 ;
        RECT 737.100 379.050 738.900 380.850 ;
        RECT 732.750 377.400 735.000 378.300 ;
        RECT 732.750 376.500 738.450 377.400 ;
        RECT 696.750 373.200 703.050 374.100 ;
        RECT 703.950 374.700 705.750 375.300 ;
        RECT 703.950 373.500 711.450 374.700 ;
        RECT 696.750 372.600 698.550 373.200 ;
        RECT 710.250 372.600 711.450 373.500 ;
        RECT 691.950 369.600 695.850 371.700 ;
        RECT 700.950 370.500 707.850 372.300 ;
        RECT 710.250 370.500 715.050 372.600 ;
        RECT 689.550 363.750 691.350 366.600 ;
        RECT 694.050 363.750 695.850 369.600 ;
        RECT 698.250 363.750 700.050 369.600 ;
        RECT 702.150 363.750 703.950 370.500 ;
        RECT 710.250 369.600 711.450 370.500 ;
        RECT 705.150 363.750 706.950 369.600 ;
        RECT 709.950 363.750 711.750 369.600 ;
        RECT 715.050 363.750 716.850 369.600 ;
        RECT 718.050 363.750 719.850 375.600 ;
        RECT 730.350 363.750 732.150 375.600 ;
        RECT 733.350 363.750 735.150 375.600 ;
        RECT 737.250 369.600 738.450 376.500 ;
        RECT 736.650 363.750 738.450 369.600 ;
        RECT 740.550 375.600 741.750 385.050 ;
        RECT 742.950 383.250 746.850 385.050 ;
        RECT 742.950 382.950 745.050 383.250 ;
        RECT 754.050 382.950 754.950 387.000 ;
        RECT 764.100 385.800 765.150 387.000 ;
        RECT 764.100 384.600 771.000 385.800 ;
        RECT 764.100 384.000 765.900 384.600 ;
        RECT 770.100 383.850 771.000 384.600 ;
        RECT 767.100 382.950 768.900 383.700 ;
        RECT 754.050 380.850 757.050 382.950 ;
        RECT 760.950 381.900 768.900 382.950 ;
        RECT 770.100 382.050 771.900 383.850 ;
        RECT 760.950 380.850 763.050 381.900 ;
        RECT 742.950 377.400 744.750 379.200 ;
        RECT 743.850 376.200 748.050 377.400 ;
        RECT 754.050 376.200 754.950 380.850 ;
        RECT 762.750 377.100 764.550 377.400 ;
        RECT 740.550 363.750 742.350 375.600 ;
        RECT 745.950 375.300 748.050 376.200 ;
        RECT 748.950 375.300 754.950 376.200 ;
        RECT 756.150 376.800 764.550 377.100 ;
        RECT 772.950 376.800 773.850 389.400 ;
        RECT 756.150 376.200 773.850 376.800 ;
        RECT 748.950 374.400 749.850 375.300 ;
        RECT 747.150 372.600 749.850 374.400 ;
        RECT 750.750 374.100 752.550 374.400 ;
        RECT 756.150 374.100 757.050 376.200 ;
        RECT 762.750 375.600 773.850 376.200 ;
        RECT 750.750 373.200 757.050 374.100 ;
        RECT 757.950 374.700 759.750 375.300 ;
        RECT 757.950 373.500 765.450 374.700 ;
        RECT 750.750 372.600 752.550 373.200 ;
        RECT 764.250 372.600 765.450 373.500 ;
        RECT 745.950 369.600 749.850 371.700 ;
        RECT 754.950 370.500 761.850 372.300 ;
        RECT 764.250 370.500 769.050 372.600 ;
        RECT 743.550 363.750 745.350 366.600 ;
        RECT 748.050 363.750 749.850 369.600 ;
        RECT 752.250 363.750 754.050 369.600 ;
        RECT 756.150 363.750 757.950 370.500 ;
        RECT 764.250 369.600 765.450 370.500 ;
        RECT 759.150 363.750 760.950 369.600 ;
        RECT 763.950 363.750 765.750 369.600 ;
        RECT 769.050 363.750 770.850 369.600 ;
        RECT 772.050 363.750 773.850 375.600 ;
        RECT 776.550 389.400 778.350 395.250 ;
        RECT 779.850 392.400 781.650 395.250 ;
        RECT 784.350 392.400 786.150 395.250 ;
        RECT 788.550 392.400 790.350 395.250 ;
        RECT 792.450 392.400 794.250 395.250 ;
        RECT 795.750 392.400 797.550 395.250 ;
        RECT 800.250 393.300 802.050 395.250 ;
        RECT 800.250 392.400 804.000 393.300 ;
        RECT 805.050 392.400 806.850 395.250 ;
        RECT 784.650 391.500 785.700 392.400 ;
        RECT 781.950 390.300 785.700 391.500 ;
        RECT 793.200 390.600 794.250 392.400 ;
        RECT 802.950 391.500 804.000 392.400 ;
        RECT 781.950 389.400 784.050 390.300 ;
        RECT 776.550 387.150 777.750 389.400 ;
        RECT 789.150 388.200 790.950 390.000 ;
        RECT 793.200 389.550 798.150 390.600 ;
        RECT 796.350 388.800 798.150 389.550 ;
        RECT 799.650 388.800 801.450 390.600 ;
        RECT 802.950 389.400 805.050 391.500 ;
        RECT 808.050 389.400 809.850 395.250 ;
        RECT 820.650 389.400 822.450 395.250 ;
        RECT 790.050 387.900 790.950 388.200 ;
        RECT 800.100 387.900 801.150 388.800 ;
        RECT 776.550 385.050 781.050 387.150 ;
        RECT 790.050 387.000 801.150 387.900 ;
        RECT 776.550 375.600 777.750 385.050 ;
        RECT 778.950 383.250 782.850 385.050 ;
        RECT 778.950 382.950 781.050 383.250 ;
        RECT 790.050 382.950 790.950 387.000 ;
        RECT 800.100 385.800 801.150 387.000 ;
        RECT 800.100 384.600 807.000 385.800 ;
        RECT 800.100 384.000 801.900 384.600 ;
        RECT 806.100 383.850 807.000 384.600 ;
        RECT 803.100 382.950 804.900 383.700 ;
        RECT 790.050 380.850 793.050 382.950 ;
        RECT 796.950 381.900 804.900 382.950 ;
        RECT 806.100 382.050 807.900 383.850 ;
        RECT 796.950 380.850 799.050 381.900 ;
        RECT 778.950 377.400 780.750 379.200 ;
        RECT 779.850 376.200 784.050 377.400 ;
        RECT 790.050 376.200 790.950 380.850 ;
        RECT 798.750 377.100 800.550 377.400 ;
        RECT 776.550 363.750 778.350 375.600 ;
        RECT 781.950 375.300 784.050 376.200 ;
        RECT 784.950 375.300 790.950 376.200 ;
        RECT 792.150 376.800 800.550 377.100 ;
        RECT 808.950 376.800 809.850 389.400 ;
        RECT 821.250 387.300 822.450 389.400 ;
        RECT 823.650 390.300 825.450 395.250 ;
        RECT 826.650 391.200 828.450 395.250 ;
        RECT 829.650 390.300 831.450 395.250 ;
        RECT 841.650 392.400 843.450 395.250 ;
        RECT 844.650 392.400 846.450 395.250 ;
        RECT 823.650 388.950 831.450 390.300 ;
        RECT 821.250 386.250 825.000 387.300 ;
        RECT 823.950 382.950 825.150 386.250 ;
        RECT 827.100 384.150 828.900 385.950 ;
        RECT 842.400 384.150 843.600 392.400 ;
        RECT 848.550 389.400 850.350 395.250 ;
        RECT 851.850 392.400 853.650 395.250 ;
        RECT 856.350 392.400 858.150 395.250 ;
        RECT 860.550 392.400 862.350 395.250 ;
        RECT 864.450 392.400 866.250 395.250 ;
        RECT 867.750 392.400 869.550 395.250 ;
        RECT 872.250 393.300 874.050 395.250 ;
        RECT 872.250 392.400 876.000 393.300 ;
        RECT 877.050 392.400 878.850 395.250 ;
        RECT 856.650 391.500 857.700 392.400 ;
        RECT 853.950 390.300 857.700 391.500 ;
        RECT 865.200 390.600 866.250 392.400 ;
        RECT 874.950 391.500 876.000 392.400 ;
        RECT 853.950 389.400 856.050 390.300 ;
        RECT 848.550 387.150 849.750 389.400 ;
        RECT 861.150 388.200 862.950 390.000 ;
        RECT 865.200 389.550 870.150 390.600 ;
        RECT 868.350 388.800 870.150 389.550 ;
        RECT 871.650 388.800 873.450 390.600 ;
        RECT 874.950 389.400 877.050 391.500 ;
        RECT 880.050 389.400 881.850 395.250 ;
        RECT 862.050 387.900 862.950 388.200 ;
        RECT 872.100 387.900 873.150 388.800 ;
        RECT 823.950 380.850 826.050 382.950 ;
        RECT 826.950 382.050 829.050 384.150 ;
        RECT 829.950 380.850 832.050 382.950 ;
        RECT 841.950 382.050 844.050 384.150 ;
        RECT 844.950 383.850 847.050 385.950 ;
        RECT 848.550 385.050 853.050 387.150 ;
        RECT 862.050 387.000 873.150 387.900 ;
        RECT 845.100 382.050 846.900 383.850 ;
        RECT 820.950 377.850 823.050 379.950 ;
        RECT 792.150 376.200 809.850 376.800 ;
        RECT 784.950 374.400 785.850 375.300 ;
        RECT 783.150 372.600 785.850 374.400 ;
        RECT 786.750 374.100 788.550 374.400 ;
        RECT 792.150 374.100 793.050 376.200 ;
        RECT 798.750 375.600 809.850 376.200 ;
        RECT 821.250 376.050 823.050 377.850 ;
        RECT 824.850 375.600 826.050 380.850 ;
        RECT 830.100 379.050 831.900 380.850 ;
        RECT 786.750 373.200 793.050 374.100 ;
        RECT 793.950 374.700 795.750 375.300 ;
        RECT 793.950 373.500 801.450 374.700 ;
        RECT 786.750 372.600 788.550 373.200 ;
        RECT 800.250 372.600 801.450 373.500 ;
        RECT 781.950 369.600 785.850 371.700 ;
        RECT 790.950 370.500 797.850 372.300 ;
        RECT 800.250 370.500 805.050 372.600 ;
        RECT 779.550 363.750 781.350 366.600 ;
        RECT 784.050 363.750 785.850 369.600 ;
        RECT 788.250 363.750 790.050 369.600 ;
        RECT 792.150 363.750 793.950 370.500 ;
        RECT 800.250 369.600 801.450 370.500 ;
        RECT 795.150 363.750 796.950 369.600 ;
        RECT 799.950 363.750 801.750 369.600 ;
        RECT 805.050 363.750 806.850 369.600 ;
        RECT 808.050 363.750 809.850 375.600 ;
        RECT 821.400 363.750 823.200 369.600 ;
        RECT 824.700 363.750 826.500 375.600 ;
        RECT 828.900 363.750 830.700 375.600 ;
        RECT 842.400 369.600 843.600 382.050 ;
        RECT 848.550 375.600 849.750 385.050 ;
        RECT 850.950 383.250 854.850 385.050 ;
        RECT 850.950 382.950 853.050 383.250 ;
        RECT 862.050 382.950 862.950 387.000 ;
        RECT 872.100 385.800 873.150 387.000 ;
        RECT 872.100 384.600 879.000 385.800 ;
        RECT 872.100 384.000 873.900 384.600 ;
        RECT 878.100 383.850 879.000 384.600 ;
        RECT 875.100 382.950 876.900 383.700 ;
        RECT 862.050 380.850 865.050 382.950 ;
        RECT 868.950 381.900 876.900 382.950 ;
        RECT 878.100 382.050 879.900 383.850 ;
        RECT 868.950 380.850 871.050 381.900 ;
        RECT 850.950 377.400 852.750 379.200 ;
        RECT 851.850 376.200 856.050 377.400 ;
        RECT 862.050 376.200 862.950 380.850 ;
        RECT 870.750 377.100 872.550 377.400 ;
        RECT 841.650 363.750 843.450 369.600 ;
        RECT 844.650 363.750 846.450 369.600 ;
        RECT 848.550 363.750 850.350 375.600 ;
        RECT 853.950 375.300 856.050 376.200 ;
        RECT 856.950 375.300 862.950 376.200 ;
        RECT 864.150 376.800 872.550 377.100 ;
        RECT 880.950 376.800 881.850 389.400 ;
        RECT 864.150 376.200 881.850 376.800 ;
        RECT 856.950 374.400 857.850 375.300 ;
        RECT 855.150 372.600 857.850 374.400 ;
        RECT 858.750 374.100 860.550 374.400 ;
        RECT 864.150 374.100 865.050 376.200 ;
        RECT 870.750 375.600 881.850 376.200 ;
        RECT 858.750 373.200 865.050 374.100 ;
        RECT 865.950 374.700 867.750 375.300 ;
        RECT 865.950 373.500 873.450 374.700 ;
        RECT 858.750 372.600 860.550 373.200 ;
        RECT 872.250 372.600 873.450 373.500 ;
        RECT 853.950 369.600 857.850 371.700 ;
        RECT 862.950 370.500 869.850 372.300 ;
        RECT 872.250 370.500 877.050 372.600 ;
        RECT 851.550 363.750 853.350 366.600 ;
        RECT 856.050 363.750 857.850 369.600 ;
        RECT 860.250 363.750 862.050 369.600 ;
        RECT 864.150 363.750 865.950 370.500 ;
        RECT 872.250 369.600 873.450 370.500 ;
        RECT 867.150 363.750 868.950 369.600 ;
        RECT 871.950 363.750 873.750 369.600 ;
        RECT 877.050 363.750 878.850 369.600 ;
        RECT 880.050 363.750 881.850 375.600 ;
        RECT 13.650 353.400 15.450 359.250 ;
        RECT 16.650 353.400 18.450 359.250 ;
        RECT 14.400 340.950 15.600 353.400 ;
        RECT 31.650 347.400 33.450 359.250 ;
        RECT 34.650 348.300 36.450 359.250 ;
        RECT 37.650 349.200 39.450 359.250 ;
        RECT 40.650 348.300 42.450 359.250 ;
        RECT 34.650 347.400 42.450 348.300 ;
        RECT 52.650 347.400 54.450 359.250 ;
        RECT 55.650 348.300 57.450 359.250 ;
        RECT 58.650 349.200 60.450 359.250 ;
        RECT 61.650 348.300 63.450 359.250 ;
        RECT 75.150 348.900 76.950 359.250 ;
        RECT 55.650 347.400 63.450 348.300 ;
        RECT 74.550 347.550 76.950 348.900 ;
        RECT 78.150 347.550 79.950 359.250 ;
        RECT 32.100 342.150 33.300 347.400 ;
        RECT 53.100 342.150 54.300 347.400 ;
        RECT 13.950 338.850 16.050 340.950 ;
        RECT 17.100 339.150 18.900 340.950 ;
        RECT 31.950 340.050 34.050 342.150 ;
        RECT 14.400 330.600 15.600 338.850 ;
        RECT 16.950 337.050 19.050 339.150 ;
        RECT 32.100 333.600 33.300 340.050 ;
        RECT 34.950 338.850 37.050 340.950 ;
        RECT 38.100 339.150 39.900 340.950 ;
        RECT 35.100 337.050 36.900 338.850 ;
        RECT 37.950 337.050 40.050 339.150 ;
        RECT 40.950 338.850 43.050 340.950 ;
        RECT 52.950 340.050 55.050 342.150 ;
        RECT 74.550 340.950 75.900 347.550 ;
        RECT 82.650 347.400 84.450 359.250 ;
        RECT 93.300 347.400 95.100 359.250 ;
        RECT 97.500 347.400 99.300 359.250 ;
        RECT 100.800 353.400 102.600 359.250 ;
        RECT 117.300 347.400 119.100 359.250 ;
        RECT 121.500 347.400 123.300 359.250 ;
        RECT 124.800 353.400 126.600 359.250 ;
        RECT 141.450 347.400 143.250 359.250 ;
        RECT 145.650 347.400 147.450 359.250 ;
        RECT 158.400 353.400 160.200 359.250 ;
        RECT 161.700 347.400 163.500 359.250 ;
        RECT 165.900 347.400 167.700 359.250 ;
        RECT 176.550 353.400 178.350 359.250 ;
        RECT 77.250 346.200 79.050 346.650 ;
        RECT 83.250 346.200 84.450 347.400 ;
        RECT 77.250 345.000 84.450 346.200 ;
        RECT 77.250 344.850 79.050 345.000 ;
        RECT 41.100 337.050 42.900 338.850 ;
        RECT 53.100 333.600 54.300 340.050 ;
        RECT 55.950 338.850 58.050 340.950 ;
        RECT 59.100 339.150 60.900 340.950 ;
        RECT 56.100 337.050 57.900 338.850 ;
        RECT 58.950 337.050 61.050 339.150 ;
        RECT 61.950 338.850 64.050 340.950 ;
        RECT 73.950 338.850 76.050 340.950 ;
        RECT 62.100 337.050 63.900 338.850 ;
        RECT 73.950 333.600 75.000 338.850 ;
        RECT 77.400 336.600 78.300 344.850 ;
        RECT 80.100 342.150 81.900 343.950 ;
        RECT 92.100 342.150 93.900 343.950 ;
        RECT 97.950 342.150 99.150 347.400 ;
        RECT 100.950 345.150 102.750 346.950 ;
        RECT 100.950 343.050 103.050 345.150 ;
        RECT 116.100 342.150 117.900 343.950 ;
        RECT 121.950 342.150 123.150 347.400 ;
        RECT 124.950 345.150 126.750 346.950 ;
        RECT 141.450 346.350 144.000 347.400 ;
        RECT 124.950 343.050 127.050 345.150 ;
        RECT 140.100 342.150 141.900 343.950 ;
        RECT 79.950 340.050 82.050 342.150 ;
        RECT 83.100 339.150 84.900 340.950 ;
        RECT 91.950 340.050 94.050 342.150 ;
        RECT 82.950 337.050 85.050 339.150 ;
        RECT 94.950 338.850 97.050 340.950 ;
        RECT 97.950 340.050 100.050 342.150 ;
        RECT 115.950 340.050 118.050 342.150 ;
        RECT 95.100 337.050 96.900 338.850 ;
        RECT 98.850 336.750 100.050 340.050 ;
        RECT 118.950 338.850 121.050 340.950 ;
        RECT 121.950 340.050 124.050 342.150 ;
        RECT 139.950 340.050 142.050 342.150 ;
        RECT 119.100 337.050 120.900 338.850 ;
        RECT 122.850 336.750 124.050 340.050 ;
        RECT 142.950 339.150 144.000 346.350 ;
        RECT 158.250 345.150 160.050 346.950 ;
        RECT 146.100 342.150 147.900 343.950 ;
        RECT 157.950 343.050 160.050 345.150 ;
        RECT 161.850 342.150 163.050 347.400 ;
        RECT 176.550 346.500 177.750 353.400 ;
        RECT 179.850 347.400 181.650 359.250 ;
        RECT 182.850 347.400 184.650 359.250 ;
        RECT 199.350 347.400 201.150 359.250 ;
        RECT 202.350 347.400 204.150 359.250 ;
        RECT 205.650 353.400 207.450 359.250 ;
        RECT 176.550 345.600 182.250 346.500 ;
        RECT 180.000 344.700 182.250 345.600 ;
        RECT 167.100 342.150 168.900 343.950 ;
        RECT 176.100 342.150 177.900 343.950 ;
        RECT 145.950 340.050 148.050 342.150 ;
        RECT 160.950 340.050 163.050 342.150 ;
        RECT 142.950 337.050 145.050 339.150 ;
        RECT 77.250 335.700 79.050 336.600 ;
        RECT 99.000 335.700 102.750 336.750 ;
        RECT 123.000 335.700 126.750 336.750 ;
        RECT 77.250 334.800 80.550 335.700 ;
        RECT 32.100 331.950 37.800 333.600 ;
        RECT 13.650 327.750 15.450 330.600 ;
        RECT 16.650 327.750 18.450 330.600 ;
        RECT 32.700 327.750 34.500 330.600 ;
        RECT 36.000 327.750 37.800 331.950 ;
        RECT 40.200 327.750 42.000 333.600 ;
        RECT 53.100 331.950 58.800 333.600 ;
        RECT 53.700 327.750 55.500 330.600 ;
        RECT 57.000 327.750 58.800 331.950 ;
        RECT 61.200 327.750 63.000 333.600 ;
        RECT 73.650 327.750 75.450 333.600 ;
        RECT 79.650 330.600 80.550 334.800 ;
        RECT 92.550 332.700 100.350 334.050 ;
        RECT 76.650 327.750 78.450 330.600 ;
        RECT 79.650 327.750 81.450 330.600 ;
        RECT 82.650 327.750 84.450 330.600 ;
        RECT 92.550 327.750 94.350 332.700 ;
        RECT 95.550 327.750 97.350 331.800 ;
        RECT 98.550 327.750 100.350 332.700 ;
        RECT 101.550 333.600 102.750 335.700 ;
        RECT 101.550 327.750 103.350 333.600 ;
        RECT 116.550 332.700 124.350 334.050 ;
        RECT 116.550 327.750 118.350 332.700 ;
        RECT 119.550 327.750 121.350 331.800 ;
        RECT 122.550 327.750 124.350 332.700 ;
        RECT 125.550 333.600 126.750 335.700 ;
        RECT 125.550 327.750 127.350 333.600 ;
        RECT 142.950 330.600 144.000 337.050 ;
        RECT 160.950 336.750 162.150 340.050 ;
        RECT 163.950 338.850 166.050 340.950 ;
        RECT 166.950 340.050 169.050 342.150 ;
        RECT 175.950 340.050 178.050 342.150 ;
        RECT 164.100 337.050 165.900 338.850 ;
        RECT 158.250 335.700 162.000 336.750 ;
        RECT 180.000 336.300 181.050 344.700 ;
        RECT 183.150 342.150 184.350 347.400 ;
        RECT 181.950 340.050 184.350 342.150 ;
        RECT 158.250 333.600 159.450 335.700 ;
        RECT 180.000 335.400 182.250 336.300 ;
        RECT 177.150 334.500 182.250 335.400 ;
        RECT 139.650 327.750 141.450 330.600 ;
        RECT 142.650 327.750 144.450 330.600 ;
        RECT 145.650 327.750 147.450 330.600 ;
        RECT 157.650 327.750 159.450 333.600 ;
        RECT 160.650 332.700 168.450 334.050 ;
        RECT 160.650 327.750 162.450 332.700 ;
        RECT 163.650 327.750 165.450 331.800 ;
        RECT 166.650 327.750 168.450 332.700 ;
        RECT 177.150 330.600 178.350 334.500 ;
        RECT 183.150 333.600 184.350 340.050 ;
        RECT 199.650 342.150 200.850 347.400 ;
        RECT 206.250 346.500 207.450 353.400 ;
        RECT 215.550 352.200 217.350 358.200 ;
        RECT 218.550 352.200 220.350 359.250 ;
        RECT 201.750 345.600 207.450 346.500 ;
        RECT 216.450 347.100 217.350 352.200 ;
        RECT 223.050 348.900 224.850 358.200 ;
        RECT 223.050 348.000 225.150 348.900 ;
        RECT 216.450 346.200 222.600 347.100 ;
        RECT 201.750 344.700 204.000 345.600 ;
        RECT 199.650 340.050 202.050 342.150 ;
        RECT 199.650 333.600 200.850 340.050 ;
        RECT 202.950 336.300 204.000 344.700 ;
        RECT 206.100 342.150 207.900 343.950 ;
        RECT 218.250 342.150 220.050 343.950 ;
        RECT 205.950 340.050 208.050 342.150 ;
        RECT 214.950 338.850 217.050 340.950 ;
        RECT 217.950 340.050 220.050 342.150 ;
        RECT 221.250 343.500 222.600 346.200 ;
        RECT 221.250 341.700 223.050 343.500 ;
        RECT 215.250 337.050 217.050 338.850 ;
        RECT 201.750 335.400 204.000 336.300 ;
        RECT 221.250 336.000 222.600 341.700 ;
        RECT 224.250 340.950 225.150 348.000 ;
        RECT 227.550 347.400 229.350 359.250 ;
        RECT 242.550 353.400 244.350 359.250 ;
        RECT 242.550 346.500 243.750 353.400 ;
        RECT 245.850 347.400 247.650 359.250 ;
        RECT 248.850 347.400 250.650 359.250 ;
        RECT 260.550 353.400 262.350 359.250 ;
        RECT 263.550 353.400 265.350 359.250 ;
        RECT 266.550 353.400 268.350 359.250 ;
        RECT 242.550 345.600 248.250 346.500 ;
        RECT 246.000 344.700 248.250 345.600 ;
        RECT 227.100 342.150 228.900 343.950 ;
        RECT 242.100 342.150 243.900 343.950 ;
        RECT 223.950 338.850 226.050 340.950 ;
        RECT 226.950 340.050 229.050 342.150 ;
        RECT 241.950 340.050 244.050 342.150 ;
        RECT 201.750 334.500 206.850 335.400 ;
        RECT 176.550 327.750 178.350 330.600 ;
        RECT 179.850 327.750 181.650 333.600 ;
        RECT 182.850 327.750 184.650 333.600 ;
        RECT 199.350 327.750 201.150 333.600 ;
        RECT 202.350 327.750 204.150 333.600 ;
        RECT 205.650 330.600 206.850 334.500 ;
        RECT 216.300 335.100 222.600 336.000 ;
        RECT 216.300 331.800 217.350 335.100 ;
        RECT 224.250 334.200 225.150 338.850 ;
        RECT 246.000 336.300 247.050 344.700 ;
        RECT 249.150 342.150 250.350 347.400 ;
        RECT 263.550 345.150 264.750 353.400 ;
        RECT 280.350 347.400 282.150 359.250 ;
        RECT 283.350 347.400 285.150 359.250 ;
        RECT 286.650 353.400 288.450 359.250 ;
        RECT 247.950 340.050 250.350 342.150 ;
        RECT 259.950 341.850 262.050 343.950 ;
        RECT 262.950 343.050 265.050 345.150 ;
        RECT 260.100 340.050 261.900 341.850 ;
        RECT 246.000 335.400 248.250 336.300 ;
        RECT 223.050 333.300 225.150 334.200 ;
        RECT 205.650 327.750 207.450 330.600 ;
        RECT 215.550 328.800 217.350 331.800 ;
        RECT 218.550 327.750 220.350 331.800 ;
        RECT 223.050 328.800 224.850 333.300 ;
        RECT 227.550 327.750 229.350 334.800 ;
        RECT 243.150 334.500 248.250 335.400 ;
        RECT 243.150 330.600 244.350 334.500 ;
        RECT 249.150 333.600 250.350 340.050 ;
        RECT 263.550 335.700 264.750 343.050 ;
        RECT 265.950 341.850 268.050 343.950 ;
        RECT 280.650 342.150 281.850 347.400 ;
        RECT 287.250 346.500 288.450 353.400 ;
        RECT 303.150 347.400 304.950 359.250 ;
        RECT 307.650 347.400 310.950 359.250 ;
        RECT 313.650 347.400 315.450 359.250 ;
        RECT 327.150 347.400 328.950 359.250 ;
        RECT 331.650 347.400 334.950 359.250 ;
        RECT 337.650 347.400 339.450 359.250 ;
        RECT 349.650 353.400 351.450 359.250 ;
        RECT 352.650 353.400 354.450 359.250 ;
        RECT 355.650 353.400 357.450 359.250 ;
        RECT 365.550 353.400 367.350 359.250 ;
        RECT 282.750 345.600 288.450 346.500 ;
        RECT 282.750 344.700 285.000 345.600 ;
        RECT 266.100 340.050 267.900 341.850 ;
        RECT 280.650 340.050 283.050 342.150 ;
        RECT 263.550 334.800 267.150 335.700 ;
        RECT 242.550 327.750 244.350 330.600 ;
        RECT 245.850 327.750 247.650 333.600 ;
        RECT 248.850 327.750 250.650 333.600 ;
        RECT 260.850 327.750 262.650 333.600 ;
        RECT 265.350 327.750 267.150 334.800 ;
        RECT 280.650 333.600 281.850 340.050 ;
        RECT 283.950 336.300 285.000 344.700 ;
        RECT 287.100 342.150 288.900 343.950 ;
        RECT 302.250 342.150 304.050 343.950 ;
        RECT 308.250 342.150 309.450 347.400 ;
        RECT 314.100 342.150 315.900 343.950 ;
        RECT 326.250 342.150 328.050 343.950 ;
        RECT 332.250 342.150 333.450 347.400 ;
        RECT 353.250 345.150 354.450 353.400 ;
        RECT 365.550 346.500 366.750 353.400 ;
        RECT 368.850 347.400 370.650 359.250 ;
        RECT 371.850 347.400 373.650 359.250 ;
        RECT 383.550 353.400 385.350 359.250 ;
        RECT 365.550 345.600 371.250 346.500 ;
        RECT 338.100 342.150 339.900 343.950 ;
        RECT 286.950 340.050 289.050 342.150 ;
        RECT 301.950 340.050 304.050 342.150 ;
        RECT 304.950 338.850 307.050 340.950 ;
        RECT 307.950 340.050 310.050 342.150 ;
        RECT 305.700 337.050 307.500 338.850 ;
        RECT 282.750 335.400 285.000 336.300 ;
        RECT 308.400 336.150 309.600 340.050 ;
        RECT 310.950 338.850 313.050 340.950 ;
        RECT 313.950 340.050 316.050 342.150 ;
        RECT 325.950 340.050 328.050 342.150 ;
        RECT 328.950 338.850 331.050 340.950 ;
        RECT 331.950 340.050 334.050 342.150 ;
        RECT 311.100 337.050 312.900 338.850 ;
        RECT 329.700 337.050 331.500 338.850 ;
        RECT 332.400 336.150 333.600 340.050 ;
        RECT 334.950 338.850 337.050 340.950 ;
        RECT 337.950 340.050 340.050 342.150 ;
        RECT 349.950 341.850 352.050 343.950 ;
        RECT 352.950 343.050 355.050 345.150 ;
        RECT 369.000 344.700 371.250 345.600 ;
        RECT 350.100 340.050 351.900 341.850 ;
        RECT 335.100 337.050 336.900 338.850 ;
        RECT 282.750 334.500 287.850 335.400 ;
        RECT 280.350 327.750 282.150 333.600 ;
        RECT 283.350 327.750 285.150 333.600 ;
        RECT 286.650 330.600 287.850 334.500 ;
        RECT 305.250 335.100 309.600 336.150 ;
        RECT 329.250 335.100 333.600 336.150 ;
        RECT 353.250 335.700 354.450 343.050 ;
        RECT 355.950 341.850 358.050 343.950 ;
        RECT 365.100 342.150 366.900 343.950 ;
        RECT 356.100 340.050 357.900 341.850 ;
        RECT 364.950 340.050 367.050 342.150 ;
        RECT 305.250 333.600 306.150 335.100 ;
        RECT 286.650 327.750 288.450 330.600 ;
        RECT 301.650 328.500 303.450 333.600 ;
        RECT 304.650 329.400 306.450 333.600 ;
        RECT 307.650 333.000 315.450 333.900 ;
        RECT 329.250 333.600 330.150 335.100 ;
        RECT 350.850 334.800 354.450 335.700 ;
        RECT 369.000 336.300 370.050 344.700 ;
        RECT 372.150 342.150 373.350 347.400 ;
        RECT 383.550 346.500 384.750 353.400 ;
        RECT 386.850 347.400 388.650 359.250 ;
        RECT 389.850 347.400 391.650 359.250 ;
        RECT 401.550 348.300 403.350 359.250 ;
        RECT 404.550 349.200 406.350 359.250 ;
        RECT 407.550 348.300 409.350 359.250 ;
        RECT 401.550 347.400 409.350 348.300 ;
        RECT 410.550 347.400 412.350 359.250 ;
        RECT 427.650 347.400 429.450 359.250 ;
        RECT 432.150 348.900 433.950 358.200 ;
        RECT 436.650 352.200 438.450 359.250 ;
        RECT 439.650 352.200 441.450 358.200 ;
        RECT 431.850 348.000 433.950 348.900 ;
        RECT 383.550 345.600 389.250 346.500 ;
        RECT 387.000 344.700 389.250 345.600 ;
        RECT 383.100 342.150 384.900 343.950 ;
        RECT 370.950 340.050 373.350 342.150 ;
        RECT 382.950 340.050 385.050 342.150 ;
        RECT 369.000 335.400 371.250 336.300 ;
        RECT 307.650 328.500 309.450 333.000 ;
        RECT 301.650 327.750 309.450 328.500 ;
        RECT 310.650 327.750 312.450 332.100 ;
        RECT 313.650 327.750 315.450 333.000 ;
        RECT 325.650 328.500 327.450 333.600 ;
        RECT 328.650 329.400 330.450 333.600 ;
        RECT 331.650 333.000 339.450 333.900 ;
        RECT 331.650 328.500 333.450 333.000 ;
        RECT 325.650 327.750 333.450 328.500 ;
        RECT 334.650 327.750 336.450 332.100 ;
        RECT 337.650 327.750 339.450 333.000 ;
        RECT 350.850 327.750 352.650 334.800 ;
        RECT 366.150 334.500 371.250 335.400 ;
        RECT 355.350 327.750 357.150 333.600 ;
        RECT 366.150 330.600 367.350 334.500 ;
        RECT 372.150 333.600 373.350 340.050 ;
        RECT 387.000 336.300 388.050 344.700 ;
        RECT 390.150 342.150 391.350 347.400 ;
        RECT 410.700 342.150 411.900 347.400 ;
        RECT 428.100 342.150 429.900 343.950 ;
        RECT 388.950 340.050 391.350 342.150 ;
        RECT 387.000 335.400 389.250 336.300 ;
        RECT 384.150 334.500 389.250 335.400 ;
        RECT 365.550 327.750 367.350 330.600 ;
        RECT 368.850 327.750 370.650 333.600 ;
        RECT 371.850 327.750 373.650 333.600 ;
        RECT 384.150 330.600 385.350 334.500 ;
        RECT 390.150 333.600 391.350 340.050 ;
        RECT 400.950 338.850 403.050 340.950 ;
        RECT 404.100 339.150 405.900 340.950 ;
        RECT 401.100 337.050 402.900 338.850 ;
        RECT 403.950 337.050 406.050 339.150 ;
        RECT 406.950 338.850 409.050 340.950 ;
        RECT 409.950 340.050 412.050 342.150 ;
        RECT 427.950 340.050 430.050 342.150 ;
        RECT 431.850 340.950 432.750 348.000 ;
        RECT 439.650 347.100 440.550 352.200 ;
        RECT 451.650 347.400 453.450 359.250 ;
        RECT 456.150 348.900 457.950 358.200 ;
        RECT 460.650 352.200 462.450 359.250 ;
        RECT 463.650 352.200 465.450 358.200 ;
        RECT 473.550 353.400 475.350 359.250 ;
        RECT 455.850 348.000 457.950 348.900 ;
        RECT 434.400 346.200 440.550 347.100 ;
        RECT 434.400 343.500 435.750 346.200 ;
        RECT 433.950 341.700 435.750 343.500 ;
        RECT 407.100 337.050 408.900 338.850 ;
        RECT 410.700 333.600 411.900 340.050 ;
        RECT 430.950 338.850 433.050 340.950 ;
        RECT 383.550 327.750 385.350 330.600 ;
        RECT 386.850 327.750 388.650 333.600 ;
        RECT 389.850 327.750 391.650 333.600 ;
        RECT 402.000 327.750 403.800 333.600 ;
        RECT 406.200 331.950 411.900 333.600 ;
        RECT 406.200 327.750 408.000 331.950 ;
        RECT 409.500 327.750 411.300 330.600 ;
        RECT 427.650 327.750 429.450 334.800 ;
        RECT 431.850 334.200 432.750 338.850 ;
        RECT 434.400 336.000 435.750 341.700 ;
        RECT 436.950 342.150 438.750 343.950 ;
        RECT 452.100 342.150 453.900 343.950 ;
        RECT 436.950 340.050 439.050 342.150 ;
        RECT 439.950 338.850 442.050 340.950 ;
        RECT 451.950 340.050 454.050 342.150 ;
        RECT 455.850 340.950 456.750 348.000 ;
        RECT 463.650 347.100 464.550 352.200 ;
        RECT 458.400 346.200 464.550 347.100 ;
        RECT 473.550 346.500 474.750 353.400 ;
        RECT 476.850 347.400 478.650 359.250 ;
        RECT 479.850 347.400 481.650 359.250 ;
        RECT 491.550 353.400 493.350 359.250 ;
        RECT 494.550 353.400 496.350 359.250 ;
        RECT 497.550 354.000 499.350 359.250 ;
        RECT 494.700 353.100 496.350 353.400 ;
        RECT 500.550 353.400 502.350 359.250 ;
        RECT 500.550 353.100 501.750 353.400 ;
        RECT 494.700 352.200 501.750 353.100 ;
        RECT 494.100 348.150 495.900 349.950 ;
        RECT 458.400 343.500 459.750 346.200 ;
        RECT 473.550 345.600 479.250 346.500 ;
        RECT 477.000 344.700 479.250 345.600 ;
        RECT 457.950 341.700 459.750 343.500 ;
        RECT 454.950 338.850 457.050 340.950 ;
        RECT 439.950 337.050 441.750 338.850 ;
        RECT 434.400 335.100 440.700 336.000 ;
        RECT 431.850 333.300 433.950 334.200 ;
        RECT 432.150 328.800 433.950 333.300 ;
        RECT 439.650 331.800 440.700 335.100 ;
        RECT 436.650 327.750 438.450 331.800 ;
        RECT 439.650 328.800 441.450 331.800 ;
        RECT 451.650 327.750 453.450 334.800 ;
        RECT 455.850 334.200 456.750 338.850 ;
        RECT 458.400 336.000 459.750 341.700 ;
        RECT 460.950 342.150 462.750 343.950 ;
        RECT 473.100 342.150 474.900 343.950 ;
        RECT 460.950 340.050 463.050 342.150 ;
        RECT 463.950 338.850 466.050 340.950 ;
        RECT 472.950 340.050 475.050 342.150 ;
        RECT 463.950 337.050 465.750 338.850 ;
        RECT 477.000 336.300 478.050 344.700 ;
        RECT 480.150 342.150 481.350 347.400 ;
        RECT 491.100 345.150 492.900 346.950 ;
        RECT 493.950 346.050 496.050 348.150 ;
        RECT 497.250 345.150 499.050 346.950 ;
        RECT 490.950 343.050 493.050 345.150 ;
        RECT 496.950 343.050 499.050 345.150 ;
        RECT 500.700 343.950 501.750 352.200 ;
        RECT 517.650 347.400 519.450 359.250 ;
        RECT 522.150 348.900 523.950 358.200 ;
        RECT 526.650 352.200 528.450 359.250 ;
        RECT 529.650 352.200 531.450 358.200 ;
        RECT 539.550 353.400 541.350 359.250 ;
        RECT 521.850 348.000 523.950 348.900 ;
        RECT 478.950 340.050 481.350 342.150 ;
        RECT 499.950 341.850 502.050 343.950 ;
        RECT 518.100 342.150 519.900 343.950 ;
        RECT 458.400 335.100 464.700 336.000 ;
        RECT 477.000 335.400 479.250 336.300 ;
        RECT 455.850 333.300 457.950 334.200 ;
        RECT 456.150 328.800 457.950 333.300 ;
        RECT 463.650 331.800 464.700 335.100 ;
        RECT 474.150 334.500 479.250 335.400 ;
        RECT 460.650 327.750 462.450 331.800 ;
        RECT 463.650 328.800 465.450 331.800 ;
        RECT 474.150 330.600 475.350 334.500 ;
        RECT 480.150 333.600 481.350 340.050 ;
        RECT 500.400 337.650 501.600 341.850 ;
        RECT 517.950 340.050 520.050 342.150 ;
        RECT 521.850 340.950 522.750 348.000 ;
        RECT 529.650 347.100 530.550 352.200 ;
        RECT 524.400 346.200 530.550 347.100 ;
        RECT 539.550 346.500 540.750 353.400 ;
        RECT 542.850 347.400 544.650 359.250 ;
        RECT 545.850 347.400 547.650 359.250 ;
        RECT 557.550 353.400 559.350 359.250 ;
        RECT 560.550 353.400 562.350 359.250 ;
        RECT 563.550 353.400 565.350 359.250 ;
        RECT 524.400 343.500 525.750 346.200 ;
        RECT 539.550 345.600 545.250 346.500 ;
        RECT 543.000 344.700 545.250 345.600 ;
        RECT 523.950 341.700 525.750 343.500 ;
        RECT 520.950 338.850 523.050 340.950 ;
        RECT 473.550 327.750 475.350 330.600 ;
        RECT 476.850 327.750 478.650 333.600 ;
        RECT 479.850 327.750 481.650 333.600 ;
        RECT 491.700 327.750 493.500 336.600 ;
        RECT 497.100 336.000 501.600 337.650 ;
        RECT 497.100 327.750 498.900 336.000 ;
        RECT 517.650 327.750 519.450 334.800 ;
        RECT 521.850 334.200 522.750 338.850 ;
        RECT 524.400 336.000 525.750 341.700 ;
        RECT 526.950 342.150 528.750 343.950 ;
        RECT 539.100 342.150 540.900 343.950 ;
        RECT 526.950 340.050 529.050 342.150 ;
        RECT 529.950 338.850 532.050 340.950 ;
        RECT 538.950 340.050 541.050 342.150 ;
        RECT 529.950 337.050 531.750 338.850 ;
        RECT 543.000 336.300 544.050 344.700 ;
        RECT 546.150 342.150 547.350 347.400 ;
        RECT 560.550 345.150 561.750 353.400 ;
        RECT 579.300 347.400 581.100 359.250 ;
        RECT 583.500 347.400 585.300 359.250 ;
        RECT 586.800 353.400 588.600 359.250 ;
        RECT 602.550 347.400 604.350 359.250 ;
        RECT 606.750 347.400 608.550 359.250 ;
        RECT 625.650 353.400 627.450 359.250 ;
        RECT 628.650 353.400 630.450 359.250 ;
        RECT 631.650 353.400 633.450 359.250 ;
        RECT 544.950 340.050 547.350 342.150 ;
        RECT 556.950 341.850 559.050 343.950 ;
        RECT 559.950 343.050 562.050 345.150 ;
        RECT 557.100 340.050 558.900 341.850 ;
        RECT 524.400 335.100 530.700 336.000 ;
        RECT 543.000 335.400 545.250 336.300 ;
        RECT 521.850 333.300 523.950 334.200 ;
        RECT 522.150 328.800 523.950 333.300 ;
        RECT 529.650 331.800 530.700 335.100 ;
        RECT 540.150 334.500 545.250 335.400 ;
        RECT 526.650 327.750 528.450 331.800 ;
        RECT 529.650 328.800 531.450 331.800 ;
        RECT 540.150 330.600 541.350 334.500 ;
        RECT 546.150 333.600 547.350 340.050 ;
        RECT 560.550 335.700 561.750 343.050 ;
        RECT 562.950 341.850 565.050 343.950 ;
        RECT 578.100 342.150 579.900 343.950 ;
        RECT 583.950 342.150 585.150 347.400 ;
        RECT 586.950 345.150 588.750 346.950 ;
        RECT 606.000 346.350 608.550 347.400 ;
        RECT 586.950 343.050 589.050 345.150 ;
        RECT 602.100 342.150 603.900 343.950 ;
        RECT 563.100 340.050 564.900 341.850 ;
        RECT 577.950 340.050 580.050 342.150 ;
        RECT 580.950 338.850 583.050 340.950 ;
        RECT 583.950 340.050 586.050 342.150 ;
        RECT 601.950 340.050 604.050 342.150 ;
        RECT 581.100 337.050 582.900 338.850 ;
        RECT 584.850 336.750 586.050 340.050 ;
        RECT 606.000 339.150 607.050 346.350 ;
        RECT 629.250 345.150 630.450 353.400 ;
        RECT 645.450 347.400 647.250 359.250 ;
        RECT 649.650 347.400 651.450 359.250 ;
        RECT 660.300 347.400 662.100 359.250 ;
        RECT 664.500 347.400 666.300 359.250 ;
        RECT 667.800 353.400 669.600 359.250 ;
        RECT 682.650 353.400 684.450 359.250 ;
        RECT 685.650 353.400 687.450 359.250 ;
        RECT 695.550 353.400 697.350 359.250 ;
        RECT 645.450 346.350 648.000 347.400 ;
        RECT 608.100 342.150 609.900 343.950 ;
        RECT 607.950 340.050 610.050 342.150 ;
        RECT 625.950 341.850 628.050 343.950 ;
        RECT 628.950 343.050 631.050 345.150 ;
        RECT 626.100 340.050 627.900 341.850 ;
        RECT 604.950 337.050 607.050 339.150 ;
        RECT 585.000 335.700 588.750 336.750 ;
        RECT 560.550 334.800 564.150 335.700 ;
        RECT 539.550 327.750 541.350 330.600 ;
        RECT 542.850 327.750 544.650 333.600 ;
        RECT 545.850 327.750 547.650 333.600 ;
        RECT 557.850 327.750 559.650 333.600 ;
        RECT 562.350 327.750 564.150 334.800 ;
        RECT 578.550 332.700 586.350 334.050 ;
        RECT 578.550 327.750 580.350 332.700 ;
        RECT 581.550 327.750 583.350 331.800 ;
        RECT 584.550 327.750 586.350 332.700 ;
        RECT 587.550 333.600 588.750 335.700 ;
        RECT 587.550 327.750 589.350 333.600 ;
        RECT 606.000 330.600 607.050 337.050 ;
        RECT 629.250 335.700 630.450 343.050 ;
        RECT 631.950 341.850 634.050 343.950 ;
        RECT 644.100 342.150 645.900 343.950 ;
        RECT 632.100 340.050 633.900 341.850 ;
        RECT 643.950 340.050 646.050 342.150 ;
        RECT 626.850 334.800 630.450 335.700 ;
        RECT 646.950 339.150 648.000 346.350 ;
        RECT 650.100 342.150 651.900 343.950 ;
        RECT 659.100 342.150 660.900 343.950 ;
        RECT 664.950 342.150 666.150 347.400 ;
        RECT 667.950 345.150 669.750 346.950 ;
        RECT 667.950 343.050 670.050 345.150 ;
        RECT 649.950 340.050 652.050 342.150 ;
        RECT 658.950 340.050 661.050 342.150 ;
        RECT 646.950 337.050 649.050 339.150 ;
        RECT 661.950 338.850 664.050 340.950 ;
        RECT 664.950 340.050 667.050 342.150 ;
        RECT 683.400 340.950 684.600 353.400 ;
        RECT 695.550 346.500 696.750 353.400 ;
        RECT 698.850 347.400 700.650 359.250 ;
        RECT 701.850 347.400 703.650 359.250 ;
        RECT 713.550 347.400 715.350 359.250 ;
        RECT 717.750 347.400 719.550 359.250 ;
        RECT 736.650 353.400 738.450 359.250 ;
        RECT 739.650 354.000 741.450 359.250 ;
        RECT 695.550 345.600 701.250 346.500 ;
        RECT 699.000 344.700 701.250 345.600 ;
        RECT 695.100 342.150 696.900 343.950 ;
        RECT 662.100 337.050 663.900 338.850 ;
        RECT 602.550 327.750 604.350 330.600 ;
        RECT 605.550 327.750 607.350 330.600 ;
        RECT 608.550 327.750 610.350 330.600 ;
        RECT 626.850 327.750 628.650 334.800 ;
        RECT 631.350 327.750 633.150 333.600 ;
        RECT 646.950 330.600 648.000 337.050 ;
        RECT 665.850 336.750 667.050 340.050 ;
        RECT 682.950 338.850 685.050 340.950 ;
        RECT 686.100 339.150 687.900 340.950 ;
        RECT 694.950 340.050 697.050 342.150 ;
        RECT 666.000 335.700 669.750 336.750 ;
        RECT 659.550 332.700 667.350 334.050 ;
        RECT 643.650 327.750 645.450 330.600 ;
        RECT 646.650 327.750 648.450 330.600 ;
        RECT 649.650 327.750 651.450 330.600 ;
        RECT 659.550 327.750 661.350 332.700 ;
        RECT 662.550 327.750 664.350 331.800 ;
        RECT 665.550 327.750 667.350 332.700 ;
        RECT 668.550 333.600 669.750 335.700 ;
        RECT 668.550 327.750 670.350 333.600 ;
        RECT 683.400 330.600 684.600 338.850 ;
        RECT 685.950 337.050 688.050 339.150 ;
        RECT 699.000 336.300 700.050 344.700 ;
        RECT 702.150 342.150 703.350 347.400 ;
        RECT 717.000 346.350 719.550 347.400 ;
        RECT 737.250 353.100 738.450 353.400 ;
        RECT 742.650 353.400 744.450 359.250 ;
        RECT 745.650 353.400 747.450 359.250 ;
        RECT 757.650 353.400 759.450 359.250 ;
        RECT 760.650 353.400 762.450 359.250 ;
        RECT 763.650 353.400 765.450 359.250 ;
        RECT 776.400 353.400 778.200 359.250 ;
        RECT 742.650 353.100 744.300 353.400 ;
        RECT 737.250 352.200 744.300 353.100 ;
        RECT 713.100 342.150 714.900 343.950 ;
        RECT 700.950 340.050 703.350 342.150 ;
        RECT 712.950 340.050 715.050 342.150 ;
        RECT 699.000 335.400 701.250 336.300 ;
        RECT 696.150 334.500 701.250 335.400 ;
        RECT 696.150 330.600 697.350 334.500 ;
        RECT 702.150 333.600 703.350 340.050 ;
        RECT 717.000 339.150 718.050 346.350 ;
        RECT 737.250 343.950 738.300 352.200 ;
        RECT 743.100 348.150 744.900 349.950 ;
        RECT 739.950 345.150 741.750 346.950 ;
        RECT 742.950 346.050 745.050 348.150 ;
        RECT 746.100 345.150 747.900 346.950 ;
        RECT 761.250 345.150 762.450 353.400 ;
        RECT 779.700 347.400 781.500 359.250 ;
        RECT 783.900 347.400 785.700 359.250 ;
        RECT 789.150 347.400 790.950 359.250 ;
        RECT 792.150 353.400 793.950 359.250 ;
        RECT 797.250 353.400 799.050 359.250 ;
        RECT 802.050 353.400 803.850 359.250 ;
        RECT 797.550 352.500 798.750 353.400 ;
        RECT 805.050 352.500 806.850 359.250 ;
        RECT 808.950 353.400 810.750 359.250 ;
        RECT 813.150 353.400 814.950 359.250 ;
        RECT 817.650 356.400 819.450 359.250 ;
        RECT 793.950 350.400 798.750 352.500 ;
        RECT 801.150 350.700 808.050 352.500 ;
        RECT 813.150 351.300 817.050 353.400 ;
        RECT 797.550 349.500 798.750 350.400 ;
        RECT 810.450 349.800 812.250 350.400 ;
        RECT 797.550 348.300 805.050 349.500 ;
        RECT 803.250 347.700 805.050 348.300 ;
        RECT 805.950 348.900 812.250 349.800 ;
        RECT 776.250 345.150 778.050 346.950 ;
        RECT 719.100 342.150 720.900 343.950 ;
        RECT 718.950 340.050 721.050 342.150 ;
        RECT 736.950 341.850 739.050 343.950 ;
        RECT 739.950 343.050 742.050 345.150 ;
        RECT 745.950 343.050 748.050 345.150 ;
        RECT 757.950 341.850 760.050 343.950 ;
        RECT 760.950 343.050 763.050 345.150 ;
        RECT 715.950 337.050 718.050 339.150 ;
        RECT 682.650 327.750 684.450 330.600 ;
        RECT 685.650 327.750 687.450 330.600 ;
        RECT 695.550 327.750 697.350 330.600 ;
        RECT 698.850 327.750 700.650 333.600 ;
        RECT 701.850 327.750 703.650 333.600 ;
        RECT 717.000 330.600 718.050 337.050 ;
        RECT 737.400 337.650 738.600 341.850 ;
        RECT 758.100 340.050 759.900 341.850 ;
        RECT 737.400 336.000 741.900 337.650 ;
        RECT 713.550 327.750 715.350 330.600 ;
        RECT 716.550 327.750 718.350 330.600 ;
        RECT 719.550 327.750 721.350 330.600 ;
        RECT 740.100 327.750 741.900 336.000 ;
        RECT 745.500 327.750 747.300 336.600 ;
        RECT 761.250 335.700 762.450 343.050 ;
        RECT 763.950 341.850 766.050 343.950 ;
        RECT 775.950 343.050 778.050 345.150 ;
        RECT 779.850 342.150 781.050 347.400 ;
        RECT 789.150 346.800 800.250 347.400 ;
        RECT 805.950 346.800 806.850 348.900 ;
        RECT 810.450 348.600 812.250 348.900 ;
        RECT 813.150 348.600 815.850 350.400 ;
        RECT 813.150 347.700 814.050 348.600 ;
        RECT 789.150 346.200 806.850 346.800 ;
        RECT 785.100 342.150 786.900 343.950 ;
        RECT 764.100 340.050 765.900 341.850 ;
        RECT 778.950 340.050 781.050 342.150 ;
        RECT 778.950 336.750 780.150 340.050 ;
        RECT 781.950 338.850 784.050 340.950 ;
        RECT 784.950 340.050 787.050 342.150 ;
        RECT 782.100 337.050 783.900 338.850 ;
        RECT 758.850 334.800 762.450 335.700 ;
        RECT 776.250 335.700 780.000 336.750 ;
        RECT 758.850 327.750 760.650 334.800 ;
        RECT 776.250 333.600 777.450 335.700 ;
        RECT 763.350 327.750 765.150 333.600 ;
        RECT 775.650 327.750 777.450 333.600 ;
        RECT 778.650 332.700 786.450 334.050 ;
        RECT 778.650 327.750 780.450 332.700 ;
        RECT 781.650 327.750 783.450 331.800 ;
        RECT 784.650 327.750 786.450 332.700 ;
        RECT 789.150 333.600 790.050 346.200 ;
        RECT 798.450 345.900 806.850 346.200 ;
        RECT 808.050 346.800 814.050 347.700 ;
        RECT 814.950 346.800 817.050 347.700 ;
        RECT 820.650 347.400 822.450 359.250 ;
        RECT 832.650 358.500 840.450 359.250 ;
        RECT 832.650 347.400 834.450 358.500 ;
        RECT 835.650 347.400 837.450 357.600 ;
        RECT 838.650 348.600 840.450 358.500 ;
        RECT 841.650 349.500 843.450 359.250 ;
        RECT 844.650 348.600 846.450 359.250 ;
        RECT 838.650 347.700 846.450 348.600 ;
        RECT 855.300 347.400 857.100 359.250 ;
        RECT 859.500 347.400 861.300 359.250 ;
        RECT 862.800 353.400 864.600 359.250 ;
        RECT 875.550 353.400 877.350 359.250 ;
        RECT 798.450 345.600 800.250 345.900 ;
        RECT 808.050 342.150 808.950 346.800 ;
        RECT 814.950 345.600 819.150 346.800 ;
        RECT 818.250 343.800 820.050 345.600 ;
        RECT 799.950 341.100 802.050 342.150 ;
        RECT 791.100 339.150 792.900 340.950 ;
        RECT 794.100 340.050 802.050 341.100 ;
        RECT 805.950 340.050 808.950 342.150 ;
        RECT 794.100 339.300 795.900 340.050 ;
        RECT 792.000 338.400 792.900 339.150 ;
        RECT 797.100 338.400 798.900 339.000 ;
        RECT 792.000 337.200 798.900 338.400 ;
        RECT 797.850 336.000 798.900 337.200 ;
        RECT 808.050 336.000 808.950 340.050 ;
        RECT 817.950 339.750 820.050 340.050 ;
        RECT 816.150 337.950 820.050 339.750 ;
        RECT 821.250 337.950 822.450 347.400 ;
        RECT 835.800 346.500 837.600 347.400 ;
        RECT 835.800 345.600 839.850 346.500 ;
        RECT 833.100 342.150 834.900 343.950 ;
        RECT 838.950 342.150 839.850 345.600 ;
        RECT 844.950 342.150 846.750 343.950 ;
        RECT 854.100 342.150 855.900 343.950 ;
        RECT 859.950 342.150 861.150 347.400 ;
        RECT 862.950 345.150 864.750 346.950 ;
        RECT 875.550 346.500 876.750 353.400 ;
        RECT 878.850 347.400 880.650 359.250 ;
        RECT 881.850 347.400 883.650 359.250 ;
        RECT 875.550 345.600 881.250 346.500 ;
        RECT 862.950 343.050 865.050 345.150 ;
        RECT 879.000 344.700 881.250 345.600 ;
        RECT 875.100 342.150 876.900 343.950 ;
        RECT 832.950 340.050 835.050 342.150 ;
        RECT 835.950 338.850 838.050 340.950 ;
        RECT 838.950 340.050 841.050 342.150 ;
        RECT 797.850 335.100 808.950 336.000 ;
        RECT 817.950 335.850 822.450 337.950 ;
        RECT 836.250 337.050 838.050 338.850 ;
        RECT 797.850 334.200 798.900 335.100 ;
        RECT 808.050 334.800 808.950 335.100 ;
        RECT 789.150 327.750 790.950 333.600 ;
        RECT 793.950 331.500 796.050 333.600 ;
        RECT 797.550 332.400 799.350 334.200 ;
        RECT 800.850 333.450 802.650 334.200 ;
        RECT 800.850 332.400 805.800 333.450 ;
        RECT 808.050 333.000 809.850 334.800 ;
        RECT 821.250 333.600 822.450 335.850 ;
        RECT 840.000 333.600 841.050 340.050 ;
        RECT 841.950 338.850 844.050 340.950 ;
        RECT 844.950 340.050 847.050 342.150 ;
        RECT 853.950 340.050 856.050 342.150 ;
        RECT 856.950 338.850 859.050 340.950 ;
        RECT 859.950 340.050 862.050 342.150 ;
        RECT 874.950 340.050 877.050 342.150 ;
        RECT 841.950 337.050 843.750 338.850 ;
        RECT 857.100 337.050 858.900 338.850 ;
        RECT 860.850 336.750 862.050 340.050 ;
        RECT 861.000 335.700 864.750 336.750 ;
        RECT 814.950 332.700 817.050 333.600 ;
        RECT 795.000 330.600 796.050 331.500 ;
        RECT 804.750 330.600 805.800 332.400 ;
        RECT 813.300 331.500 817.050 332.700 ;
        RECT 813.300 330.600 814.350 331.500 ;
        RECT 792.150 327.750 793.950 330.600 ;
        RECT 795.000 329.700 798.750 330.600 ;
        RECT 796.950 327.750 798.750 329.700 ;
        RECT 801.450 327.750 803.250 330.600 ;
        RECT 804.750 327.750 806.550 330.600 ;
        RECT 808.650 327.750 810.450 330.600 ;
        RECT 812.850 327.750 814.650 330.600 ;
        RECT 817.350 327.750 819.150 330.600 ;
        RECT 820.650 327.750 822.450 333.600 ;
        RECT 835.800 327.750 837.600 333.600 ;
        RECT 840.000 327.750 841.800 333.600 ;
        RECT 844.200 327.750 846.000 333.600 ;
        RECT 854.550 332.700 862.350 334.050 ;
        RECT 854.550 327.750 856.350 332.700 ;
        RECT 857.550 327.750 859.350 331.800 ;
        RECT 860.550 327.750 862.350 332.700 ;
        RECT 863.550 333.600 864.750 335.700 ;
        RECT 879.000 336.300 880.050 344.700 ;
        RECT 882.150 342.150 883.350 347.400 ;
        RECT 880.950 340.050 883.350 342.150 ;
        RECT 879.000 335.400 881.250 336.300 ;
        RECT 876.150 334.500 881.250 335.400 ;
        RECT 863.550 327.750 865.350 333.600 ;
        RECT 876.150 330.600 877.350 334.500 ;
        RECT 882.150 333.600 883.350 340.050 ;
        RECT 875.550 327.750 877.350 330.600 ;
        RECT 878.850 327.750 880.650 333.600 ;
        RECT 881.850 327.750 883.650 333.600 ;
        RECT 14.850 316.200 16.650 323.250 ;
        RECT 19.350 317.400 21.150 323.250 ;
        RECT 32.850 316.200 34.650 323.250 ;
        RECT 37.350 317.400 39.150 323.250 ;
        RECT 47.550 320.400 49.350 323.250 ;
        RECT 50.550 320.400 52.350 323.250 ;
        RECT 53.550 320.400 55.350 323.250 ;
        RECT 65.550 320.400 67.350 323.250 ;
        RECT 68.550 320.400 70.350 323.250 ;
        RECT 85.650 320.400 87.450 323.250 ;
        RECT 88.650 320.400 90.450 323.250 ;
        RECT 91.650 320.400 93.450 323.250 ;
        RECT 40.950 318.450 43.050 319.050 ;
        RECT 46.950 318.450 49.050 319.050 ;
        RECT 40.950 317.550 49.050 318.450 ;
        RECT 40.950 316.950 43.050 317.550 ;
        RECT 46.950 316.950 49.050 317.550 ;
        RECT 14.850 315.300 18.450 316.200 ;
        RECT 32.850 315.300 36.450 316.200 ;
        RECT 14.100 309.150 15.900 310.950 ;
        RECT 13.950 307.050 16.050 309.150 ;
        RECT 17.250 307.950 18.450 315.300 ;
        RECT 20.100 309.150 21.900 310.950 ;
        RECT 32.100 309.150 33.900 310.950 ;
        RECT 16.950 305.850 19.050 307.950 ;
        RECT 19.950 307.050 22.050 309.150 ;
        RECT 31.950 307.050 34.050 309.150 ;
        RECT 35.250 307.950 36.450 315.300 ;
        RECT 51.000 313.950 52.050 320.400 ;
        RECT 49.950 311.850 52.050 313.950 ;
        RECT 64.950 311.850 67.050 313.950 ;
        RECT 68.400 312.150 69.600 320.400 ;
        RECT 88.950 313.950 90.000 320.400 ;
        RECT 105.000 317.400 106.800 323.250 ;
        RECT 109.200 319.050 111.000 323.250 ;
        RECT 112.500 320.400 114.300 323.250 ;
        RECT 109.200 317.400 114.900 319.050 ;
        RECT 38.100 309.150 39.900 310.950 ;
        RECT 34.950 305.850 37.050 307.950 ;
        RECT 37.950 307.050 40.050 309.150 ;
        RECT 46.950 308.850 49.050 310.950 ;
        RECT 47.100 307.050 48.900 308.850 ;
        RECT 17.250 297.600 18.450 305.850 ;
        RECT 19.950 303.450 22.050 304.050 ;
        RECT 31.950 303.450 34.050 304.050 ;
        RECT 19.950 302.550 34.050 303.450 ;
        RECT 19.950 301.950 22.050 302.550 ;
        RECT 31.950 301.950 34.050 302.550 ;
        RECT 35.250 297.600 36.450 305.850 ;
        RECT 51.000 304.650 52.050 311.850 ;
        RECT 52.950 308.850 55.050 310.950 ;
        RECT 65.100 310.050 66.900 311.850 ;
        RECT 67.950 310.050 70.050 312.150 ;
        RECT 88.950 311.850 91.050 313.950 ;
        RECT 104.100 312.150 105.900 313.950 ;
        RECT 53.100 307.050 54.900 308.850 ;
        RECT 51.000 303.600 53.550 304.650 ;
        RECT 13.650 291.750 15.450 297.600 ;
        RECT 16.650 291.750 18.450 297.600 ;
        RECT 19.650 291.750 21.450 297.600 ;
        RECT 31.650 291.750 33.450 297.600 ;
        RECT 34.650 291.750 36.450 297.600 ;
        RECT 37.650 291.750 39.450 297.600 ;
        RECT 47.550 291.750 49.350 303.600 ;
        RECT 51.750 291.750 53.550 303.600 ;
        RECT 68.400 297.600 69.600 310.050 ;
        RECT 85.950 308.850 88.050 310.950 ;
        RECT 86.100 307.050 87.900 308.850 ;
        RECT 88.950 304.650 90.000 311.850 ;
        RECT 91.950 308.850 94.050 310.950 ;
        RECT 103.950 310.050 106.050 312.150 ;
        RECT 106.950 311.850 109.050 313.950 ;
        RECT 110.100 312.150 111.900 313.950 ;
        RECT 107.100 310.050 108.900 311.850 ;
        RECT 109.950 310.050 112.050 312.150 ;
        RECT 113.700 310.950 114.900 317.400 ;
        RECT 128.850 316.200 130.650 323.250 ;
        RECT 133.350 317.400 135.150 323.250 ;
        RECT 143.550 318.300 145.350 323.250 ;
        RECT 146.550 319.200 148.350 323.250 ;
        RECT 149.550 318.300 151.350 323.250 ;
        RECT 143.550 316.950 151.350 318.300 ;
        RECT 152.550 317.400 154.350 323.250 ;
        RECT 169.650 317.400 171.450 323.250 ;
        RECT 128.850 315.300 132.450 316.200 ;
        RECT 152.550 315.300 153.750 317.400 ;
        RECT 112.950 308.850 115.050 310.950 ;
        RECT 128.100 309.150 129.900 310.950 ;
        RECT 92.100 307.050 93.900 308.850 ;
        RECT 87.450 303.600 90.000 304.650 ;
        RECT 113.700 303.600 114.900 308.850 ;
        RECT 127.950 307.050 130.050 309.150 ;
        RECT 131.250 307.950 132.450 315.300 ;
        RECT 150.000 314.250 153.750 315.300 ;
        RECT 170.250 315.300 171.450 317.400 ;
        RECT 172.650 318.300 174.450 323.250 ;
        RECT 175.650 319.200 177.450 323.250 ;
        RECT 178.650 318.300 180.450 323.250 ;
        RECT 172.650 316.950 180.450 318.300 ;
        RECT 190.350 317.400 192.150 323.250 ;
        RECT 193.350 317.400 195.150 323.250 ;
        RECT 196.650 320.400 198.450 323.250 ;
        RECT 170.250 314.250 174.000 315.300 ;
        RECT 146.100 312.150 147.900 313.950 ;
        RECT 134.100 309.150 135.900 310.950 ;
        RECT 130.950 305.850 133.050 307.950 ;
        RECT 133.950 307.050 136.050 309.150 ;
        RECT 142.950 308.850 145.050 310.950 ;
        RECT 145.950 310.050 148.050 312.150 ;
        RECT 149.850 310.950 151.050 314.250 ;
        RECT 148.950 308.850 151.050 310.950 ;
        RECT 172.950 310.950 174.150 314.250 ;
        RECT 176.100 312.150 177.900 313.950 ;
        RECT 172.950 308.850 175.050 310.950 ;
        RECT 175.950 310.050 178.050 312.150 ;
        RECT 190.650 310.950 191.850 317.400 ;
        RECT 196.650 316.500 197.850 320.400 ;
        RECT 209.850 317.400 211.650 323.250 ;
        RECT 192.750 315.600 197.850 316.500 ;
        RECT 214.350 316.200 216.150 323.250 ;
        RECT 192.750 314.700 195.000 315.600 ;
        RECT 178.950 308.850 181.050 310.950 ;
        RECT 190.650 308.850 193.050 310.950 ;
        RECT 143.100 307.050 144.900 308.850 ;
        RECT 65.550 291.750 67.350 297.600 ;
        RECT 68.550 291.750 70.350 297.600 ;
        RECT 87.450 291.750 89.250 303.600 ;
        RECT 91.650 291.750 93.450 303.600 ;
        RECT 104.550 302.700 112.350 303.600 ;
        RECT 104.550 291.750 106.350 302.700 ;
        RECT 107.550 291.750 109.350 301.800 ;
        RECT 110.550 291.750 112.350 302.700 ;
        RECT 113.550 291.750 115.350 303.600 ;
        RECT 131.250 297.600 132.450 305.850 ;
        RECT 148.950 303.600 150.150 308.850 ;
        RECT 151.950 305.850 154.050 307.950 ;
        RECT 169.950 305.850 172.050 307.950 ;
        RECT 151.950 304.050 153.750 305.850 ;
        RECT 170.250 304.050 172.050 305.850 ;
        RECT 173.850 303.600 175.050 308.850 ;
        RECT 179.100 307.050 180.900 308.850 ;
        RECT 190.650 303.600 191.850 308.850 ;
        RECT 193.950 306.300 195.000 314.700 ;
        RECT 212.550 315.300 216.150 316.200 ;
        RECT 230.850 316.200 232.650 323.250 ;
        RECT 235.350 317.400 237.150 323.250 ;
        RECT 245.550 319.200 247.350 322.200 ;
        RECT 248.550 319.200 250.350 323.250 ;
        RECT 230.850 315.300 234.450 316.200 ;
        RECT 196.950 308.850 199.050 310.950 ;
        RECT 209.100 309.150 210.900 310.950 ;
        RECT 197.100 307.050 198.900 308.850 ;
        RECT 208.950 307.050 211.050 309.150 ;
        RECT 212.550 307.950 213.750 315.300 ;
        RECT 215.100 309.150 216.900 310.950 ;
        RECT 230.100 309.150 231.900 310.950 ;
        RECT 192.750 305.400 195.000 306.300 ;
        RECT 211.950 305.850 214.050 307.950 ;
        RECT 214.950 307.050 217.050 309.150 ;
        RECT 229.950 307.050 232.050 309.150 ;
        RECT 233.250 307.950 234.450 315.300 ;
        RECT 246.300 315.900 247.350 319.200 ;
        RECT 253.050 317.700 254.850 322.200 ;
        RECT 253.050 316.800 255.150 317.700 ;
        RECT 246.300 315.000 252.600 315.900 ;
        RECT 245.250 312.150 247.050 313.950 ;
        RECT 236.100 309.150 237.900 310.950 ;
        RECT 244.950 310.050 247.050 312.150 ;
        RECT 232.950 305.850 235.050 307.950 ;
        RECT 235.950 307.050 238.050 309.150 ;
        RECT 247.950 308.850 250.050 310.950 ;
        RECT 248.250 307.050 250.050 308.850 ;
        RECT 251.250 309.300 252.600 315.000 ;
        RECT 254.250 312.150 255.150 316.800 ;
        RECT 257.550 316.200 259.350 323.250 ;
        RECT 272.550 318.300 274.350 323.250 ;
        RECT 275.550 319.200 277.350 323.250 ;
        RECT 278.550 318.300 280.350 323.250 ;
        RECT 272.550 316.950 280.350 318.300 ;
        RECT 281.550 317.400 283.350 323.250 ;
        RECT 293.550 319.200 295.350 322.200 ;
        RECT 296.550 319.200 298.350 323.250 ;
        RECT 281.550 315.300 282.750 317.400 ;
        RECT 279.000 314.250 282.750 315.300 ;
        RECT 294.300 315.900 295.350 319.200 ;
        RECT 301.050 317.700 302.850 322.200 ;
        RECT 301.050 316.800 303.150 317.700 ;
        RECT 294.300 315.000 300.600 315.900 ;
        RECT 275.100 312.150 276.900 313.950 ;
        RECT 253.950 310.050 256.050 312.150 ;
        RECT 251.250 307.500 253.050 309.300 ;
        RECT 192.750 304.500 198.450 305.400 ;
        RECT 127.650 291.750 129.450 297.600 ;
        RECT 130.650 291.750 132.450 297.600 ;
        RECT 133.650 291.750 135.450 297.600 ;
        RECT 144.300 291.750 146.100 303.600 ;
        RECT 148.500 291.750 150.300 303.600 ;
        RECT 151.800 291.750 153.600 297.600 ;
        RECT 170.400 291.750 172.200 297.600 ;
        RECT 173.700 291.750 175.500 303.600 ;
        RECT 177.900 291.750 179.700 303.600 ;
        RECT 190.350 291.750 192.150 303.600 ;
        RECT 193.350 291.750 195.150 303.600 ;
        RECT 197.250 297.600 198.450 304.500 ;
        RECT 212.550 297.600 213.750 305.850 ;
        RECT 233.250 297.600 234.450 305.850 ;
        RECT 251.250 304.800 252.600 307.500 ;
        RECT 246.450 303.900 252.600 304.800 ;
        RECT 246.450 298.800 247.350 303.900 ;
        RECT 254.250 303.000 255.150 310.050 ;
        RECT 256.950 308.850 259.050 310.950 ;
        RECT 271.950 308.850 274.050 310.950 ;
        RECT 274.950 310.050 277.050 312.150 ;
        RECT 278.850 310.950 280.050 314.250 ;
        RECT 293.250 312.150 295.050 313.950 ;
        RECT 277.950 308.850 280.050 310.950 ;
        RECT 292.950 310.050 295.050 312.150 ;
        RECT 295.950 308.850 298.050 310.950 ;
        RECT 257.100 307.050 258.900 308.850 ;
        RECT 272.100 307.050 273.900 308.850 ;
        RECT 277.950 303.600 279.150 308.850 ;
        RECT 280.950 305.850 283.050 307.950 ;
        RECT 296.250 307.050 298.050 308.850 ;
        RECT 299.250 309.300 300.600 315.000 ;
        RECT 302.250 312.150 303.150 316.800 ;
        RECT 305.550 316.200 307.350 323.250 ;
        RECT 320.550 320.400 322.350 323.250 ;
        RECT 321.150 316.500 322.350 320.400 ;
        RECT 323.850 317.400 325.650 323.250 ;
        RECT 326.850 317.400 328.650 323.250 ;
        RECT 339.000 317.400 340.800 323.250 ;
        RECT 343.200 319.050 345.000 323.250 ;
        RECT 346.500 320.400 348.300 323.250 ;
        RECT 362.550 320.400 364.350 323.250 ;
        RECT 365.550 320.400 367.350 323.250 ;
        RECT 343.200 317.400 348.900 319.050 ;
        RECT 321.150 315.600 326.250 316.500 ;
        RECT 324.000 314.700 326.250 315.600 ;
        RECT 301.950 310.050 304.050 312.150 ;
        RECT 299.250 307.500 301.050 309.300 ;
        RECT 280.950 304.050 282.750 305.850 ;
        RECT 299.250 304.800 300.600 307.500 ;
        RECT 294.450 303.900 300.600 304.800 ;
        RECT 253.050 302.100 255.150 303.000 ;
        RECT 196.650 291.750 198.450 297.600 ;
        RECT 209.550 291.750 211.350 297.600 ;
        RECT 212.550 291.750 214.350 297.600 ;
        RECT 215.550 291.750 217.350 297.600 ;
        RECT 229.650 291.750 231.450 297.600 ;
        RECT 232.650 291.750 234.450 297.600 ;
        RECT 235.650 291.750 237.450 297.600 ;
        RECT 245.550 292.800 247.350 298.800 ;
        RECT 248.550 291.750 250.350 298.800 ;
        RECT 253.050 292.800 254.850 302.100 ;
        RECT 257.550 291.750 259.350 303.600 ;
        RECT 273.300 291.750 275.100 303.600 ;
        RECT 277.500 291.750 279.300 303.600 ;
        RECT 294.450 298.800 295.350 303.900 ;
        RECT 302.250 303.000 303.150 310.050 ;
        RECT 304.950 308.850 307.050 310.950 ;
        RECT 319.950 308.850 322.050 310.950 ;
        RECT 305.100 307.050 306.900 308.850 ;
        RECT 320.100 307.050 321.900 308.850 ;
        RECT 324.000 306.300 325.050 314.700 ;
        RECT 327.150 310.950 328.350 317.400 ;
        RECT 338.100 312.150 339.900 313.950 ;
        RECT 325.950 308.850 328.350 310.950 ;
        RECT 337.950 310.050 340.050 312.150 ;
        RECT 340.950 311.850 343.050 313.950 ;
        RECT 344.100 312.150 345.900 313.950 ;
        RECT 341.100 310.050 342.900 311.850 ;
        RECT 343.950 310.050 346.050 312.150 ;
        RECT 347.700 310.950 348.900 317.400 ;
        RECT 361.950 311.850 364.050 313.950 ;
        RECT 365.400 312.150 366.600 320.400 ;
        RECT 380.850 316.200 382.650 323.250 ;
        RECT 385.350 317.400 387.150 323.250 ;
        RECT 395.850 317.400 397.650 323.250 ;
        RECT 400.350 316.200 402.150 323.250 ;
        RECT 413.850 317.400 415.650 323.250 ;
        RECT 418.350 316.200 420.150 323.250 ;
        RECT 431.550 320.400 433.350 323.250 ;
        RECT 434.550 320.400 436.350 323.250 ;
        RECT 446.550 320.400 448.350 323.250 ;
        RECT 380.850 315.300 384.450 316.200 ;
        RECT 346.950 308.850 349.050 310.950 ;
        RECT 362.100 310.050 363.900 311.850 ;
        RECT 364.950 310.050 367.050 312.150 ;
        RECT 324.000 305.400 326.250 306.300 ;
        RECT 320.550 304.500 326.250 305.400 ;
        RECT 301.050 302.100 303.150 303.000 ;
        RECT 280.800 291.750 282.600 297.600 ;
        RECT 293.550 292.800 295.350 298.800 ;
        RECT 296.550 291.750 298.350 298.800 ;
        RECT 301.050 292.800 302.850 302.100 ;
        RECT 305.550 291.750 307.350 303.600 ;
        RECT 320.550 297.600 321.750 304.500 ;
        RECT 327.150 303.600 328.350 308.850 ;
        RECT 347.700 303.600 348.900 308.850 ;
        RECT 320.550 291.750 322.350 297.600 ;
        RECT 323.850 291.750 325.650 303.600 ;
        RECT 326.850 291.750 328.650 303.600 ;
        RECT 338.550 302.700 346.350 303.600 ;
        RECT 338.550 291.750 340.350 302.700 ;
        RECT 341.550 291.750 343.350 301.800 ;
        RECT 344.550 291.750 346.350 302.700 ;
        RECT 347.550 291.750 349.350 303.600 ;
        RECT 365.400 297.600 366.600 310.050 ;
        RECT 380.100 309.150 381.900 310.950 ;
        RECT 379.950 307.050 382.050 309.150 ;
        RECT 383.250 307.950 384.450 315.300 ;
        RECT 398.550 315.300 402.150 316.200 ;
        RECT 416.550 315.300 420.150 316.200 ;
        RECT 386.100 309.150 387.900 310.950 ;
        RECT 395.100 309.150 396.900 310.950 ;
        RECT 382.950 305.850 385.050 307.950 ;
        RECT 385.950 307.050 388.050 309.150 ;
        RECT 394.950 307.050 397.050 309.150 ;
        RECT 398.550 307.950 399.750 315.300 ;
        RECT 401.100 309.150 402.900 310.950 ;
        RECT 413.100 309.150 414.900 310.950 ;
        RECT 397.950 305.850 400.050 307.950 ;
        RECT 400.950 307.050 403.050 309.150 ;
        RECT 412.950 307.050 415.050 309.150 ;
        RECT 416.550 307.950 417.750 315.300 ;
        RECT 430.950 311.850 433.050 313.950 ;
        RECT 434.400 312.150 435.600 320.400 ;
        RECT 447.150 316.500 448.350 320.400 ;
        RECT 449.850 317.400 451.650 323.250 ;
        RECT 452.850 317.400 454.650 323.250 ;
        RECT 447.150 315.600 452.250 316.500 ;
        RECT 450.000 314.700 452.250 315.600 ;
        RECT 419.100 309.150 420.900 310.950 ;
        RECT 431.100 310.050 432.900 311.850 ;
        RECT 433.950 310.050 436.050 312.150 ;
        RECT 415.950 305.850 418.050 307.950 ;
        RECT 418.950 307.050 421.050 309.150 ;
        RECT 383.250 297.600 384.450 305.850 ;
        RECT 398.550 297.600 399.750 305.850 ;
        RECT 416.550 297.600 417.750 305.850 ;
        RECT 434.400 297.600 435.600 310.050 ;
        RECT 445.950 308.850 448.050 310.950 ;
        RECT 446.100 307.050 447.900 308.850 ;
        RECT 450.000 306.300 451.050 314.700 ;
        RECT 453.150 310.950 454.350 317.400 ;
        RECT 470.850 316.200 472.650 323.250 ;
        RECT 475.350 317.400 477.150 323.250 ;
        RECT 491.850 316.200 493.650 323.250 ;
        RECT 496.350 317.400 498.150 323.250 ;
        RECT 509.550 320.400 511.350 323.250 ;
        RECT 510.150 316.500 511.350 320.400 ;
        RECT 512.850 317.400 514.650 323.250 ;
        RECT 515.850 317.400 517.650 323.250 ;
        RECT 530.550 319.200 532.350 322.200 ;
        RECT 533.550 319.200 535.350 323.250 ;
        RECT 470.850 315.300 474.450 316.200 ;
        RECT 491.850 315.300 495.450 316.200 ;
        RECT 510.150 315.600 515.250 316.500 ;
        RECT 451.950 308.850 454.350 310.950 ;
        RECT 470.100 309.150 471.900 310.950 ;
        RECT 450.000 305.400 452.250 306.300 ;
        RECT 446.550 304.500 452.250 305.400 ;
        RECT 446.550 297.600 447.750 304.500 ;
        RECT 453.150 303.600 454.350 308.850 ;
        RECT 469.950 307.050 472.050 309.150 ;
        RECT 473.250 307.950 474.450 315.300 ;
        RECT 476.100 309.150 477.900 310.950 ;
        RECT 491.100 309.150 492.900 310.950 ;
        RECT 472.950 305.850 475.050 307.950 ;
        RECT 475.950 307.050 478.050 309.150 ;
        RECT 490.950 307.050 493.050 309.150 ;
        RECT 494.250 307.950 495.450 315.300 ;
        RECT 513.000 314.700 515.250 315.600 ;
        RECT 497.100 309.150 498.900 310.950 ;
        RECT 493.950 305.850 496.050 307.950 ;
        RECT 496.950 307.050 499.050 309.150 ;
        RECT 508.950 308.850 511.050 310.950 ;
        RECT 509.100 307.050 510.900 308.850 ;
        RECT 513.000 306.300 514.050 314.700 ;
        RECT 516.150 310.950 517.350 317.400 ;
        RECT 531.300 315.900 532.350 319.200 ;
        RECT 538.050 317.700 539.850 322.200 ;
        RECT 538.050 316.800 540.150 317.700 ;
        RECT 531.300 315.000 537.600 315.900 ;
        RECT 530.250 312.150 532.050 313.950 ;
        RECT 514.950 308.850 517.350 310.950 ;
        RECT 529.950 310.050 532.050 312.150 ;
        RECT 532.950 308.850 535.050 310.950 ;
        RECT 362.550 291.750 364.350 297.600 ;
        RECT 365.550 291.750 367.350 297.600 ;
        RECT 379.650 291.750 381.450 297.600 ;
        RECT 382.650 291.750 384.450 297.600 ;
        RECT 385.650 291.750 387.450 297.600 ;
        RECT 395.550 291.750 397.350 297.600 ;
        RECT 398.550 291.750 400.350 297.600 ;
        RECT 401.550 291.750 403.350 297.600 ;
        RECT 413.550 291.750 415.350 297.600 ;
        RECT 416.550 291.750 418.350 297.600 ;
        RECT 419.550 291.750 421.350 297.600 ;
        RECT 431.550 291.750 433.350 297.600 ;
        RECT 434.550 291.750 436.350 297.600 ;
        RECT 446.550 291.750 448.350 297.600 ;
        RECT 449.850 291.750 451.650 303.600 ;
        RECT 452.850 291.750 454.650 303.600 ;
        RECT 473.250 297.600 474.450 305.850 ;
        RECT 494.250 297.600 495.450 305.850 ;
        RECT 513.000 305.400 515.250 306.300 ;
        RECT 509.550 304.500 515.250 305.400 ;
        RECT 509.550 297.600 510.750 304.500 ;
        RECT 516.150 303.600 517.350 308.850 ;
        RECT 533.250 307.050 535.050 308.850 ;
        RECT 536.250 309.300 537.600 315.000 ;
        RECT 539.250 312.150 540.150 316.800 ;
        RECT 542.550 316.200 544.350 323.250 ;
        RECT 557.550 319.200 559.350 322.200 ;
        RECT 560.550 319.200 562.350 323.250 ;
        RECT 558.300 315.900 559.350 319.200 ;
        RECT 565.050 317.700 566.850 322.200 ;
        RECT 565.050 316.800 567.150 317.700 ;
        RECT 558.300 315.000 564.600 315.900 ;
        RECT 557.250 312.150 559.050 313.950 ;
        RECT 538.950 310.050 541.050 312.150 ;
        RECT 536.250 307.500 538.050 309.300 ;
        RECT 536.250 304.800 537.600 307.500 ;
        RECT 531.450 303.900 537.600 304.800 ;
        RECT 469.650 291.750 471.450 297.600 ;
        RECT 472.650 291.750 474.450 297.600 ;
        RECT 475.650 291.750 477.450 297.600 ;
        RECT 490.650 291.750 492.450 297.600 ;
        RECT 493.650 291.750 495.450 297.600 ;
        RECT 496.650 291.750 498.450 297.600 ;
        RECT 509.550 291.750 511.350 297.600 ;
        RECT 512.850 291.750 514.650 303.600 ;
        RECT 515.850 291.750 517.650 303.600 ;
        RECT 531.450 298.800 532.350 303.900 ;
        RECT 539.250 303.000 540.150 310.050 ;
        RECT 541.950 308.850 544.050 310.950 ;
        RECT 556.950 310.050 559.050 312.150 ;
        RECT 559.950 308.850 562.050 310.950 ;
        RECT 542.100 307.050 543.900 308.850 ;
        RECT 560.250 307.050 562.050 308.850 ;
        RECT 563.250 309.300 564.600 315.000 ;
        RECT 566.250 312.150 567.150 316.800 ;
        RECT 569.550 316.200 571.350 323.250 ;
        RECT 583.650 317.400 585.450 323.250 ;
        RECT 584.250 315.300 585.450 317.400 ;
        RECT 586.650 318.300 588.450 323.250 ;
        RECT 589.650 319.200 591.450 323.250 ;
        RECT 592.650 318.300 594.450 323.250 ;
        RECT 586.650 316.950 594.450 318.300 ;
        RECT 605.850 316.200 607.650 323.250 ;
        RECT 610.350 317.400 612.150 323.250 ;
        RECT 620.550 318.300 622.350 323.250 ;
        RECT 623.550 319.200 625.350 323.250 ;
        RECT 626.550 318.300 628.350 323.250 ;
        RECT 620.550 316.950 628.350 318.300 ;
        RECT 629.550 317.400 631.350 323.250 ;
        RECT 642.000 317.400 643.800 323.250 ;
        RECT 646.200 319.050 648.000 323.250 ;
        RECT 649.500 320.400 651.300 323.250 ;
        RECT 646.200 317.400 651.900 319.050 ;
        RECT 605.850 315.300 609.450 316.200 ;
        RECT 629.550 315.300 630.750 317.400 ;
        RECT 584.250 314.250 588.000 315.300 ;
        RECT 565.950 310.050 568.050 312.150 ;
        RECT 586.950 310.950 588.150 314.250 ;
        RECT 590.100 312.150 591.900 313.950 ;
        RECT 563.250 307.500 565.050 309.300 ;
        RECT 563.250 304.800 564.600 307.500 ;
        RECT 558.450 303.900 564.600 304.800 ;
        RECT 538.050 302.100 540.150 303.000 ;
        RECT 530.550 292.800 532.350 298.800 ;
        RECT 533.550 291.750 535.350 298.800 ;
        RECT 538.050 292.800 539.850 302.100 ;
        RECT 542.550 291.750 544.350 303.600 ;
        RECT 558.450 298.800 559.350 303.900 ;
        RECT 566.250 303.000 567.150 310.050 ;
        RECT 568.950 308.850 571.050 310.950 ;
        RECT 586.950 308.850 589.050 310.950 ;
        RECT 589.950 310.050 592.050 312.150 ;
        RECT 592.950 308.850 595.050 310.950 ;
        RECT 605.100 309.150 606.900 310.950 ;
        RECT 569.100 307.050 570.900 308.850 ;
        RECT 583.950 305.850 586.050 307.950 ;
        RECT 584.250 304.050 586.050 305.850 ;
        RECT 587.850 303.600 589.050 308.850 ;
        RECT 593.100 307.050 594.900 308.850 ;
        RECT 604.950 307.050 607.050 309.150 ;
        RECT 608.250 307.950 609.450 315.300 ;
        RECT 627.000 314.250 630.750 315.300 ;
        RECT 623.100 312.150 624.900 313.950 ;
        RECT 611.100 309.150 612.900 310.950 ;
        RECT 607.950 305.850 610.050 307.950 ;
        RECT 610.950 307.050 613.050 309.150 ;
        RECT 619.950 308.850 622.050 310.950 ;
        RECT 622.950 310.050 625.050 312.150 ;
        RECT 626.850 310.950 628.050 314.250 ;
        RECT 641.100 312.150 642.900 313.950 ;
        RECT 625.950 308.850 628.050 310.950 ;
        RECT 640.950 310.050 643.050 312.150 ;
        RECT 643.950 311.850 646.050 313.950 ;
        RECT 647.100 312.150 648.900 313.950 ;
        RECT 644.100 310.050 645.900 311.850 ;
        RECT 646.950 310.050 649.050 312.150 ;
        RECT 650.700 310.950 651.900 317.400 ;
        RECT 662.700 314.400 664.500 323.250 ;
        RECT 668.100 315.000 669.900 323.250 ;
        RECT 684.000 317.400 685.800 323.250 ;
        RECT 688.200 319.050 690.000 323.250 ;
        RECT 691.500 320.400 693.300 323.250 ;
        RECT 707.550 320.400 709.350 323.250 ;
        RECT 710.550 320.400 712.350 323.250 ;
        RECT 688.200 317.400 693.900 319.050 ;
        RECT 668.100 313.350 672.600 315.000 ;
        RECT 649.950 308.850 652.050 310.950 ;
        RECT 671.400 309.150 672.600 313.350 ;
        RECT 683.100 312.150 684.900 313.950 ;
        RECT 682.950 310.050 685.050 312.150 ;
        RECT 685.950 311.850 688.050 313.950 ;
        RECT 689.100 312.150 690.900 313.950 ;
        RECT 686.100 310.050 687.900 311.850 ;
        RECT 688.950 310.050 691.050 312.150 ;
        RECT 692.700 310.950 693.900 317.400 ;
        RECT 706.950 311.850 709.050 313.950 ;
        RECT 710.400 312.150 711.600 320.400 ;
        RECT 722.550 315.900 724.350 323.250 ;
        RECT 727.050 317.400 728.850 323.250 ;
        RECT 730.050 318.900 731.850 323.250 ;
        RECT 743.550 320.400 745.350 323.250 ;
        RECT 746.550 320.400 748.350 323.250 ;
        RECT 749.550 320.400 751.350 323.250 ;
        RECT 730.050 317.400 733.350 318.900 ;
        RECT 728.250 315.900 730.050 316.500 ;
        RECT 722.550 314.700 730.050 315.900 ;
        RECT 620.100 307.050 621.900 308.850 ;
        RECT 565.050 302.100 567.150 303.000 ;
        RECT 557.550 292.800 559.350 298.800 ;
        RECT 560.550 291.750 562.350 298.800 ;
        RECT 565.050 292.800 566.850 302.100 ;
        RECT 569.550 291.750 571.350 303.600 ;
        RECT 584.400 291.750 586.200 297.600 ;
        RECT 587.700 291.750 589.500 303.600 ;
        RECT 591.900 291.750 593.700 303.600 ;
        RECT 608.250 297.600 609.450 305.850 ;
        RECT 625.950 303.600 627.150 308.850 ;
        RECT 628.950 305.850 631.050 307.950 ;
        RECT 628.950 304.050 630.750 305.850 ;
        RECT 650.700 303.600 651.900 308.850 ;
        RECT 661.950 305.850 664.050 307.950 ;
        RECT 667.950 305.850 670.050 307.950 ;
        RECT 670.950 307.050 673.050 309.150 ;
        RECT 691.950 308.850 694.050 310.950 ;
        RECT 707.100 310.050 708.900 311.850 ;
        RECT 709.950 310.050 712.050 312.150 ;
        RECT 662.100 304.050 663.900 305.850 ;
        RECT 604.650 291.750 606.450 297.600 ;
        RECT 607.650 291.750 609.450 297.600 ;
        RECT 610.650 291.750 612.450 297.600 ;
        RECT 621.300 291.750 623.100 303.600 ;
        RECT 625.500 291.750 627.300 303.600 ;
        RECT 641.550 302.700 649.350 303.600 ;
        RECT 628.800 291.750 630.600 297.600 ;
        RECT 641.550 291.750 643.350 302.700 ;
        RECT 644.550 291.750 646.350 301.800 ;
        RECT 647.550 291.750 649.350 302.700 ;
        RECT 650.550 291.750 652.350 303.600 ;
        RECT 664.950 302.850 667.050 304.950 ;
        RECT 668.250 304.050 670.050 305.850 ;
        RECT 665.100 301.050 666.900 302.850 ;
        RECT 671.700 298.800 672.750 307.050 ;
        RECT 692.700 303.600 693.900 308.850 ;
        RECT 665.700 297.900 672.750 298.800 ;
        RECT 665.700 297.600 667.350 297.900 ;
        RECT 662.550 291.750 664.350 297.600 ;
        RECT 665.550 291.750 667.350 297.600 ;
        RECT 671.550 297.600 672.750 297.900 ;
        RECT 683.550 302.700 691.350 303.600 ;
        RECT 668.550 291.750 670.350 297.000 ;
        RECT 671.550 291.750 673.350 297.600 ;
        RECT 683.550 291.750 685.350 302.700 ;
        RECT 686.550 291.750 688.350 301.800 ;
        RECT 689.550 291.750 691.350 302.700 ;
        RECT 692.550 291.750 694.350 303.600 ;
        RECT 710.400 297.600 711.600 310.050 ;
        RECT 721.950 308.850 724.050 310.950 ;
        RECT 722.100 307.050 723.900 308.850 ;
        RECT 725.700 297.600 726.900 314.700 ;
        RECT 732.150 310.950 733.350 317.400 ;
        RECT 747.450 316.200 748.350 320.400 ;
        RECT 752.550 317.400 754.350 323.250 ;
        RECT 766.650 320.400 768.450 323.250 ;
        RECT 769.650 320.400 771.450 323.250 ;
        RECT 772.650 320.400 774.450 323.250 ;
        RECT 785.700 320.400 787.500 323.250 ;
        RECT 747.450 315.300 750.750 316.200 ;
        RECT 748.950 314.400 750.750 315.300 ;
        RECT 742.950 311.850 745.050 313.950 ;
        RECT 728.100 309.150 729.900 310.950 ;
        RECT 727.950 307.050 730.050 309.150 ;
        RECT 730.950 308.850 733.350 310.950 ;
        RECT 743.100 310.050 744.900 311.850 ;
        RECT 745.950 308.850 748.050 310.950 ;
        RECT 732.150 303.600 733.350 308.850 ;
        RECT 746.100 307.050 747.900 308.850 ;
        RECT 749.700 306.150 750.600 314.400 ;
        RECT 753.000 312.150 754.050 317.400 ;
        RECT 751.950 310.050 754.050 312.150 ;
        RECT 769.950 313.950 771.000 320.400 ;
        RECT 789.000 319.050 790.800 323.250 ;
        RECT 785.100 317.400 790.800 319.050 ;
        RECT 793.200 317.400 795.000 323.250 ;
        RECT 806.550 320.400 808.350 323.250 ;
        RECT 809.550 320.400 811.350 323.250 ;
        RECT 824.550 320.400 826.350 323.250 ;
        RECT 827.550 320.400 829.350 323.250 ;
        RECT 839.550 320.400 841.350 323.250 ;
        RECT 769.950 311.850 772.050 313.950 ;
        RECT 748.950 306.000 750.750 306.150 ;
        RECT 743.550 304.800 750.750 306.000 ;
        RECT 743.550 303.600 744.750 304.800 ;
        RECT 748.950 304.350 750.750 304.800 ;
        RECT 707.550 291.750 709.350 297.600 ;
        RECT 710.550 291.750 712.350 297.600 ;
        RECT 722.550 291.750 724.350 297.600 ;
        RECT 725.550 291.750 727.350 297.600 ;
        RECT 729.150 291.750 730.950 303.600 ;
        RECT 732.150 291.750 733.950 303.600 ;
        RECT 743.550 291.750 745.350 303.600 ;
        RECT 752.100 303.450 753.450 310.050 ;
        RECT 766.950 308.850 769.050 310.950 ;
        RECT 767.100 307.050 768.900 308.850 ;
        RECT 769.950 304.650 771.000 311.850 ;
        RECT 785.100 310.950 786.300 317.400 ;
        RECT 788.100 312.150 789.900 313.950 ;
        RECT 772.950 308.850 775.050 310.950 ;
        RECT 784.950 308.850 787.050 310.950 ;
        RECT 787.950 310.050 790.050 312.150 ;
        RECT 790.950 311.850 793.050 313.950 ;
        RECT 794.100 312.150 795.900 313.950 ;
        RECT 791.100 310.050 792.900 311.850 ;
        RECT 793.950 310.050 796.050 312.150 ;
        RECT 805.950 311.850 808.050 313.950 ;
        RECT 809.400 312.150 810.600 320.400 ;
        RECT 814.950 318.450 817.050 319.050 ;
        RECT 823.950 318.450 826.050 319.050 ;
        RECT 814.950 317.550 826.050 318.450 ;
        RECT 814.950 316.950 817.050 317.550 ;
        RECT 823.950 316.950 826.050 317.550 ;
        RECT 806.100 310.050 807.900 311.850 ;
        RECT 808.950 310.050 811.050 312.150 ;
        RECT 823.950 311.850 826.050 313.950 ;
        RECT 827.400 312.150 828.600 320.400 ;
        RECT 840.150 316.500 841.350 320.400 ;
        RECT 842.850 317.400 844.650 323.250 ;
        RECT 845.850 317.400 847.650 323.250 ;
        RECT 859.650 317.400 861.450 323.250 ;
        RECT 840.150 315.600 845.250 316.500 ;
        RECT 843.000 314.700 845.250 315.600 ;
        RECT 824.100 310.050 825.900 311.850 ;
        RECT 826.950 310.050 829.050 312.150 ;
        RECT 773.100 307.050 774.900 308.850 ;
        RECT 748.050 291.750 749.850 303.450 ;
        RECT 751.050 302.100 753.450 303.450 ;
        RECT 768.450 303.600 771.000 304.650 ;
        RECT 785.100 303.600 786.300 308.850 ;
        RECT 751.050 291.750 752.850 302.100 ;
        RECT 768.450 291.750 770.250 303.600 ;
        RECT 772.650 291.750 774.450 303.600 ;
        RECT 784.650 291.750 786.450 303.600 ;
        RECT 787.650 302.700 795.450 303.600 ;
        RECT 787.650 291.750 789.450 302.700 ;
        RECT 790.650 291.750 792.450 301.800 ;
        RECT 793.650 291.750 795.450 302.700 ;
        RECT 809.400 297.600 810.600 310.050 ;
        RECT 827.400 297.600 828.600 310.050 ;
        RECT 838.950 308.850 841.050 310.950 ;
        RECT 839.100 307.050 840.900 308.850 ;
        RECT 843.000 306.300 844.050 314.700 ;
        RECT 846.150 310.950 847.350 317.400 ;
        RECT 860.250 315.300 861.450 317.400 ;
        RECT 862.650 318.300 864.450 323.250 ;
        RECT 865.650 319.200 867.450 323.250 ;
        RECT 868.650 318.300 870.450 323.250 ;
        RECT 878.550 320.400 880.350 323.250 ;
        RECT 862.650 316.950 870.450 318.300 ;
        RECT 879.150 316.500 880.350 320.400 ;
        RECT 881.850 317.400 883.650 323.250 ;
        RECT 884.850 317.400 886.650 323.250 ;
        RECT 879.150 315.600 884.250 316.500 ;
        RECT 860.250 314.250 864.000 315.300 ;
        RECT 882.000 314.700 884.250 315.600 ;
        RECT 859.950 312.450 862.050 313.050 ;
        RECT 844.950 308.850 847.350 310.950 ;
        RECT 843.000 305.400 845.250 306.300 ;
        RECT 839.550 304.500 845.250 305.400 ;
        RECT 839.550 297.600 840.750 304.500 ;
        RECT 846.150 303.600 847.350 308.850 ;
        RECT 857.550 311.550 862.050 312.450 ;
        RECT 806.550 291.750 808.350 297.600 ;
        RECT 809.550 291.750 811.350 297.600 ;
        RECT 824.550 291.750 826.350 297.600 ;
        RECT 827.550 291.750 829.350 297.600 ;
        RECT 839.550 291.750 841.350 297.600 ;
        RECT 842.850 291.750 844.650 303.600 ;
        RECT 845.850 291.750 847.650 303.600 ;
        RECT 857.550 300.450 858.450 311.550 ;
        RECT 859.950 310.950 862.050 311.550 ;
        RECT 862.950 310.950 864.150 314.250 ;
        RECT 866.100 312.150 867.900 313.950 ;
        RECT 862.950 308.850 865.050 310.950 ;
        RECT 865.950 310.050 868.050 312.150 ;
        RECT 868.950 308.850 871.050 310.950 ;
        RECT 877.950 308.850 880.050 310.950 ;
        RECT 859.950 305.850 862.050 307.950 ;
        RECT 860.250 304.050 862.050 305.850 ;
        RECT 863.850 303.600 865.050 308.850 ;
        RECT 869.100 307.050 870.900 308.850 ;
        RECT 878.100 307.050 879.900 308.850 ;
        RECT 882.000 306.300 883.050 314.700 ;
        RECT 885.150 310.950 886.350 317.400 ;
        RECT 883.950 308.850 886.350 310.950 ;
        RECT 882.000 305.400 884.250 306.300 ;
        RECT 878.550 304.500 884.250 305.400 ;
        RECT 859.950 300.450 862.050 301.050 ;
        RECT 857.550 299.550 862.050 300.450 ;
        RECT 859.950 298.950 862.050 299.550 ;
        RECT 860.400 291.750 862.200 297.600 ;
        RECT 863.700 291.750 865.500 303.600 ;
        RECT 867.900 291.750 869.700 303.600 ;
        RECT 878.550 297.600 879.750 304.500 ;
        RECT 885.150 303.600 886.350 308.850 ;
        RECT 878.550 291.750 880.350 297.600 ;
        RECT 881.850 291.750 883.650 303.600 ;
        RECT 884.850 291.750 886.650 303.600 ;
        RECT 3.150 275.400 4.950 287.250 ;
        RECT 6.150 281.400 7.950 287.250 ;
        RECT 11.250 281.400 13.050 287.250 ;
        RECT 16.050 281.400 17.850 287.250 ;
        RECT 11.550 280.500 12.750 281.400 ;
        RECT 19.050 280.500 20.850 287.250 ;
        RECT 22.950 281.400 24.750 287.250 ;
        RECT 27.150 281.400 28.950 287.250 ;
        RECT 31.650 284.400 33.450 287.250 ;
        RECT 7.950 278.400 12.750 280.500 ;
        RECT 15.150 278.700 22.050 280.500 ;
        RECT 27.150 279.300 31.050 281.400 ;
        RECT 11.550 277.500 12.750 278.400 ;
        RECT 24.450 277.800 26.250 278.400 ;
        RECT 11.550 276.300 19.050 277.500 ;
        RECT 17.250 275.700 19.050 276.300 ;
        RECT 19.950 276.900 26.250 277.800 ;
        RECT 3.150 274.800 14.250 275.400 ;
        RECT 19.950 274.800 20.850 276.900 ;
        RECT 24.450 276.600 26.250 276.900 ;
        RECT 27.150 276.600 29.850 278.400 ;
        RECT 27.150 275.700 28.050 276.600 ;
        RECT 3.150 274.200 20.850 274.800 ;
        RECT 3.150 261.600 4.050 274.200 ;
        RECT 12.450 273.900 20.850 274.200 ;
        RECT 22.050 274.800 28.050 275.700 ;
        RECT 28.950 274.800 31.050 275.700 ;
        RECT 34.650 275.400 36.450 287.250 ;
        RECT 47.550 281.400 49.350 287.250 ;
        RECT 50.550 281.400 52.350 287.250 ;
        RECT 67.650 281.400 69.450 287.250 ;
        RECT 70.650 281.400 72.450 287.250 ;
        RECT 73.650 281.400 75.450 287.250 ;
        RECT 86.400 281.400 88.200 287.250 ;
        RECT 12.450 273.600 14.250 273.900 ;
        RECT 22.050 270.150 22.950 274.800 ;
        RECT 28.950 273.600 33.150 274.800 ;
        RECT 32.250 271.800 34.050 273.600 ;
        RECT 13.950 269.100 16.050 270.150 ;
        RECT 5.100 267.150 6.900 268.950 ;
        RECT 8.100 268.050 16.050 269.100 ;
        RECT 19.950 268.050 22.950 270.150 ;
        RECT 8.100 267.300 9.900 268.050 ;
        RECT 6.000 266.400 6.900 267.150 ;
        RECT 11.100 266.400 12.900 267.000 ;
        RECT 6.000 265.200 12.900 266.400 ;
        RECT 11.850 264.000 12.900 265.200 ;
        RECT 22.050 264.000 22.950 268.050 ;
        RECT 31.950 267.750 34.050 268.050 ;
        RECT 30.150 265.950 34.050 267.750 ;
        RECT 35.250 265.950 36.450 275.400 ;
        RECT 50.400 268.950 51.600 281.400 ;
        RECT 71.250 273.150 72.450 281.400 ;
        RECT 89.700 275.400 91.500 287.250 ;
        RECT 93.900 275.400 95.700 287.250 ;
        RECT 111.450 275.400 113.250 287.250 ;
        RECT 115.650 275.400 117.450 287.250 ;
        RECT 128.550 276.300 130.350 287.250 ;
        RECT 131.550 277.200 133.350 287.250 ;
        RECT 134.550 276.300 136.350 287.250 ;
        RECT 128.550 275.400 136.350 276.300 ;
        RECT 137.550 275.400 139.350 287.250 ;
        RECT 149.550 276.300 151.350 287.250 ;
        RECT 152.550 277.200 154.350 287.250 ;
        RECT 155.550 276.300 157.350 287.250 ;
        RECT 149.550 275.400 157.350 276.300 ;
        RECT 158.550 275.400 160.350 287.250 ;
        RECT 175.650 275.400 177.450 287.250 ;
        RECT 180.150 276.900 181.950 286.200 ;
        RECT 184.650 280.200 186.450 287.250 ;
        RECT 187.650 280.200 189.450 286.200 ;
        RECT 179.850 276.000 181.950 276.900 ;
        RECT 86.250 273.150 88.050 274.950 ;
        RECT 67.950 269.850 70.050 271.950 ;
        RECT 70.950 271.050 73.050 273.150 ;
        RECT 47.100 267.150 48.900 268.950 ;
        RECT 11.850 263.100 22.950 264.000 ;
        RECT 31.950 263.850 36.450 265.950 ;
        RECT 46.950 265.050 49.050 267.150 ;
        RECT 49.950 266.850 52.050 268.950 ;
        RECT 68.100 268.050 69.900 269.850 ;
        RECT 11.850 262.200 12.900 263.100 ;
        RECT 22.050 262.800 22.950 263.100 ;
        RECT 3.150 255.750 4.950 261.600 ;
        RECT 7.950 259.500 10.050 261.600 ;
        RECT 11.550 260.400 13.350 262.200 ;
        RECT 14.850 261.450 16.650 262.200 ;
        RECT 14.850 260.400 19.800 261.450 ;
        RECT 22.050 261.000 23.850 262.800 ;
        RECT 35.250 261.600 36.450 263.850 ;
        RECT 28.950 260.700 31.050 261.600 ;
        RECT 9.000 258.600 10.050 259.500 ;
        RECT 18.750 258.600 19.800 260.400 ;
        RECT 27.300 259.500 31.050 260.700 ;
        RECT 27.300 258.600 28.350 259.500 ;
        RECT 6.150 255.750 7.950 258.600 ;
        RECT 9.000 257.700 12.750 258.600 ;
        RECT 10.950 255.750 12.750 257.700 ;
        RECT 15.450 255.750 17.250 258.600 ;
        RECT 18.750 255.750 20.550 258.600 ;
        RECT 22.650 255.750 24.450 258.600 ;
        RECT 26.850 255.750 28.650 258.600 ;
        RECT 31.350 255.750 33.150 258.600 ;
        RECT 34.650 255.750 36.450 261.600 ;
        RECT 50.400 258.600 51.600 266.850 ;
        RECT 71.250 263.700 72.450 271.050 ;
        RECT 73.950 269.850 76.050 271.950 ;
        RECT 85.950 271.050 88.050 273.150 ;
        RECT 89.850 270.150 91.050 275.400 ;
        RECT 111.450 274.350 114.000 275.400 ;
        RECT 95.100 270.150 96.900 271.950 ;
        RECT 110.100 270.150 111.900 271.950 ;
        RECT 74.100 268.050 75.900 269.850 ;
        RECT 88.950 268.050 91.050 270.150 ;
        RECT 88.950 264.750 90.150 268.050 ;
        RECT 91.950 266.850 94.050 268.950 ;
        RECT 94.950 268.050 97.050 270.150 ;
        RECT 109.950 268.050 112.050 270.150 ;
        RECT 112.950 267.150 114.000 274.350 ;
        RECT 116.100 270.150 117.900 271.950 ;
        RECT 137.700 270.150 138.900 275.400 ;
        RECT 158.700 270.150 159.900 275.400 ;
        RECT 176.100 270.150 177.900 271.950 ;
        RECT 115.950 268.050 118.050 270.150 ;
        RECT 92.100 265.050 93.900 266.850 ;
        RECT 112.950 265.050 115.050 267.150 ;
        RECT 127.950 266.850 130.050 268.950 ;
        RECT 131.100 267.150 132.900 268.950 ;
        RECT 128.100 265.050 129.900 266.850 ;
        RECT 130.950 265.050 133.050 267.150 ;
        RECT 133.950 266.850 136.050 268.950 ;
        RECT 136.950 268.050 139.050 270.150 ;
        RECT 134.100 265.050 135.900 266.850 ;
        RECT 68.850 262.800 72.450 263.700 ;
        RECT 86.250 263.700 90.000 264.750 ;
        RECT 47.550 255.750 49.350 258.600 ;
        RECT 50.550 255.750 52.350 258.600 ;
        RECT 68.850 255.750 70.650 262.800 ;
        RECT 86.250 261.600 87.450 263.700 ;
        RECT 73.350 255.750 75.150 261.600 ;
        RECT 85.650 255.750 87.450 261.600 ;
        RECT 88.650 260.700 96.450 262.050 ;
        RECT 88.650 255.750 90.450 260.700 ;
        RECT 91.650 255.750 93.450 259.800 ;
        RECT 94.650 255.750 96.450 260.700 ;
        RECT 112.950 258.600 114.000 265.050 ;
        RECT 137.700 261.600 138.900 268.050 ;
        RECT 148.950 266.850 151.050 268.950 ;
        RECT 152.100 267.150 153.900 268.950 ;
        RECT 149.100 265.050 150.900 266.850 ;
        RECT 151.950 265.050 154.050 267.150 ;
        RECT 154.950 266.850 157.050 268.950 ;
        RECT 157.950 268.050 160.050 270.150 ;
        RECT 175.950 268.050 178.050 270.150 ;
        RECT 179.850 268.950 180.750 276.000 ;
        RECT 187.650 275.100 188.550 280.200 ;
        RECT 202.350 275.400 204.150 287.250 ;
        RECT 205.350 275.400 207.150 287.250 ;
        RECT 208.650 281.400 210.450 287.250 ;
        RECT 182.400 274.200 188.550 275.100 ;
        RECT 182.400 271.500 183.750 274.200 ;
        RECT 181.950 269.700 183.750 271.500 ;
        RECT 155.100 265.050 156.900 266.850 ;
        RECT 158.700 261.600 159.900 268.050 ;
        RECT 178.950 266.850 181.050 268.950 ;
        RECT 109.650 255.750 111.450 258.600 ;
        RECT 112.650 255.750 114.450 258.600 ;
        RECT 115.650 255.750 117.450 258.600 ;
        RECT 129.000 255.750 130.800 261.600 ;
        RECT 133.200 259.950 138.900 261.600 ;
        RECT 133.200 255.750 135.000 259.950 ;
        RECT 136.500 255.750 138.300 258.600 ;
        RECT 150.000 255.750 151.800 261.600 ;
        RECT 154.200 259.950 159.900 261.600 ;
        RECT 154.200 255.750 156.000 259.950 ;
        RECT 157.500 255.750 159.300 258.600 ;
        RECT 175.650 255.750 177.450 262.800 ;
        RECT 179.850 262.200 180.750 266.850 ;
        RECT 182.400 264.000 183.750 269.700 ;
        RECT 184.950 270.150 186.750 271.950 ;
        RECT 202.650 270.150 203.850 275.400 ;
        RECT 209.250 274.500 210.450 281.400 ;
        RECT 220.350 275.400 222.150 287.250 ;
        RECT 223.350 275.400 225.150 287.250 ;
        RECT 226.650 281.400 228.450 287.250 ;
        RECT 239.400 281.400 241.200 287.250 ;
        RECT 204.750 273.600 210.450 274.500 ;
        RECT 204.750 272.700 207.000 273.600 ;
        RECT 184.950 268.050 187.050 270.150 ;
        RECT 187.950 266.850 190.050 268.950 ;
        RECT 202.650 268.050 205.050 270.150 ;
        RECT 187.950 265.050 189.750 266.850 ;
        RECT 182.400 263.100 188.700 264.000 ;
        RECT 179.850 261.300 181.950 262.200 ;
        RECT 180.150 256.800 181.950 261.300 ;
        RECT 187.650 259.800 188.700 263.100 ;
        RECT 202.650 261.600 203.850 268.050 ;
        RECT 205.950 264.300 207.000 272.700 ;
        RECT 209.100 270.150 210.900 271.950 ;
        RECT 220.650 270.150 221.850 275.400 ;
        RECT 227.250 274.500 228.450 281.400 ;
        RECT 242.700 275.400 244.500 287.250 ;
        RECT 246.900 275.400 248.700 287.250 ;
        RECT 259.350 275.400 261.150 287.250 ;
        RECT 262.350 275.400 264.150 287.250 ;
        RECT 265.650 281.400 267.450 287.250 ;
        RECT 222.750 273.600 228.450 274.500 ;
        RECT 222.750 272.700 225.000 273.600 ;
        RECT 239.250 273.150 241.050 274.950 ;
        RECT 208.950 268.050 211.050 270.150 ;
        RECT 220.650 268.050 223.050 270.150 ;
        RECT 204.750 263.400 207.000 264.300 ;
        RECT 204.750 262.500 209.850 263.400 ;
        RECT 184.650 255.750 186.450 259.800 ;
        RECT 187.650 256.800 189.450 259.800 ;
        RECT 202.350 255.750 204.150 261.600 ;
        RECT 205.350 255.750 207.150 261.600 ;
        RECT 208.650 258.600 209.850 262.500 ;
        RECT 220.650 261.600 221.850 268.050 ;
        RECT 223.950 264.300 225.000 272.700 ;
        RECT 227.100 270.150 228.900 271.950 ;
        RECT 238.950 271.050 241.050 273.150 ;
        RECT 242.850 270.150 244.050 275.400 ;
        RECT 248.100 270.150 249.900 271.950 ;
        RECT 259.650 270.150 260.850 275.400 ;
        RECT 266.250 274.500 267.450 281.400 ;
        RECT 275.550 275.400 277.350 287.250 ;
        RECT 278.550 275.400 280.350 287.250 ;
        RECT 281.550 275.400 283.350 287.250 ;
        RECT 293.550 281.400 295.350 287.250 ;
        RECT 296.550 281.400 298.350 287.250 ;
        RECT 299.550 281.400 301.350 287.250 ;
        RECT 261.750 273.600 267.450 274.500 ;
        RECT 261.750 272.700 264.000 273.600 ;
        RECT 226.950 268.050 229.050 270.150 ;
        RECT 241.950 268.050 244.050 270.150 ;
        RECT 232.950 267.450 235.050 268.050 ;
        RECT 238.950 267.450 241.050 268.050 ;
        RECT 232.950 266.550 241.050 267.450 ;
        RECT 232.950 265.950 235.050 266.550 ;
        RECT 238.950 265.950 241.050 266.550 ;
        RECT 241.950 264.750 243.150 268.050 ;
        RECT 244.950 266.850 247.050 268.950 ;
        RECT 247.950 268.050 250.050 270.150 ;
        RECT 259.650 268.050 262.050 270.150 ;
        RECT 245.100 265.050 246.900 266.850 ;
        RECT 222.750 263.400 225.000 264.300 ;
        RECT 239.250 263.700 243.000 264.750 ;
        RECT 222.750 262.500 227.850 263.400 ;
        RECT 208.650 255.750 210.450 258.600 ;
        RECT 220.350 255.750 222.150 261.600 ;
        RECT 223.350 255.750 225.150 261.600 ;
        RECT 226.650 258.600 227.850 262.500 ;
        RECT 239.250 261.600 240.450 263.700 ;
        RECT 226.650 255.750 228.450 258.600 ;
        RECT 238.650 255.750 240.450 261.600 ;
        RECT 241.650 260.700 249.450 262.050 ;
        RECT 259.650 261.600 260.850 268.050 ;
        RECT 262.950 264.300 264.000 272.700 ;
        RECT 266.100 270.150 267.900 271.950 ;
        RECT 265.950 268.050 268.050 270.150 ;
        RECT 278.850 268.950 280.200 275.400 ;
        RECT 296.550 273.150 297.750 281.400 ;
        RECT 313.650 275.400 315.450 287.250 ;
        RECT 316.650 276.300 318.450 287.250 ;
        RECT 319.650 277.200 321.450 287.250 ;
        RECT 322.650 276.300 324.450 287.250 ;
        RECT 332.550 280.200 334.350 286.200 ;
        RECT 335.550 280.200 337.350 287.250 ;
        RECT 316.650 275.400 324.450 276.300 ;
        RECT 292.950 269.850 295.050 271.950 ;
        RECT 295.950 271.050 298.050 273.150 ;
        RECT 274.950 266.850 277.050 268.950 ;
        RECT 278.850 266.850 283.050 268.950 ;
        RECT 293.100 268.050 294.900 269.850 ;
        RECT 275.100 265.050 276.900 266.850 ;
        RECT 261.750 263.400 264.000 264.300 ;
        RECT 261.750 262.500 266.850 263.400 ;
        RECT 241.650 255.750 243.450 260.700 ;
        RECT 244.650 255.750 246.450 259.800 ;
        RECT 247.650 255.750 249.450 260.700 ;
        RECT 259.350 255.750 261.150 261.600 ;
        RECT 262.350 255.750 264.150 261.600 ;
        RECT 265.650 258.600 266.850 262.500 ;
        RECT 278.850 261.600 280.200 266.850 ;
        RECT 296.550 263.700 297.750 271.050 ;
        RECT 298.950 269.850 301.050 271.950 ;
        RECT 314.100 270.150 315.300 275.400 ;
        RECT 333.450 275.100 334.350 280.200 ;
        RECT 340.050 276.900 341.850 286.200 ;
        RECT 340.050 276.000 342.150 276.900 ;
        RECT 333.450 274.200 339.600 275.100 ;
        RECT 335.250 270.150 337.050 271.950 ;
        RECT 299.100 268.050 300.900 269.850 ;
        RECT 313.950 268.050 316.050 270.150 ;
        RECT 296.550 262.800 300.150 263.700 ;
        RECT 265.650 255.750 267.450 258.600 ;
        RECT 275.550 255.750 277.350 261.600 ;
        RECT 278.550 255.750 280.350 261.600 ;
        RECT 281.550 255.750 283.350 261.600 ;
        RECT 293.850 255.750 295.650 261.600 ;
        RECT 298.350 255.750 300.150 262.800 ;
        RECT 314.100 261.600 315.300 268.050 ;
        RECT 316.950 266.850 319.050 268.950 ;
        RECT 320.100 267.150 321.900 268.950 ;
        RECT 317.100 265.050 318.900 266.850 ;
        RECT 319.950 265.050 322.050 267.150 ;
        RECT 322.950 266.850 325.050 268.950 ;
        RECT 331.950 266.850 334.050 268.950 ;
        RECT 334.950 268.050 337.050 270.150 ;
        RECT 338.250 271.500 339.600 274.200 ;
        RECT 338.250 269.700 340.050 271.500 ;
        RECT 323.100 265.050 324.900 266.850 ;
        RECT 332.250 265.050 334.050 266.850 ;
        RECT 338.250 264.000 339.600 269.700 ;
        RECT 341.250 268.950 342.150 276.000 ;
        RECT 344.550 275.400 346.350 287.250 ;
        RECT 361.350 275.400 363.150 287.250 ;
        RECT 364.350 275.400 366.150 287.250 ;
        RECT 367.650 281.400 369.450 287.250 ;
        RECT 344.100 270.150 345.900 271.950 ;
        RECT 361.650 270.150 362.850 275.400 ;
        RECT 368.250 274.500 369.450 281.400 ;
        RECT 382.650 275.400 384.450 287.250 ;
        RECT 387.150 276.900 388.950 286.200 ;
        RECT 391.650 280.200 393.450 287.250 ;
        RECT 394.650 280.200 396.450 286.200 ;
        RECT 404.550 281.400 406.350 287.250 ;
        RECT 407.550 281.400 409.350 287.250 ;
        RECT 410.550 281.400 412.350 287.250 ;
        RECT 425.550 281.400 427.350 287.250 ;
        RECT 386.850 276.000 388.950 276.900 ;
        RECT 363.750 273.600 369.450 274.500 ;
        RECT 363.750 272.700 366.000 273.600 ;
        RECT 340.950 266.850 343.050 268.950 ;
        RECT 343.950 268.050 346.050 270.150 ;
        RECT 361.650 268.050 364.050 270.150 ;
        RECT 333.300 263.100 339.600 264.000 ;
        RECT 314.100 259.950 319.800 261.600 ;
        RECT 314.700 255.750 316.500 258.600 ;
        RECT 318.000 255.750 319.800 259.950 ;
        RECT 322.200 255.750 324.000 261.600 ;
        RECT 333.300 259.800 334.350 263.100 ;
        RECT 341.250 262.200 342.150 266.850 ;
        RECT 340.050 261.300 342.150 262.200 ;
        RECT 332.550 256.800 334.350 259.800 ;
        RECT 335.550 255.750 337.350 259.800 ;
        RECT 340.050 256.800 341.850 261.300 ;
        RECT 344.550 255.750 346.350 262.800 ;
        RECT 361.650 261.600 362.850 268.050 ;
        RECT 364.950 264.300 366.000 272.700 ;
        RECT 368.100 270.150 369.900 271.950 ;
        RECT 383.100 270.150 384.900 271.950 ;
        RECT 367.950 268.050 370.050 270.150 ;
        RECT 382.950 268.050 385.050 270.150 ;
        RECT 386.850 268.950 387.750 276.000 ;
        RECT 394.650 275.100 395.550 280.200 ;
        RECT 389.400 274.200 395.550 275.100 ;
        RECT 389.400 271.500 390.750 274.200 ;
        RECT 407.550 273.150 408.750 281.400 ;
        RECT 425.550 274.500 426.750 281.400 ;
        RECT 428.850 275.400 430.650 287.250 ;
        RECT 431.850 275.400 433.650 287.250 ;
        RECT 448.650 275.400 450.450 287.250 ;
        RECT 425.550 273.600 431.250 274.500 ;
        RECT 388.950 269.700 390.750 271.500 ;
        RECT 385.950 266.850 388.050 268.950 ;
        RECT 363.750 263.400 366.000 264.300 ;
        RECT 363.750 262.500 368.850 263.400 ;
        RECT 361.350 255.750 363.150 261.600 ;
        RECT 364.350 255.750 366.150 261.600 ;
        RECT 367.650 258.600 368.850 262.500 ;
        RECT 367.650 255.750 369.450 258.600 ;
        RECT 382.650 255.750 384.450 262.800 ;
        RECT 386.850 262.200 387.750 266.850 ;
        RECT 389.400 264.000 390.750 269.700 ;
        RECT 391.950 270.150 393.750 271.950 ;
        RECT 391.950 268.050 394.050 270.150 ;
        RECT 403.950 269.850 406.050 271.950 ;
        RECT 406.950 271.050 409.050 273.150 ;
        RECT 429.000 272.700 431.250 273.600 ;
        RECT 394.950 266.850 397.050 268.950 ;
        RECT 404.100 268.050 405.900 269.850 ;
        RECT 394.950 265.050 396.750 266.850 ;
        RECT 389.400 263.100 395.700 264.000 ;
        RECT 386.850 261.300 388.950 262.200 ;
        RECT 387.150 256.800 388.950 261.300 ;
        RECT 394.650 259.800 395.700 263.100 ;
        RECT 407.550 263.700 408.750 271.050 ;
        RECT 409.950 269.850 412.050 271.950 ;
        RECT 425.100 270.150 426.900 271.950 ;
        RECT 410.100 268.050 411.900 269.850 ;
        RECT 424.950 268.050 427.050 270.150 ;
        RECT 429.000 264.300 430.050 272.700 ;
        RECT 432.150 270.150 433.350 275.400 ;
        RECT 451.650 274.500 453.450 287.250 ;
        RECT 454.650 275.400 456.450 287.250 ;
        RECT 457.650 274.500 459.450 287.250 ;
        RECT 460.650 275.400 462.450 287.250 ;
        RECT 463.650 274.500 465.450 287.250 ;
        RECT 466.650 275.400 468.450 287.250 ;
        RECT 469.650 274.500 471.450 287.250 ;
        RECT 472.650 275.400 474.450 287.250 ;
        RECT 482.550 281.400 484.350 287.250 ;
        RECT 485.550 281.400 487.350 287.250 ;
        RECT 500.400 281.400 502.200 287.250 ;
        RECT 430.950 268.050 433.350 270.150 ;
        RECT 450.750 273.300 453.450 274.500 ;
        RECT 455.700 273.300 459.450 274.500 ;
        RECT 461.700 273.300 465.450 274.500 ;
        RECT 467.550 273.300 471.450 274.500 ;
        RECT 450.750 268.950 451.800 273.300 ;
        RECT 407.550 262.800 411.150 263.700 ;
        RECT 429.000 263.400 431.250 264.300 ;
        RECT 391.650 255.750 393.450 259.800 ;
        RECT 394.650 256.800 396.450 259.800 ;
        RECT 404.850 255.750 406.650 261.600 ;
        RECT 409.350 255.750 411.150 262.800 ;
        RECT 426.150 262.500 431.250 263.400 ;
        RECT 426.150 258.600 427.350 262.500 ;
        RECT 432.150 261.600 433.350 268.050 ;
        RECT 448.950 266.850 451.800 268.950 ;
        RECT 450.750 263.700 451.800 266.850 ;
        RECT 455.700 266.400 456.900 273.300 ;
        RECT 461.700 266.400 462.900 273.300 ;
        RECT 467.550 266.400 468.750 273.300 ;
        RECT 485.400 268.950 486.600 281.400 ;
        RECT 503.700 275.400 505.500 287.250 ;
        RECT 507.900 275.400 509.700 287.250 ;
        RECT 521.400 281.400 523.200 287.250 ;
        RECT 524.700 275.400 526.500 287.250 ;
        RECT 528.900 275.400 530.700 287.250 ;
        RECT 542.400 281.400 544.200 287.250 ;
        RECT 545.700 275.400 547.500 287.250 ;
        RECT 549.900 275.400 551.700 287.250 ;
        RECT 563.550 281.400 565.350 287.250 ;
        RECT 566.550 281.400 568.350 287.250 ;
        RECT 569.550 281.400 571.350 287.250 ;
        RECT 500.250 273.150 502.050 274.950 ;
        RECT 499.950 271.050 502.050 273.150 ;
        RECT 503.850 270.150 505.050 275.400 ;
        RECT 521.250 273.150 523.050 274.950 ;
        RECT 509.100 270.150 510.900 271.950 ;
        RECT 520.950 271.050 523.050 273.150 ;
        RECT 524.850 270.150 526.050 275.400 ;
        RECT 542.250 273.150 544.050 274.950 ;
        RECT 530.100 270.150 531.900 271.950 ;
        RECT 541.950 271.050 544.050 273.150 ;
        RECT 545.850 270.150 547.050 275.400 ;
        RECT 566.550 273.150 567.750 281.400 ;
        RECT 575.550 275.400 577.350 287.250 ;
        RECT 578.550 284.400 580.350 287.250 ;
        RECT 583.050 281.400 584.850 287.250 ;
        RECT 587.250 281.400 589.050 287.250 ;
        RECT 580.950 279.300 584.850 281.400 ;
        RECT 591.150 280.500 592.950 287.250 ;
        RECT 594.150 281.400 595.950 287.250 ;
        RECT 598.950 281.400 600.750 287.250 ;
        RECT 604.050 281.400 605.850 287.250 ;
        RECT 599.250 280.500 600.450 281.400 ;
        RECT 589.950 278.700 596.850 280.500 ;
        RECT 599.250 278.400 604.050 280.500 ;
        RECT 582.150 276.600 584.850 278.400 ;
        RECT 585.750 277.800 587.550 278.400 ;
        RECT 585.750 276.900 592.050 277.800 ;
        RECT 599.250 277.500 600.450 278.400 ;
        RECT 585.750 276.600 587.550 276.900 ;
        RECT 583.950 275.700 584.850 276.600 ;
        RECT 551.100 270.150 552.900 271.950 ;
        RECT 469.950 266.850 472.050 268.950 ;
        RECT 482.100 267.150 483.900 268.950 ;
        RECT 452.700 264.600 456.900 266.400 ;
        RECT 458.700 264.600 462.900 266.400 ;
        RECT 464.700 264.600 468.750 266.400 ;
        RECT 470.100 265.050 471.900 266.850 ;
        RECT 481.950 265.050 484.050 267.150 ;
        RECT 484.950 266.850 487.050 268.950 ;
        RECT 502.950 268.050 505.050 270.150 ;
        RECT 455.700 263.700 456.900 264.600 ;
        RECT 461.700 263.700 462.900 264.600 ;
        RECT 467.550 263.700 468.750 264.600 ;
        RECT 450.750 262.650 453.600 263.700 ;
        RECT 450.900 262.500 453.600 262.650 ;
        RECT 455.700 262.500 459.600 263.700 ;
        RECT 461.700 262.500 465.450 263.700 ;
        RECT 467.550 262.500 471.600 263.700 ;
        RECT 451.800 261.600 453.600 262.500 ;
        RECT 457.800 261.600 459.600 262.500 ;
        RECT 425.550 255.750 427.350 258.600 ;
        RECT 428.850 255.750 430.650 261.600 ;
        RECT 431.850 255.750 433.650 261.600 ;
        RECT 448.650 255.750 450.450 261.600 ;
        RECT 451.650 255.750 453.450 261.600 ;
        RECT 454.650 255.750 456.450 261.600 ;
        RECT 457.650 255.750 459.450 261.600 ;
        RECT 460.650 255.750 462.450 261.600 ;
        RECT 463.650 255.750 465.450 262.500 ;
        RECT 469.800 261.600 471.600 262.500 ;
        RECT 466.650 255.750 468.450 261.600 ;
        RECT 469.650 255.750 471.450 261.600 ;
        RECT 472.650 255.750 474.450 261.600 ;
        RECT 485.400 258.600 486.600 266.850 ;
        RECT 502.950 264.750 504.150 268.050 ;
        RECT 505.950 266.850 508.050 268.950 ;
        RECT 508.950 268.050 511.050 270.150 ;
        RECT 523.950 268.050 526.050 270.150 ;
        RECT 506.100 265.050 507.900 266.850 ;
        RECT 523.950 264.750 525.150 268.050 ;
        RECT 526.950 266.850 529.050 268.950 ;
        RECT 529.950 268.050 532.050 270.150 ;
        RECT 544.950 268.050 547.050 270.150 ;
        RECT 527.100 265.050 528.900 266.850 ;
        RECT 544.950 264.750 546.150 268.050 ;
        RECT 547.950 266.850 550.050 268.950 ;
        RECT 550.950 268.050 553.050 270.150 ;
        RECT 562.950 269.850 565.050 271.950 ;
        RECT 565.950 271.050 568.050 273.150 ;
        RECT 563.100 268.050 564.900 269.850 ;
        RECT 548.100 265.050 549.900 266.850 ;
        RECT 500.250 263.700 504.000 264.750 ;
        RECT 521.250 263.700 525.000 264.750 ;
        RECT 542.250 263.700 546.000 264.750 ;
        RECT 566.550 263.700 567.750 271.050 ;
        RECT 568.950 269.850 571.050 271.950 ;
        RECT 569.100 268.050 570.900 269.850 ;
        RECT 575.550 265.950 576.750 275.400 ;
        RECT 580.950 274.800 583.050 275.700 ;
        RECT 583.950 274.800 589.950 275.700 ;
        RECT 578.850 273.600 583.050 274.800 ;
        RECT 577.950 271.800 579.750 273.600 ;
        RECT 589.050 270.150 589.950 274.800 ;
        RECT 591.150 274.800 592.050 276.900 ;
        RECT 592.950 276.300 600.450 277.500 ;
        RECT 592.950 275.700 594.750 276.300 ;
        RECT 607.050 275.400 608.850 287.250 ;
        RECT 617.550 281.400 619.350 287.250 ;
        RECT 620.550 281.400 622.350 287.250 ;
        RECT 635.400 281.400 637.200 287.250 ;
        RECT 597.750 274.800 608.850 275.400 ;
        RECT 591.150 274.200 608.850 274.800 ;
        RECT 591.150 273.900 599.550 274.200 ;
        RECT 597.750 273.600 599.550 273.900 ;
        RECT 589.050 268.050 592.050 270.150 ;
        RECT 595.950 269.100 598.050 270.150 ;
        RECT 595.950 268.050 603.900 269.100 ;
        RECT 577.950 267.750 580.050 268.050 ;
        RECT 577.950 265.950 581.850 267.750 ;
        RECT 575.550 263.850 580.050 265.950 ;
        RECT 589.050 264.000 589.950 268.050 ;
        RECT 602.100 267.300 603.900 268.050 ;
        RECT 605.100 267.150 606.900 268.950 ;
        RECT 599.100 266.400 600.900 267.000 ;
        RECT 605.100 266.400 606.000 267.150 ;
        RECT 599.100 265.200 606.000 266.400 ;
        RECT 599.100 264.000 600.150 265.200 ;
        RECT 500.250 261.600 501.450 263.700 ;
        RECT 482.550 255.750 484.350 258.600 ;
        RECT 485.550 255.750 487.350 258.600 ;
        RECT 499.650 255.750 501.450 261.600 ;
        RECT 502.650 260.700 510.450 262.050 ;
        RECT 521.250 261.600 522.450 263.700 ;
        RECT 502.650 255.750 504.450 260.700 ;
        RECT 505.650 255.750 507.450 259.800 ;
        RECT 508.650 255.750 510.450 260.700 ;
        RECT 520.650 255.750 522.450 261.600 ;
        RECT 523.650 260.700 531.450 262.050 ;
        RECT 542.250 261.600 543.450 263.700 ;
        RECT 566.550 262.800 570.150 263.700 ;
        RECT 523.650 255.750 525.450 260.700 ;
        RECT 526.650 255.750 528.450 259.800 ;
        RECT 529.650 255.750 531.450 260.700 ;
        RECT 541.650 255.750 543.450 261.600 ;
        RECT 544.650 260.700 552.450 262.050 ;
        RECT 544.650 255.750 546.450 260.700 ;
        RECT 547.650 255.750 549.450 259.800 ;
        RECT 550.650 255.750 552.450 260.700 ;
        RECT 563.850 255.750 565.650 261.600 ;
        RECT 568.350 255.750 570.150 262.800 ;
        RECT 575.550 261.600 576.750 263.850 ;
        RECT 589.050 263.100 600.150 264.000 ;
        RECT 589.050 262.800 589.950 263.100 ;
        RECT 575.550 255.750 577.350 261.600 ;
        RECT 580.950 260.700 583.050 261.600 ;
        RECT 588.150 261.000 589.950 262.800 ;
        RECT 599.100 262.200 600.150 263.100 ;
        RECT 595.350 261.450 597.150 262.200 ;
        RECT 580.950 259.500 584.700 260.700 ;
        RECT 583.650 258.600 584.700 259.500 ;
        RECT 592.200 260.400 597.150 261.450 ;
        RECT 598.650 260.400 600.450 262.200 ;
        RECT 607.950 261.600 608.850 274.200 ;
        RECT 620.400 268.950 621.600 281.400 ;
        RECT 638.700 275.400 640.500 287.250 ;
        RECT 642.900 275.400 644.700 287.250 ;
        RECT 655.650 281.400 657.450 287.250 ;
        RECT 658.650 281.400 660.450 287.250 ;
        RECT 635.250 273.150 637.050 274.950 ;
        RECT 634.950 271.050 637.050 273.150 ;
        RECT 638.850 270.150 640.050 275.400 ;
        RECT 644.100 270.150 645.900 271.950 ;
        RECT 617.100 267.150 618.900 268.950 ;
        RECT 616.950 265.050 619.050 267.150 ;
        RECT 619.950 266.850 622.050 268.950 ;
        RECT 637.950 268.050 640.050 270.150 ;
        RECT 592.200 258.600 593.250 260.400 ;
        RECT 601.950 259.500 604.050 261.600 ;
        RECT 601.950 258.600 603.000 259.500 ;
        RECT 578.850 255.750 580.650 258.600 ;
        RECT 583.350 255.750 585.150 258.600 ;
        RECT 587.550 255.750 589.350 258.600 ;
        RECT 591.450 255.750 593.250 258.600 ;
        RECT 594.750 255.750 596.550 258.600 ;
        RECT 599.250 257.700 603.000 258.600 ;
        RECT 599.250 255.750 601.050 257.700 ;
        RECT 604.050 255.750 605.850 258.600 ;
        RECT 607.050 255.750 608.850 261.600 ;
        RECT 620.400 258.600 621.600 266.850 ;
        RECT 637.950 264.750 639.150 268.050 ;
        RECT 640.950 266.850 643.050 268.950 ;
        RECT 643.950 268.050 646.050 270.150 ;
        RECT 656.400 268.950 657.600 281.400 ;
        RECT 669.300 275.400 671.100 287.250 ;
        RECT 673.500 275.400 675.300 287.250 ;
        RECT 676.800 281.400 678.600 287.250 ;
        RECT 684.150 275.400 685.950 287.250 ;
        RECT 687.150 281.400 688.950 287.250 ;
        RECT 692.250 281.400 694.050 287.250 ;
        RECT 697.050 281.400 698.850 287.250 ;
        RECT 692.550 280.500 693.750 281.400 ;
        RECT 700.050 280.500 701.850 287.250 ;
        RECT 703.950 281.400 705.750 287.250 ;
        RECT 708.150 281.400 709.950 287.250 ;
        RECT 712.650 284.400 714.450 287.250 ;
        RECT 688.950 278.400 693.750 280.500 ;
        RECT 696.150 278.700 703.050 280.500 ;
        RECT 708.150 279.300 712.050 281.400 ;
        RECT 692.550 277.500 693.750 278.400 ;
        RECT 705.450 277.800 707.250 278.400 ;
        RECT 692.550 276.300 700.050 277.500 ;
        RECT 698.250 275.700 700.050 276.300 ;
        RECT 700.950 276.900 707.250 277.800 ;
        RECT 668.100 270.150 669.900 271.950 ;
        RECT 673.950 270.150 675.150 275.400 ;
        RECT 676.950 273.150 678.750 274.950 ;
        RECT 684.150 274.800 695.250 275.400 ;
        RECT 700.950 274.800 701.850 276.900 ;
        RECT 705.450 276.600 707.250 276.900 ;
        RECT 708.150 276.600 710.850 278.400 ;
        RECT 708.150 275.700 709.050 276.600 ;
        RECT 684.150 274.200 701.850 274.800 ;
        RECT 676.950 271.050 679.050 273.150 ;
        RECT 655.950 266.850 658.050 268.950 ;
        RECT 659.100 267.150 660.900 268.950 ;
        RECT 667.950 268.050 670.050 270.150 ;
        RECT 641.100 265.050 642.900 266.850 ;
        RECT 635.250 263.700 639.000 264.750 ;
        RECT 635.250 261.600 636.450 263.700 ;
        RECT 617.550 255.750 619.350 258.600 ;
        RECT 620.550 255.750 622.350 258.600 ;
        RECT 634.650 255.750 636.450 261.600 ;
        RECT 637.650 260.700 645.450 262.050 ;
        RECT 637.650 255.750 639.450 260.700 ;
        RECT 640.650 255.750 642.450 259.800 ;
        RECT 643.650 255.750 645.450 260.700 ;
        RECT 656.400 258.600 657.600 266.850 ;
        RECT 658.950 265.050 661.050 267.150 ;
        RECT 670.950 266.850 673.050 268.950 ;
        RECT 673.950 268.050 676.050 270.150 ;
        RECT 671.100 265.050 672.900 266.850 ;
        RECT 674.850 264.750 676.050 268.050 ;
        RECT 675.000 263.700 678.750 264.750 ;
        RECT 668.550 260.700 676.350 262.050 ;
        RECT 655.650 255.750 657.450 258.600 ;
        RECT 658.650 255.750 660.450 258.600 ;
        RECT 668.550 255.750 670.350 260.700 ;
        RECT 671.550 255.750 673.350 259.800 ;
        RECT 674.550 255.750 676.350 260.700 ;
        RECT 677.550 261.600 678.750 263.700 ;
        RECT 684.150 261.600 685.050 274.200 ;
        RECT 693.450 273.900 701.850 274.200 ;
        RECT 703.050 274.800 709.050 275.700 ;
        RECT 709.950 274.800 712.050 275.700 ;
        RECT 715.650 275.400 717.450 287.250 ;
        RECT 729.300 275.400 731.100 287.250 ;
        RECT 733.500 275.400 735.300 287.250 ;
        RECT 736.800 281.400 738.600 287.250 ;
        RECT 749.550 276.300 751.350 287.250 ;
        RECT 752.550 277.200 754.350 287.250 ;
        RECT 755.550 276.300 757.350 287.250 ;
        RECT 749.550 275.400 757.350 276.300 ;
        RECT 758.550 275.400 760.350 287.250 ;
        RECT 773.550 275.400 775.350 287.250 ;
        RECT 776.550 275.400 778.350 287.250 ;
        RECT 792.300 275.400 794.100 287.250 ;
        RECT 796.500 275.400 798.300 287.250 ;
        RECT 799.800 281.400 801.600 287.250 ;
        RECT 807.150 275.400 808.950 287.250 ;
        RECT 810.150 281.400 811.950 287.250 ;
        RECT 815.250 281.400 817.050 287.250 ;
        RECT 820.050 281.400 821.850 287.250 ;
        RECT 815.550 280.500 816.750 281.400 ;
        RECT 823.050 280.500 824.850 287.250 ;
        RECT 826.950 281.400 828.750 287.250 ;
        RECT 831.150 281.400 832.950 287.250 ;
        RECT 835.650 284.400 837.450 287.250 ;
        RECT 811.950 278.400 816.750 280.500 ;
        RECT 819.150 278.700 826.050 280.500 ;
        RECT 831.150 279.300 835.050 281.400 ;
        RECT 815.550 277.500 816.750 278.400 ;
        RECT 828.450 277.800 830.250 278.400 ;
        RECT 815.550 276.300 823.050 277.500 ;
        RECT 821.250 275.700 823.050 276.300 ;
        RECT 823.950 276.900 830.250 277.800 ;
        RECT 693.450 273.600 695.250 273.900 ;
        RECT 703.050 270.150 703.950 274.800 ;
        RECT 709.950 273.600 714.150 274.800 ;
        RECT 713.250 271.800 715.050 273.600 ;
        RECT 694.950 269.100 697.050 270.150 ;
        RECT 686.100 267.150 687.900 268.950 ;
        RECT 689.100 268.050 697.050 269.100 ;
        RECT 700.950 268.050 703.950 270.150 ;
        RECT 689.100 267.300 690.900 268.050 ;
        RECT 687.000 266.400 687.900 267.150 ;
        RECT 692.100 266.400 693.900 267.000 ;
        RECT 687.000 265.200 693.900 266.400 ;
        RECT 692.850 264.000 693.900 265.200 ;
        RECT 703.050 264.000 703.950 268.050 ;
        RECT 712.950 267.750 715.050 268.050 ;
        RECT 711.150 265.950 715.050 267.750 ;
        RECT 716.250 265.950 717.450 275.400 ;
        RECT 728.100 270.150 729.900 271.950 ;
        RECT 733.950 270.150 735.150 275.400 ;
        RECT 736.950 273.150 738.750 274.950 ;
        RECT 736.950 271.050 739.050 273.150 ;
        RECT 758.700 270.150 759.900 275.400 ;
        RECT 776.400 270.150 777.600 275.400 ;
        RECT 791.100 270.150 792.900 271.950 ;
        RECT 796.950 270.150 798.150 275.400 ;
        RECT 799.950 273.150 801.750 274.950 ;
        RECT 807.150 274.800 818.250 275.400 ;
        RECT 823.950 274.800 824.850 276.900 ;
        RECT 828.450 276.600 830.250 276.900 ;
        RECT 831.150 276.600 833.850 278.400 ;
        RECT 831.150 275.700 832.050 276.600 ;
        RECT 807.150 274.200 824.850 274.800 ;
        RECT 799.950 271.050 802.050 273.150 ;
        RECT 727.950 268.050 730.050 270.150 ;
        RECT 730.950 266.850 733.050 268.950 ;
        RECT 733.950 268.050 736.050 270.150 ;
        RECT 692.850 263.100 703.950 264.000 ;
        RECT 712.950 263.850 717.450 265.950 ;
        RECT 731.100 265.050 732.900 266.850 ;
        RECT 734.850 264.750 736.050 268.050 ;
        RECT 748.950 266.850 751.050 268.950 ;
        RECT 752.100 267.150 753.900 268.950 ;
        RECT 749.100 265.050 750.900 266.850 ;
        RECT 751.950 265.050 754.050 267.150 ;
        RECT 754.950 266.850 757.050 268.950 ;
        RECT 757.950 268.050 760.050 270.150 ;
        RECT 755.100 265.050 756.900 266.850 ;
        RECT 692.850 262.200 693.900 263.100 ;
        RECT 703.050 262.800 703.950 263.100 ;
        RECT 677.550 255.750 679.350 261.600 ;
        RECT 684.150 255.750 685.950 261.600 ;
        RECT 688.950 259.500 691.050 261.600 ;
        RECT 692.550 260.400 694.350 262.200 ;
        RECT 695.850 261.450 697.650 262.200 ;
        RECT 695.850 260.400 700.800 261.450 ;
        RECT 703.050 261.000 704.850 262.800 ;
        RECT 716.250 261.600 717.450 263.850 ;
        RECT 735.000 263.700 738.750 264.750 ;
        RECT 709.950 260.700 712.050 261.600 ;
        RECT 690.000 258.600 691.050 259.500 ;
        RECT 699.750 258.600 700.800 260.400 ;
        RECT 708.300 259.500 712.050 260.700 ;
        RECT 708.300 258.600 709.350 259.500 ;
        RECT 687.150 255.750 688.950 258.600 ;
        RECT 690.000 257.700 693.750 258.600 ;
        RECT 691.950 255.750 693.750 257.700 ;
        RECT 696.450 255.750 698.250 258.600 ;
        RECT 699.750 255.750 701.550 258.600 ;
        RECT 703.650 255.750 705.450 258.600 ;
        RECT 707.850 255.750 709.650 258.600 ;
        RECT 712.350 255.750 714.150 258.600 ;
        RECT 715.650 255.750 717.450 261.600 ;
        RECT 728.550 260.700 736.350 262.050 ;
        RECT 728.550 255.750 730.350 260.700 ;
        RECT 731.550 255.750 733.350 259.800 ;
        RECT 734.550 255.750 736.350 260.700 ;
        RECT 737.550 261.600 738.750 263.700 ;
        RECT 758.700 261.600 759.900 268.050 ;
        RECT 772.950 266.850 775.050 268.950 ;
        RECT 775.950 268.050 778.050 270.150 ;
        RECT 790.950 268.050 793.050 270.150 ;
        RECT 773.100 265.050 774.900 266.850 ;
        RECT 776.400 261.600 777.600 268.050 ;
        RECT 793.950 266.850 796.050 268.950 ;
        RECT 796.950 268.050 799.050 270.150 ;
        RECT 794.100 265.050 795.900 266.850 ;
        RECT 797.850 264.750 799.050 268.050 ;
        RECT 798.000 263.700 801.750 264.750 ;
        RECT 737.550 255.750 739.350 261.600 ;
        RECT 750.000 255.750 751.800 261.600 ;
        RECT 754.200 259.950 759.900 261.600 ;
        RECT 754.200 255.750 756.000 259.950 ;
        RECT 757.500 255.750 759.300 258.600 ;
        RECT 773.550 255.750 775.350 261.600 ;
        RECT 776.550 255.750 778.350 261.600 ;
        RECT 791.550 260.700 799.350 262.050 ;
        RECT 791.550 255.750 793.350 260.700 ;
        RECT 794.550 255.750 796.350 259.800 ;
        RECT 797.550 255.750 799.350 260.700 ;
        RECT 800.550 261.600 801.750 263.700 ;
        RECT 807.150 261.600 808.050 274.200 ;
        RECT 816.450 273.900 824.850 274.200 ;
        RECT 826.050 274.800 832.050 275.700 ;
        RECT 832.950 274.800 835.050 275.700 ;
        RECT 838.650 275.400 840.450 287.250 ;
        RECT 853.650 275.400 855.450 287.250 ;
        RECT 816.450 273.600 818.250 273.900 ;
        RECT 826.050 270.150 826.950 274.800 ;
        RECT 832.950 273.600 837.150 274.800 ;
        RECT 836.250 271.800 838.050 273.600 ;
        RECT 817.950 269.100 820.050 270.150 ;
        RECT 809.100 267.150 810.900 268.950 ;
        RECT 812.100 268.050 820.050 269.100 ;
        RECT 823.950 268.050 826.950 270.150 ;
        RECT 812.100 267.300 813.900 268.050 ;
        RECT 810.000 266.400 810.900 267.150 ;
        RECT 815.100 266.400 816.900 267.000 ;
        RECT 810.000 265.200 816.900 266.400 ;
        RECT 815.850 264.000 816.900 265.200 ;
        RECT 826.050 264.000 826.950 268.050 ;
        RECT 835.950 267.750 838.050 268.050 ;
        RECT 834.150 265.950 838.050 267.750 ;
        RECT 839.250 265.950 840.450 275.400 ;
        RECT 856.650 274.500 858.450 287.250 ;
        RECT 859.650 275.400 861.450 287.250 ;
        RECT 862.650 274.500 864.450 287.250 ;
        RECT 865.650 275.400 867.450 287.250 ;
        RECT 868.650 274.500 870.450 287.250 ;
        RECT 871.650 275.400 873.450 287.250 ;
        RECT 874.650 274.500 876.450 287.250 ;
        RECT 877.650 275.400 879.450 287.250 ;
        RECT 855.750 273.300 858.450 274.500 ;
        RECT 860.700 273.300 864.450 274.500 ;
        RECT 866.700 273.300 870.450 274.500 ;
        RECT 872.550 273.300 876.450 274.500 ;
        RECT 855.750 268.950 856.800 273.300 ;
        RECT 853.950 266.850 856.800 268.950 ;
        RECT 815.850 263.100 826.950 264.000 ;
        RECT 835.950 263.850 840.450 265.950 ;
        RECT 815.850 262.200 816.900 263.100 ;
        RECT 826.050 262.800 826.950 263.100 ;
        RECT 800.550 255.750 802.350 261.600 ;
        RECT 807.150 255.750 808.950 261.600 ;
        RECT 811.950 259.500 814.050 261.600 ;
        RECT 815.550 260.400 817.350 262.200 ;
        RECT 818.850 261.450 820.650 262.200 ;
        RECT 818.850 260.400 823.800 261.450 ;
        RECT 826.050 261.000 827.850 262.800 ;
        RECT 839.250 261.600 840.450 263.850 ;
        RECT 855.750 263.700 856.800 266.850 ;
        RECT 860.700 266.400 861.900 273.300 ;
        RECT 866.700 266.400 867.900 273.300 ;
        RECT 872.550 266.400 873.750 273.300 ;
        RECT 874.950 266.850 877.050 268.950 ;
        RECT 857.700 264.600 861.900 266.400 ;
        RECT 863.700 264.600 867.900 266.400 ;
        RECT 869.700 264.600 873.750 266.400 ;
        RECT 875.100 265.050 876.900 266.850 ;
        RECT 860.700 263.700 861.900 264.600 ;
        RECT 866.700 263.700 867.900 264.600 ;
        RECT 872.550 263.700 873.750 264.600 ;
        RECT 855.750 262.650 858.600 263.700 ;
        RECT 855.900 262.500 858.600 262.650 ;
        RECT 860.700 262.500 864.600 263.700 ;
        RECT 866.700 262.500 870.450 263.700 ;
        RECT 872.550 262.500 876.600 263.700 ;
        RECT 856.800 261.600 858.600 262.500 ;
        RECT 862.800 261.600 864.600 262.500 ;
        RECT 832.950 260.700 835.050 261.600 ;
        RECT 813.000 258.600 814.050 259.500 ;
        RECT 822.750 258.600 823.800 260.400 ;
        RECT 831.300 259.500 835.050 260.700 ;
        RECT 831.300 258.600 832.350 259.500 ;
        RECT 810.150 255.750 811.950 258.600 ;
        RECT 813.000 257.700 816.750 258.600 ;
        RECT 814.950 255.750 816.750 257.700 ;
        RECT 819.450 255.750 821.250 258.600 ;
        RECT 822.750 255.750 824.550 258.600 ;
        RECT 826.650 255.750 828.450 258.600 ;
        RECT 830.850 255.750 832.650 258.600 ;
        RECT 835.350 255.750 837.150 258.600 ;
        RECT 838.650 255.750 840.450 261.600 ;
        RECT 853.650 255.750 855.450 261.600 ;
        RECT 856.650 255.750 858.450 261.600 ;
        RECT 859.650 255.750 861.450 261.600 ;
        RECT 862.650 255.750 864.450 261.600 ;
        RECT 865.650 255.750 867.450 261.600 ;
        RECT 868.650 255.750 870.450 262.500 ;
        RECT 874.800 261.600 876.600 262.500 ;
        RECT 871.650 255.750 873.450 261.600 ;
        RECT 874.650 255.750 876.450 261.600 ;
        RECT 877.650 255.750 879.450 261.600 ;
        RECT 10.650 245.400 12.450 251.250 ;
        RECT 11.250 243.300 12.450 245.400 ;
        RECT 13.650 246.300 15.450 251.250 ;
        RECT 16.650 247.200 18.450 251.250 ;
        RECT 19.650 246.300 21.450 251.250 ;
        RECT 13.650 244.950 21.450 246.300 ;
        RECT 32.850 244.200 34.650 251.250 ;
        RECT 37.350 245.400 39.150 251.250 ;
        RECT 53.850 244.200 55.650 251.250 ;
        RECT 58.350 245.400 60.150 251.250 ;
        RECT 70.650 245.400 72.450 251.250 ;
        RECT 32.850 243.300 36.450 244.200 ;
        RECT 53.850 243.300 57.450 244.200 ;
        RECT 11.250 242.250 15.000 243.300 ;
        RECT 13.950 238.950 15.150 242.250 ;
        RECT 17.100 240.150 18.900 241.950 ;
        RECT 13.950 236.850 16.050 238.950 ;
        RECT 16.950 238.050 19.050 240.150 ;
        RECT 19.950 236.850 22.050 238.950 ;
        RECT 32.100 237.150 33.900 238.950 ;
        RECT 10.950 233.850 13.050 235.950 ;
        RECT 11.250 232.050 13.050 233.850 ;
        RECT 14.850 231.600 16.050 236.850 ;
        RECT 20.100 235.050 21.900 236.850 ;
        RECT 31.950 235.050 34.050 237.150 ;
        RECT 35.250 235.950 36.450 243.300 ;
        RECT 38.100 237.150 39.900 238.950 ;
        RECT 53.100 237.150 54.900 238.950 ;
        RECT 34.950 233.850 37.050 235.950 ;
        RECT 37.950 235.050 40.050 237.150 ;
        RECT 52.950 235.050 55.050 237.150 ;
        RECT 56.250 235.950 57.450 243.300 ;
        RECT 71.250 243.300 72.450 245.400 ;
        RECT 73.650 246.300 75.450 251.250 ;
        RECT 76.650 247.200 78.450 251.250 ;
        RECT 79.650 246.300 81.450 251.250 ;
        RECT 91.650 248.400 93.450 251.250 ;
        RECT 94.650 248.400 96.450 251.250 ;
        RECT 97.650 248.400 99.450 251.250 ;
        RECT 73.650 244.950 81.450 246.300 ;
        RECT 71.250 242.250 75.000 243.300 ;
        RECT 73.950 238.950 75.150 242.250 ;
        RECT 94.950 241.950 96.000 248.400 ;
        RECT 113.850 244.200 115.650 251.250 ;
        RECT 118.350 245.400 120.150 251.250 ;
        RECT 130.650 245.400 132.450 251.250 ;
        RECT 113.850 243.300 117.450 244.200 ;
        RECT 77.100 240.150 78.900 241.950 ;
        RECT 59.100 237.150 60.900 238.950 ;
        RECT 55.950 233.850 58.050 235.950 ;
        RECT 58.950 235.050 61.050 237.150 ;
        RECT 73.950 236.850 76.050 238.950 ;
        RECT 76.950 238.050 79.050 240.150 ;
        RECT 94.950 239.850 97.050 241.950 ;
        RECT 79.950 236.850 82.050 238.950 ;
        RECT 91.950 236.850 94.050 238.950 ;
        RECT 70.950 233.850 73.050 235.950 ;
        RECT 11.400 219.750 13.200 225.600 ;
        RECT 14.700 219.750 16.500 231.600 ;
        RECT 18.900 219.750 20.700 231.600 ;
        RECT 35.250 225.600 36.450 233.850 ;
        RECT 56.250 225.600 57.450 233.850 ;
        RECT 71.250 232.050 73.050 233.850 ;
        RECT 74.850 231.600 76.050 236.850 ;
        RECT 80.100 235.050 81.900 236.850 ;
        RECT 92.100 235.050 93.900 236.850 ;
        RECT 94.950 232.650 96.000 239.850 ;
        RECT 97.950 236.850 100.050 238.950 ;
        RECT 113.100 237.150 114.900 238.950 ;
        RECT 98.100 235.050 99.900 236.850 ;
        RECT 112.950 235.050 115.050 237.150 ;
        RECT 116.250 235.950 117.450 243.300 ;
        RECT 131.250 243.300 132.450 245.400 ;
        RECT 133.650 246.300 135.450 251.250 ;
        RECT 136.650 247.200 138.450 251.250 ;
        RECT 139.650 246.300 141.450 251.250 ;
        RECT 133.650 244.950 141.450 246.300 ;
        RECT 152.850 244.200 154.650 251.250 ;
        RECT 157.350 245.400 159.150 251.250 ;
        RECT 167.550 248.400 169.350 251.250 ;
        RECT 170.550 248.400 172.350 251.250 ;
        RECT 185.700 248.400 187.500 251.250 ;
        RECT 152.850 243.300 156.450 244.200 ;
        RECT 131.250 242.250 135.000 243.300 ;
        RECT 133.950 238.950 135.150 242.250 ;
        RECT 137.100 240.150 138.900 241.950 ;
        RECT 119.100 237.150 120.900 238.950 ;
        RECT 115.950 233.850 118.050 235.950 ;
        RECT 118.950 235.050 121.050 237.150 ;
        RECT 133.950 236.850 136.050 238.950 ;
        RECT 136.950 238.050 139.050 240.150 ;
        RECT 139.950 236.850 142.050 238.950 ;
        RECT 152.100 237.150 153.900 238.950 ;
        RECT 130.950 233.850 133.050 235.950 ;
        RECT 93.450 231.600 96.000 232.650 ;
        RECT 31.650 219.750 33.450 225.600 ;
        RECT 34.650 219.750 36.450 225.600 ;
        RECT 37.650 219.750 39.450 225.600 ;
        RECT 52.650 219.750 54.450 225.600 ;
        RECT 55.650 219.750 57.450 225.600 ;
        RECT 58.650 219.750 60.450 225.600 ;
        RECT 71.400 219.750 73.200 225.600 ;
        RECT 74.700 219.750 76.500 231.600 ;
        RECT 78.900 219.750 80.700 231.600 ;
        RECT 93.450 219.750 95.250 231.600 ;
        RECT 97.650 219.750 99.450 231.600 ;
        RECT 116.250 225.600 117.450 233.850 ;
        RECT 131.250 232.050 133.050 233.850 ;
        RECT 134.850 231.600 136.050 236.850 ;
        RECT 140.100 235.050 141.900 236.850 ;
        RECT 151.950 235.050 154.050 237.150 ;
        RECT 155.250 235.950 156.450 243.300 ;
        RECT 157.950 243.450 160.050 244.050 ;
        RECT 163.950 243.450 166.050 244.050 ;
        RECT 157.950 242.550 166.050 243.450 ;
        RECT 157.950 241.950 160.050 242.550 ;
        RECT 163.950 241.950 166.050 242.550 ;
        RECT 166.950 239.850 169.050 241.950 ;
        RECT 170.400 240.150 171.600 248.400 ;
        RECT 189.000 247.050 190.800 251.250 ;
        RECT 185.100 245.400 190.800 247.050 ;
        RECT 193.200 245.400 195.000 251.250 ;
        RECT 158.100 237.150 159.900 238.950 ;
        RECT 167.100 238.050 168.900 239.850 ;
        RECT 169.950 238.050 172.050 240.150 ;
        RECT 185.100 238.950 186.300 245.400 ;
        RECT 206.850 244.200 208.650 251.250 ;
        RECT 211.350 245.400 213.150 251.250 ;
        RECT 226.650 245.400 228.450 251.250 ;
        RECT 206.850 243.300 210.450 244.200 ;
        RECT 188.100 240.150 189.900 241.950 ;
        RECT 154.950 233.850 157.050 235.950 ;
        RECT 157.950 235.050 160.050 237.150 ;
        RECT 112.650 219.750 114.450 225.600 ;
        RECT 115.650 219.750 117.450 225.600 ;
        RECT 118.650 219.750 120.450 225.600 ;
        RECT 131.400 219.750 133.200 225.600 ;
        RECT 134.700 219.750 136.500 231.600 ;
        RECT 138.900 219.750 140.700 231.600 ;
        RECT 155.250 225.600 156.450 233.850 ;
        RECT 170.400 225.600 171.600 238.050 ;
        RECT 184.950 236.850 187.050 238.950 ;
        RECT 187.950 238.050 190.050 240.150 ;
        RECT 190.950 239.850 193.050 241.950 ;
        RECT 194.100 240.150 195.900 241.950 ;
        RECT 191.100 238.050 192.900 239.850 ;
        RECT 193.950 238.050 196.050 240.150 ;
        RECT 206.100 237.150 207.900 238.950 ;
        RECT 185.100 231.600 186.300 236.850 ;
        RECT 205.950 235.050 208.050 237.150 ;
        RECT 209.250 235.950 210.450 243.300 ;
        RECT 227.250 243.300 228.450 245.400 ;
        RECT 229.650 246.300 231.450 251.250 ;
        RECT 232.650 247.200 234.450 251.250 ;
        RECT 235.650 246.300 237.450 251.250 ;
        RECT 229.650 244.950 237.450 246.300 ;
        RECT 245.550 246.300 247.350 251.250 ;
        RECT 248.550 247.200 250.350 251.250 ;
        RECT 251.550 246.300 253.350 251.250 ;
        RECT 245.550 244.950 253.350 246.300 ;
        RECT 254.550 245.400 256.350 251.250 ;
        RECT 268.650 248.400 270.450 251.250 ;
        RECT 271.650 248.400 273.450 251.250 ;
        RECT 254.550 243.300 255.750 245.400 ;
        RECT 227.250 242.250 231.000 243.300 ;
        RECT 252.000 242.250 255.750 243.300 ;
        RECT 229.950 238.950 231.150 242.250 ;
        RECT 233.100 240.150 234.900 241.950 ;
        RECT 248.100 240.150 249.900 241.950 ;
        RECT 212.100 237.150 213.900 238.950 ;
        RECT 208.950 233.850 211.050 235.950 ;
        RECT 211.950 235.050 214.050 237.150 ;
        RECT 229.950 236.850 232.050 238.950 ;
        RECT 232.950 238.050 235.050 240.150 ;
        RECT 235.950 236.850 238.050 238.950 ;
        RECT 244.950 236.850 247.050 238.950 ;
        RECT 247.950 238.050 250.050 240.150 ;
        RECT 251.850 238.950 253.050 242.250 ;
        RECT 269.400 240.150 270.600 248.400 ;
        RECT 285.000 245.400 286.800 251.250 ;
        RECT 289.200 247.050 291.000 251.250 ;
        RECT 292.500 248.400 294.300 251.250 ;
        RECT 289.200 245.400 294.900 247.050 ;
        RECT 250.950 236.850 253.050 238.950 ;
        RECT 268.950 238.050 271.050 240.150 ;
        RECT 271.950 239.850 274.050 241.950 ;
        RECT 284.100 240.150 285.900 241.950 ;
        RECT 272.100 238.050 273.900 239.850 ;
        RECT 283.950 238.050 286.050 240.150 ;
        RECT 286.950 239.850 289.050 241.950 ;
        RECT 290.100 240.150 291.900 241.950 ;
        RECT 287.100 238.050 288.900 239.850 ;
        RECT 289.950 238.050 292.050 240.150 ;
        RECT 293.700 238.950 294.900 245.400 ;
        RECT 311.100 243.000 312.900 251.250 ;
        RECT 308.400 241.350 312.900 243.000 ;
        RECT 316.500 242.400 318.300 251.250 ;
        RECT 328.650 245.400 330.450 251.250 ;
        RECT 329.250 243.300 330.450 245.400 ;
        RECT 331.650 246.300 333.450 251.250 ;
        RECT 334.650 247.200 336.450 251.250 ;
        RECT 337.650 246.300 339.450 251.250 ;
        RECT 349.650 248.400 351.450 251.250 ;
        RECT 352.650 248.400 354.450 251.250 ;
        RECT 364.650 248.400 366.450 251.250 ;
        RECT 367.650 248.400 369.450 251.250 ;
        RECT 370.650 248.400 372.450 251.250 ;
        RECT 331.650 244.950 339.450 246.300 ;
        RECT 329.250 242.250 333.000 243.300 ;
        RECT 226.950 233.850 229.050 235.950 ;
        RECT 151.650 219.750 153.450 225.600 ;
        RECT 154.650 219.750 156.450 225.600 ;
        RECT 157.650 219.750 159.450 225.600 ;
        RECT 167.550 219.750 169.350 225.600 ;
        RECT 170.550 219.750 172.350 225.600 ;
        RECT 184.650 219.750 186.450 231.600 ;
        RECT 187.650 230.700 195.450 231.600 ;
        RECT 187.650 219.750 189.450 230.700 ;
        RECT 190.650 219.750 192.450 229.800 ;
        RECT 193.650 219.750 195.450 230.700 ;
        RECT 209.250 225.600 210.450 233.850 ;
        RECT 227.250 232.050 229.050 233.850 ;
        RECT 230.850 231.600 232.050 236.850 ;
        RECT 236.100 235.050 237.900 236.850 ;
        RECT 245.100 235.050 246.900 236.850 ;
        RECT 250.950 231.600 252.150 236.850 ;
        RECT 253.950 233.850 256.050 235.950 ;
        RECT 253.950 232.050 255.750 233.850 ;
        RECT 205.650 219.750 207.450 225.600 ;
        RECT 208.650 219.750 210.450 225.600 ;
        RECT 211.650 219.750 213.450 225.600 ;
        RECT 227.400 219.750 229.200 225.600 ;
        RECT 230.700 219.750 232.500 231.600 ;
        RECT 234.900 219.750 236.700 231.600 ;
        RECT 246.300 219.750 248.100 231.600 ;
        RECT 250.500 219.750 252.300 231.600 ;
        RECT 269.400 225.600 270.600 238.050 ;
        RECT 292.950 236.850 295.050 238.950 ;
        RECT 308.400 237.150 309.600 241.350 ;
        RECT 331.950 238.950 333.150 242.250 ;
        RECT 335.100 240.150 336.900 241.950 ;
        RECT 350.400 240.150 351.600 248.400 ;
        RECT 367.950 241.950 369.000 248.400 ;
        RECT 383.700 242.400 385.500 251.250 ;
        RECT 389.100 243.000 390.900 251.250 ;
        RECT 407.850 245.400 409.650 251.250 ;
        RECT 412.350 244.200 414.150 251.250 ;
        RECT 410.550 243.300 414.150 244.200 ;
        RECT 293.700 231.600 294.900 236.850 ;
        RECT 307.950 235.050 310.050 237.150 ;
        RECT 331.950 236.850 334.050 238.950 ;
        RECT 334.950 238.050 337.050 240.150 ;
        RECT 337.950 236.850 340.050 238.950 ;
        RECT 349.950 238.050 352.050 240.150 ;
        RECT 352.950 239.850 355.050 241.950 ;
        RECT 367.950 239.850 370.050 241.950 ;
        RECT 389.100 241.350 393.600 243.000 ;
        RECT 353.100 238.050 354.900 239.850 ;
        RECT 284.550 230.700 292.350 231.600 ;
        RECT 253.800 219.750 255.600 225.600 ;
        RECT 268.650 219.750 270.450 225.600 ;
        RECT 271.650 219.750 273.450 225.600 ;
        RECT 284.550 219.750 286.350 230.700 ;
        RECT 287.550 219.750 289.350 229.800 ;
        RECT 290.550 219.750 292.350 230.700 ;
        RECT 293.550 219.750 295.350 231.600 ;
        RECT 308.250 226.800 309.300 235.050 ;
        RECT 310.950 233.850 313.050 235.950 ;
        RECT 316.950 233.850 319.050 235.950 ;
        RECT 328.950 233.850 331.050 235.950 ;
        RECT 310.950 232.050 312.750 233.850 ;
        RECT 313.950 230.850 316.050 232.950 ;
        RECT 317.100 232.050 318.900 233.850 ;
        RECT 329.250 232.050 331.050 233.850 ;
        RECT 332.850 231.600 334.050 236.850 ;
        RECT 338.100 235.050 339.900 236.850 ;
        RECT 314.100 229.050 315.900 230.850 ;
        RECT 308.250 225.900 315.300 226.800 ;
        RECT 308.250 225.600 309.450 225.900 ;
        RECT 307.650 219.750 309.450 225.600 ;
        RECT 313.650 225.600 315.300 225.900 ;
        RECT 310.650 219.750 312.450 225.000 ;
        RECT 313.650 219.750 315.450 225.600 ;
        RECT 316.650 219.750 318.450 225.600 ;
        RECT 329.400 219.750 331.200 225.600 ;
        RECT 332.700 219.750 334.500 231.600 ;
        RECT 336.900 219.750 338.700 231.600 ;
        RECT 350.400 225.600 351.600 238.050 ;
        RECT 364.950 236.850 367.050 238.950 ;
        RECT 365.100 235.050 366.900 236.850 ;
        RECT 367.950 232.650 369.000 239.850 ;
        RECT 370.950 236.850 373.050 238.950 ;
        RECT 392.400 237.150 393.600 241.350 ;
        RECT 407.100 237.150 408.900 238.950 ;
        RECT 371.100 235.050 372.900 236.850 ;
        RECT 382.950 233.850 385.050 235.950 ;
        RECT 388.950 233.850 391.050 235.950 ;
        RECT 391.950 235.050 394.050 237.150 ;
        RECT 406.950 235.050 409.050 237.150 ;
        RECT 410.550 235.950 411.750 243.300 ;
        RECT 434.100 243.000 435.900 251.250 ;
        RECT 431.400 241.350 435.900 243.000 ;
        RECT 439.500 242.400 441.300 251.250 ;
        RECT 455.850 244.200 457.650 251.250 ;
        RECT 460.350 245.400 462.150 251.250 ;
        RECT 455.850 243.300 459.450 244.200 ;
        RECT 413.100 237.150 414.900 238.950 ;
        RECT 431.400 237.150 432.600 241.350 ;
        RECT 455.100 237.150 456.900 238.950 ;
        RECT 366.450 231.600 369.000 232.650 ;
        RECT 383.100 232.050 384.900 233.850 ;
        RECT 349.650 219.750 351.450 225.600 ;
        RECT 352.650 219.750 354.450 225.600 ;
        RECT 366.450 219.750 368.250 231.600 ;
        RECT 370.650 219.750 372.450 231.600 ;
        RECT 385.950 230.850 388.050 232.950 ;
        RECT 389.250 232.050 391.050 233.850 ;
        RECT 386.100 229.050 387.900 230.850 ;
        RECT 392.700 226.800 393.750 235.050 ;
        RECT 409.950 233.850 412.050 235.950 ;
        RECT 412.950 235.050 415.050 237.150 ;
        RECT 430.950 235.050 433.050 237.150 ;
        RECT 386.700 225.900 393.750 226.800 ;
        RECT 386.700 225.600 388.350 225.900 ;
        RECT 383.550 219.750 385.350 225.600 ;
        RECT 386.550 219.750 388.350 225.600 ;
        RECT 392.550 225.600 393.750 225.900 ;
        RECT 410.550 225.600 411.750 233.850 ;
        RECT 431.250 226.800 432.300 235.050 ;
        RECT 433.950 233.850 436.050 235.950 ;
        RECT 439.950 233.850 442.050 235.950 ;
        RECT 454.950 235.050 457.050 237.150 ;
        RECT 458.250 235.950 459.450 243.300 ;
        RECT 473.700 242.400 475.500 251.250 ;
        RECT 479.100 243.000 480.900 251.250 ;
        RECT 494.550 248.400 496.350 251.250 ;
        RECT 495.150 244.500 496.350 248.400 ;
        RECT 497.850 245.400 499.650 251.250 ;
        RECT 500.850 245.400 502.650 251.250 ;
        RECT 495.150 243.600 500.250 244.500 ;
        RECT 479.100 241.350 483.600 243.000 ;
        RECT 461.100 237.150 462.900 238.950 ;
        RECT 482.400 237.150 483.600 241.350 ;
        RECT 498.000 242.700 500.250 243.600 ;
        RECT 457.950 233.850 460.050 235.950 ;
        RECT 460.950 235.050 463.050 237.150 ;
        RECT 472.950 233.850 475.050 235.950 ;
        RECT 478.950 233.850 481.050 235.950 ;
        RECT 481.950 235.050 484.050 237.150 ;
        RECT 493.950 236.850 496.050 238.950 ;
        RECT 494.100 235.050 495.900 236.850 ;
        RECT 433.950 232.050 435.750 233.850 ;
        RECT 436.950 230.850 439.050 232.950 ;
        RECT 440.100 232.050 441.900 233.850 ;
        RECT 437.100 229.050 438.900 230.850 ;
        RECT 431.250 225.900 438.300 226.800 ;
        RECT 431.250 225.600 432.450 225.900 ;
        RECT 389.550 219.750 391.350 225.000 ;
        RECT 392.550 219.750 394.350 225.600 ;
        RECT 407.550 219.750 409.350 225.600 ;
        RECT 410.550 219.750 412.350 225.600 ;
        RECT 413.550 219.750 415.350 225.600 ;
        RECT 430.650 219.750 432.450 225.600 ;
        RECT 436.650 225.600 438.300 225.900 ;
        RECT 458.250 225.600 459.450 233.850 ;
        RECT 473.100 232.050 474.900 233.850 ;
        RECT 475.950 230.850 478.050 232.950 ;
        RECT 479.250 232.050 481.050 233.850 ;
        RECT 476.100 229.050 477.900 230.850 ;
        RECT 482.700 226.800 483.750 235.050 ;
        RECT 498.000 234.300 499.050 242.700 ;
        RECT 501.150 238.950 502.350 245.400 ;
        RECT 515.850 244.200 517.650 251.250 ;
        RECT 520.350 245.400 522.150 251.250 ;
        RECT 535.650 245.400 537.450 251.250 ;
        RECT 515.850 243.300 519.450 244.200 ;
        RECT 499.950 236.850 502.350 238.950 ;
        RECT 515.100 237.150 516.900 238.950 ;
        RECT 498.000 233.400 500.250 234.300 ;
        RECT 476.700 225.900 483.750 226.800 ;
        RECT 476.700 225.600 478.350 225.900 ;
        RECT 433.650 219.750 435.450 225.000 ;
        RECT 436.650 219.750 438.450 225.600 ;
        RECT 439.650 219.750 441.450 225.600 ;
        RECT 454.650 219.750 456.450 225.600 ;
        RECT 457.650 219.750 459.450 225.600 ;
        RECT 460.650 219.750 462.450 225.600 ;
        RECT 473.550 219.750 475.350 225.600 ;
        RECT 476.550 219.750 478.350 225.600 ;
        RECT 482.550 225.600 483.750 225.900 ;
        RECT 494.550 232.500 500.250 233.400 ;
        RECT 494.550 225.600 495.750 232.500 ;
        RECT 501.150 231.600 502.350 236.850 ;
        RECT 514.950 235.050 517.050 237.150 ;
        RECT 518.250 235.950 519.450 243.300 ;
        RECT 536.250 243.300 537.450 245.400 ;
        RECT 538.650 246.300 540.450 251.250 ;
        RECT 541.650 247.200 543.450 251.250 ;
        RECT 544.650 246.300 546.450 251.250 ;
        RECT 538.650 244.950 546.450 246.300 ;
        RECT 536.250 242.250 540.000 243.300 ;
        RECT 560.100 243.000 561.900 251.250 ;
        RECT 538.950 238.950 540.150 242.250 ;
        RECT 542.100 240.150 543.900 241.950 ;
        RECT 557.400 241.350 561.900 243.000 ;
        RECT 565.500 242.400 567.300 251.250 ;
        RECT 579.000 245.400 580.800 251.250 ;
        RECT 583.200 247.050 585.000 251.250 ;
        RECT 586.500 248.400 588.300 251.250 ;
        RECT 601.650 248.400 603.450 251.250 ;
        RECT 604.650 248.400 606.450 251.250 ;
        RECT 583.200 245.400 588.900 247.050 ;
        RECT 521.100 237.150 522.900 238.950 ;
        RECT 517.950 233.850 520.050 235.950 ;
        RECT 520.950 235.050 523.050 237.150 ;
        RECT 538.950 236.850 541.050 238.950 ;
        RECT 541.950 238.050 544.050 240.150 ;
        RECT 544.950 236.850 547.050 238.950 ;
        RECT 557.400 237.150 558.600 241.350 ;
        RECT 578.100 240.150 579.900 241.950 ;
        RECT 577.950 238.050 580.050 240.150 ;
        RECT 580.950 239.850 583.050 241.950 ;
        RECT 584.100 240.150 585.900 241.950 ;
        RECT 581.100 238.050 582.900 239.850 ;
        RECT 583.950 238.050 586.050 240.150 ;
        RECT 587.700 238.950 588.900 245.400 ;
        RECT 602.400 240.150 603.600 248.400 ;
        RECT 608.550 245.400 610.350 251.250 ;
        RECT 611.850 248.400 613.650 251.250 ;
        RECT 616.350 248.400 618.150 251.250 ;
        RECT 620.550 248.400 622.350 251.250 ;
        RECT 624.450 248.400 626.250 251.250 ;
        RECT 627.750 248.400 629.550 251.250 ;
        RECT 632.250 249.300 634.050 251.250 ;
        RECT 632.250 248.400 636.000 249.300 ;
        RECT 637.050 248.400 638.850 251.250 ;
        RECT 616.650 247.500 617.700 248.400 ;
        RECT 613.950 246.300 617.700 247.500 ;
        RECT 625.200 246.600 626.250 248.400 ;
        RECT 634.950 247.500 636.000 248.400 ;
        RECT 613.950 245.400 616.050 246.300 ;
        RECT 608.550 243.150 609.750 245.400 ;
        RECT 621.150 244.200 622.950 246.000 ;
        RECT 625.200 245.550 630.150 246.600 ;
        RECT 628.350 244.800 630.150 245.550 ;
        RECT 631.650 244.800 633.450 246.600 ;
        RECT 634.950 245.400 637.050 247.500 ;
        RECT 640.050 245.400 641.850 251.250 ;
        RECT 622.050 243.900 622.950 244.200 ;
        RECT 632.100 243.900 633.150 244.800 ;
        RECT 535.950 233.850 538.050 235.950 ;
        RECT 479.550 219.750 481.350 225.000 ;
        RECT 482.550 219.750 484.350 225.600 ;
        RECT 494.550 219.750 496.350 225.600 ;
        RECT 497.850 219.750 499.650 231.600 ;
        RECT 500.850 219.750 502.650 231.600 ;
        RECT 518.250 225.600 519.450 233.850 ;
        RECT 536.250 232.050 538.050 233.850 ;
        RECT 539.850 231.600 541.050 236.850 ;
        RECT 545.100 235.050 546.900 236.850 ;
        RECT 556.950 235.050 559.050 237.150 ;
        RECT 586.950 236.850 589.050 238.950 ;
        RECT 601.950 238.050 604.050 240.150 ;
        RECT 604.950 239.850 607.050 241.950 ;
        RECT 608.550 241.050 613.050 243.150 ;
        RECT 622.050 243.000 633.150 243.900 ;
        RECT 605.100 238.050 606.900 239.850 ;
        RECT 514.650 219.750 516.450 225.600 ;
        RECT 517.650 219.750 519.450 225.600 ;
        RECT 520.650 219.750 522.450 225.600 ;
        RECT 536.400 219.750 538.200 225.600 ;
        RECT 539.700 219.750 541.500 231.600 ;
        RECT 543.900 219.750 545.700 231.600 ;
        RECT 557.250 226.800 558.300 235.050 ;
        RECT 559.950 233.850 562.050 235.950 ;
        RECT 565.950 233.850 568.050 235.950 ;
        RECT 559.950 232.050 561.750 233.850 ;
        RECT 562.950 230.850 565.050 232.950 ;
        RECT 566.100 232.050 567.900 233.850 ;
        RECT 587.700 231.600 588.900 236.850 ;
        RECT 563.100 229.050 564.900 230.850 ;
        RECT 578.550 230.700 586.350 231.600 ;
        RECT 557.250 225.900 564.300 226.800 ;
        RECT 557.250 225.600 558.450 225.900 ;
        RECT 556.650 219.750 558.450 225.600 ;
        RECT 562.650 225.600 564.300 225.900 ;
        RECT 559.650 219.750 561.450 225.000 ;
        RECT 562.650 219.750 564.450 225.600 ;
        RECT 565.650 219.750 567.450 225.600 ;
        RECT 578.550 219.750 580.350 230.700 ;
        RECT 581.550 219.750 583.350 229.800 ;
        RECT 584.550 219.750 586.350 230.700 ;
        RECT 587.550 219.750 589.350 231.600 ;
        RECT 602.400 225.600 603.600 238.050 ;
        RECT 608.550 231.600 609.750 241.050 ;
        RECT 610.950 239.250 614.850 241.050 ;
        RECT 610.950 238.950 613.050 239.250 ;
        RECT 622.050 238.950 622.950 243.000 ;
        RECT 632.100 241.800 633.150 243.000 ;
        RECT 632.100 240.600 639.000 241.800 ;
        RECT 632.100 240.000 633.900 240.600 ;
        RECT 638.100 239.850 639.000 240.600 ;
        RECT 635.100 238.950 636.900 239.700 ;
        RECT 622.050 236.850 625.050 238.950 ;
        RECT 628.950 237.900 636.900 238.950 ;
        RECT 638.100 238.050 639.900 239.850 ;
        RECT 628.950 236.850 631.050 237.900 ;
        RECT 610.950 233.400 612.750 235.200 ;
        RECT 611.850 232.200 616.050 233.400 ;
        RECT 622.050 232.200 622.950 236.850 ;
        RECT 630.750 233.100 632.550 233.400 ;
        RECT 601.650 219.750 603.450 225.600 ;
        RECT 604.650 219.750 606.450 225.600 ;
        RECT 608.550 219.750 610.350 231.600 ;
        RECT 613.950 231.300 616.050 232.200 ;
        RECT 616.950 231.300 622.950 232.200 ;
        RECT 624.150 232.800 632.550 233.100 ;
        RECT 640.950 232.800 641.850 245.400 ;
        RECT 653.550 246.300 655.350 251.250 ;
        RECT 656.550 247.200 658.350 251.250 ;
        RECT 659.550 246.300 661.350 251.250 ;
        RECT 653.550 244.950 661.350 246.300 ;
        RECT 662.550 245.400 664.350 251.250 ;
        RECT 677.850 245.400 679.650 251.250 ;
        RECT 662.550 243.300 663.750 245.400 ;
        RECT 682.350 244.200 684.150 251.250 ;
        RECT 695.850 245.400 697.650 251.250 ;
        RECT 700.350 244.200 702.150 251.250 ;
        RECT 713.550 246.300 715.350 251.250 ;
        RECT 716.550 247.200 718.350 251.250 ;
        RECT 719.550 246.300 721.350 251.250 ;
        RECT 713.550 244.950 721.350 246.300 ;
        RECT 722.550 245.400 724.350 251.250 ;
        RECT 734.550 248.400 736.350 251.250 ;
        RECT 737.550 248.400 739.350 251.250 ;
        RECT 752.550 248.400 754.350 251.250 ;
        RECT 755.550 248.400 757.350 251.250 ;
        RECT 758.550 248.400 760.350 251.250 ;
        RECT 660.000 242.250 663.750 243.300 ;
        RECT 680.550 243.300 684.150 244.200 ;
        RECT 698.550 243.300 702.150 244.200 ;
        RECT 722.550 243.300 723.750 245.400 ;
        RECT 656.100 240.150 657.900 241.950 ;
        RECT 652.950 236.850 655.050 238.950 ;
        RECT 655.950 238.050 658.050 240.150 ;
        RECT 659.850 238.950 661.050 242.250 ;
        RECT 658.950 236.850 661.050 238.950 ;
        RECT 677.100 237.150 678.900 238.950 ;
        RECT 653.100 235.050 654.900 236.850 ;
        RECT 624.150 232.200 641.850 232.800 ;
        RECT 616.950 230.400 617.850 231.300 ;
        RECT 615.150 228.600 617.850 230.400 ;
        RECT 618.750 230.100 620.550 230.400 ;
        RECT 624.150 230.100 625.050 232.200 ;
        RECT 630.750 231.600 641.850 232.200 ;
        RECT 658.950 231.600 660.150 236.850 ;
        RECT 661.950 233.850 664.050 235.950 ;
        RECT 676.950 235.050 679.050 237.150 ;
        RECT 680.550 235.950 681.750 243.300 ;
        RECT 683.100 237.150 684.900 238.950 ;
        RECT 695.100 237.150 696.900 238.950 ;
        RECT 679.950 233.850 682.050 235.950 ;
        RECT 682.950 235.050 685.050 237.150 ;
        RECT 694.950 235.050 697.050 237.150 ;
        RECT 698.550 235.950 699.750 243.300 ;
        RECT 720.000 242.250 723.750 243.300 ;
        RECT 716.100 240.150 717.900 241.950 ;
        RECT 701.100 237.150 702.900 238.950 ;
        RECT 697.950 233.850 700.050 235.950 ;
        RECT 700.950 235.050 703.050 237.150 ;
        RECT 712.950 236.850 715.050 238.950 ;
        RECT 715.950 238.050 718.050 240.150 ;
        RECT 719.850 238.950 721.050 242.250 ;
        RECT 733.950 239.850 736.050 241.950 ;
        RECT 737.400 240.150 738.600 248.400 ;
        RECT 756.450 244.200 757.350 248.400 ;
        RECT 761.550 245.400 763.350 251.250 ;
        RECT 773.550 246.300 775.350 251.250 ;
        RECT 776.550 247.200 778.350 251.250 ;
        RECT 779.550 246.300 781.350 251.250 ;
        RECT 756.450 243.300 759.750 244.200 ;
        RECT 757.950 242.400 759.750 243.300 ;
        RECT 718.950 236.850 721.050 238.950 ;
        RECT 734.100 238.050 735.900 239.850 ;
        RECT 736.950 238.050 739.050 240.150 ;
        RECT 751.950 239.850 754.050 241.950 ;
        RECT 752.100 238.050 753.900 239.850 ;
        RECT 713.100 235.050 714.900 236.850 ;
        RECT 661.950 232.050 663.750 233.850 ;
        RECT 618.750 229.200 625.050 230.100 ;
        RECT 625.950 230.700 627.750 231.300 ;
        RECT 625.950 229.500 633.450 230.700 ;
        RECT 618.750 228.600 620.550 229.200 ;
        RECT 632.250 228.600 633.450 229.500 ;
        RECT 613.950 225.600 617.850 227.700 ;
        RECT 622.950 226.500 629.850 228.300 ;
        RECT 632.250 226.500 637.050 228.600 ;
        RECT 611.550 219.750 613.350 222.600 ;
        RECT 616.050 219.750 617.850 225.600 ;
        RECT 620.250 219.750 622.050 225.600 ;
        RECT 624.150 219.750 625.950 226.500 ;
        RECT 632.250 225.600 633.450 226.500 ;
        RECT 627.150 219.750 628.950 225.600 ;
        RECT 631.950 219.750 633.750 225.600 ;
        RECT 637.050 219.750 638.850 225.600 ;
        RECT 640.050 219.750 641.850 231.600 ;
        RECT 654.300 219.750 656.100 231.600 ;
        RECT 658.500 219.750 660.300 231.600 ;
        RECT 680.550 225.600 681.750 233.850 ;
        RECT 698.550 225.600 699.750 233.850 ;
        RECT 718.950 231.600 720.150 236.850 ;
        RECT 721.950 233.850 724.050 235.950 ;
        RECT 721.950 232.050 723.750 233.850 ;
        RECT 661.800 219.750 663.600 225.600 ;
        RECT 677.550 219.750 679.350 225.600 ;
        RECT 680.550 219.750 682.350 225.600 ;
        RECT 683.550 219.750 685.350 225.600 ;
        RECT 695.550 219.750 697.350 225.600 ;
        RECT 698.550 219.750 700.350 225.600 ;
        RECT 701.550 219.750 703.350 225.600 ;
        RECT 714.300 219.750 716.100 231.600 ;
        RECT 718.500 219.750 720.300 231.600 ;
        RECT 737.400 225.600 738.600 238.050 ;
        RECT 754.950 236.850 757.050 238.950 ;
        RECT 755.100 235.050 756.900 236.850 ;
        RECT 758.700 234.150 759.600 242.400 ;
        RECT 762.000 240.150 763.050 245.400 ;
        RECT 773.550 244.950 781.350 246.300 ;
        RECT 782.550 245.400 784.350 251.250 ;
        RECT 798.150 246.900 799.950 251.250 ;
        RECT 796.650 245.400 799.950 246.900 ;
        RECT 801.150 245.400 802.950 251.250 ;
        RECT 782.550 243.300 783.750 245.400 ;
        RECT 780.000 242.250 783.750 243.300 ;
        RECT 776.100 240.150 777.900 241.950 ;
        RECT 760.950 238.050 763.050 240.150 ;
        RECT 757.950 234.000 759.750 234.150 ;
        RECT 752.550 232.800 759.750 234.000 ;
        RECT 752.550 231.600 753.750 232.800 ;
        RECT 757.950 232.350 759.750 232.800 ;
        RECT 721.800 219.750 723.600 225.600 ;
        RECT 734.550 219.750 736.350 225.600 ;
        RECT 737.550 219.750 739.350 225.600 ;
        RECT 752.550 219.750 754.350 231.600 ;
        RECT 761.100 231.450 762.450 238.050 ;
        RECT 772.950 236.850 775.050 238.950 ;
        RECT 775.950 238.050 778.050 240.150 ;
        RECT 779.850 238.950 781.050 242.250 ;
        RECT 778.950 236.850 781.050 238.950 ;
        RECT 796.650 238.950 797.850 245.400 ;
        RECT 799.950 243.900 801.750 244.500 ;
        RECT 805.650 243.900 807.450 251.250 ;
        RECT 818.550 248.400 820.350 251.250 ;
        RECT 821.550 248.400 823.350 251.250 ;
        RECT 824.550 248.400 826.350 251.250 ;
        RECT 799.950 242.700 807.450 243.900 ;
        RECT 796.650 236.850 799.050 238.950 ;
        RECT 800.100 237.150 801.900 238.950 ;
        RECT 773.100 235.050 774.900 236.850 ;
        RECT 778.950 231.600 780.150 236.850 ;
        RECT 781.950 233.850 784.050 235.950 ;
        RECT 781.950 232.050 783.750 233.850 ;
        RECT 796.650 231.600 797.850 236.850 ;
        RECT 799.950 235.050 802.050 237.150 ;
        RECT 757.050 219.750 758.850 231.450 ;
        RECT 760.050 230.100 762.450 231.450 ;
        RECT 760.050 219.750 761.850 230.100 ;
        RECT 774.300 219.750 776.100 231.600 ;
        RECT 778.500 219.750 780.300 231.600 ;
        RECT 781.800 219.750 783.600 225.600 ;
        RECT 796.050 219.750 797.850 231.600 ;
        RECT 799.050 219.750 800.850 231.600 ;
        RECT 803.100 225.600 804.300 242.700 ;
        RECT 822.000 241.950 823.050 248.400 ;
        RECT 836.850 245.400 838.650 251.250 ;
        RECT 841.350 244.200 843.150 251.250 ;
        RECT 858.000 245.400 859.800 251.250 ;
        RECT 862.200 245.400 864.000 251.250 ;
        RECT 866.400 245.400 868.200 251.250 ;
        RECT 820.950 239.850 823.050 241.950 ;
        RECT 805.950 236.850 808.050 238.950 ;
        RECT 817.950 236.850 820.050 238.950 ;
        RECT 806.100 235.050 807.900 236.850 ;
        RECT 818.100 235.050 819.900 236.850 ;
        RECT 822.000 232.650 823.050 239.850 ;
        RECT 839.550 243.300 843.150 244.200 ;
        RECT 823.950 236.850 826.050 238.950 ;
        RECT 836.100 237.150 837.900 238.950 ;
        RECT 824.100 235.050 825.900 236.850 ;
        RECT 835.950 235.050 838.050 237.150 ;
        RECT 839.550 235.950 840.750 243.300 ;
        RECT 860.250 240.150 862.050 241.950 ;
        RECT 842.100 237.150 843.900 238.950 ;
        RECT 838.950 233.850 841.050 235.950 ;
        RECT 841.950 235.050 844.050 237.150 ;
        RECT 856.950 236.850 859.050 238.950 ;
        RECT 859.950 238.050 862.050 240.150 ;
        RECT 862.950 238.950 864.000 245.400 ;
        RECT 865.950 240.150 867.750 241.950 ;
        RECT 862.950 236.850 865.050 238.950 ;
        RECT 865.950 238.050 868.050 240.150 ;
        RECT 868.950 236.850 871.050 238.950 ;
        RECT 857.250 235.050 859.050 236.850 ;
        RECT 822.000 231.600 824.550 232.650 ;
        RECT 802.650 219.750 804.450 225.600 ;
        RECT 805.650 219.750 807.450 225.600 ;
        RECT 818.550 219.750 820.350 231.600 ;
        RECT 822.750 219.750 824.550 231.600 ;
        RECT 839.550 225.600 840.750 233.850 ;
        RECT 864.150 233.400 865.050 236.850 ;
        RECT 869.100 235.050 870.900 236.850 ;
        RECT 864.150 232.500 868.200 233.400 ;
        RECT 866.400 231.600 868.200 232.500 ;
        RECT 857.550 230.400 865.350 231.300 ;
        RECT 836.550 219.750 838.350 225.600 ;
        RECT 839.550 219.750 841.350 225.600 ;
        RECT 842.550 219.750 844.350 225.600 ;
        RECT 857.550 219.750 859.350 230.400 ;
        RECT 860.550 219.750 862.350 229.500 ;
        RECT 863.550 220.500 865.350 230.400 ;
        RECT 866.550 221.400 868.350 231.600 ;
        RECT 869.550 220.500 871.350 231.600 ;
        RECT 863.550 219.750 871.350 220.500 ;
        RECT 10.650 209.400 12.450 215.250 ;
        RECT 13.650 209.400 15.450 215.250 ;
        RECT 16.650 209.400 18.450 215.250 ;
        RECT 14.250 201.150 15.450 209.400 ;
        RECT 28.650 203.400 30.450 215.250 ;
        RECT 31.650 202.500 33.450 215.250 ;
        RECT 34.650 203.400 36.450 215.250 ;
        RECT 37.650 202.500 39.450 215.250 ;
        RECT 40.650 203.400 42.450 215.250 ;
        RECT 43.650 202.500 45.450 215.250 ;
        RECT 46.650 203.400 48.450 215.250 ;
        RECT 49.650 202.500 51.450 215.250 ;
        RECT 52.650 203.400 54.450 215.250 ;
        RECT 64.650 209.400 66.450 215.250 ;
        RECT 67.650 209.400 69.450 215.250 ;
        RECT 30.750 201.300 33.450 202.500 ;
        RECT 35.700 201.300 39.450 202.500 ;
        RECT 41.700 201.300 45.450 202.500 ;
        RECT 47.550 201.300 51.450 202.500 ;
        RECT 10.950 197.850 13.050 199.950 ;
        RECT 13.950 199.050 16.050 201.150 ;
        RECT 11.100 196.050 12.900 197.850 ;
        RECT 14.250 191.700 15.450 199.050 ;
        RECT 16.950 197.850 19.050 199.950 ;
        RECT 17.100 196.050 18.900 197.850 ;
        RECT 30.750 196.950 31.800 201.300 ;
        RECT 28.950 194.850 31.800 196.950 ;
        RECT 11.850 190.800 15.450 191.700 ;
        RECT 30.750 191.700 31.800 194.850 ;
        RECT 35.700 194.400 36.900 201.300 ;
        RECT 41.700 194.400 42.900 201.300 ;
        RECT 47.550 194.400 48.750 201.300 ;
        RECT 65.400 196.950 66.600 209.400 ;
        RECT 71.550 203.400 73.350 215.250 ;
        RECT 74.550 212.400 76.350 215.250 ;
        RECT 79.050 209.400 80.850 215.250 ;
        RECT 83.250 209.400 85.050 215.250 ;
        RECT 76.950 207.300 80.850 209.400 ;
        RECT 87.150 208.500 88.950 215.250 ;
        RECT 90.150 209.400 91.950 215.250 ;
        RECT 94.950 209.400 96.750 215.250 ;
        RECT 100.050 209.400 101.850 215.250 ;
        RECT 95.250 208.500 96.450 209.400 ;
        RECT 85.950 206.700 92.850 208.500 ;
        RECT 95.250 206.400 100.050 208.500 ;
        RECT 78.150 204.600 80.850 206.400 ;
        RECT 81.750 205.800 83.550 206.400 ;
        RECT 81.750 204.900 88.050 205.800 ;
        RECT 95.250 205.500 96.450 206.400 ;
        RECT 81.750 204.600 83.550 204.900 ;
        RECT 79.950 203.700 80.850 204.600 ;
        RECT 49.950 194.850 52.050 196.950 ;
        RECT 64.950 194.850 67.050 196.950 ;
        RECT 68.100 195.150 69.900 196.950 ;
        RECT 32.700 192.600 36.900 194.400 ;
        RECT 38.700 192.600 42.900 194.400 ;
        RECT 44.700 192.600 48.750 194.400 ;
        RECT 50.100 193.050 51.900 194.850 ;
        RECT 35.700 191.700 36.900 192.600 ;
        RECT 41.700 191.700 42.900 192.600 ;
        RECT 47.550 191.700 48.750 192.600 ;
        RECT 11.850 183.750 13.650 190.800 ;
        RECT 30.750 190.650 33.600 191.700 ;
        RECT 30.900 190.500 33.600 190.650 ;
        RECT 35.700 190.500 39.600 191.700 ;
        RECT 41.700 190.500 45.450 191.700 ;
        RECT 47.550 190.500 51.600 191.700 ;
        RECT 31.800 189.600 33.600 190.500 ;
        RECT 37.800 189.600 39.600 190.500 ;
        RECT 16.350 183.750 18.150 189.600 ;
        RECT 28.650 183.750 30.450 189.600 ;
        RECT 31.650 183.750 33.450 189.600 ;
        RECT 34.650 183.750 36.450 189.600 ;
        RECT 37.650 183.750 39.450 189.600 ;
        RECT 40.650 183.750 42.450 189.600 ;
        RECT 43.650 183.750 45.450 190.500 ;
        RECT 49.800 189.600 51.600 190.500 ;
        RECT 46.650 183.750 48.450 189.600 ;
        RECT 49.650 183.750 51.450 189.600 ;
        RECT 52.650 183.750 54.450 189.600 ;
        RECT 65.400 186.600 66.600 194.850 ;
        RECT 67.950 193.050 70.050 195.150 ;
        RECT 71.550 193.950 72.750 203.400 ;
        RECT 76.950 202.800 79.050 203.700 ;
        RECT 79.950 202.800 85.950 203.700 ;
        RECT 74.850 201.600 79.050 202.800 ;
        RECT 73.950 199.800 75.750 201.600 ;
        RECT 85.050 198.150 85.950 202.800 ;
        RECT 87.150 202.800 88.050 204.900 ;
        RECT 88.950 204.300 96.450 205.500 ;
        RECT 88.950 203.700 90.750 204.300 ;
        RECT 103.050 203.400 104.850 215.250 ;
        RECT 118.650 209.400 120.450 215.250 ;
        RECT 121.650 209.400 123.450 215.250 ;
        RECT 124.650 209.400 126.450 215.250 ;
        RECT 137.400 209.400 139.200 215.250 ;
        RECT 93.750 202.800 104.850 203.400 ;
        RECT 87.150 202.200 104.850 202.800 ;
        RECT 87.150 201.900 95.550 202.200 ;
        RECT 93.750 201.600 95.550 201.900 ;
        RECT 85.050 196.050 88.050 198.150 ;
        RECT 91.950 197.100 94.050 198.150 ;
        RECT 91.950 196.050 99.900 197.100 ;
        RECT 73.950 195.750 76.050 196.050 ;
        RECT 73.950 193.950 77.850 195.750 ;
        RECT 71.550 191.850 76.050 193.950 ;
        RECT 85.050 192.000 85.950 196.050 ;
        RECT 98.100 195.300 99.900 196.050 ;
        RECT 101.100 195.150 102.900 196.950 ;
        RECT 95.100 194.400 96.900 195.000 ;
        RECT 101.100 194.400 102.000 195.150 ;
        RECT 95.100 193.200 102.000 194.400 ;
        RECT 95.100 192.000 96.150 193.200 ;
        RECT 71.550 189.600 72.750 191.850 ;
        RECT 85.050 191.100 96.150 192.000 ;
        RECT 85.050 190.800 85.950 191.100 ;
        RECT 64.650 183.750 66.450 186.600 ;
        RECT 67.650 183.750 69.450 186.600 ;
        RECT 71.550 183.750 73.350 189.600 ;
        RECT 76.950 188.700 79.050 189.600 ;
        RECT 84.150 189.000 85.950 190.800 ;
        RECT 95.100 190.200 96.150 191.100 ;
        RECT 91.350 189.450 93.150 190.200 ;
        RECT 76.950 187.500 80.700 188.700 ;
        RECT 79.650 186.600 80.700 187.500 ;
        RECT 88.200 188.400 93.150 189.450 ;
        RECT 94.650 188.400 96.450 190.200 ;
        RECT 103.950 189.600 104.850 202.200 ;
        RECT 122.250 201.150 123.450 209.400 ;
        RECT 140.700 203.400 142.500 215.250 ;
        RECT 144.900 203.400 146.700 215.250 ;
        RECT 158.400 209.400 160.200 215.250 ;
        RECT 161.700 203.400 163.500 215.250 ;
        RECT 165.900 203.400 167.700 215.250 ;
        RECT 177.300 203.400 179.100 215.250 ;
        RECT 181.500 203.400 183.300 215.250 ;
        RECT 184.800 209.400 186.600 215.250 ;
        RECT 200.550 209.400 202.350 215.250 ;
        RECT 203.550 209.400 205.350 215.250 ;
        RECT 137.250 201.150 139.050 202.950 ;
        RECT 118.950 197.850 121.050 199.950 ;
        RECT 121.950 199.050 124.050 201.150 ;
        RECT 119.100 196.050 120.900 197.850 ;
        RECT 122.250 191.700 123.450 199.050 ;
        RECT 124.950 197.850 127.050 199.950 ;
        RECT 136.950 199.050 139.050 201.150 ;
        RECT 140.850 198.150 142.050 203.400 ;
        RECT 158.250 201.150 160.050 202.950 ;
        RECT 146.100 198.150 147.900 199.950 ;
        RECT 157.950 199.050 160.050 201.150 ;
        RECT 161.850 198.150 163.050 203.400 ;
        RECT 167.100 198.150 168.900 199.950 ;
        RECT 176.100 198.150 177.900 199.950 ;
        RECT 181.950 198.150 183.150 203.400 ;
        RECT 184.950 201.150 186.750 202.950 ;
        RECT 184.950 199.050 187.050 201.150 ;
        RECT 125.100 196.050 126.900 197.850 ;
        RECT 139.950 196.050 142.050 198.150 ;
        RECT 139.950 192.750 141.150 196.050 ;
        RECT 142.950 194.850 145.050 196.950 ;
        RECT 145.950 196.050 148.050 198.150 ;
        RECT 160.950 196.050 163.050 198.150 ;
        RECT 143.100 193.050 144.900 194.850 ;
        RECT 160.950 192.750 162.150 196.050 ;
        RECT 163.950 194.850 166.050 196.950 ;
        RECT 166.950 196.050 169.050 198.150 ;
        RECT 175.950 196.050 178.050 198.150 ;
        RECT 178.950 194.850 181.050 196.950 ;
        RECT 181.950 196.050 184.050 198.150 ;
        RECT 203.400 196.950 204.600 209.400 ;
        RECT 216.300 203.400 218.100 215.250 ;
        RECT 220.500 203.400 222.300 215.250 ;
        RECT 223.800 209.400 225.600 215.250 ;
        RECT 240.300 203.400 242.100 215.250 ;
        RECT 244.500 203.400 246.300 215.250 ;
        RECT 247.800 209.400 249.600 215.250 ;
        RECT 260.550 209.400 262.350 215.250 ;
        RECT 263.550 209.400 265.350 215.250 ;
        RECT 266.550 209.400 268.350 215.250 ;
        RECT 215.100 198.150 216.900 199.950 ;
        RECT 220.950 198.150 222.150 203.400 ;
        RECT 223.950 201.150 225.750 202.950 ;
        RECT 223.950 199.050 226.050 201.150 ;
        RECT 239.100 198.150 240.900 199.950 ;
        RECT 244.950 198.150 246.150 203.400 ;
        RECT 247.950 201.150 249.750 202.950 ;
        RECT 263.550 201.150 264.750 209.400 ;
        RECT 283.350 203.400 285.150 215.250 ;
        RECT 286.350 203.400 288.150 215.250 ;
        RECT 289.650 209.400 291.450 215.250 ;
        RECT 304.650 209.400 306.450 215.250 ;
        RECT 307.650 209.400 309.450 215.250 ;
        RECT 310.650 209.400 312.450 215.250 ;
        RECT 323.400 209.400 325.200 215.250 ;
        RECT 247.950 199.050 250.050 201.150 ;
        RECT 164.100 193.050 165.900 194.850 ;
        RECT 179.100 193.050 180.900 194.850 ;
        RECT 182.850 192.750 184.050 196.050 ;
        RECT 200.100 195.150 201.900 196.950 ;
        RECT 199.950 193.050 202.050 195.150 ;
        RECT 202.950 194.850 205.050 196.950 ;
        RECT 214.950 196.050 217.050 198.150 ;
        RECT 217.950 194.850 220.050 196.950 ;
        RECT 220.950 196.050 223.050 198.150 ;
        RECT 238.950 196.050 241.050 198.150 ;
        RECT 88.200 186.600 89.250 188.400 ;
        RECT 97.950 187.500 100.050 189.600 ;
        RECT 97.950 186.600 99.000 187.500 ;
        RECT 74.850 183.750 76.650 186.600 ;
        RECT 79.350 183.750 81.150 186.600 ;
        RECT 83.550 183.750 85.350 186.600 ;
        RECT 87.450 183.750 89.250 186.600 ;
        RECT 90.750 183.750 92.550 186.600 ;
        RECT 95.250 185.700 99.000 186.600 ;
        RECT 95.250 183.750 97.050 185.700 ;
        RECT 100.050 183.750 101.850 186.600 ;
        RECT 103.050 183.750 104.850 189.600 ;
        RECT 119.850 190.800 123.450 191.700 ;
        RECT 137.250 191.700 141.000 192.750 ;
        RECT 158.250 191.700 162.000 192.750 ;
        RECT 183.000 191.700 186.750 192.750 ;
        RECT 119.850 183.750 121.650 190.800 ;
        RECT 137.250 189.600 138.450 191.700 ;
        RECT 124.350 183.750 126.150 189.600 ;
        RECT 136.650 183.750 138.450 189.600 ;
        RECT 139.650 188.700 147.450 190.050 ;
        RECT 158.250 189.600 159.450 191.700 ;
        RECT 139.650 183.750 141.450 188.700 ;
        RECT 142.650 183.750 144.450 187.800 ;
        RECT 145.650 183.750 147.450 188.700 ;
        RECT 157.650 183.750 159.450 189.600 ;
        RECT 160.650 188.700 168.450 190.050 ;
        RECT 160.650 183.750 162.450 188.700 ;
        RECT 163.650 183.750 165.450 187.800 ;
        RECT 166.650 183.750 168.450 188.700 ;
        RECT 176.550 188.700 184.350 190.050 ;
        RECT 176.550 183.750 178.350 188.700 ;
        RECT 179.550 183.750 181.350 187.800 ;
        RECT 182.550 183.750 184.350 188.700 ;
        RECT 185.550 189.600 186.750 191.700 ;
        RECT 185.550 183.750 187.350 189.600 ;
        RECT 203.400 186.600 204.600 194.850 ;
        RECT 218.100 193.050 219.900 194.850 ;
        RECT 221.850 192.750 223.050 196.050 ;
        RECT 241.950 194.850 244.050 196.950 ;
        RECT 244.950 196.050 247.050 198.150 ;
        RECT 259.950 197.850 262.050 199.950 ;
        RECT 262.950 199.050 265.050 201.150 ;
        RECT 260.100 196.050 261.900 197.850 ;
        RECT 242.100 193.050 243.900 194.850 ;
        RECT 245.850 192.750 247.050 196.050 ;
        RECT 222.000 191.700 225.750 192.750 ;
        RECT 246.000 191.700 249.750 192.750 ;
        RECT 215.550 188.700 223.350 190.050 ;
        RECT 200.550 183.750 202.350 186.600 ;
        RECT 203.550 183.750 205.350 186.600 ;
        RECT 215.550 183.750 217.350 188.700 ;
        RECT 218.550 183.750 220.350 187.800 ;
        RECT 221.550 183.750 223.350 188.700 ;
        RECT 224.550 189.600 225.750 191.700 ;
        RECT 224.550 183.750 226.350 189.600 ;
        RECT 239.550 188.700 247.350 190.050 ;
        RECT 239.550 183.750 241.350 188.700 ;
        RECT 242.550 183.750 244.350 187.800 ;
        RECT 245.550 183.750 247.350 188.700 ;
        RECT 248.550 189.600 249.750 191.700 ;
        RECT 263.550 191.700 264.750 199.050 ;
        RECT 265.950 197.850 268.050 199.950 ;
        RECT 283.650 198.150 284.850 203.400 ;
        RECT 290.250 202.500 291.450 209.400 ;
        RECT 285.750 201.600 291.450 202.500 ;
        RECT 285.750 200.700 288.000 201.600 ;
        RECT 308.250 201.150 309.450 209.400 ;
        RECT 326.700 203.400 328.500 215.250 ;
        RECT 330.900 203.400 332.700 215.250 ;
        RECT 336.150 203.400 337.950 215.250 ;
        RECT 339.150 209.400 340.950 215.250 ;
        RECT 344.250 209.400 346.050 215.250 ;
        RECT 349.050 209.400 350.850 215.250 ;
        RECT 344.550 208.500 345.750 209.400 ;
        RECT 352.050 208.500 353.850 215.250 ;
        RECT 355.950 209.400 357.750 215.250 ;
        RECT 360.150 209.400 361.950 215.250 ;
        RECT 364.650 212.400 366.450 215.250 ;
        RECT 340.950 206.400 345.750 208.500 ;
        RECT 348.150 206.700 355.050 208.500 ;
        RECT 360.150 207.300 364.050 209.400 ;
        RECT 344.550 205.500 345.750 206.400 ;
        RECT 357.450 205.800 359.250 206.400 ;
        RECT 344.550 204.300 352.050 205.500 ;
        RECT 350.250 203.700 352.050 204.300 ;
        RECT 352.950 204.900 359.250 205.800 ;
        RECT 323.250 201.150 325.050 202.950 ;
        RECT 266.100 196.050 267.900 197.850 ;
        RECT 283.650 196.050 286.050 198.150 ;
        RECT 263.550 190.800 267.150 191.700 ;
        RECT 248.550 183.750 250.350 189.600 ;
        RECT 260.850 183.750 262.650 189.600 ;
        RECT 265.350 183.750 267.150 190.800 ;
        RECT 283.650 189.600 284.850 196.050 ;
        RECT 286.950 192.300 288.000 200.700 ;
        RECT 290.100 198.150 291.900 199.950 ;
        RECT 289.950 196.050 292.050 198.150 ;
        RECT 304.950 197.850 307.050 199.950 ;
        RECT 307.950 199.050 310.050 201.150 ;
        RECT 305.100 196.050 306.900 197.850 ;
        RECT 285.750 191.400 288.000 192.300 ;
        RECT 308.250 191.700 309.450 199.050 ;
        RECT 310.950 197.850 313.050 199.950 ;
        RECT 322.950 199.050 325.050 201.150 ;
        RECT 326.850 198.150 328.050 203.400 ;
        RECT 336.150 202.800 347.250 203.400 ;
        RECT 352.950 202.800 353.850 204.900 ;
        RECT 357.450 204.600 359.250 204.900 ;
        RECT 360.150 204.600 362.850 206.400 ;
        RECT 360.150 203.700 361.050 204.600 ;
        RECT 336.150 202.200 353.850 202.800 ;
        RECT 332.100 198.150 333.900 199.950 ;
        RECT 311.100 196.050 312.900 197.850 ;
        RECT 325.950 196.050 328.050 198.150 ;
        RECT 325.950 192.750 327.150 196.050 ;
        RECT 328.950 194.850 331.050 196.950 ;
        RECT 331.950 196.050 334.050 198.150 ;
        RECT 329.100 193.050 330.900 194.850 ;
        RECT 285.750 190.500 290.850 191.400 ;
        RECT 283.350 183.750 285.150 189.600 ;
        RECT 286.350 183.750 288.150 189.600 ;
        RECT 289.650 186.600 290.850 190.500 ;
        RECT 305.850 190.800 309.450 191.700 ;
        RECT 323.250 191.700 327.000 192.750 ;
        RECT 289.650 183.750 291.450 186.600 ;
        RECT 305.850 183.750 307.650 190.800 ;
        RECT 323.250 189.600 324.450 191.700 ;
        RECT 310.350 183.750 312.150 189.600 ;
        RECT 322.650 183.750 324.450 189.600 ;
        RECT 325.650 188.700 333.450 190.050 ;
        RECT 325.650 183.750 327.450 188.700 ;
        RECT 328.650 183.750 330.450 187.800 ;
        RECT 331.650 183.750 333.450 188.700 ;
        RECT 336.150 189.600 337.050 202.200 ;
        RECT 345.450 201.900 353.850 202.200 ;
        RECT 355.050 202.800 361.050 203.700 ;
        RECT 361.950 202.800 364.050 203.700 ;
        RECT 367.650 203.400 369.450 215.250 ;
        RECT 382.650 209.400 384.450 215.250 ;
        RECT 385.650 209.400 387.450 215.250 ;
        RECT 388.650 209.400 390.450 215.250 ;
        RECT 401.400 209.400 403.200 215.250 ;
        RECT 345.450 201.600 347.250 201.900 ;
        RECT 355.050 198.150 355.950 202.800 ;
        RECT 361.950 201.600 366.150 202.800 ;
        RECT 365.250 199.800 367.050 201.600 ;
        RECT 346.950 197.100 349.050 198.150 ;
        RECT 338.100 195.150 339.900 196.950 ;
        RECT 341.100 196.050 349.050 197.100 ;
        RECT 352.950 196.050 355.950 198.150 ;
        RECT 341.100 195.300 342.900 196.050 ;
        RECT 339.000 194.400 339.900 195.150 ;
        RECT 344.100 194.400 345.900 195.000 ;
        RECT 339.000 193.200 345.900 194.400 ;
        RECT 344.850 192.000 345.900 193.200 ;
        RECT 355.050 192.000 355.950 196.050 ;
        RECT 364.950 195.750 367.050 196.050 ;
        RECT 363.150 193.950 367.050 195.750 ;
        RECT 368.250 193.950 369.450 203.400 ;
        RECT 386.250 201.150 387.450 209.400 ;
        RECT 404.700 203.400 406.500 215.250 ;
        RECT 408.900 203.400 410.700 215.250 ;
        RECT 423.300 203.400 425.100 215.250 ;
        RECT 427.500 203.400 429.300 215.250 ;
        RECT 430.800 209.400 432.600 215.250 ;
        RECT 443.550 209.400 445.350 215.250 ;
        RECT 446.550 209.400 448.350 215.250 ;
        RECT 449.550 209.400 451.350 215.250 ;
        RECT 401.250 201.150 403.050 202.950 ;
        RECT 382.950 197.850 385.050 199.950 ;
        RECT 385.950 199.050 388.050 201.150 ;
        RECT 383.100 196.050 384.900 197.850 ;
        RECT 344.850 191.100 355.950 192.000 ;
        RECT 364.950 191.850 369.450 193.950 ;
        RECT 344.850 190.200 345.900 191.100 ;
        RECT 355.050 190.800 355.950 191.100 ;
        RECT 336.150 183.750 337.950 189.600 ;
        RECT 340.950 187.500 343.050 189.600 ;
        RECT 344.550 188.400 346.350 190.200 ;
        RECT 347.850 189.450 349.650 190.200 ;
        RECT 347.850 188.400 352.800 189.450 ;
        RECT 355.050 189.000 356.850 190.800 ;
        RECT 368.250 189.600 369.450 191.850 ;
        RECT 386.250 191.700 387.450 199.050 ;
        RECT 388.950 197.850 391.050 199.950 ;
        RECT 400.950 199.050 403.050 201.150 ;
        RECT 404.850 198.150 406.050 203.400 ;
        RECT 410.100 198.150 411.900 199.950 ;
        RECT 422.100 198.150 423.900 199.950 ;
        RECT 427.950 198.150 429.150 203.400 ;
        RECT 430.950 201.150 432.750 202.950 ;
        RECT 446.550 201.150 447.750 209.400 ;
        RECT 462.300 203.400 464.100 215.250 ;
        RECT 466.500 203.400 468.300 215.250 ;
        RECT 469.800 209.400 471.600 215.250 ;
        RECT 487.650 209.400 489.450 215.250 ;
        RECT 490.650 209.400 492.450 215.250 ;
        RECT 493.650 209.400 495.450 215.250 ;
        RECT 430.950 199.050 433.050 201.150 ;
        RECT 389.100 196.050 390.900 197.850 ;
        RECT 403.950 196.050 406.050 198.150 ;
        RECT 403.950 192.750 405.150 196.050 ;
        RECT 406.950 194.850 409.050 196.950 ;
        RECT 409.950 196.050 412.050 198.150 ;
        RECT 421.950 196.050 424.050 198.150 ;
        RECT 424.950 194.850 427.050 196.950 ;
        RECT 427.950 196.050 430.050 198.150 ;
        RECT 442.950 197.850 445.050 199.950 ;
        RECT 445.950 199.050 448.050 201.150 ;
        RECT 443.100 196.050 444.900 197.850 ;
        RECT 407.100 193.050 408.900 194.850 ;
        RECT 425.100 193.050 426.900 194.850 ;
        RECT 428.850 192.750 430.050 196.050 ;
        RECT 361.950 188.700 364.050 189.600 ;
        RECT 342.000 186.600 343.050 187.500 ;
        RECT 351.750 186.600 352.800 188.400 ;
        RECT 360.300 187.500 364.050 188.700 ;
        RECT 360.300 186.600 361.350 187.500 ;
        RECT 339.150 183.750 340.950 186.600 ;
        RECT 342.000 185.700 345.750 186.600 ;
        RECT 343.950 183.750 345.750 185.700 ;
        RECT 348.450 183.750 350.250 186.600 ;
        RECT 351.750 183.750 353.550 186.600 ;
        RECT 355.650 183.750 357.450 186.600 ;
        RECT 359.850 183.750 361.650 186.600 ;
        RECT 364.350 183.750 366.150 186.600 ;
        RECT 367.650 183.750 369.450 189.600 ;
        RECT 383.850 190.800 387.450 191.700 ;
        RECT 401.250 191.700 405.000 192.750 ;
        RECT 429.000 191.700 432.750 192.750 ;
        RECT 383.850 183.750 385.650 190.800 ;
        RECT 401.250 189.600 402.450 191.700 ;
        RECT 388.350 183.750 390.150 189.600 ;
        RECT 400.650 183.750 402.450 189.600 ;
        RECT 403.650 188.700 411.450 190.050 ;
        RECT 403.650 183.750 405.450 188.700 ;
        RECT 406.650 183.750 408.450 187.800 ;
        RECT 409.650 183.750 411.450 188.700 ;
        RECT 422.550 188.700 430.350 190.050 ;
        RECT 422.550 183.750 424.350 188.700 ;
        RECT 425.550 183.750 427.350 187.800 ;
        RECT 428.550 183.750 430.350 188.700 ;
        RECT 431.550 189.600 432.750 191.700 ;
        RECT 446.550 191.700 447.750 199.050 ;
        RECT 448.950 197.850 451.050 199.950 ;
        RECT 461.100 198.150 462.900 199.950 ;
        RECT 466.950 198.150 468.150 203.400 ;
        RECT 469.950 201.150 471.750 202.950 ;
        RECT 491.250 201.150 492.450 209.400 ;
        RECT 504.300 203.400 506.100 215.250 ;
        RECT 508.500 203.400 510.300 215.250 ;
        RECT 511.800 209.400 513.600 215.250 ;
        RECT 526.650 209.400 528.450 215.250 ;
        RECT 529.650 209.400 531.450 215.250 ;
        RECT 532.650 209.400 534.450 215.250 ;
        RECT 469.950 199.050 472.050 201.150 ;
        RECT 449.100 196.050 450.900 197.850 ;
        RECT 460.950 196.050 463.050 198.150 ;
        RECT 463.950 194.850 466.050 196.950 ;
        RECT 466.950 196.050 469.050 198.150 ;
        RECT 487.950 197.850 490.050 199.950 ;
        RECT 490.950 199.050 493.050 201.150 ;
        RECT 488.100 196.050 489.900 197.850 ;
        RECT 464.100 193.050 465.900 194.850 ;
        RECT 467.850 192.750 469.050 196.050 ;
        RECT 468.000 191.700 471.750 192.750 ;
        RECT 491.250 191.700 492.450 199.050 ;
        RECT 493.950 197.850 496.050 199.950 ;
        RECT 503.100 198.150 504.900 199.950 ;
        RECT 508.950 198.150 510.150 203.400 ;
        RECT 511.950 201.150 513.750 202.950 ;
        RECT 530.250 201.150 531.450 209.400 ;
        RECT 536.550 203.400 538.350 215.250 ;
        RECT 539.550 212.400 541.350 215.250 ;
        RECT 544.050 209.400 545.850 215.250 ;
        RECT 548.250 209.400 550.050 215.250 ;
        RECT 541.950 207.300 545.850 209.400 ;
        RECT 552.150 208.500 553.950 215.250 ;
        RECT 555.150 209.400 556.950 215.250 ;
        RECT 559.950 209.400 561.750 215.250 ;
        RECT 565.050 209.400 566.850 215.250 ;
        RECT 560.250 208.500 561.450 209.400 ;
        RECT 550.950 206.700 557.850 208.500 ;
        RECT 560.250 206.400 565.050 208.500 ;
        RECT 543.150 204.600 545.850 206.400 ;
        RECT 546.750 205.800 548.550 206.400 ;
        RECT 546.750 204.900 553.050 205.800 ;
        RECT 560.250 205.500 561.450 206.400 ;
        RECT 546.750 204.600 548.550 204.900 ;
        RECT 544.950 203.700 545.850 204.600 ;
        RECT 511.950 199.050 514.050 201.150 ;
        RECT 494.100 196.050 495.900 197.850 ;
        RECT 502.950 196.050 505.050 198.150 ;
        RECT 505.950 194.850 508.050 196.950 ;
        RECT 508.950 196.050 511.050 198.150 ;
        RECT 526.950 197.850 529.050 199.950 ;
        RECT 529.950 199.050 532.050 201.150 ;
        RECT 527.100 196.050 528.900 197.850 ;
        RECT 506.100 193.050 507.900 194.850 ;
        RECT 509.850 192.750 511.050 196.050 ;
        RECT 510.000 191.700 513.750 192.750 ;
        RECT 530.250 191.700 531.450 199.050 ;
        RECT 532.950 197.850 535.050 199.950 ;
        RECT 533.100 196.050 534.900 197.850 ;
        RECT 446.550 190.800 450.150 191.700 ;
        RECT 431.550 183.750 433.350 189.600 ;
        RECT 443.850 183.750 445.650 189.600 ;
        RECT 448.350 183.750 450.150 190.800 ;
        RECT 461.550 188.700 469.350 190.050 ;
        RECT 461.550 183.750 463.350 188.700 ;
        RECT 464.550 183.750 466.350 187.800 ;
        RECT 467.550 183.750 469.350 188.700 ;
        RECT 470.550 189.600 471.750 191.700 ;
        RECT 488.850 190.800 492.450 191.700 ;
        RECT 470.550 183.750 472.350 189.600 ;
        RECT 488.850 183.750 490.650 190.800 ;
        RECT 493.350 183.750 495.150 189.600 ;
        RECT 503.550 188.700 511.350 190.050 ;
        RECT 503.550 183.750 505.350 188.700 ;
        RECT 506.550 183.750 508.350 187.800 ;
        RECT 509.550 183.750 511.350 188.700 ;
        RECT 512.550 189.600 513.750 191.700 ;
        RECT 527.850 190.800 531.450 191.700 ;
        RECT 536.550 193.950 537.750 203.400 ;
        RECT 541.950 202.800 544.050 203.700 ;
        RECT 544.950 202.800 550.950 203.700 ;
        RECT 539.850 201.600 544.050 202.800 ;
        RECT 538.950 199.800 540.750 201.600 ;
        RECT 550.050 198.150 550.950 202.800 ;
        RECT 552.150 202.800 553.050 204.900 ;
        RECT 553.950 204.300 561.450 205.500 ;
        RECT 553.950 203.700 555.750 204.300 ;
        RECT 568.050 203.400 569.850 215.250 ;
        RECT 579.300 203.400 581.100 215.250 ;
        RECT 583.500 203.400 585.300 215.250 ;
        RECT 586.800 209.400 588.600 215.250 ;
        RECT 602.550 209.400 604.350 215.250 ;
        RECT 605.550 209.400 607.350 215.250 ;
        RECT 608.550 209.400 610.350 215.250 ;
        RECT 620.550 209.400 622.350 215.250 ;
        RECT 623.550 209.400 625.350 215.250 ;
        RECT 626.550 209.400 628.350 215.250 ;
        RECT 643.650 209.400 645.450 215.250 ;
        RECT 646.650 209.400 648.450 215.250 ;
        RECT 649.650 209.400 651.450 215.250 ;
        RECT 659.550 209.400 661.350 215.250 ;
        RECT 662.550 209.400 664.350 215.250 ;
        RECT 558.750 202.800 569.850 203.400 ;
        RECT 552.150 202.200 569.850 202.800 ;
        RECT 552.150 201.900 560.550 202.200 ;
        RECT 558.750 201.600 560.550 201.900 ;
        RECT 550.050 196.050 553.050 198.150 ;
        RECT 556.950 197.100 559.050 198.150 ;
        RECT 556.950 196.050 564.900 197.100 ;
        RECT 538.950 195.750 541.050 196.050 ;
        RECT 538.950 193.950 542.850 195.750 ;
        RECT 536.550 191.850 541.050 193.950 ;
        RECT 550.050 192.000 550.950 196.050 ;
        RECT 563.100 195.300 564.900 196.050 ;
        RECT 566.100 195.150 567.900 196.950 ;
        RECT 560.100 194.400 561.900 195.000 ;
        RECT 566.100 194.400 567.000 195.150 ;
        RECT 560.100 193.200 567.000 194.400 ;
        RECT 560.100 192.000 561.150 193.200 ;
        RECT 512.550 183.750 514.350 189.600 ;
        RECT 527.850 183.750 529.650 190.800 ;
        RECT 536.550 189.600 537.750 191.850 ;
        RECT 550.050 191.100 561.150 192.000 ;
        RECT 550.050 190.800 550.950 191.100 ;
        RECT 532.350 183.750 534.150 189.600 ;
        RECT 536.550 183.750 538.350 189.600 ;
        RECT 541.950 188.700 544.050 189.600 ;
        RECT 549.150 189.000 550.950 190.800 ;
        RECT 560.100 190.200 561.150 191.100 ;
        RECT 556.350 189.450 558.150 190.200 ;
        RECT 541.950 187.500 545.700 188.700 ;
        RECT 544.650 186.600 545.700 187.500 ;
        RECT 553.200 188.400 558.150 189.450 ;
        RECT 559.650 188.400 561.450 190.200 ;
        RECT 568.950 189.600 569.850 202.200 ;
        RECT 578.100 198.150 579.900 199.950 ;
        RECT 583.950 198.150 585.150 203.400 ;
        RECT 586.950 201.150 588.750 202.950 ;
        RECT 605.550 201.150 606.750 209.400 ;
        RECT 623.550 201.150 624.750 209.400 ;
        RECT 647.250 201.150 648.450 209.400 ;
        RECT 586.950 199.050 589.050 201.150 ;
        RECT 577.950 196.050 580.050 198.150 ;
        RECT 580.950 194.850 583.050 196.950 ;
        RECT 583.950 196.050 586.050 198.150 ;
        RECT 601.950 197.850 604.050 199.950 ;
        RECT 604.950 199.050 607.050 201.150 ;
        RECT 602.100 196.050 603.900 197.850 ;
        RECT 581.100 193.050 582.900 194.850 ;
        RECT 584.850 192.750 586.050 196.050 ;
        RECT 585.000 191.700 588.750 192.750 ;
        RECT 553.200 186.600 554.250 188.400 ;
        RECT 562.950 187.500 565.050 189.600 ;
        RECT 562.950 186.600 564.000 187.500 ;
        RECT 539.850 183.750 541.650 186.600 ;
        RECT 544.350 183.750 546.150 186.600 ;
        RECT 548.550 183.750 550.350 186.600 ;
        RECT 552.450 183.750 554.250 186.600 ;
        RECT 555.750 183.750 557.550 186.600 ;
        RECT 560.250 185.700 564.000 186.600 ;
        RECT 560.250 183.750 562.050 185.700 ;
        RECT 565.050 183.750 566.850 186.600 ;
        RECT 568.050 183.750 569.850 189.600 ;
        RECT 578.550 188.700 586.350 190.050 ;
        RECT 578.550 183.750 580.350 188.700 ;
        RECT 581.550 183.750 583.350 187.800 ;
        RECT 584.550 183.750 586.350 188.700 ;
        RECT 587.550 189.600 588.750 191.700 ;
        RECT 605.550 191.700 606.750 199.050 ;
        RECT 607.950 197.850 610.050 199.950 ;
        RECT 619.950 197.850 622.050 199.950 ;
        RECT 622.950 199.050 625.050 201.150 ;
        RECT 608.100 196.050 609.900 197.850 ;
        RECT 620.100 196.050 621.900 197.850 ;
        RECT 623.550 191.700 624.750 199.050 ;
        RECT 625.950 197.850 628.050 199.950 ;
        RECT 643.950 197.850 646.050 199.950 ;
        RECT 646.950 199.050 649.050 201.150 ;
        RECT 626.100 196.050 627.900 197.850 ;
        RECT 644.100 196.050 645.900 197.850 ;
        RECT 647.250 191.700 648.450 199.050 ;
        RECT 649.950 197.850 652.050 199.950 ;
        RECT 650.100 196.050 651.900 197.850 ;
        RECT 662.400 196.950 663.600 209.400 ;
        RECT 675.300 203.400 677.100 215.250 ;
        RECT 679.500 203.400 681.300 215.250 ;
        RECT 682.800 209.400 684.600 215.250 ;
        RECT 695.550 209.400 697.350 215.250 ;
        RECT 698.550 209.400 700.350 215.250 ;
        RECT 701.550 209.400 703.350 215.250 ;
        RECT 713.550 209.400 715.350 215.250 ;
        RECT 716.550 209.400 718.350 215.250 ;
        RECT 730.650 209.400 732.450 215.250 ;
        RECT 733.650 209.400 735.450 215.250 ;
        RECT 736.650 209.400 738.450 215.250 ;
        RECT 749.400 209.400 751.200 215.250 ;
        RECT 674.100 198.150 675.900 199.950 ;
        RECT 679.950 198.150 681.150 203.400 ;
        RECT 682.950 201.150 684.750 202.950 ;
        RECT 698.550 201.150 699.750 209.400 ;
        RECT 682.950 199.050 685.050 201.150 ;
        RECT 659.100 195.150 660.900 196.950 ;
        RECT 658.950 193.050 661.050 195.150 ;
        RECT 661.950 194.850 664.050 196.950 ;
        RECT 673.950 196.050 676.050 198.150 ;
        RECT 676.950 194.850 679.050 196.950 ;
        RECT 679.950 196.050 682.050 198.150 ;
        RECT 694.950 197.850 697.050 199.950 ;
        RECT 697.950 199.050 700.050 201.150 ;
        RECT 695.100 196.050 696.900 197.850 ;
        RECT 605.550 190.800 609.150 191.700 ;
        RECT 623.550 190.800 627.150 191.700 ;
        RECT 587.550 183.750 589.350 189.600 ;
        RECT 602.850 183.750 604.650 189.600 ;
        RECT 607.350 183.750 609.150 190.800 ;
        RECT 620.850 183.750 622.650 189.600 ;
        RECT 625.350 183.750 627.150 190.800 ;
        RECT 644.850 190.800 648.450 191.700 ;
        RECT 644.850 183.750 646.650 190.800 ;
        RECT 649.350 183.750 651.150 189.600 ;
        RECT 662.400 186.600 663.600 194.850 ;
        RECT 677.100 193.050 678.900 194.850 ;
        RECT 680.850 192.750 682.050 196.050 ;
        RECT 681.000 191.700 684.750 192.750 ;
        RECT 674.550 188.700 682.350 190.050 ;
        RECT 659.550 183.750 661.350 186.600 ;
        RECT 662.550 183.750 664.350 186.600 ;
        RECT 674.550 183.750 676.350 188.700 ;
        RECT 677.550 183.750 679.350 187.800 ;
        RECT 680.550 183.750 682.350 188.700 ;
        RECT 683.550 189.600 684.750 191.700 ;
        RECT 698.550 191.700 699.750 199.050 ;
        RECT 700.950 197.850 703.050 199.950 ;
        RECT 701.100 196.050 702.900 197.850 ;
        RECT 716.400 196.950 717.600 209.400 ;
        RECT 734.250 201.150 735.450 209.400 ;
        RECT 752.700 203.400 754.500 215.250 ;
        RECT 756.900 203.400 758.700 215.250 ;
        RECT 768.300 203.400 770.100 215.250 ;
        RECT 772.500 203.400 774.300 215.250 ;
        RECT 775.800 209.400 777.600 215.250 ;
        RECT 791.550 209.400 793.350 215.250 ;
        RECT 794.550 209.400 796.350 215.250 ;
        RECT 797.550 209.400 799.350 215.250 ;
        RECT 749.250 201.150 751.050 202.950 ;
        RECT 730.950 197.850 733.050 199.950 ;
        RECT 733.950 199.050 736.050 201.150 ;
        RECT 713.100 195.150 714.900 196.950 ;
        RECT 712.950 193.050 715.050 195.150 ;
        RECT 715.950 194.850 718.050 196.950 ;
        RECT 731.100 196.050 732.900 197.850 ;
        RECT 698.550 190.800 702.150 191.700 ;
        RECT 683.550 183.750 685.350 189.600 ;
        RECT 695.850 183.750 697.650 189.600 ;
        RECT 700.350 183.750 702.150 190.800 ;
        RECT 716.400 186.600 717.600 194.850 ;
        RECT 734.250 191.700 735.450 199.050 ;
        RECT 736.950 197.850 739.050 199.950 ;
        RECT 748.950 199.050 751.050 201.150 ;
        RECT 752.850 198.150 754.050 203.400 ;
        RECT 758.100 198.150 759.900 199.950 ;
        RECT 767.100 198.150 768.900 199.950 ;
        RECT 772.950 198.150 774.150 203.400 ;
        RECT 775.950 201.150 777.750 202.950 ;
        RECT 794.550 201.150 795.750 209.400 ;
        RECT 812.550 204.300 814.350 215.250 ;
        RECT 815.550 205.200 817.350 215.250 ;
        RECT 818.550 204.300 820.350 215.250 ;
        RECT 812.550 203.400 820.350 204.300 ;
        RECT 821.550 203.400 823.350 215.250 ;
        RECT 833.550 204.300 835.350 215.250 ;
        RECT 836.550 205.200 838.350 215.250 ;
        RECT 839.550 204.300 841.350 215.250 ;
        RECT 833.550 203.400 841.350 204.300 ;
        RECT 842.550 203.400 844.350 215.250 ;
        RECT 856.650 203.400 858.450 215.250 ;
        RECT 775.950 199.050 778.050 201.150 ;
        RECT 737.100 196.050 738.900 197.850 ;
        RECT 751.950 196.050 754.050 198.150 ;
        RECT 751.950 192.750 753.150 196.050 ;
        RECT 754.950 194.850 757.050 196.950 ;
        RECT 757.950 196.050 760.050 198.150 ;
        RECT 766.950 196.050 769.050 198.150 ;
        RECT 769.950 194.850 772.050 196.950 ;
        RECT 772.950 196.050 775.050 198.150 ;
        RECT 790.950 197.850 793.050 199.950 ;
        RECT 793.950 199.050 796.050 201.150 ;
        RECT 791.100 196.050 792.900 197.850 ;
        RECT 755.100 193.050 756.900 194.850 ;
        RECT 770.100 193.050 771.900 194.850 ;
        RECT 773.850 192.750 775.050 196.050 ;
        RECT 731.850 190.800 735.450 191.700 ;
        RECT 749.250 191.700 753.000 192.750 ;
        RECT 774.000 191.700 777.750 192.750 ;
        RECT 713.550 183.750 715.350 186.600 ;
        RECT 716.550 183.750 718.350 186.600 ;
        RECT 731.850 183.750 733.650 190.800 ;
        RECT 749.250 189.600 750.450 191.700 ;
        RECT 736.350 183.750 738.150 189.600 ;
        RECT 748.650 183.750 750.450 189.600 ;
        RECT 751.650 188.700 759.450 190.050 ;
        RECT 751.650 183.750 753.450 188.700 ;
        RECT 754.650 183.750 756.450 187.800 ;
        RECT 757.650 183.750 759.450 188.700 ;
        RECT 767.550 188.700 775.350 190.050 ;
        RECT 767.550 183.750 769.350 188.700 ;
        RECT 770.550 183.750 772.350 187.800 ;
        RECT 773.550 183.750 775.350 188.700 ;
        RECT 776.550 189.600 777.750 191.700 ;
        RECT 794.550 191.700 795.750 199.050 ;
        RECT 796.950 197.850 799.050 199.950 ;
        RECT 821.700 198.150 822.900 203.400 ;
        RECT 842.700 198.150 843.900 203.400 ;
        RECT 859.650 202.500 861.450 215.250 ;
        RECT 862.650 203.400 864.450 215.250 ;
        RECT 865.650 202.500 867.450 215.250 ;
        RECT 868.650 203.400 870.450 215.250 ;
        RECT 871.650 202.500 873.450 215.250 ;
        RECT 874.650 203.400 876.450 215.250 ;
        RECT 877.650 202.500 879.450 215.250 ;
        RECT 880.650 203.400 882.450 215.250 ;
        RECT 858.750 201.300 861.450 202.500 ;
        RECT 863.700 201.300 867.450 202.500 ;
        RECT 869.700 201.300 873.450 202.500 ;
        RECT 875.550 201.300 879.450 202.500 ;
        RECT 797.100 196.050 798.900 197.850 ;
        RECT 811.950 194.850 814.050 196.950 ;
        RECT 815.100 195.150 816.900 196.950 ;
        RECT 812.100 193.050 813.900 194.850 ;
        RECT 814.950 193.050 817.050 195.150 ;
        RECT 817.950 194.850 820.050 196.950 ;
        RECT 820.950 196.050 823.050 198.150 ;
        RECT 818.100 193.050 819.900 194.850 ;
        RECT 794.550 190.800 798.150 191.700 ;
        RECT 776.550 183.750 778.350 189.600 ;
        RECT 791.850 183.750 793.650 189.600 ;
        RECT 796.350 183.750 798.150 190.800 ;
        RECT 821.700 189.600 822.900 196.050 ;
        RECT 832.950 194.850 835.050 196.950 ;
        RECT 836.100 195.150 837.900 196.950 ;
        RECT 833.100 193.050 834.900 194.850 ;
        RECT 835.950 193.050 838.050 195.150 ;
        RECT 838.950 194.850 841.050 196.950 ;
        RECT 841.950 196.050 844.050 198.150 ;
        RECT 858.750 196.950 859.800 201.300 ;
        RECT 839.100 193.050 840.900 194.850 ;
        RECT 842.700 189.600 843.900 196.050 ;
        RECT 856.950 194.850 859.800 196.950 ;
        RECT 858.750 191.700 859.800 194.850 ;
        RECT 863.700 194.400 864.900 201.300 ;
        RECT 869.700 194.400 870.900 201.300 ;
        RECT 875.550 194.400 876.750 201.300 ;
        RECT 877.950 194.850 880.050 196.950 ;
        RECT 860.700 192.600 864.900 194.400 ;
        RECT 866.700 192.600 870.900 194.400 ;
        RECT 872.700 192.600 876.750 194.400 ;
        RECT 878.100 193.050 879.900 194.850 ;
        RECT 863.700 191.700 864.900 192.600 ;
        RECT 869.700 191.700 870.900 192.600 ;
        RECT 875.550 191.700 876.750 192.600 ;
        RECT 858.750 190.650 861.600 191.700 ;
        RECT 858.900 190.500 861.600 190.650 ;
        RECT 863.700 190.500 867.600 191.700 ;
        RECT 869.700 190.500 873.450 191.700 ;
        RECT 875.550 190.500 879.600 191.700 ;
        RECT 859.800 189.600 861.600 190.500 ;
        RECT 865.800 189.600 867.600 190.500 ;
        RECT 813.000 183.750 814.800 189.600 ;
        RECT 817.200 187.950 822.900 189.600 ;
        RECT 817.200 183.750 819.000 187.950 ;
        RECT 820.500 183.750 822.300 186.600 ;
        RECT 834.000 183.750 835.800 189.600 ;
        RECT 838.200 187.950 843.900 189.600 ;
        RECT 838.200 183.750 840.000 187.950 ;
        RECT 841.500 183.750 843.300 186.600 ;
        RECT 856.650 183.750 858.450 189.600 ;
        RECT 859.650 183.750 861.450 189.600 ;
        RECT 862.650 183.750 864.450 189.600 ;
        RECT 865.650 183.750 867.450 189.600 ;
        RECT 868.650 183.750 870.450 189.600 ;
        RECT 871.650 183.750 873.450 190.500 ;
        RECT 877.800 189.600 879.600 190.500 ;
        RECT 874.650 183.750 876.450 189.600 ;
        RECT 877.650 183.750 879.450 189.600 ;
        RECT 880.650 183.750 882.450 189.600 ;
        RECT 11.550 174.300 13.350 179.250 ;
        RECT 14.550 175.200 16.350 179.250 ;
        RECT 17.550 174.300 19.350 179.250 ;
        RECT 11.550 172.950 19.350 174.300 ;
        RECT 20.550 173.400 22.350 179.250 ;
        RECT 20.550 171.300 21.750 173.400 ;
        RECT 35.850 172.200 37.650 179.250 ;
        RECT 40.350 173.400 42.150 179.250 ;
        RECT 50.550 174.300 52.350 179.250 ;
        RECT 53.550 175.200 55.350 179.250 ;
        RECT 56.550 174.300 58.350 179.250 ;
        RECT 50.550 172.950 58.350 174.300 ;
        RECT 59.550 173.400 61.350 179.250 ;
        RECT 35.850 171.300 39.450 172.200 ;
        RECT 59.550 171.300 60.750 173.400 ;
        RECT 74.850 172.200 76.650 179.250 ;
        RECT 79.350 173.400 81.150 179.250 ;
        RECT 94.650 173.400 96.450 179.250 ;
        RECT 74.850 171.300 78.450 172.200 ;
        RECT 18.000 170.250 21.750 171.300 ;
        RECT 14.100 168.150 15.900 169.950 ;
        RECT 10.950 164.850 13.050 166.950 ;
        RECT 13.950 166.050 16.050 168.150 ;
        RECT 17.850 166.950 19.050 170.250 ;
        RECT 16.950 164.850 19.050 166.950 ;
        RECT 35.100 165.150 36.900 166.950 ;
        RECT 11.100 163.050 12.900 164.850 ;
        RECT 16.950 159.600 18.150 164.850 ;
        RECT 19.950 161.850 22.050 163.950 ;
        RECT 34.950 163.050 37.050 165.150 ;
        RECT 38.250 163.950 39.450 171.300 ;
        RECT 57.000 170.250 60.750 171.300 ;
        RECT 53.100 168.150 54.900 169.950 ;
        RECT 41.100 165.150 42.900 166.950 ;
        RECT 37.950 161.850 40.050 163.950 ;
        RECT 40.950 163.050 43.050 165.150 ;
        RECT 49.950 164.850 52.050 166.950 ;
        RECT 52.950 166.050 55.050 168.150 ;
        RECT 56.850 166.950 58.050 170.250 ;
        RECT 55.950 164.850 58.050 166.950 ;
        RECT 74.100 165.150 75.900 166.950 ;
        RECT 50.100 163.050 51.900 164.850 ;
        RECT 19.950 160.050 21.750 161.850 ;
        RECT 12.300 147.750 14.100 159.600 ;
        RECT 16.500 147.750 18.300 159.600 ;
        RECT 38.250 153.600 39.450 161.850 ;
        RECT 55.950 159.600 57.150 164.850 ;
        RECT 58.950 161.850 61.050 163.950 ;
        RECT 73.950 163.050 76.050 165.150 ;
        RECT 77.250 163.950 78.450 171.300 ;
        RECT 95.250 171.300 96.450 173.400 ;
        RECT 97.650 174.300 99.450 179.250 ;
        RECT 100.650 175.200 102.450 179.250 ;
        RECT 103.650 174.300 105.450 179.250 ;
        RECT 113.550 176.400 115.350 179.250 ;
        RECT 116.550 176.400 118.350 179.250 ;
        RECT 97.650 172.950 105.450 174.300 ;
        RECT 95.250 170.250 99.000 171.300 ;
        RECT 97.950 166.950 99.150 170.250 ;
        RECT 101.100 168.150 102.900 169.950 ;
        RECT 80.100 165.150 81.900 166.950 ;
        RECT 76.950 161.850 79.050 163.950 ;
        RECT 79.950 163.050 82.050 165.150 ;
        RECT 97.950 164.850 100.050 166.950 ;
        RECT 100.950 166.050 103.050 168.150 ;
        RECT 112.950 167.850 115.050 169.950 ;
        RECT 116.400 168.150 117.600 176.400 ;
        RECT 123.150 173.400 124.950 179.250 ;
        RECT 126.150 176.400 127.950 179.250 ;
        RECT 130.950 177.300 132.750 179.250 ;
        RECT 129.000 176.400 132.750 177.300 ;
        RECT 135.450 176.400 137.250 179.250 ;
        RECT 138.750 176.400 140.550 179.250 ;
        RECT 142.650 176.400 144.450 179.250 ;
        RECT 146.850 176.400 148.650 179.250 ;
        RECT 151.350 176.400 153.150 179.250 ;
        RECT 129.000 175.500 130.050 176.400 ;
        RECT 127.950 173.400 130.050 175.500 ;
        RECT 138.750 174.600 139.800 176.400 ;
        RECT 103.950 164.850 106.050 166.950 ;
        RECT 113.100 166.050 114.900 167.850 ;
        RECT 115.950 166.050 118.050 168.150 ;
        RECT 94.950 161.850 97.050 163.950 ;
        RECT 58.950 160.050 60.750 161.850 ;
        RECT 19.800 147.750 21.600 153.600 ;
        RECT 34.650 147.750 36.450 153.600 ;
        RECT 37.650 147.750 39.450 153.600 ;
        RECT 40.650 147.750 42.450 153.600 ;
        RECT 51.300 147.750 53.100 159.600 ;
        RECT 55.500 147.750 57.300 159.600 ;
        RECT 77.250 153.600 78.450 161.850 ;
        RECT 95.250 160.050 97.050 161.850 ;
        RECT 98.850 159.600 100.050 164.850 ;
        RECT 104.100 163.050 105.900 164.850 ;
        RECT 58.800 147.750 60.600 153.600 ;
        RECT 73.650 147.750 75.450 153.600 ;
        RECT 76.650 147.750 78.450 153.600 ;
        RECT 79.650 147.750 81.450 153.600 ;
        RECT 95.400 147.750 97.200 153.600 ;
        RECT 98.700 147.750 100.500 159.600 ;
        RECT 102.900 147.750 104.700 159.600 ;
        RECT 116.400 153.600 117.600 166.050 ;
        RECT 123.150 160.800 124.050 173.400 ;
        RECT 131.550 172.800 133.350 174.600 ;
        RECT 134.850 173.550 139.800 174.600 ;
        RECT 147.300 175.500 148.350 176.400 ;
        RECT 147.300 174.300 151.050 175.500 ;
        RECT 134.850 172.800 136.650 173.550 ;
        RECT 131.850 171.900 132.900 172.800 ;
        RECT 142.050 172.200 143.850 174.000 ;
        RECT 148.950 173.400 151.050 174.300 ;
        RECT 154.650 173.400 156.450 179.250 ;
        RECT 166.650 173.400 168.450 179.250 ;
        RECT 142.050 171.900 142.950 172.200 ;
        RECT 131.850 171.000 142.950 171.900 ;
        RECT 155.250 171.150 156.450 173.400 ;
        RECT 131.850 169.800 132.900 171.000 ;
        RECT 126.000 168.600 132.900 169.800 ;
        RECT 126.000 167.850 126.900 168.600 ;
        RECT 131.100 168.000 132.900 168.600 ;
        RECT 125.100 166.050 126.900 167.850 ;
        RECT 128.100 166.950 129.900 167.700 ;
        RECT 142.050 166.950 142.950 171.000 ;
        RECT 151.950 169.050 156.450 171.150 ;
        RECT 167.250 171.300 168.450 173.400 ;
        RECT 169.650 174.300 171.450 179.250 ;
        RECT 172.650 175.200 174.450 179.250 ;
        RECT 175.650 174.300 177.450 179.250 ;
        RECT 169.650 172.950 177.450 174.300 ;
        RECT 191.850 172.200 193.650 179.250 ;
        RECT 196.350 173.400 198.150 179.250 ;
        RECT 208.650 173.400 210.450 179.250 ;
        RECT 191.850 171.300 195.450 172.200 ;
        RECT 167.250 170.250 171.000 171.300 ;
        RECT 150.150 167.250 154.050 169.050 ;
        RECT 151.950 166.950 154.050 167.250 ;
        RECT 128.100 165.900 136.050 166.950 ;
        RECT 133.950 164.850 136.050 165.900 ;
        RECT 139.950 164.850 142.950 166.950 ;
        RECT 132.450 161.100 134.250 161.400 ;
        RECT 132.450 160.800 140.850 161.100 ;
        RECT 123.150 160.200 140.850 160.800 ;
        RECT 123.150 159.600 134.250 160.200 ;
        RECT 113.550 147.750 115.350 153.600 ;
        RECT 116.550 147.750 118.350 153.600 ;
        RECT 123.150 147.750 124.950 159.600 ;
        RECT 137.250 158.700 139.050 159.300 ;
        RECT 131.550 157.500 139.050 158.700 ;
        RECT 139.950 158.100 140.850 160.200 ;
        RECT 142.050 160.200 142.950 164.850 ;
        RECT 152.250 161.400 154.050 163.200 ;
        RECT 148.950 160.200 153.150 161.400 ;
        RECT 142.050 159.300 148.050 160.200 ;
        RECT 148.950 159.300 151.050 160.200 ;
        RECT 155.250 159.600 156.450 169.050 ;
        RECT 169.950 166.950 171.150 170.250 ;
        RECT 173.100 168.150 174.900 169.950 ;
        RECT 169.950 164.850 172.050 166.950 ;
        RECT 172.950 166.050 175.050 168.150 ;
        RECT 175.950 164.850 178.050 166.950 ;
        RECT 191.100 165.150 192.900 166.950 ;
        RECT 166.950 161.850 169.050 163.950 ;
        RECT 167.250 160.050 169.050 161.850 ;
        RECT 170.850 159.600 172.050 164.850 ;
        RECT 176.100 163.050 177.900 164.850 ;
        RECT 190.950 163.050 193.050 165.150 ;
        RECT 194.250 163.950 195.450 171.300 ;
        RECT 209.250 171.300 210.450 173.400 ;
        RECT 211.650 174.300 213.450 179.250 ;
        RECT 214.650 175.200 216.450 179.250 ;
        RECT 217.650 174.300 219.450 179.250 ;
        RECT 211.650 172.950 219.450 174.300 ;
        RECT 230.850 172.200 232.650 179.250 ;
        RECT 235.350 173.400 237.150 179.250 ;
        RECT 250.350 173.400 252.150 179.250 ;
        RECT 253.350 173.400 255.150 179.250 ;
        RECT 256.650 176.400 258.450 179.250 ;
        RECT 230.850 171.300 234.450 172.200 ;
        RECT 209.250 170.250 213.000 171.300 ;
        RECT 211.950 166.950 213.150 170.250 ;
        RECT 215.100 168.150 216.900 169.950 ;
        RECT 197.100 165.150 198.900 166.950 ;
        RECT 193.950 161.850 196.050 163.950 ;
        RECT 196.950 163.050 199.050 165.150 ;
        RECT 211.950 164.850 214.050 166.950 ;
        RECT 214.950 166.050 217.050 168.150 ;
        RECT 217.950 164.850 220.050 166.950 ;
        RECT 230.100 165.150 231.900 166.950 ;
        RECT 208.950 161.850 211.050 163.950 ;
        RECT 147.150 158.400 148.050 159.300 ;
        RECT 144.450 158.100 146.250 158.400 ;
        RECT 131.550 156.600 132.750 157.500 ;
        RECT 139.950 157.200 146.250 158.100 ;
        RECT 144.450 156.600 146.250 157.200 ;
        RECT 147.150 156.600 149.850 158.400 ;
        RECT 127.950 154.500 132.750 156.600 ;
        RECT 135.150 154.500 142.050 156.300 ;
        RECT 131.550 153.600 132.750 154.500 ;
        RECT 126.150 147.750 127.950 153.600 ;
        RECT 131.250 147.750 133.050 153.600 ;
        RECT 136.050 147.750 137.850 153.600 ;
        RECT 139.050 147.750 140.850 154.500 ;
        RECT 147.150 153.600 151.050 155.700 ;
        RECT 142.950 147.750 144.750 153.600 ;
        RECT 147.150 147.750 148.950 153.600 ;
        RECT 151.650 147.750 153.450 150.600 ;
        RECT 154.650 147.750 156.450 159.600 ;
        RECT 167.400 147.750 169.200 153.600 ;
        RECT 170.700 147.750 172.500 159.600 ;
        RECT 174.900 147.750 176.700 159.600 ;
        RECT 194.250 153.600 195.450 161.850 ;
        RECT 209.250 160.050 211.050 161.850 ;
        RECT 212.850 159.600 214.050 164.850 ;
        RECT 218.100 163.050 219.900 164.850 ;
        RECT 229.950 163.050 232.050 165.150 ;
        RECT 233.250 163.950 234.450 171.300 ;
        RECT 250.650 166.950 251.850 173.400 ;
        RECT 256.650 172.500 257.850 176.400 ;
        RECT 271.650 173.400 273.450 179.250 ;
        RECT 252.750 171.600 257.850 172.500 ;
        RECT 252.750 170.700 255.000 171.600 ;
        RECT 236.100 165.150 237.900 166.950 ;
        RECT 232.950 161.850 235.050 163.950 ;
        RECT 235.950 163.050 238.050 165.150 ;
        RECT 250.650 164.850 253.050 166.950 ;
        RECT 190.650 147.750 192.450 153.600 ;
        RECT 193.650 147.750 195.450 153.600 ;
        RECT 196.650 147.750 198.450 153.600 ;
        RECT 209.400 147.750 211.200 153.600 ;
        RECT 212.700 147.750 214.500 159.600 ;
        RECT 216.900 147.750 218.700 159.600 ;
        RECT 233.250 153.600 234.450 161.850 ;
        RECT 250.650 159.600 251.850 164.850 ;
        RECT 253.950 162.300 255.000 170.700 ;
        RECT 272.250 171.300 273.450 173.400 ;
        RECT 274.650 174.300 276.450 179.250 ;
        RECT 277.650 175.200 279.450 179.250 ;
        RECT 280.650 174.300 282.450 179.250 ;
        RECT 293.250 176.400 295.350 179.250 ;
        RECT 296.550 176.400 298.350 179.250 ;
        RECT 299.550 176.400 301.350 179.250 ;
        RECT 302.550 176.400 304.350 179.250 ;
        RECT 323.550 176.400 325.350 179.250 ;
        RECT 326.550 176.400 328.350 179.250 ;
        RECT 297.300 175.500 298.350 176.400 ;
        RECT 303.300 175.500 304.350 176.400 ;
        RECT 297.300 174.600 308.100 175.500 ;
        RECT 274.650 172.950 282.450 174.300 ;
        RECT 272.250 170.250 276.000 171.300 ;
        RECT 274.950 166.950 276.150 170.250 ;
        RECT 278.100 168.150 279.900 169.950 ;
        RECT 299.100 168.150 300.900 169.950 ;
        RECT 306.900 168.150 308.100 174.600 ;
        RECT 256.950 164.850 259.050 166.950 ;
        RECT 274.950 164.850 277.050 166.950 ;
        RECT 277.950 166.050 280.050 168.150 ;
        RECT 280.950 164.850 283.050 166.950 ;
        RECT 292.950 164.850 295.050 166.950 ;
        RECT 298.950 166.050 301.050 168.150 ;
        RECT 301.950 164.850 304.050 166.950 ;
        RECT 306.900 166.050 310.050 168.150 ;
        RECT 322.950 167.850 325.050 169.950 ;
        RECT 326.400 168.150 327.600 176.400 ;
        RECT 338.550 174.300 340.350 179.250 ;
        RECT 341.550 175.200 343.350 179.250 ;
        RECT 344.550 174.300 346.350 179.250 ;
        RECT 338.550 172.950 346.350 174.300 ;
        RECT 347.550 173.400 349.350 179.250 ;
        RECT 362.850 173.400 364.650 179.250 ;
        RECT 347.550 171.300 348.750 173.400 ;
        RECT 367.350 172.200 369.150 179.250 ;
        RECT 380.550 176.400 382.350 179.250 ;
        RECT 383.550 176.400 385.350 179.250 ;
        RECT 395.550 176.400 397.350 179.250 ;
        RECT 345.000 170.250 348.750 171.300 ;
        RECT 365.550 171.300 369.150 172.200 ;
        RECT 341.100 168.150 342.900 169.950 ;
        RECT 323.100 166.050 324.900 167.850 ;
        RECT 325.950 166.050 328.050 168.150 ;
        RECT 257.100 163.050 258.900 164.850 ;
        RECT 252.750 161.400 255.000 162.300 ;
        RECT 271.950 161.850 274.050 163.950 ;
        RECT 252.750 160.500 258.450 161.400 ;
        RECT 229.650 147.750 231.450 153.600 ;
        RECT 232.650 147.750 234.450 153.600 ;
        RECT 235.650 147.750 237.450 153.600 ;
        RECT 250.350 147.750 252.150 159.600 ;
        RECT 253.350 147.750 255.150 159.600 ;
        RECT 257.250 153.600 258.450 160.500 ;
        RECT 272.250 160.050 274.050 161.850 ;
        RECT 275.850 159.600 277.050 164.850 ;
        RECT 281.100 163.050 282.900 164.850 ;
        RECT 293.100 163.050 294.900 164.850 ;
        RECT 302.100 163.050 303.900 164.850 ;
        RECT 306.900 160.800 308.100 166.050 ;
        RECT 306.900 159.600 310.350 160.800 ;
        RECT 256.650 147.750 258.450 153.600 ;
        RECT 272.400 147.750 274.200 153.600 ;
        RECT 275.700 147.750 277.500 159.600 ;
        RECT 279.900 147.750 281.700 159.600 ;
        RECT 290.550 157.500 298.350 158.400 ;
        RECT 290.550 147.750 292.350 157.500 ;
        RECT 293.550 147.750 295.350 156.600 ;
        RECT 296.550 148.500 298.350 157.500 ;
        RECT 299.550 157.200 307.950 158.100 ;
        RECT 299.550 149.400 301.350 157.200 ;
        RECT 302.550 148.500 304.350 156.300 ;
        RECT 296.550 147.750 304.350 148.500 ;
        RECT 306.150 148.500 307.950 157.200 ;
        RECT 309.150 157.200 310.350 159.600 ;
        RECT 309.150 149.400 310.950 157.200 ;
        RECT 312.150 148.500 313.950 157.800 ;
        RECT 326.400 153.600 327.600 166.050 ;
        RECT 337.950 164.850 340.050 166.950 ;
        RECT 340.950 166.050 343.050 168.150 ;
        RECT 344.850 166.950 346.050 170.250 ;
        RECT 343.950 164.850 346.050 166.950 ;
        RECT 362.100 165.150 363.900 166.950 ;
        RECT 338.100 163.050 339.900 164.850 ;
        RECT 343.950 159.600 345.150 164.850 ;
        RECT 346.950 161.850 349.050 163.950 ;
        RECT 361.950 163.050 364.050 165.150 ;
        RECT 365.550 163.950 366.750 171.300 ;
        RECT 379.950 167.850 382.050 169.950 ;
        RECT 383.400 168.150 384.600 176.400 ;
        RECT 396.150 172.500 397.350 176.400 ;
        RECT 398.850 173.400 400.650 179.250 ;
        RECT 401.850 173.400 403.650 179.250 ;
        RECT 407.550 173.400 409.350 179.250 ;
        RECT 410.850 176.400 412.650 179.250 ;
        RECT 415.350 176.400 417.150 179.250 ;
        RECT 419.550 176.400 421.350 179.250 ;
        RECT 423.450 176.400 425.250 179.250 ;
        RECT 426.750 176.400 428.550 179.250 ;
        RECT 431.250 177.300 433.050 179.250 ;
        RECT 431.250 176.400 435.000 177.300 ;
        RECT 436.050 176.400 437.850 179.250 ;
        RECT 415.650 175.500 416.700 176.400 ;
        RECT 412.950 174.300 416.700 175.500 ;
        RECT 424.200 174.600 425.250 176.400 ;
        RECT 433.950 175.500 435.000 176.400 ;
        RECT 412.950 173.400 415.050 174.300 ;
        RECT 396.150 171.600 401.250 172.500 ;
        RECT 399.000 170.700 401.250 171.600 ;
        RECT 368.100 165.150 369.900 166.950 ;
        RECT 380.100 166.050 381.900 167.850 ;
        RECT 382.950 166.050 385.050 168.150 ;
        RECT 364.950 161.850 367.050 163.950 ;
        RECT 367.950 163.050 370.050 165.150 ;
        RECT 346.950 160.050 348.750 161.850 ;
        RECT 306.150 147.750 313.950 148.500 ;
        RECT 323.550 147.750 325.350 153.600 ;
        RECT 326.550 147.750 328.350 153.600 ;
        RECT 339.300 147.750 341.100 159.600 ;
        RECT 343.500 147.750 345.300 159.600 ;
        RECT 365.550 153.600 366.750 161.850 ;
        RECT 383.400 153.600 384.600 166.050 ;
        RECT 394.950 164.850 397.050 166.950 ;
        RECT 395.100 163.050 396.900 164.850 ;
        RECT 399.000 162.300 400.050 170.700 ;
        RECT 402.150 166.950 403.350 173.400 ;
        RECT 400.950 164.850 403.350 166.950 ;
        RECT 399.000 161.400 401.250 162.300 ;
        RECT 395.550 160.500 401.250 161.400 ;
        RECT 395.550 153.600 396.750 160.500 ;
        RECT 402.150 159.600 403.350 164.850 ;
        RECT 407.550 171.150 408.750 173.400 ;
        RECT 420.150 172.200 421.950 174.000 ;
        RECT 424.200 173.550 429.150 174.600 ;
        RECT 427.350 172.800 429.150 173.550 ;
        RECT 430.650 172.800 432.450 174.600 ;
        RECT 433.950 173.400 436.050 175.500 ;
        RECT 439.050 173.400 440.850 179.250 ;
        RECT 421.050 171.900 421.950 172.200 ;
        RECT 431.100 171.900 432.150 172.800 ;
        RECT 407.550 169.050 412.050 171.150 ;
        RECT 421.050 171.000 432.150 171.900 ;
        RECT 407.550 159.600 408.750 169.050 ;
        RECT 409.950 167.250 413.850 169.050 ;
        RECT 409.950 166.950 412.050 167.250 ;
        RECT 421.050 166.950 421.950 171.000 ;
        RECT 431.100 169.800 432.150 171.000 ;
        RECT 431.100 168.600 438.000 169.800 ;
        RECT 431.100 168.000 432.900 168.600 ;
        RECT 437.100 167.850 438.000 168.600 ;
        RECT 434.100 166.950 435.900 167.700 ;
        RECT 421.050 164.850 424.050 166.950 ;
        RECT 427.950 165.900 435.900 166.950 ;
        RECT 437.100 166.050 438.900 167.850 ;
        RECT 427.950 164.850 430.050 165.900 ;
        RECT 409.950 161.400 411.750 163.200 ;
        RECT 410.850 160.200 415.050 161.400 ;
        RECT 421.050 160.200 421.950 164.850 ;
        RECT 429.750 161.100 431.550 161.400 ;
        RECT 346.800 147.750 348.600 153.600 ;
        RECT 362.550 147.750 364.350 153.600 ;
        RECT 365.550 147.750 367.350 153.600 ;
        RECT 368.550 147.750 370.350 153.600 ;
        RECT 380.550 147.750 382.350 153.600 ;
        RECT 383.550 147.750 385.350 153.600 ;
        RECT 395.550 147.750 397.350 153.600 ;
        RECT 398.850 147.750 400.650 159.600 ;
        RECT 401.850 147.750 403.650 159.600 ;
        RECT 407.550 147.750 409.350 159.600 ;
        RECT 412.950 159.300 415.050 160.200 ;
        RECT 415.950 159.300 421.950 160.200 ;
        RECT 423.150 160.800 431.550 161.100 ;
        RECT 439.950 160.800 440.850 173.400 ;
        RECT 449.700 170.400 451.500 179.250 ;
        RECT 455.100 171.000 456.900 179.250 ;
        RECT 472.650 176.400 474.450 179.250 ;
        RECT 475.650 176.400 477.450 179.250 ;
        RECT 455.100 169.350 459.600 171.000 ;
        RECT 458.400 165.150 459.600 169.350 ;
        RECT 473.400 168.150 474.600 176.400 ;
        RECT 479.550 173.400 481.350 179.250 ;
        RECT 482.850 176.400 484.650 179.250 ;
        RECT 487.350 176.400 489.150 179.250 ;
        RECT 491.550 176.400 493.350 179.250 ;
        RECT 495.450 176.400 497.250 179.250 ;
        RECT 498.750 176.400 500.550 179.250 ;
        RECT 503.250 177.300 505.050 179.250 ;
        RECT 503.250 176.400 507.000 177.300 ;
        RECT 508.050 176.400 509.850 179.250 ;
        RECT 487.650 175.500 488.700 176.400 ;
        RECT 484.950 174.300 488.700 175.500 ;
        RECT 496.200 174.600 497.250 176.400 ;
        RECT 505.950 175.500 507.000 176.400 ;
        RECT 484.950 173.400 487.050 174.300 ;
        RECT 479.550 171.150 480.750 173.400 ;
        RECT 492.150 172.200 493.950 174.000 ;
        RECT 496.200 173.550 501.150 174.600 ;
        RECT 499.350 172.800 501.150 173.550 ;
        RECT 502.650 172.800 504.450 174.600 ;
        RECT 505.950 173.400 508.050 175.500 ;
        RECT 511.050 173.400 512.850 179.250 ;
        RECT 523.650 176.400 525.450 179.250 ;
        RECT 526.650 176.400 528.450 179.250 ;
        RECT 493.050 171.900 493.950 172.200 ;
        RECT 503.100 171.900 504.150 172.800 ;
        RECT 472.950 166.050 475.050 168.150 ;
        RECT 475.950 167.850 478.050 169.950 ;
        RECT 479.550 169.050 484.050 171.150 ;
        RECT 493.050 171.000 504.150 171.900 ;
        RECT 476.100 166.050 477.900 167.850 ;
        RECT 448.950 161.850 451.050 163.950 ;
        RECT 454.950 161.850 457.050 163.950 ;
        RECT 457.950 163.050 460.050 165.150 ;
        RECT 423.150 160.200 440.850 160.800 ;
        RECT 415.950 158.400 416.850 159.300 ;
        RECT 414.150 156.600 416.850 158.400 ;
        RECT 417.750 158.100 419.550 158.400 ;
        RECT 423.150 158.100 424.050 160.200 ;
        RECT 429.750 159.600 440.850 160.200 ;
        RECT 449.100 160.050 450.900 161.850 ;
        RECT 417.750 157.200 424.050 158.100 ;
        RECT 424.950 158.700 426.750 159.300 ;
        RECT 424.950 157.500 432.450 158.700 ;
        RECT 417.750 156.600 419.550 157.200 ;
        RECT 431.250 156.600 432.450 157.500 ;
        RECT 412.950 153.600 416.850 155.700 ;
        RECT 421.950 154.500 428.850 156.300 ;
        RECT 431.250 154.500 436.050 156.600 ;
        RECT 410.550 147.750 412.350 150.600 ;
        RECT 415.050 147.750 416.850 153.600 ;
        RECT 419.250 147.750 421.050 153.600 ;
        RECT 423.150 147.750 424.950 154.500 ;
        RECT 431.250 153.600 432.450 154.500 ;
        RECT 426.150 147.750 427.950 153.600 ;
        RECT 430.950 147.750 432.750 153.600 ;
        RECT 436.050 147.750 437.850 153.600 ;
        RECT 439.050 147.750 440.850 159.600 ;
        RECT 451.950 158.850 454.050 160.950 ;
        RECT 455.250 160.050 457.050 161.850 ;
        RECT 452.100 157.050 453.900 158.850 ;
        RECT 458.700 154.800 459.750 163.050 ;
        RECT 452.700 153.900 459.750 154.800 ;
        RECT 452.700 153.600 454.350 153.900 ;
        RECT 449.550 147.750 451.350 153.600 ;
        RECT 452.550 147.750 454.350 153.600 ;
        RECT 458.550 153.600 459.750 153.900 ;
        RECT 473.400 153.600 474.600 166.050 ;
        RECT 479.550 159.600 480.750 169.050 ;
        RECT 481.950 167.250 485.850 169.050 ;
        RECT 481.950 166.950 484.050 167.250 ;
        RECT 493.050 166.950 493.950 171.000 ;
        RECT 503.100 169.800 504.150 171.000 ;
        RECT 503.100 168.600 510.000 169.800 ;
        RECT 503.100 168.000 504.900 168.600 ;
        RECT 509.100 167.850 510.000 168.600 ;
        RECT 506.100 166.950 507.900 167.700 ;
        RECT 493.050 164.850 496.050 166.950 ;
        RECT 499.950 165.900 507.900 166.950 ;
        RECT 509.100 166.050 510.900 167.850 ;
        RECT 499.950 164.850 502.050 165.900 ;
        RECT 481.950 161.400 483.750 163.200 ;
        RECT 482.850 160.200 487.050 161.400 ;
        RECT 493.050 160.200 493.950 164.850 ;
        RECT 501.750 161.100 503.550 161.400 ;
        RECT 455.550 147.750 457.350 153.000 ;
        RECT 458.550 147.750 460.350 153.600 ;
        RECT 472.650 147.750 474.450 153.600 ;
        RECT 475.650 147.750 477.450 153.600 ;
        RECT 479.550 147.750 481.350 159.600 ;
        RECT 484.950 159.300 487.050 160.200 ;
        RECT 487.950 159.300 493.950 160.200 ;
        RECT 495.150 160.800 503.550 161.100 ;
        RECT 511.950 160.800 512.850 173.400 ;
        RECT 524.400 168.150 525.600 176.400 ;
        RECT 536.550 174.300 538.350 179.250 ;
        RECT 539.550 175.200 541.350 179.250 ;
        RECT 542.550 174.300 544.350 179.250 ;
        RECT 536.550 172.950 544.350 174.300 ;
        RECT 545.550 173.400 547.350 179.250 ;
        RECT 557.550 176.400 559.350 179.250 ;
        RECT 560.550 176.400 562.350 179.250 ;
        RECT 545.550 171.300 546.750 173.400 ;
        RECT 543.000 170.250 546.750 171.300 ;
        RECT 523.950 166.050 526.050 168.150 ;
        RECT 526.950 167.850 529.050 169.950 ;
        RECT 539.100 168.150 540.900 169.950 ;
        RECT 527.100 166.050 528.900 167.850 ;
        RECT 495.150 160.200 512.850 160.800 ;
        RECT 487.950 158.400 488.850 159.300 ;
        RECT 486.150 156.600 488.850 158.400 ;
        RECT 489.750 158.100 491.550 158.400 ;
        RECT 495.150 158.100 496.050 160.200 ;
        RECT 501.750 159.600 512.850 160.200 ;
        RECT 489.750 157.200 496.050 158.100 ;
        RECT 496.950 158.700 498.750 159.300 ;
        RECT 496.950 157.500 504.450 158.700 ;
        RECT 489.750 156.600 491.550 157.200 ;
        RECT 503.250 156.600 504.450 157.500 ;
        RECT 484.950 153.600 488.850 155.700 ;
        RECT 493.950 154.500 500.850 156.300 ;
        RECT 503.250 154.500 508.050 156.600 ;
        RECT 482.550 147.750 484.350 150.600 ;
        RECT 487.050 147.750 488.850 153.600 ;
        RECT 491.250 147.750 493.050 153.600 ;
        RECT 495.150 147.750 496.950 154.500 ;
        RECT 503.250 153.600 504.450 154.500 ;
        RECT 498.150 147.750 499.950 153.600 ;
        RECT 502.950 147.750 504.750 153.600 ;
        RECT 508.050 147.750 509.850 153.600 ;
        RECT 511.050 147.750 512.850 159.600 ;
        RECT 524.400 153.600 525.600 166.050 ;
        RECT 535.950 164.850 538.050 166.950 ;
        RECT 538.950 166.050 541.050 168.150 ;
        RECT 542.850 166.950 544.050 170.250 ;
        RECT 556.950 167.850 559.050 169.950 ;
        RECT 560.400 168.150 561.600 176.400 ;
        RECT 580.800 173.400 582.600 179.250 ;
        RECT 585.000 173.400 586.800 179.250 ;
        RECT 589.200 173.400 591.000 179.250 ;
        RECT 594.150 173.400 595.950 179.250 ;
        RECT 597.150 176.400 598.950 179.250 ;
        RECT 601.950 177.300 603.750 179.250 ;
        RECT 600.000 176.400 603.750 177.300 ;
        RECT 606.450 176.400 608.250 179.250 ;
        RECT 609.750 176.400 611.550 179.250 ;
        RECT 613.650 176.400 615.450 179.250 ;
        RECT 617.850 176.400 619.650 179.250 ;
        RECT 622.350 176.400 624.150 179.250 ;
        RECT 600.000 175.500 601.050 176.400 ;
        RECT 598.950 173.400 601.050 175.500 ;
        RECT 609.750 174.600 610.800 176.400 ;
        RECT 581.250 168.150 583.050 169.950 ;
        RECT 541.950 164.850 544.050 166.950 ;
        RECT 557.100 166.050 558.900 167.850 ;
        RECT 559.950 166.050 562.050 168.150 ;
        RECT 536.100 163.050 537.900 164.850 ;
        RECT 541.950 159.600 543.150 164.850 ;
        RECT 544.950 161.850 547.050 163.950 ;
        RECT 544.950 160.050 546.750 161.850 ;
        RECT 523.650 147.750 525.450 153.600 ;
        RECT 526.650 147.750 528.450 153.600 ;
        RECT 537.300 147.750 539.100 159.600 ;
        RECT 541.500 147.750 543.300 159.600 ;
        RECT 560.400 153.600 561.600 166.050 ;
        RECT 577.950 164.850 580.050 166.950 ;
        RECT 580.950 166.050 583.050 168.150 ;
        RECT 585.000 166.950 586.050 173.400 ;
        RECT 583.950 164.850 586.050 166.950 ;
        RECT 586.950 168.150 588.750 169.950 ;
        RECT 586.950 166.050 589.050 168.150 ;
        RECT 589.950 164.850 592.050 166.950 ;
        RECT 578.100 163.050 579.900 164.850 ;
        RECT 583.950 161.400 584.850 164.850 ;
        RECT 589.950 163.050 591.750 164.850 ;
        RECT 580.800 160.500 584.850 161.400 ;
        RECT 594.150 160.800 595.050 173.400 ;
        RECT 602.550 172.800 604.350 174.600 ;
        RECT 605.850 173.550 610.800 174.600 ;
        RECT 618.300 175.500 619.350 176.400 ;
        RECT 618.300 174.300 622.050 175.500 ;
        RECT 605.850 172.800 607.650 173.550 ;
        RECT 602.850 171.900 603.900 172.800 ;
        RECT 613.050 172.200 614.850 174.000 ;
        RECT 619.950 173.400 622.050 174.300 ;
        RECT 625.650 173.400 627.450 179.250 ;
        RECT 640.650 173.400 642.450 179.250 ;
        RECT 613.050 171.900 613.950 172.200 ;
        RECT 602.850 171.000 613.950 171.900 ;
        RECT 626.250 171.150 627.450 173.400 ;
        RECT 602.850 169.800 603.900 171.000 ;
        RECT 597.000 168.600 603.900 169.800 ;
        RECT 597.000 167.850 597.900 168.600 ;
        RECT 602.100 168.000 603.900 168.600 ;
        RECT 596.100 166.050 597.900 167.850 ;
        RECT 599.100 166.950 600.900 167.700 ;
        RECT 613.050 166.950 613.950 171.000 ;
        RECT 622.950 169.050 627.450 171.150 ;
        RECT 641.250 171.300 642.450 173.400 ;
        RECT 643.650 174.300 645.450 179.250 ;
        RECT 646.650 175.200 648.450 179.250 ;
        RECT 649.650 174.300 651.450 179.250 ;
        RECT 643.650 172.950 651.450 174.300 ;
        RECT 654.150 173.400 655.950 179.250 ;
        RECT 657.150 176.400 658.950 179.250 ;
        RECT 661.950 177.300 663.750 179.250 ;
        RECT 660.000 176.400 663.750 177.300 ;
        RECT 666.450 176.400 668.250 179.250 ;
        RECT 669.750 176.400 671.550 179.250 ;
        RECT 673.650 176.400 675.450 179.250 ;
        RECT 677.850 176.400 679.650 179.250 ;
        RECT 682.350 176.400 684.150 179.250 ;
        RECT 660.000 175.500 661.050 176.400 ;
        RECT 658.950 173.400 661.050 175.500 ;
        RECT 669.750 174.600 670.800 176.400 ;
        RECT 641.250 170.250 645.000 171.300 ;
        RECT 621.150 167.250 625.050 169.050 ;
        RECT 622.950 166.950 625.050 167.250 ;
        RECT 599.100 165.900 607.050 166.950 ;
        RECT 604.950 164.850 607.050 165.900 ;
        RECT 610.950 164.850 613.950 166.950 ;
        RECT 603.450 161.100 605.250 161.400 ;
        RECT 603.450 160.800 611.850 161.100 ;
        RECT 580.800 159.600 582.600 160.500 ;
        RECT 594.150 160.200 611.850 160.800 ;
        RECT 594.150 159.600 605.250 160.200 ;
        RECT 544.800 147.750 546.600 153.600 ;
        RECT 557.550 147.750 559.350 153.600 ;
        RECT 560.550 147.750 562.350 153.600 ;
        RECT 577.650 148.500 579.450 159.600 ;
        RECT 580.650 149.400 582.450 159.600 ;
        RECT 583.650 158.400 591.450 159.300 ;
        RECT 583.650 148.500 585.450 158.400 ;
        RECT 577.650 147.750 585.450 148.500 ;
        RECT 586.650 147.750 588.450 157.500 ;
        RECT 589.650 147.750 591.450 158.400 ;
        RECT 594.150 147.750 595.950 159.600 ;
        RECT 608.250 158.700 610.050 159.300 ;
        RECT 602.550 157.500 610.050 158.700 ;
        RECT 610.950 158.100 611.850 160.200 ;
        RECT 613.050 160.200 613.950 164.850 ;
        RECT 623.250 161.400 625.050 163.200 ;
        RECT 619.950 160.200 624.150 161.400 ;
        RECT 613.050 159.300 619.050 160.200 ;
        RECT 619.950 159.300 622.050 160.200 ;
        RECT 626.250 159.600 627.450 169.050 ;
        RECT 643.950 166.950 645.150 170.250 ;
        RECT 647.100 168.150 648.900 169.950 ;
        RECT 643.950 164.850 646.050 166.950 ;
        RECT 646.950 166.050 649.050 168.150 ;
        RECT 649.950 164.850 652.050 166.950 ;
        RECT 640.950 161.850 643.050 163.950 ;
        RECT 641.250 160.050 643.050 161.850 ;
        RECT 644.850 159.600 646.050 164.850 ;
        RECT 650.100 163.050 651.900 164.850 ;
        RECT 654.150 160.800 655.050 173.400 ;
        RECT 662.550 172.800 664.350 174.600 ;
        RECT 665.850 173.550 670.800 174.600 ;
        RECT 678.300 175.500 679.350 176.400 ;
        RECT 678.300 174.300 682.050 175.500 ;
        RECT 665.850 172.800 667.650 173.550 ;
        RECT 662.850 171.900 663.900 172.800 ;
        RECT 673.050 172.200 674.850 174.000 ;
        RECT 679.950 173.400 682.050 174.300 ;
        RECT 685.650 173.400 687.450 179.250 ;
        RECT 703.800 173.400 705.600 179.250 ;
        RECT 708.000 173.400 709.800 179.250 ;
        RECT 712.200 173.400 714.000 179.250 ;
        RECT 724.650 176.400 726.450 179.250 ;
        RECT 727.650 176.400 729.450 179.250 ;
        RECT 673.050 171.900 673.950 172.200 ;
        RECT 662.850 171.000 673.950 171.900 ;
        RECT 686.250 171.150 687.450 173.400 ;
        RECT 662.850 169.800 663.900 171.000 ;
        RECT 657.000 168.600 663.900 169.800 ;
        RECT 657.000 167.850 657.900 168.600 ;
        RECT 662.100 168.000 663.900 168.600 ;
        RECT 656.100 166.050 657.900 167.850 ;
        RECT 659.100 166.950 660.900 167.700 ;
        RECT 673.050 166.950 673.950 171.000 ;
        RECT 682.950 169.050 687.450 171.150 ;
        RECT 681.150 167.250 685.050 169.050 ;
        RECT 682.950 166.950 685.050 167.250 ;
        RECT 659.100 165.900 667.050 166.950 ;
        RECT 664.950 164.850 667.050 165.900 ;
        RECT 670.950 164.850 673.950 166.950 ;
        RECT 663.450 161.100 665.250 161.400 ;
        RECT 663.450 160.800 671.850 161.100 ;
        RECT 654.150 160.200 671.850 160.800 ;
        RECT 654.150 159.600 665.250 160.200 ;
        RECT 618.150 158.400 619.050 159.300 ;
        RECT 615.450 158.100 617.250 158.400 ;
        RECT 602.550 156.600 603.750 157.500 ;
        RECT 610.950 157.200 617.250 158.100 ;
        RECT 615.450 156.600 617.250 157.200 ;
        RECT 618.150 156.600 620.850 158.400 ;
        RECT 598.950 154.500 603.750 156.600 ;
        RECT 606.150 154.500 613.050 156.300 ;
        RECT 602.550 153.600 603.750 154.500 ;
        RECT 597.150 147.750 598.950 153.600 ;
        RECT 602.250 147.750 604.050 153.600 ;
        RECT 607.050 147.750 608.850 153.600 ;
        RECT 610.050 147.750 611.850 154.500 ;
        RECT 618.150 153.600 622.050 155.700 ;
        RECT 613.950 147.750 615.750 153.600 ;
        RECT 618.150 147.750 619.950 153.600 ;
        RECT 622.650 147.750 624.450 150.600 ;
        RECT 625.650 147.750 627.450 159.600 ;
        RECT 641.400 147.750 643.200 153.600 ;
        RECT 644.700 147.750 646.500 159.600 ;
        RECT 648.900 147.750 650.700 159.600 ;
        RECT 654.150 147.750 655.950 159.600 ;
        RECT 668.250 158.700 670.050 159.300 ;
        RECT 662.550 157.500 670.050 158.700 ;
        RECT 670.950 158.100 671.850 160.200 ;
        RECT 673.050 160.200 673.950 164.850 ;
        RECT 683.250 161.400 685.050 163.200 ;
        RECT 679.950 160.200 684.150 161.400 ;
        RECT 673.050 159.300 679.050 160.200 ;
        RECT 679.950 159.300 682.050 160.200 ;
        RECT 686.250 159.600 687.450 169.050 ;
        RECT 704.250 168.150 706.050 169.950 ;
        RECT 700.950 164.850 703.050 166.950 ;
        RECT 703.950 166.050 706.050 168.150 ;
        RECT 708.000 166.950 709.050 173.400 ;
        RECT 706.950 164.850 709.050 166.950 ;
        RECT 709.950 168.150 711.750 169.950 ;
        RECT 725.400 168.150 726.600 176.400 ;
        RECT 731.550 173.400 733.350 179.250 ;
        RECT 734.850 176.400 736.650 179.250 ;
        RECT 739.350 176.400 741.150 179.250 ;
        RECT 743.550 176.400 745.350 179.250 ;
        RECT 747.450 176.400 749.250 179.250 ;
        RECT 750.750 176.400 752.550 179.250 ;
        RECT 755.250 177.300 757.050 179.250 ;
        RECT 755.250 176.400 759.000 177.300 ;
        RECT 760.050 176.400 761.850 179.250 ;
        RECT 739.650 175.500 740.700 176.400 ;
        RECT 736.950 174.300 740.700 175.500 ;
        RECT 748.200 174.600 749.250 176.400 ;
        RECT 757.950 175.500 759.000 176.400 ;
        RECT 736.950 173.400 739.050 174.300 ;
        RECT 731.550 171.150 732.750 173.400 ;
        RECT 744.150 172.200 745.950 174.000 ;
        RECT 748.200 173.550 753.150 174.600 ;
        RECT 751.350 172.800 753.150 173.550 ;
        RECT 754.650 172.800 756.450 174.600 ;
        RECT 757.950 173.400 760.050 175.500 ;
        RECT 763.050 173.400 764.850 179.250 ;
        RECT 745.050 171.900 745.950 172.200 ;
        RECT 755.100 171.900 756.150 172.800 ;
        RECT 709.950 166.050 712.050 168.150 ;
        RECT 712.950 164.850 715.050 166.950 ;
        RECT 724.950 166.050 727.050 168.150 ;
        RECT 727.950 167.850 730.050 169.950 ;
        RECT 731.550 169.050 736.050 171.150 ;
        RECT 745.050 171.000 756.150 171.900 ;
        RECT 728.100 166.050 729.900 167.850 ;
        RECT 701.100 163.050 702.900 164.850 ;
        RECT 706.950 161.400 707.850 164.850 ;
        RECT 712.950 163.050 714.750 164.850 ;
        RECT 703.800 160.500 707.850 161.400 ;
        RECT 703.800 159.600 705.600 160.500 ;
        RECT 678.150 158.400 679.050 159.300 ;
        RECT 675.450 158.100 677.250 158.400 ;
        RECT 662.550 156.600 663.750 157.500 ;
        RECT 670.950 157.200 677.250 158.100 ;
        RECT 675.450 156.600 677.250 157.200 ;
        RECT 678.150 156.600 680.850 158.400 ;
        RECT 658.950 154.500 663.750 156.600 ;
        RECT 666.150 154.500 673.050 156.300 ;
        RECT 662.550 153.600 663.750 154.500 ;
        RECT 657.150 147.750 658.950 153.600 ;
        RECT 662.250 147.750 664.050 153.600 ;
        RECT 667.050 147.750 668.850 153.600 ;
        RECT 670.050 147.750 671.850 154.500 ;
        RECT 678.150 153.600 682.050 155.700 ;
        RECT 673.950 147.750 675.750 153.600 ;
        RECT 678.150 147.750 679.950 153.600 ;
        RECT 682.650 147.750 684.450 150.600 ;
        RECT 685.650 147.750 687.450 159.600 ;
        RECT 700.650 148.500 702.450 159.600 ;
        RECT 703.650 149.400 705.450 159.600 ;
        RECT 706.650 158.400 714.450 159.300 ;
        RECT 706.650 148.500 708.450 158.400 ;
        RECT 700.650 147.750 708.450 148.500 ;
        RECT 709.650 147.750 711.450 157.500 ;
        RECT 712.650 147.750 714.450 158.400 ;
        RECT 725.400 153.600 726.600 166.050 ;
        RECT 731.550 159.600 732.750 169.050 ;
        RECT 733.950 167.250 737.850 169.050 ;
        RECT 733.950 166.950 736.050 167.250 ;
        RECT 745.050 166.950 745.950 171.000 ;
        RECT 755.100 169.800 756.150 171.000 ;
        RECT 755.100 168.600 762.000 169.800 ;
        RECT 755.100 168.000 756.900 168.600 ;
        RECT 761.100 167.850 762.000 168.600 ;
        RECT 758.100 166.950 759.900 167.700 ;
        RECT 745.050 164.850 748.050 166.950 ;
        RECT 751.950 165.900 759.900 166.950 ;
        RECT 761.100 166.050 762.900 167.850 ;
        RECT 751.950 164.850 754.050 165.900 ;
        RECT 733.950 161.400 735.750 163.200 ;
        RECT 734.850 160.200 739.050 161.400 ;
        RECT 745.050 160.200 745.950 164.850 ;
        RECT 753.750 161.100 755.550 161.400 ;
        RECT 724.650 147.750 726.450 153.600 ;
        RECT 727.650 147.750 729.450 153.600 ;
        RECT 731.550 147.750 733.350 159.600 ;
        RECT 736.950 159.300 739.050 160.200 ;
        RECT 739.950 159.300 745.950 160.200 ;
        RECT 747.150 160.800 755.550 161.100 ;
        RECT 763.950 160.800 764.850 173.400 ;
        RECT 773.550 174.000 775.350 179.250 ;
        RECT 776.550 174.900 778.350 179.250 ;
        RECT 779.550 178.500 787.350 179.250 ;
        RECT 779.550 174.000 781.350 178.500 ;
        RECT 773.550 173.100 781.350 174.000 ;
        RECT 782.550 173.400 784.350 177.600 ;
        RECT 785.550 173.400 787.350 178.500 ;
        RECT 799.650 173.400 801.450 179.250 ;
        RECT 782.850 171.900 783.750 173.400 ;
        RECT 779.400 170.850 783.750 171.900 ;
        RECT 784.950 171.450 787.050 172.050 ;
        RECT 776.100 168.150 777.900 169.950 ;
        RECT 772.950 164.850 775.050 166.950 ;
        RECT 775.950 166.050 778.050 168.150 ;
        RECT 779.400 166.950 780.600 170.850 ;
        RECT 784.950 170.550 789.450 171.450 ;
        RECT 784.950 169.950 787.050 170.550 ;
        RECT 781.500 168.150 783.300 169.950 ;
        RECT 788.550 169.050 789.450 170.550 ;
        RECT 800.250 171.300 801.450 173.400 ;
        RECT 802.650 174.300 804.450 179.250 ;
        RECT 805.650 175.200 807.450 179.250 ;
        RECT 808.650 174.300 810.450 179.250 ;
        RECT 802.650 172.950 810.450 174.300 ;
        RECT 818.550 174.000 820.350 179.250 ;
        RECT 821.550 174.900 823.350 179.250 ;
        RECT 824.550 178.500 832.350 179.250 ;
        RECT 824.550 174.000 826.350 178.500 ;
        RECT 818.550 173.100 826.350 174.000 ;
        RECT 827.550 173.400 829.350 177.600 ;
        RECT 830.550 173.400 832.350 178.500 ;
        RECT 844.650 176.400 846.450 179.250 ;
        RECT 847.650 176.400 849.450 179.250 ;
        RECT 827.850 171.900 828.750 173.400 ;
        RECT 800.250 170.250 804.000 171.300 ;
        RECT 824.400 170.850 828.750 171.900 ;
        RECT 778.950 164.850 781.050 166.950 ;
        RECT 781.950 166.050 784.050 168.150 ;
        RECT 787.950 166.950 790.050 169.050 ;
        RECT 802.950 166.950 804.150 170.250 ;
        RECT 806.100 168.150 807.900 169.950 ;
        RECT 821.100 168.150 822.900 169.950 ;
        RECT 784.950 164.850 787.050 166.950 ;
        RECT 802.950 164.850 805.050 166.950 ;
        RECT 805.950 166.050 808.050 168.150 ;
        RECT 808.950 164.850 811.050 166.950 ;
        RECT 817.950 164.850 820.050 166.950 ;
        RECT 820.950 166.050 823.050 168.150 ;
        RECT 824.400 166.950 825.600 170.850 ;
        RECT 826.500 168.150 828.300 169.950 ;
        RECT 845.400 168.150 846.600 176.400 ;
        RECT 851.550 173.400 853.350 179.250 ;
        RECT 854.850 176.400 856.650 179.250 ;
        RECT 859.350 176.400 861.150 179.250 ;
        RECT 863.550 176.400 865.350 179.250 ;
        RECT 867.450 176.400 869.250 179.250 ;
        RECT 870.750 176.400 872.550 179.250 ;
        RECT 875.250 177.300 877.050 179.250 ;
        RECT 875.250 176.400 879.000 177.300 ;
        RECT 880.050 176.400 881.850 179.250 ;
        RECT 859.650 175.500 860.700 176.400 ;
        RECT 856.950 174.300 860.700 175.500 ;
        RECT 868.200 174.600 869.250 176.400 ;
        RECT 877.950 175.500 879.000 176.400 ;
        RECT 856.950 173.400 859.050 174.300 ;
        RECT 851.550 171.150 852.750 173.400 ;
        RECT 864.150 172.200 865.950 174.000 ;
        RECT 868.200 173.550 873.150 174.600 ;
        RECT 871.350 172.800 873.150 173.550 ;
        RECT 874.650 172.800 876.450 174.600 ;
        RECT 877.950 173.400 880.050 175.500 ;
        RECT 883.050 173.400 884.850 179.250 ;
        RECT 865.050 171.900 865.950 172.200 ;
        RECT 875.100 171.900 876.150 172.800 ;
        RECT 823.950 164.850 826.050 166.950 ;
        RECT 826.950 166.050 829.050 168.150 ;
        RECT 829.950 164.850 832.050 166.950 ;
        RECT 844.950 166.050 847.050 168.150 ;
        RECT 847.950 167.850 850.050 169.950 ;
        RECT 851.550 169.050 856.050 171.150 ;
        RECT 865.050 171.000 876.150 171.900 ;
        RECT 848.100 166.050 849.900 167.850 ;
        RECT 773.100 163.050 774.900 164.850 ;
        RECT 747.150 160.200 764.850 160.800 ;
        RECT 739.950 158.400 740.850 159.300 ;
        RECT 738.150 156.600 740.850 158.400 ;
        RECT 741.750 158.100 743.550 158.400 ;
        RECT 747.150 158.100 748.050 160.200 ;
        RECT 753.750 159.600 764.850 160.200 ;
        RECT 779.550 159.600 780.750 164.850 ;
        RECT 784.950 163.050 786.750 164.850 ;
        RECT 799.950 161.850 802.050 163.950 ;
        RECT 800.250 160.050 802.050 161.850 ;
        RECT 803.850 159.600 805.050 164.850 ;
        RECT 809.100 163.050 810.900 164.850 ;
        RECT 818.100 163.050 819.900 164.850 ;
        RECT 824.550 159.600 825.750 164.850 ;
        RECT 829.950 163.050 831.750 164.850 ;
        RECT 741.750 157.200 748.050 158.100 ;
        RECT 748.950 158.700 750.750 159.300 ;
        RECT 748.950 157.500 756.450 158.700 ;
        RECT 741.750 156.600 743.550 157.200 ;
        RECT 755.250 156.600 756.450 157.500 ;
        RECT 736.950 153.600 740.850 155.700 ;
        RECT 745.950 154.500 752.850 156.300 ;
        RECT 755.250 154.500 760.050 156.600 ;
        RECT 734.550 147.750 736.350 150.600 ;
        RECT 739.050 147.750 740.850 153.600 ;
        RECT 743.250 147.750 745.050 153.600 ;
        RECT 747.150 147.750 748.950 154.500 ;
        RECT 755.250 153.600 756.450 154.500 ;
        RECT 750.150 147.750 751.950 153.600 ;
        RECT 754.950 147.750 756.750 153.600 ;
        RECT 760.050 147.750 761.850 153.600 ;
        RECT 763.050 147.750 764.850 159.600 ;
        RECT 773.550 147.750 775.350 159.600 ;
        RECT 778.050 147.750 781.350 159.600 ;
        RECT 784.050 147.750 785.850 159.600 ;
        RECT 800.400 147.750 802.200 153.600 ;
        RECT 803.700 147.750 805.500 159.600 ;
        RECT 807.900 147.750 809.700 159.600 ;
        RECT 818.550 147.750 820.350 159.600 ;
        RECT 823.050 147.750 826.350 159.600 ;
        RECT 829.050 147.750 830.850 159.600 ;
        RECT 845.400 153.600 846.600 166.050 ;
        RECT 851.550 159.600 852.750 169.050 ;
        RECT 853.950 167.250 857.850 169.050 ;
        RECT 853.950 166.950 856.050 167.250 ;
        RECT 865.050 166.950 865.950 171.000 ;
        RECT 875.100 169.800 876.150 171.000 ;
        RECT 875.100 168.600 882.000 169.800 ;
        RECT 875.100 168.000 876.900 168.600 ;
        RECT 881.100 167.850 882.000 168.600 ;
        RECT 878.100 166.950 879.900 167.700 ;
        RECT 865.050 164.850 868.050 166.950 ;
        RECT 871.950 165.900 879.900 166.950 ;
        RECT 881.100 166.050 882.900 167.850 ;
        RECT 871.950 164.850 874.050 165.900 ;
        RECT 853.950 161.400 855.750 163.200 ;
        RECT 854.850 160.200 859.050 161.400 ;
        RECT 865.050 160.200 865.950 164.850 ;
        RECT 873.750 161.100 875.550 161.400 ;
        RECT 844.650 147.750 846.450 153.600 ;
        RECT 847.650 147.750 849.450 153.600 ;
        RECT 851.550 147.750 853.350 159.600 ;
        RECT 856.950 159.300 859.050 160.200 ;
        RECT 859.950 159.300 865.950 160.200 ;
        RECT 867.150 160.800 875.550 161.100 ;
        RECT 883.950 160.800 884.850 173.400 ;
        RECT 867.150 160.200 884.850 160.800 ;
        RECT 859.950 158.400 860.850 159.300 ;
        RECT 858.150 156.600 860.850 158.400 ;
        RECT 861.750 158.100 863.550 158.400 ;
        RECT 867.150 158.100 868.050 160.200 ;
        RECT 873.750 159.600 884.850 160.200 ;
        RECT 861.750 157.200 868.050 158.100 ;
        RECT 868.950 158.700 870.750 159.300 ;
        RECT 868.950 157.500 876.450 158.700 ;
        RECT 861.750 156.600 863.550 157.200 ;
        RECT 875.250 156.600 876.450 157.500 ;
        RECT 856.950 153.600 860.850 155.700 ;
        RECT 865.950 154.500 872.850 156.300 ;
        RECT 875.250 154.500 880.050 156.600 ;
        RECT 854.550 147.750 856.350 150.600 ;
        RECT 859.050 147.750 860.850 153.600 ;
        RECT 863.250 147.750 865.050 153.600 ;
        RECT 867.150 147.750 868.950 154.500 ;
        RECT 875.250 153.600 876.450 154.500 ;
        RECT 870.150 147.750 871.950 153.600 ;
        RECT 874.950 147.750 876.750 153.600 ;
        RECT 880.050 147.750 881.850 153.600 ;
        RECT 883.050 147.750 884.850 159.600 ;
        RECT 2.550 131.400 4.350 143.250 ;
        RECT 5.550 140.400 7.350 143.250 ;
        RECT 10.050 137.400 11.850 143.250 ;
        RECT 14.250 137.400 16.050 143.250 ;
        RECT 7.950 135.300 11.850 137.400 ;
        RECT 18.150 136.500 19.950 143.250 ;
        RECT 21.150 137.400 22.950 143.250 ;
        RECT 25.950 137.400 27.750 143.250 ;
        RECT 31.050 137.400 32.850 143.250 ;
        RECT 26.250 136.500 27.450 137.400 ;
        RECT 16.950 134.700 23.850 136.500 ;
        RECT 26.250 134.400 31.050 136.500 ;
        RECT 9.150 132.600 11.850 134.400 ;
        RECT 12.750 133.800 14.550 134.400 ;
        RECT 12.750 132.900 19.050 133.800 ;
        RECT 26.250 133.500 27.450 134.400 ;
        RECT 12.750 132.600 14.550 132.900 ;
        RECT 10.950 131.700 11.850 132.600 ;
        RECT 2.550 121.950 3.750 131.400 ;
        RECT 7.950 130.800 10.050 131.700 ;
        RECT 10.950 130.800 16.950 131.700 ;
        RECT 5.850 129.600 10.050 130.800 ;
        RECT 4.950 127.800 6.750 129.600 ;
        RECT 16.050 126.150 16.950 130.800 ;
        RECT 18.150 130.800 19.050 132.900 ;
        RECT 19.950 132.300 27.450 133.500 ;
        RECT 19.950 131.700 21.750 132.300 ;
        RECT 34.050 131.400 35.850 143.250 ;
        RECT 48.150 132.900 49.950 143.250 ;
        RECT 24.750 130.800 35.850 131.400 ;
        RECT 18.150 130.200 35.850 130.800 ;
        RECT 18.150 129.900 26.550 130.200 ;
        RECT 24.750 129.600 26.550 129.900 ;
        RECT 16.050 124.050 19.050 126.150 ;
        RECT 22.950 125.100 25.050 126.150 ;
        RECT 22.950 124.050 30.900 125.100 ;
        RECT 4.950 123.750 7.050 124.050 ;
        RECT 4.950 121.950 8.850 123.750 ;
        RECT 2.550 119.850 7.050 121.950 ;
        RECT 16.050 120.000 16.950 124.050 ;
        RECT 29.100 123.300 30.900 124.050 ;
        RECT 32.100 123.150 33.900 124.950 ;
        RECT 26.100 122.400 27.900 123.000 ;
        RECT 32.100 122.400 33.000 123.150 ;
        RECT 26.100 121.200 33.000 122.400 ;
        RECT 26.100 120.000 27.150 121.200 ;
        RECT 2.550 117.600 3.750 119.850 ;
        RECT 16.050 119.100 27.150 120.000 ;
        RECT 16.050 118.800 16.950 119.100 ;
        RECT 2.550 111.750 4.350 117.600 ;
        RECT 7.950 116.700 10.050 117.600 ;
        RECT 15.150 117.000 16.950 118.800 ;
        RECT 26.100 118.200 27.150 119.100 ;
        RECT 22.350 117.450 24.150 118.200 ;
        RECT 7.950 115.500 11.700 116.700 ;
        RECT 10.650 114.600 11.700 115.500 ;
        RECT 19.200 116.400 24.150 117.450 ;
        RECT 25.650 116.400 27.450 118.200 ;
        RECT 34.950 117.600 35.850 130.200 ;
        RECT 47.550 131.550 49.950 132.900 ;
        RECT 51.150 131.550 52.950 143.250 ;
        RECT 47.550 124.950 48.900 131.550 ;
        RECT 55.650 131.400 57.450 143.250 ;
        RECT 70.650 137.400 72.450 143.250 ;
        RECT 73.650 137.400 75.450 143.250 ;
        RECT 76.650 137.400 78.450 143.250 ;
        RECT 50.250 130.200 52.050 130.650 ;
        RECT 56.250 130.200 57.450 131.400 ;
        RECT 50.250 129.000 57.450 130.200 ;
        RECT 74.250 129.150 75.450 137.400 ;
        RECT 81.150 131.400 82.950 143.250 ;
        RECT 84.150 137.400 85.950 143.250 ;
        RECT 89.250 137.400 91.050 143.250 ;
        RECT 94.050 137.400 95.850 143.250 ;
        RECT 89.550 136.500 90.750 137.400 ;
        RECT 97.050 136.500 98.850 143.250 ;
        RECT 100.950 137.400 102.750 143.250 ;
        RECT 105.150 137.400 106.950 143.250 ;
        RECT 109.650 140.400 111.450 143.250 ;
        RECT 85.950 134.400 90.750 136.500 ;
        RECT 93.150 134.700 100.050 136.500 ;
        RECT 105.150 135.300 109.050 137.400 ;
        RECT 89.550 133.500 90.750 134.400 ;
        RECT 102.450 133.800 104.250 134.400 ;
        RECT 89.550 132.300 97.050 133.500 ;
        RECT 95.250 131.700 97.050 132.300 ;
        RECT 97.950 132.900 104.250 133.800 ;
        RECT 81.150 130.800 92.250 131.400 ;
        RECT 97.950 130.800 98.850 132.900 ;
        RECT 102.450 132.600 104.250 132.900 ;
        RECT 105.150 132.600 107.850 134.400 ;
        RECT 105.150 131.700 106.050 132.600 ;
        RECT 81.150 130.200 98.850 130.800 ;
        RECT 50.250 128.850 52.050 129.000 ;
        RECT 46.950 122.850 49.050 124.950 ;
        RECT 46.950 117.600 48.000 122.850 ;
        RECT 50.400 120.600 51.300 128.850 ;
        RECT 53.100 126.150 54.900 127.950 ;
        RECT 52.950 124.050 55.050 126.150 ;
        RECT 70.950 125.850 73.050 127.950 ;
        RECT 73.950 127.050 76.050 129.150 ;
        RECT 56.100 123.150 57.900 124.950 ;
        RECT 71.100 124.050 72.900 125.850 ;
        RECT 55.950 121.050 58.050 123.150 ;
        RECT 50.250 119.700 52.050 120.600 ;
        RECT 74.250 119.700 75.450 127.050 ;
        RECT 76.950 125.850 79.050 127.950 ;
        RECT 77.100 124.050 78.900 125.850 ;
        RECT 50.250 118.800 53.550 119.700 ;
        RECT 19.200 114.600 20.250 116.400 ;
        RECT 28.950 115.500 31.050 117.600 ;
        RECT 28.950 114.600 30.000 115.500 ;
        RECT 5.850 111.750 7.650 114.600 ;
        RECT 10.350 111.750 12.150 114.600 ;
        RECT 14.550 111.750 16.350 114.600 ;
        RECT 18.450 111.750 20.250 114.600 ;
        RECT 21.750 111.750 23.550 114.600 ;
        RECT 26.250 113.700 30.000 114.600 ;
        RECT 26.250 111.750 28.050 113.700 ;
        RECT 31.050 111.750 32.850 114.600 ;
        RECT 34.050 111.750 35.850 117.600 ;
        RECT 46.650 111.750 48.450 117.600 ;
        RECT 52.650 114.600 53.550 118.800 ;
        RECT 71.850 118.800 75.450 119.700 ;
        RECT 49.650 111.750 51.450 114.600 ;
        RECT 52.650 111.750 54.450 114.600 ;
        RECT 55.650 111.750 57.450 114.600 ;
        RECT 71.850 111.750 73.650 118.800 ;
        RECT 81.150 117.600 82.050 130.200 ;
        RECT 90.450 129.900 98.850 130.200 ;
        RECT 100.050 130.800 106.050 131.700 ;
        RECT 106.950 130.800 109.050 131.700 ;
        RECT 112.650 131.400 114.450 143.250 ;
        RECT 123.300 131.400 125.100 143.250 ;
        RECT 127.500 131.400 129.300 143.250 ;
        RECT 130.800 137.400 132.600 143.250 ;
        RECT 146.550 137.400 148.350 143.250 ;
        RECT 149.550 137.400 151.350 143.250 ;
        RECT 152.550 137.400 154.350 143.250 ;
        RECT 164.550 137.400 166.350 143.250 ;
        RECT 167.550 137.400 169.350 143.250 ;
        RECT 170.550 137.400 172.350 143.250 ;
        RECT 185.550 137.400 187.350 143.250 ;
        RECT 188.550 137.400 190.350 143.250 ;
        RECT 90.450 129.600 92.250 129.900 ;
        RECT 100.050 126.150 100.950 130.800 ;
        RECT 106.950 129.600 111.150 130.800 ;
        RECT 110.250 127.800 112.050 129.600 ;
        RECT 91.950 125.100 94.050 126.150 ;
        RECT 83.100 123.150 84.900 124.950 ;
        RECT 86.100 124.050 94.050 125.100 ;
        RECT 97.950 124.050 100.950 126.150 ;
        RECT 86.100 123.300 87.900 124.050 ;
        RECT 84.000 122.400 84.900 123.150 ;
        RECT 89.100 122.400 90.900 123.000 ;
        RECT 84.000 121.200 90.900 122.400 ;
        RECT 89.850 120.000 90.900 121.200 ;
        RECT 100.050 120.000 100.950 124.050 ;
        RECT 109.950 123.750 112.050 124.050 ;
        RECT 108.150 121.950 112.050 123.750 ;
        RECT 113.250 121.950 114.450 131.400 ;
        RECT 122.100 126.150 123.900 127.950 ;
        RECT 127.950 126.150 129.150 131.400 ;
        RECT 130.950 129.150 132.750 130.950 ;
        RECT 149.550 129.150 150.750 137.400 ;
        RECT 167.550 129.150 168.750 137.400 ;
        RECT 130.950 127.050 133.050 129.150 ;
        RECT 121.950 124.050 124.050 126.150 ;
        RECT 124.950 122.850 127.050 124.950 ;
        RECT 127.950 124.050 130.050 126.150 ;
        RECT 145.950 125.850 148.050 127.950 ;
        RECT 148.950 127.050 151.050 129.150 ;
        RECT 146.100 124.050 147.900 125.850 ;
        RECT 89.850 119.100 100.950 120.000 ;
        RECT 109.950 119.850 114.450 121.950 ;
        RECT 125.100 121.050 126.900 122.850 ;
        RECT 128.850 120.750 130.050 124.050 ;
        RECT 89.850 118.200 90.900 119.100 ;
        RECT 100.050 118.800 100.950 119.100 ;
        RECT 76.350 111.750 78.150 117.600 ;
        RECT 81.150 111.750 82.950 117.600 ;
        RECT 85.950 115.500 88.050 117.600 ;
        RECT 89.550 116.400 91.350 118.200 ;
        RECT 92.850 117.450 94.650 118.200 ;
        RECT 92.850 116.400 97.800 117.450 ;
        RECT 100.050 117.000 101.850 118.800 ;
        RECT 113.250 117.600 114.450 119.850 ;
        RECT 129.000 119.700 132.750 120.750 ;
        RECT 106.950 116.700 109.050 117.600 ;
        RECT 87.000 114.600 88.050 115.500 ;
        RECT 96.750 114.600 97.800 116.400 ;
        RECT 105.300 115.500 109.050 116.700 ;
        RECT 105.300 114.600 106.350 115.500 ;
        RECT 84.150 111.750 85.950 114.600 ;
        RECT 87.000 113.700 90.750 114.600 ;
        RECT 88.950 111.750 90.750 113.700 ;
        RECT 93.450 111.750 95.250 114.600 ;
        RECT 96.750 111.750 98.550 114.600 ;
        RECT 100.650 111.750 102.450 114.600 ;
        RECT 104.850 111.750 106.650 114.600 ;
        RECT 109.350 111.750 111.150 114.600 ;
        RECT 112.650 111.750 114.450 117.600 ;
        RECT 122.550 116.700 130.350 118.050 ;
        RECT 122.550 111.750 124.350 116.700 ;
        RECT 125.550 111.750 127.350 115.800 ;
        RECT 128.550 111.750 130.350 116.700 ;
        RECT 131.550 117.600 132.750 119.700 ;
        RECT 149.550 119.700 150.750 127.050 ;
        RECT 151.950 125.850 154.050 127.950 ;
        RECT 163.950 125.850 166.050 127.950 ;
        RECT 166.950 127.050 169.050 129.150 ;
        RECT 152.100 124.050 153.900 125.850 ;
        RECT 164.100 124.050 165.900 125.850 ;
        RECT 167.550 119.700 168.750 127.050 ;
        RECT 169.950 125.850 172.050 127.950 ;
        RECT 170.100 124.050 171.900 125.850 ;
        RECT 188.400 124.950 189.600 137.400 ;
        RECT 200.550 132.300 202.350 143.250 ;
        RECT 203.550 133.200 205.350 143.250 ;
        RECT 206.550 132.300 208.350 143.250 ;
        RECT 200.550 131.400 208.350 132.300 ;
        RECT 209.550 131.400 211.350 143.250 ;
        RECT 227.400 137.400 229.200 143.250 ;
        RECT 230.700 131.400 232.500 143.250 ;
        RECT 234.900 131.400 236.700 143.250 ;
        RECT 245.550 137.400 247.350 143.250 ;
        RECT 248.550 137.400 250.350 143.250 ;
        RECT 265.650 137.400 267.450 143.250 ;
        RECT 268.650 138.000 270.450 143.250 ;
        RECT 209.700 126.150 210.900 131.400 ;
        RECT 227.250 129.150 229.050 130.950 ;
        RECT 226.950 127.050 229.050 129.150 ;
        RECT 230.850 126.150 232.050 131.400 ;
        RECT 236.100 126.150 237.900 127.950 ;
        RECT 185.100 123.150 186.900 124.950 ;
        RECT 184.950 121.050 187.050 123.150 ;
        RECT 187.950 122.850 190.050 124.950 ;
        RECT 199.950 122.850 202.050 124.950 ;
        RECT 203.100 123.150 204.900 124.950 ;
        RECT 149.550 118.800 153.150 119.700 ;
        RECT 167.550 118.800 171.150 119.700 ;
        RECT 131.550 111.750 133.350 117.600 ;
        RECT 146.850 111.750 148.650 117.600 ;
        RECT 151.350 111.750 153.150 118.800 ;
        RECT 164.850 111.750 166.650 117.600 ;
        RECT 169.350 111.750 171.150 118.800 ;
        RECT 188.400 114.600 189.600 122.850 ;
        RECT 200.100 121.050 201.900 122.850 ;
        RECT 202.950 121.050 205.050 123.150 ;
        RECT 205.950 122.850 208.050 124.950 ;
        RECT 208.950 124.050 211.050 126.150 ;
        RECT 229.950 124.050 232.050 126.150 ;
        RECT 206.100 121.050 207.900 122.850 ;
        RECT 209.700 117.600 210.900 124.050 ;
        RECT 229.950 120.750 231.150 124.050 ;
        RECT 232.950 122.850 235.050 124.950 ;
        RECT 235.950 124.050 238.050 126.150 ;
        RECT 248.400 124.950 249.600 137.400 ;
        RECT 266.250 137.100 267.450 137.400 ;
        RECT 271.650 137.400 273.450 143.250 ;
        RECT 274.650 137.400 276.450 143.250 ;
        RECT 271.650 137.100 273.300 137.400 ;
        RECT 266.250 136.200 273.300 137.100 ;
        RECT 266.250 127.950 267.300 136.200 ;
        RECT 272.100 132.150 273.900 133.950 ;
        RECT 268.950 129.150 270.750 130.950 ;
        RECT 271.950 130.050 274.050 132.150 ;
        RECT 289.350 131.400 291.150 143.250 ;
        RECT 292.350 131.400 294.150 143.250 ;
        RECT 295.650 137.400 297.450 143.250 ;
        RECT 305.550 137.400 307.350 143.250 ;
        RECT 308.550 137.400 310.350 143.250 ;
        RECT 311.550 138.000 313.350 143.250 ;
        RECT 275.100 129.150 276.900 130.950 ;
        RECT 265.950 125.850 268.050 127.950 ;
        RECT 268.950 127.050 271.050 129.150 ;
        RECT 274.950 127.050 277.050 129.150 ;
        RECT 289.650 126.150 290.850 131.400 ;
        RECT 296.250 130.500 297.450 137.400 ;
        RECT 308.700 137.100 310.350 137.400 ;
        RECT 314.550 137.400 316.350 143.250 ;
        RECT 326.550 137.400 328.350 143.250 ;
        RECT 329.550 137.400 331.350 143.250 ;
        RECT 314.550 137.100 315.750 137.400 ;
        RECT 308.700 136.200 315.750 137.100 ;
        RECT 308.100 132.150 309.900 133.950 ;
        RECT 291.750 129.600 297.450 130.500 ;
        RECT 291.750 128.700 294.000 129.600 ;
        RECT 305.100 129.150 306.900 130.950 ;
        RECT 307.950 130.050 310.050 132.150 ;
        RECT 311.250 129.150 313.050 130.950 ;
        RECT 245.100 123.150 246.900 124.950 ;
        RECT 233.100 121.050 234.900 122.850 ;
        RECT 244.950 121.050 247.050 123.150 ;
        RECT 247.950 122.850 250.050 124.950 ;
        RECT 227.250 119.700 231.000 120.750 ;
        RECT 227.250 117.600 228.450 119.700 ;
        RECT 185.550 111.750 187.350 114.600 ;
        RECT 188.550 111.750 190.350 114.600 ;
        RECT 201.000 111.750 202.800 117.600 ;
        RECT 205.200 115.950 210.900 117.600 ;
        RECT 205.200 111.750 207.000 115.950 ;
        RECT 208.500 111.750 210.300 114.600 ;
        RECT 226.650 111.750 228.450 117.600 ;
        RECT 229.650 116.700 237.450 118.050 ;
        RECT 229.650 111.750 231.450 116.700 ;
        RECT 232.650 111.750 234.450 115.800 ;
        RECT 235.650 111.750 237.450 116.700 ;
        RECT 248.400 114.600 249.600 122.850 ;
        RECT 266.400 121.650 267.600 125.850 ;
        RECT 289.650 124.050 292.050 126.150 ;
        RECT 266.400 120.000 270.900 121.650 ;
        RECT 245.550 111.750 247.350 114.600 ;
        RECT 248.550 111.750 250.350 114.600 ;
        RECT 269.100 111.750 270.900 120.000 ;
        RECT 274.500 111.750 276.300 120.600 ;
        RECT 289.650 117.600 290.850 124.050 ;
        RECT 292.950 120.300 294.000 128.700 ;
        RECT 296.100 126.150 297.900 127.950 ;
        RECT 304.950 127.050 307.050 129.150 ;
        RECT 310.950 127.050 313.050 129.150 ;
        RECT 314.700 127.950 315.750 136.200 ;
        RECT 295.950 124.050 298.050 126.150 ;
        RECT 313.950 125.850 316.050 127.950 ;
        RECT 314.400 121.650 315.600 125.850 ;
        RECT 329.400 124.950 330.600 137.400 ;
        RECT 345.300 131.400 347.100 143.250 ;
        RECT 349.500 131.400 351.300 143.250 ;
        RECT 352.800 137.400 354.600 143.250 ;
        RECT 365.550 137.400 367.350 143.250 ;
        RECT 368.550 137.400 370.350 143.250 ;
        RECT 371.550 138.000 373.350 143.250 ;
        RECT 368.700 137.100 370.350 137.400 ;
        RECT 374.550 137.400 376.350 143.250 ;
        RECT 386.550 137.400 388.350 143.250 ;
        RECT 389.550 137.400 391.350 143.250 ;
        RECT 392.550 138.000 394.350 143.250 ;
        RECT 374.550 137.100 375.750 137.400 ;
        RECT 368.700 136.200 375.750 137.100 ;
        RECT 389.700 137.100 391.350 137.400 ;
        RECT 395.550 137.400 397.350 143.250 ;
        RECT 409.650 137.400 411.450 143.250 ;
        RECT 412.650 138.000 414.450 143.250 ;
        RECT 395.550 137.100 396.750 137.400 ;
        RECT 389.700 136.200 396.750 137.100 ;
        RECT 368.100 132.150 369.900 133.950 ;
        RECT 344.100 126.150 345.900 127.950 ;
        RECT 349.950 126.150 351.150 131.400 ;
        RECT 352.950 129.150 354.750 130.950 ;
        RECT 365.100 129.150 366.900 130.950 ;
        RECT 367.950 130.050 370.050 132.150 ;
        RECT 371.250 129.150 373.050 130.950 ;
        RECT 352.950 127.050 355.050 129.150 ;
        RECT 364.950 127.050 367.050 129.150 ;
        RECT 370.950 127.050 373.050 129.150 ;
        RECT 374.700 127.950 375.750 136.200 ;
        RECT 389.100 132.150 390.900 133.950 ;
        RECT 386.100 129.150 387.900 130.950 ;
        RECT 388.950 130.050 391.050 132.150 ;
        RECT 392.250 129.150 394.050 130.950 ;
        RECT 326.100 123.150 327.900 124.950 ;
        RECT 291.750 119.400 294.000 120.300 ;
        RECT 291.750 118.500 296.850 119.400 ;
        RECT 289.350 111.750 291.150 117.600 ;
        RECT 292.350 111.750 294.150 117.600 ;
        RECT 295.650 114.600 296.850 118.500 ;
        RECT 295.650 111.750 297.450 114.600 ;
        RECT 305.700 111.750 307.500 120.600 ;
        RECT 311.100 120.000 315.600 121.650 ;
        RECT 325.950 121.050 328.050 123.150 ;
        RECT 328.950 122.850 331.050 124.950 ;
        RECT 343.950 124.050 346.050 126.150 ;
        RECT 346.950 122.850 349.050 124.950 ;
        RECT 349.950 124.050 352.050 126.150 ;
        RECT 373.950 125.850 376.050 127.950 ;
        RECT 385.950 127.050 388.050 129.150 ;
        RECT 391.950 127.050 394.050 129.150 ;
        RECT 395.700 127.950 396.750 136.200 ;
        RECT 410.250 137.100 411.450 137.400 ;
        RECT 415.650 137.400 417.450 143.250 ;
        RECT 418.650 137.400 420.450 143.250 ;
        RECT 415.650 137.100 417.300 137.400 ;
        RECT 410.250 136.200 417.300 137.100 ;
        RECT 410.250 127.950 411.300 136.200 ;
        RECT 416.100 132.150 417.900 133.950 ;
        RECT 412.950 129.150 414.750 130.950 ;
        RECT 415.950 130.050 418.050 132.150 ;
        RECT 429.300 131.400 431.100 143.250 ;
        RECT 433.500 131.400 435.300 143.250 ;
        RECT 436.800 137.400 438.600 143.250 ;
        RECT 454.650 137.400 456.450 143.250 ;
        RECT 457.650 137.400 459.450 143.250 ;
        RECT 470.400 137.400 472.200 143.250 ;
        RECT 419.100 129.150 420.900 130.950 ;
        RECT 394.950 125.850 397.050 127.950 ;
        RECT 409.950 125.850 412.050 127.950 ;
        RECT 412.950 127.050 415.050 129.150 ;
        RECT 418.950 127.050 421.050 129.150 ;
        RECT 428.100 126.150 429.900 127.950 ;
        RECT 433.950 126.150 435.150 131.400 ;
        RECT 436.950 129.150 438.750 130.950 ;
        RECT 436.950 127.050 439.050 129.150 ;
        RECT 311.100 111.750 312.900 120.000 ;
        RECT 329.400 114.600 330.600 122.850 ;
        RECT 347.100 121.050 348.900 122.850 ;
        RECT 350.850 120.750 352.050 124.050 ;
        RECT 374.400 121.650 375.600 125.850 ;
        RECT 395.400 121.650 396.600 125.850 ;
        RECT 351.000 119.700 354.750 120.750 ;
        RECT 344.550 116.700 352.350 118.050 ;
        RECT 326.550 111.750 328.350 114.600 ;
        RECT 329.550 111.750 331.350 114.600 ;
        RECT 344.550 111.750 346.350 116.700 ;
        RECT 347.550 111.750 349.350 115.800 ;
        RECT 350.550 111.750 352.350 116.700 ;
        RECT 353.550 117.600 354.750 119.700 ;
        RECT 353.550 111.750 355.350 117.600 ;
        RECT 365.700 111.750 367.500 120.600 ;
        RECT 371.100 120.000 375.600 121.650 ;
        RECT 371.100 111.750 372.900 120.000 ;
        RECT 386.700 111.750 388.500 120.600 ;
        RECT 392.100 120.000 396.600 121.650 ;
        RECT 410.400 121.650 411.600 125.850 ;
        RECT 427.950 124.050 430.050 126.150 ;
        RECT 430.950 122.850 433.050 124.950 ;
        RECT 433.950 124.050 436.050 126.150 ;
        RECT 455.400 124.950 456.600 137.400 ;
        RECT 473.700 131.400 475.500 143.250 ;
        RECT 477.900 131.400 479.700 143.250 ;
        RECT 488.550 132.300 490.350 143.250 ;
        RECT 491.550 133.200 493.350 143.250 ;
        RECT 494.550 132.300 496.350 143.250 ;
        RECT 488.550 131.400 496.350 132.300 ;
        RECT 497.550 131.400 499.350 143.250 ;
        RECT 509.550 137.400 511.350 143.250 ;
        RECT 512.550 137.400 514.350 143.250 ;
        RECT 515.550 138.000 517.350 143.250 ;
        RECT 512.700 137.100 514.350 137.400 ;
        RECT 518.550 137.400 520.350 143.250 ;
        RECT 535.650 137.400 537.450 143.250 ;
        RECT 538.650 137.400 540.450 143.250 ;
        RECT 518.550 137.100 519.750 137.400 ;
        RECT 512.700 136.200 519.750 137.100 ;
        RECT 512.100 132.150 513.900 133.950 ;
        RECT 470.250 129.150 472.050 130.950 ;
        RECT 469.950 127.050 472.050 129.150 ;
        RECT 473.850 126.150 475.050 131.400 ;
        RECT 479.100 126.150 480.900 127.950 ;
        RECT 497.700 126.150 498.900 131.400 ;
        RECT 509.100 129.150 510.900 130.950 ;
        RECT 511.950 130.050 514.050 132.150 ;
        RECT 515.250 129.150 517.050 130.950 ;
        RECT 508.950 127.050 511.050 129.150 ;
        RECT 514.950 127.050 517.050 129.150 ;
        RECT 518.700 127.950 519.750 136.200 ;
        RECT 410.400 120.000 414.900 121.650 ;
        RECT 431.100 121.050 432.900 122.850 ;
        RECT 434.850 120.750 436.050 124.050 ;
        RECT 454.950 122.850 457.050 124.950 ;
        RECT 458.100 123.150 459.900 124.950 ;
        RECT 472.950 124.050 475.050 126.150 ;
        RECT 392.100 111.750 393.900 120.000 ;
        RECT 413.100 111.750 414.900 120.000 ;
        RECT 418.500 111.750 420.300 120.600 ;
        RECT 435.000 119.700 438.750 120.750 ;
        RECT 428.550 116.700 436.350 118.050 ;
        RECT 428.550 111.750 430.350 116.700 ;
        RECT 431.550 111.750 433.350 115.800 ;
        RECT 434.550 111.750 436.350 116.700 ;
        RECT 437.550 117.600 438.750 119.700 ;
        RECT 437.550 111.750 439.350 117.600 ;
        RECT 455.400 114.600 456.600 122.850 ;
        RECT 457.950 121.050 460.050 123.150 ;
        RECT 472.950 120.750 474.150 124.050 ;
        RECT 475.950 122.850 478.050 124.950 ;
        RECT 478.950 124.050 481.050 126.150 ;
        RECT 487.950 122.850 490.050 124.950 ;
        RECT 491.100 123.150 492.900 124.950 ;
        RECT 476.100 121.050 477.900 122.850 ;
        RECT 488.100 121.050 489.900 122.850 ;
        RECT 490.950 121.050 493.050 123.150 ;
        RECT 493.950 122.850 496.050 124.950 ;
        RECT 496.950 124.050 499.050 126.150 ;
        RECT 517.950 125.850 520.050 127.950 ;
        RECT 494.100 121.050 495.900 122.850 ;
        RECT 470.250 119.700 474.000 120.750 ;
        RECT 470.250 117.600 471.450 119.700 ;
        RECT 454.650 111.750 456.450 114.600 ;
        RECT 457.650 111.750 459.450 114.600 ;
        RECT 469.650 111.750 471.450 117.600 ;
        RECT 472.650 116.700 480.450 118.050 ;
        RECT 497.700 117.600 498.900 124.050 ;
        RECT 518.400 121.650 519.600 125.850 ;
        RECT 536.400 124.950 537.600 137.400 ;
        RECT 549.300 131.400 551.100 143.250 ;
        RECT 553.500 131.400 555.300 143.250 ;
        RECT 556.800 137.400 558.600 143.250 ;
        RECT 569.550 137.400 571.350 143.250 ;
        RECT 572.550 137.400 574.350 143.250 ;
        RECT 548.100 126.150 549.900 127.950 ;
        RECT 553.950 126.150 555.150 131.400 ;
        RECT 556.950 129.150 558.750 130.950 ;
        RECT 556.950 127.050 559.050 129.150 ;
        RECT 535.950 122.850 538.050 124.950 ;
        RECT 539.100 123.150 540.900 124.950 ;
        RECT 547.950 124.050 550.050 126.150 ;
        RECT 472.650 111.750 474.450 116.700 ;
        RECT 475.650 111.750 477.450 115.800 ;
        RECT 478.650 111.750 480.450 116.700 ;
        RECT 489.000 111.750 490.800 117.600 ;
        RECT 493.200 115.950 498.900 117.600 ;
        RECT 493.200 111.750 495.000 115.950 ;
        RECT 496.500 111.750 498.300 114.600 ;
        RECT 509.700 111.750 511.500 120.600 ;
        RECT 515.100 120.000 519.600 121.650 ;
        RECT 515.100 111.750 516.900 120.000 ;
        RECT 536.400 114.600 537.600 122.850 ;
        RECT 538.950 121.050 541.050 123.150 ;
        RECT 550.950 122.850 553.050 124.950 ;
        RECT 553.950 124.050 556.050 126.150 ;
        RECT 572.400 124.950 573.600 137.400 ;
        RECT 584.550 132.300 586.350 143.250 ;
        RECT 587.550 133.200 589.350 143.250 ;
        RECT 590.550 132.300 592.350 143.250 ;
        RECT 584.550 131.400 592.350 132.300 ;
        RECT 593.550 131.400 595.350 143.250 ;
        RECT 607.650 131.400 609.450 143.250 ;
        RECT 610.650 132.300 612.450 143.250 ;
        RECT 613.650 133.200 615.450 143.250 ;
        RECT 616.650 132.300 618.450 143.250 ;
        RECT 631.650 137.400 633.450 143.250 ;
        RECT 634.650 137.400 636.450 143.250 ;
        RECT 650.400 137.400 652.200 143.250 ;
        RECT 610.650 131.400 618.450 132.300 ;
        RECT 574.950 129.450 577.050 130.050 ;
        RECT 589.950 129.450 592.050 130.050 ;
        RECT 574.950 128.550 592.050 129.450 ;
        RECT 574.950 127.950 577.050 128.550 ;
        RECT 589.950 127.950 592.050 128.550 ;
        RECT 593.700 126.150 594.900 131.400 ;
        RECT 608.100 126.150 609.300 131.400 ;
        RECT 551.100 121.050 552.900 122.850 ;
        RECT 554.850 120.750 556.050 124.050 ;
        RECT 569.100 123.150 570.900 124.950 ;
        RECT 568.950 121.050 571.050 123.150 ;
        RECT 571.950 122.850 574.050 124.950 ;
        RECT 583.950 122.850 586.050 124.950 ;
        RECT 587.100 123.150 588.900 124.950 ;
        RECT 555.000 119.700 558.750 120.750 ;
        RECT 548.550 116.700 556.350 118.050 ;
        RECT 535.650 111.750 537.450 114.600 ;
        RECT 538.650 111.750 540.450 114.600 ;
        RECT 548.550 111.750 550.350 116.700 ;
        RECT 551.550 111.750 553.350 115.800 ;
        RECT 554.550 111.750 556.350 116.700 ;
        RECT 557.550 117.600 558.750 119.700 ;
        RECT 557.550 111.750 559.350 117.600 ;
        RECT 572.400 114.600 573.600 122.850 ;
        RECT 584.100 121.050 585.900 122.850 ;
        RECT 586.950 121.050 589.050 123.150 ;
        RECT 589.950 122.850 592.050 124.950 ;
        RECT 592.950 124.050 595.050 126.150 ;
        RECT 607.950 124.050 610.050 126.150 ;
        RECT 632.400 124.950 633.600 137.400 ;
        RECT 653.700 131.400 655.500 143.250 ;
        RECT 657.900 131.400 659.700 143.250 ;
        RECT 668.550 137.400 670.350 143.250 ;
        RECT 671.550 137.400 673.350 143.250 ;
        RECT 650.250 129.150 652.050 130.950 ;
        RECT 649.950 127.050 652.050 129.150 ;
        RECT 653.850 126.150 655.050 131.400 ;
        RECT 659.100 126.150 660.900 127.950 ;
        RECT 668.100 126.150 669.900 127.950 ;
        RECT 590.100 121.050 591.900 122.850 ;
        RECT 593.700 117.600 594.900 124.050 ;
        RECT 569.550 111.750 571.350 114.600 ;
        RECT 572.550 111.750 574.350 114.600 ;
        RECT 585.000 111.750 586.800 117.600 ;
        RECT 589.200 115.950 594.900 117.600 ;
        RECT 608.100 117.600 609.300 124.050 ;
        RECT 610.950 122.850 613.050 124.950 ;
        RECT 614.100 123.150 615.900 124.950 ;
        RECT 611.100 121.050 612.900 122.850 ;
        RECT 613.950 121.050 616.050 123.150 ;
        RECT 616.950 122.850 619.050 124.950 ;
        RECT 631.950 122.850 634.050 124.950 ;
        RECT 635.100 123.150 636.900 124.950 ;
        RECT 652.950 124.050 655.050 126.150 ;
        RECT 617.100 121.050 618.900 122.850 ;
        RECT 608.100 115.950 613.800 117.600 ;
        RECT 589.200 111.750 591.000 115.950 ;
        RECT 592.500 111.750 594.300 114.600 ;
        RECT 608.700 111.750 610.500 114.600 ;
        RECT 612.000 111.750 613.800 115.950 ;
        RECT 616.200 111.750 618.000 117.600 ;
        RECT 632.400 114.600 633.600 122.850 ;
        RECT 634.950 121.050 637.050 123.150 ;
        RECT 652.950 120.750 654.150 124.050 ;
        RECT 655.950 122.850 658.050 124.950 ;
        RECT 658.950 124.050 661.050 126.150 ;
        RECT 667.950 124.050 670.050 126.150 ;
        RECT 656.100 121.050 657.900 122.850 ;
        RECT 650.250 119.700 654.000 120.750 ;
        RECT 671.700 120.300 672.900 137.400 ;
        RECT 675.150 131.400 676.950 143.250 ;
        RECT 678.150 131.400 679.950 143.250 ;
        RECT 692.550 137.400 694.350 143.250 ;
        RECT 695.550 137.400 697.350 143.250 ;
        RECT 698.550 138.000 700.350 143.250 ;
        RECT 695.700 137.100 697.350 137.400 ;
        RECT 701.550 137.400 703.350 143.250 ;
        RECT 701.550 137.100 702.750 137.400 ;
        RECT 695.700 136.200 702.750 137.100 ;
        RECT 695.100 132.150 696.900 133.950 ;
        RECT 673.950 125.850 676.050 127.950 ;
        RECT 678.150 126.150 679.350 131.400 ;
        RECT 692.100 129.150 693.900 130.950 ;
        RECT 694.950 130.050 697.050 132.150 ;
        RECT 698.250 129.150 700.050 130.950 ;
        RECT 691.950 127.050 694.050 129.150 ;
        RECT 697.950 127.050 700.050 129.150 ;
        RECT 701.700 127.950 702.750 136.200 ;
        RECT 713.550 132.300 715.350 143.250 ;
        RECT 716.550 133.200 718.350 143.250 ;
        RECT 719.550 132.300 721.350 143.250 ;
        RECT 713.550 131.400 721.350 132.300 ;
        RECT 722.550 131.400 724.350 143.250 ;
        RECT 735.300 131.400 737.100 143.250 ;
        RECT 739.500 131.400 741.300 143.250 ;
        RECT 742.800 137.400 744.600 143.250 ;
        RECT 756.300 131.400 758.100 143.250 ;
        RECT 760.500 131.400 762.300 143.250 ;
        RECT 763.800 137.400 765.600 143.250 ;
        RECT 777.300 131.400 779.100 143.250 ;
        RECT 781.500 131.400 783.300 143.250 ;
        RECT 784.800 137.400 786.600 143.250 ;
        RECT 800.550 137.400 802.350 143.250 ;
        RECT 803.550 137.400 805.350 143.250 ;
        RECT 821.400 137.400 823.200 143.250 ;
        RECT 706.950 129.450 709.050 130.050 ;
        RECT 715.950 129.450 718.050 130.050 ;
        RECT 706.950 128.550 718.050 129.450 ;
        RECT 706.950 127.950 709.050 128.550 ;
        RECT 715.950 127.950 718.050 128.550 ;
        RECT 674.100 124.050 675.900 125.850 ;
        RECT 676.950 124.050 679.350 126.150 ;
        RECT 700.950 125.850 703.050 127.950 ;
        RECT 722.700 126.150 723.900 131.400 ;
        RECT 734.100 126.150 735.900 127.950 ;
        RECT 739.950 126.150 741.150 131.400 ;
        RECT 742.950 129.150 744.750 130.950 ;
        RECT 742.950 127.050 745.050 129.150 ;
        RECT 755.100 126.150 756.900 127.950 ;
        RECT 760.950 126.150 762.150 131.400 ;
        RECT 763.950 129.150 765.750 130.950 ;
        RECT 763.950 127.050 766.050 129.150 ;
        RECT 776.100 126.150 777.900 127.950 ;
        RECT 781.950 126.150 783.150 131.400 ;
        RECT 784.950 129.150 786.750 130.950 ;
        RECT 784.950 127.050 787.050 129.150 ;
        RECT 650.250 117.600 651.450 119.700 ;
        RECT 668.550 119.100 676.050 120.300 ;
        RECT 631.650 111.750 633.450 114.600 ;
        RECT 634.650 111.750 636.450 114.600 ;
        RECT 649.650 111.750 651.450 117.600 ;
        RECT 652.650 116.700 660.450 118.050 ;
        RECT 652.650 111.750 654.450 116.700 ;
        RECT 655.650 111.750 657.450 115.800 ;
        RECT 658.650 111.750 660.450 116.700 ;
        RECT 668.550 111.750 670.350 119.100 ;
        RECT 674.250 118.500 676.050 119.100 ;
        RECT 678.150 117.600 679.350 124.050 ;
        RECT 701.400 121.650 702.600 125.850 ;
        RECT 712.950 122.850 715.050 124.950 ;
        RECT 716.100 123.150 717.900 124.950 ;
        RECT 673.050 111.750 674.850 117.600 ;
        RECT 676.050 116.100 679.350 117.600 ;
        RECT 676.050 111.750 677.850 116.100 ;
        RECT 692.700 111.750 694.500 120.600 ;
        RECT 698.100 120.000 702.600 121.650 ;
        RECT 713.100 121.050 714.900 122.850 ;
        RECT 715.950 121.050 718.050 123.150 ;
        RECT 718.950 122.850 721.050 124.950 ;
        RECT 721.950 124.050 724.050 126.150 ;
        RECT 733.950 124.050 736.050 126.150 ;
        RECT 719.100 121.050 720.900 122.850 ;
        RECT 698.100 111.750 699.900 120.000 ;
        RECT 722.700 117.600 723.900 124.050 ;
        RECT 736.950 122.850 739.050 124.950 ;
        RECT 739.950 124.050 742.050 126.150 ;
        RECT 754.950 124.050 757.050 126.150 ;
        RECT 737.100 121.050 738.900 122.850 ;
        RECT 740.850 120.750 742.050 124.050 ;
        RECT 757.950 122.850 760.050 124.950 ;
        RECT 760.950 124.050 763.050 126.150 ;
        RECT 775.950 124.050 778.050 126.150 ;
        RECT 758.100 121.050 759.900 122.850 ;
        RECT 761.850 120.750 763.050 124.050 ;
        RECT 778.950 122.850 781.050 124.950 ;
        RECT 781.950 124.050 784.050 126.150 ;
        RECT 803.400 124.950 804.600 137.400 ;
        RECT 824.700 131.400 826.500 143.250 ;
        RECT 828.900 131.400 830.700 143.250 ;
        RECT 834.150 131.400 835.950 143.250 ;
        RECT 837.150 137.400 838.950 143.250 ;
        RECT 842.250 137.400 844.050 143.250 ;
        RECT 847.050 137.400 848.850 143.250 ;
        RECT 842.550 136.500 843.750 137.400 ;
        RECT 850.050 136.500 851.850 143.250 ;
        RECT 853.950 137.400 855.750 143.250 ;
        RECT 858.150 137.400 859.950 143.250 ;
        RECT 862.650 140.400 864.450 143.250 ;
        RECT 838.950 134.400 843.750 136.500 ;
        RECT 846.150 134.700 853.050 136.500 ;
        RECT 858.150 135.300 862.050 137.400 ;
        RECT 842.550 133.500 843.750 134.400 ;
        RECT 855.450 133.800 857.250 134.400 ;
        RECT 842.550 132.300 850.050 133.500 ;
        RECT 848.250 131.700 850.050 132.300 ;
        RECT 850.950 132.900 857.250 133.800 ;
        RECT 821.250 129.150 823.050 130.950 ;
        RECT 820.950 127.050 823.050 129.150 ;
        RECT 824.850 126.150 826.050 131.400 ;
        RECT 834.150 130.800 845.250 131.400 ;
        RECT 850.950 130.800 851.850 132.900 ;
        RECT 855.450 132.600 857.250 132.900 ;
        RECT 858.150 132.600 860.850 134.400 ;
        RECT 858.150 131.700 859.050 132.600 ;
        RECT 834.150 130.200 851.850 130.800 ;
        RECT 830.100 126.150 831.900 127.950 ;
        RECT 779.100 121.050 780.900 122.850 ;
        RECT 782.850 120.750 784.050 124.050 ;
        RECT 800.100 123.150 801.900 124.950 ;
        RECT 799.950 121.050 802.050 123.150 ;
        RECT 802.950 122.850 805.050 124.950 ;
        RECT 823.950 124.050 826.050 126.150 ;
        RECT 741.000 119.700 744.750 120.750 ;
        RECT 762.000 119.700 765.750 120.750 ;
        RECT 783.000 119.700 786.750 120.750 ;
        RECT 714.000 111.750 715.800 117.600 ;
        RECT 718.200 115.950 723.900 117.600 ;
        RECT 734.550 116.700 742.350 118.050 ;
        RECT 718.200 111.750 720.000 115.950 ;
        RECT 721.500 111.750 723.300 114.600 ;
        RECT 734.550 111.750 736.350 116.700 ;
        RECT 737.550 111.750 739.350 115.800 ;
        RECT 740.550 111.750 742.350 116.700 ;
        RECT 743.550 117.600 744.750 119.700 ;
        RECT 743.550 111.750 745.350 117.600 ;
        RECT 755.550 116.700 763.350 118.050 ;
        RECT 755.550 111.750 757.350 116.700 ;
        RECT 758.550 111.750 760.350 115.800 ;
        RECT 761.550 111.750 763.350 116.700 ;
        RECT 764.550 117.600 765.750 119.700 ;
        RECT 764.550 111.750 766.350 117.600 ;
        RECT 776.550 116.700 784.350 118.050 ;
        RECT 776.550 111.750 778.350 116.700 ;
        RECT 779.550 111.750 781.350 115.800 ;
        RECT 782.550 111.750 784.350 116.700 ;
        RECT 785.550 117.600 786.750 119.700 ;
        RECT 785.550 111.750 787.350 117.600 ;
        RECT 803.400 114.600 804.600 122.850 ;
        RECT 823.950 120.750 825.150 124.050 ;
        RECT 826.950 122.850 829.050 124.950 ;
        RECT 829.950 124.050 832.050 126.150 ;
        RECT 827.100 121.050 828.900 122.850 ;
        RECT 821.250 119.700 825.000 120.750 ;
        RECT 821.250 117.600 822.450 119.700 ;
        RECT 800.550 111.750 802.350 114.600 ;
        RECT 803.550 111.750 805.350 114.600 ;
        RECT 820.650 111.750 822.450 117.600 ;
        RECT 823.650 116.700 831.450 118.050 ;
        RECT 823.650 111.750 825.450 116.700 ;
        RECT 826.650 111.750 828.450 115.800 ;
        RECT 829.650 111.750 831.450 116.700 ;
        RECT 834.150 117.600 835.050 130.200 ;
        RECT 843.450 129.900 851.850 130.200 ;
        RECT 853.050 130.800 859.050 131.700 ;
        RECT 859.950 130.800 862.050 131.700 ;
        RECT 865.650 131.400 867.450 143.250 ;
        RECT 878.550 137.400 880.350 143.250 ;
        RECT 881.550 137.400 883.350 143.250 ;
        RECT 843.450 129.600 845.250 129.900 ;
        RECT 853.050 126.150 853.950 130.800 ;
        RECT 859.950 129.600 864.150 130.800 ;
        RECT 863.250 127.800 865.050 129.600 ;
        RECT 844.950 125.100 847.050 126.150 ;
        RECT 836.100 123.150 837.900 124.950 ;
        RECT 839.100 124.050 847.050 125.100 ;
        RECT 850.950 124.050 853.950 126.150 ;
        RECT 839.100 123.300 840.900 124.050 ;
        RECT 837.000 122.400 837.900 123.150 ;
        RECT 842.100 122.400 843.900 123.000 ;
        RECT 837.000 121.200 843.900 122.400 ;
        RECT 842.850 120.000 843.900 121.200 ;
        RECT 853.050 120.000 853.950 124.050 ;
        RECT 862.950 123.750 865.050 124.050 ;
        RECT 861.150 121.950 865.050 123.750 ;
        RECT 866.250 121.950 867.450 131.400 ;
        RECT 881.400 124.950 882.600 137.400 ;
        RECT 878.100 123.150 879.900 124.950 ;
        RECT 842.850 119.100 853.950 120.000 ;
        RECT 862.950 119.850 867.450 121.950 ;
        RECT 877.950 121.050 880.050 123.150 ;
        RECT 880.950 122.850 883.050 124.950 ;
        RECT 842.850 118.200 843.900 119.100 ;
        RECT 853.050 118.800 853.950 119.100 ;
        RECT 834.150 111.750 835.950 117.600 ;
        RECT 838.950 115.500 841.050 117.600 ;
        RECT 842.550 116.400 844.350 118.200 ;
        RECT 845.850 117.450 847.650 118.200 ;
        RECT 845.850 116.400 850.800 117.450 ;
        RECT 853.050 117.000 854.850 118.800 ;
        RECT 866.250 117.600 867.450 119.850 ;
        RECT 859.950 116.700 862.050 117.600 ;
        RECT 840.000 114.600 841.050 115.500 ;
        RECT 849.750 114.600 850.800 116.400 ;
        RECT 858.300 115.500 862.050 116.700 ;
        RECT 858.300 114.600 859.350 115.500 ;
        RECT 837.150 111.750 838.950 114.600 ;
        RECT 840.000 113.700 843.750 114.600 ;
        RECT 841.950 111.750 843.750 113.700 ;
        RECT 846.450 111.750 848.250 114.600 ;
        RECT 849.750 111.750 851.550 114.600 ;
        RECT 853.650 111.750 855.450 114.600 ;
        RECT 857.850 111.750 859.650 114.600 ;
        RECT 862.350 111.750 864.150 114.600 ;
        RECT 865.650 111.750 867.450 117.600 ;
        RECT 881.400 114.600 882.600 122.850 ;
        RECT 878.550 111.750 880.350 114.600 ;
        RECT 881.550 111.750 883.350 114.600 ;
        RECT 8.550 104.400 10.350 107.250 ;
        RECT 11.550 104.400 13.350 107.250 ;
        RECT 29.700 104.400 31.500 107.250 ;
        RECT 7.950 95.850 10.050 97.950 ;
        RECT 11.400 96.150 12.600 104.400 ;
        RECT 33.000 103.050 34.800 107.250 ;
        RECT 29.100 101.400 34.800 103.050 ;
        RECT 37.200 101.400 39.000 107.250 ;
        RECT 47.550 102.300 49.350 107.250 ;
        RECT 50.550 103.200 52.350 107.250 ;
        RECT 53.550 102.300 55.350 107.250 ;
        RECT 8.100 94.050 9.900 95.850 ;
        RECT 10.950 94.050 13.050 96.150 ;
        RECT 29.100 94.950 30.300 101.400 ;
        RECT 47.550 100.950 55.350 102.300 ;
        RECT 56.550 101.400 58.350 107.250 ;
        RECT 56.550 99.300 57.750 101.400 ;
        RECT 71.850 100.200 73.650 107.250 ;
        RECT 76.350 101.400 78.150 107.250 ;
        RECT 91.350 101.400 93.150 107.250 ;
        RECT 94.350 101.400 96.150 107.250 ;
        RECT 97.650 104.400 99.450 107.250 ;
        RECT 71.850 99.300 75.450 100.200 ;
        RECT 54.000 98.250 57.750 99.300 ;
        RECT 32.100 96.150 33.900 97.950 ;
        RECT 11.400 81.600 12.600 94.050 ;
        RECT 28.950 92.850 31.050 94.950 ;
        RECT 31.950 94.050 34.050 96.150 ;
        RECT 34.950 95.850 37.050 97.950 ;
        RECT 38.100 96.150 39.900 97.950 ;
        RECT 50.100 96.150 51.900 97.950 ;
        RECT 35.100 94.050 36.900 95.850 ;
        RECT 37.950 94.050 40.050 96.150 ;
        RECT 46.950 92.850 49.050 94.950 ;
        RECT 49.950 94.050 52.050 96.150 ;
        RECT 53.850 94.950 55.050 98.250 ;
        RECT 52.950 92.850 55.050 94.950 ;
        RECT 71.100 93.150 72.900 94.950 ;
        RECT 29.100 87.600 30.300 92.850 ;
        RECT 47.100 91.050 48.900 92.850 ;
        RECT 52.950 87.600 54.150 92.850 ;
        RECT 55.950 89.850 58.050 91.950 ;
        RECT 70.950 91.050 73.050 93.150 ;
        RECT 74.250 91.950 75.450 99.300 ;
        RECT 91.650 94.950 92.850 101.400 ;
        RECT 97.650 100.500 98.850 104.400 ;
        RECT 107.850 101.400 109.650 107.250 ;
        RECT 93.750 99.600 98.850 100.500 ;
        RECT 112.350 100.200 114.150 107.250 ;
        RECT 127.650 101.400 129.450 107.250 ;
        RECT 93.750 98.700 96.000 99.600 ;
        RECT 77.100 93.150 78.900 94.950 ;
        RECT 73.950 89.850 76.050 91.950 ;
        RECT 76.950 91.050 79.050 93.150 ;
        RECT 91.650 92.850 94.050 94.950 ;
        RECT 55.950 88.050 57.750 89.850 ;
        RECT 8.550 75.750 10.350 81.600 ;
        RECT 11.550 75.750 13.350 81.600 ;
        RECT 28.650 75.750 30.450 87.600 ;
        RECT 31.650 86.700 39.450 87.600 ;
        RECT 31.650 75.750 33.450 86.700 ;
        RECT 34.650 75.750 36.450 85.800 ;
        RECT 37.650 75.750 39.450 86.700 ;
        RECT 48.300 75.750 50.100 87.600 ;
        RECT 52.500 75.750 54.300 87.600 ;
        RECT 74.250 81.600 75.450 89.850 ;
        RECT 91.650 87.600 92.850 92.850 ;
        RECT 94.950 90.300 96.000 98.700 ;
        RECT 110.550 99.300 114.150 100.200 ;
        RECT 128.250 99.300 129.450 101.400 ;
        RECT 130.650 102.300 132.450 107.250 ;
        RECT 133.650 103.200 135.450 107.250 ;
        RECT 136.650 102.300 138.450 107.250 ;
        RECT 149.550 104.400 151.350 107.250 ;
        RECT 152.550 104.400 154.350 107.250 ;
        RECT 155.550 104.400 157.350 107.250 ;
        RECT 169.650 104.400 171.450 107.250 ;
        RECT 172.650 104.400 174.450 107.250 ;
        RECT 130.650 100.950 138.450 102.300 ;
        RECT 97.950 92.850 100.050 94.950 ;
        RECT 107.100 93.150 108.900 94.950 ;
        RECT 98.100 91.050 99.900 92.850 ;
        RECT 106.950 91.050 109.050 93.150 ;
        RECT 110.550 91.950 111.750 99.300 ;
        RECT 128.250 98.250 132.000 99.300 ;
        RECT 130.950 94.950 132.150 98.250 ;
        RECT 153.000 97.950 154.050 104.400 ;
        RECT 134.100 96.150 135.900 97.950 ;
        RECT 113.100 93.150 114.900 94.950 ;
        RECT 93.750 89.400 96.000 90.300 ;
        RECT 109.950 89.850 112.050 91.950 ;
        RECT 112.950 91.050 115.050 93.150 ;
        RECT 130.950 92.850 133.050 94.950 ;
        RECT 133.950 94.050 136.050 96.150 ;
        RECT 151.950 95.850 154.050 97.950 ;
        RECT 170.400 96.150 171.600 104.400 ;
        RECT 188.100 99.000 189.900 107.250 ;
        RECT 136.950 92.850 139.050 94.950 ;
        RECT 148.950 92.850 151.050 94.950 ;
        RECT 127.950 89.850 130.050 91.950 ;
        RECT 93.750 88.500 99.450 89.400 ;
        RECT 55.800 75.750 57.600 81.600 ;
        RECT 70.650 75.750 72.450 81.600 ;
        RECT 73.650 75.750 75.450 81.600 ;
        RECT 76.650 75.750 78.450 81.600 ;
        RECT 91.350 75.750 93.150 87.600 ;
        RECT 94.350 75.750 96.150 87.600 ;
        RECT 98.250 81.600 99.450 88.500 ;
        RECT 110.550 81.600 111.750 89.850 ;
        RECT 128.250 88.050 130.050 89.850 ;
        RECT 131.850 87.600 133.050 92.850 ;
        RECT 137.100 91.050 138.900 92.850 ;
        RECT 149.100 91.050 150.900 92.850 ;
        RECT 153.000 88.650 154.050 95.850 ;
        RECT 154.950 92.850 157.050 94.950 ;
        RECT 169.950 94.050 172.050 96.150 ;
        RECT 172.950 95.850 175.050 97.950 ;
        RECT 185.400 97.350 189.900 99.000 ;
        RECT 193.500 98.400 195.300 107.250 ;
        RECT 212.100 99.000 213.900 107.250 ;
        RECT 209.400 97.350 213.900 99.000 ;
        RECT 217.500 98.400 219.300 107.250 ;
        RECT 227.550 99.900 229.350 107.250 ;
        RECT 232.050 101.400 233.850 107.250 ;
        RECT 235.050 102.900 236.850 107.250 ;
        RECT 235.050 101.400 238.350 102.900 ;
        RECT 248.850 101.400 250.650 107.250 ;
        RECT 233.250 99.900 235.050 100.500 ;
        RECT 227.550 98.700 235.050 99.900 ;
        RECT 173.100 94.050 174.900 95.850 ;
        RECT 155.100 91.050 156.900 92.850 ;
        RECT 153.000 87.600 155.550 88.650 ;
        RECT 97.650 75.750 99.450 81.600 ;
        RECT 107.550 75.750 109.350 81.600 ;
        RECT 110.550 75.750 112.350 81.600 ;
        RECT 113.550 75.750 115.350 81.600 ;
        RECT 128.400 75.750 130.200 81.600 ;
        RECT 131.700 75.750 133.500 87.600 ;
        RECT 135.900 75.750 137.700 87.600 ;
        RECT 149.550 75.750 151.350 87.600 ;
        RECT 153.750 75.750 155.550 87.600 ;
        RECT 170.400 81.600 171.600 94.050 ;
        RECT 185.400 93.150 186.600 97.350 ;
        RECT 209.400 93.150 210.600 97.350 ;
        RECT 184.950 91.050 187.050 93.150 ;
        RECT 185.250 82.800 186.300 91.050 ;
        RECT 187.950 89.850 190.050 91.950 ;
        RECT 193.950 89.850 196.050 91.950 ;
        RECT 208.950 91.050 211.050 93.150 ;
        RECT 226.950 92.850 229.050 94.950 ;
        RECT 187.950 88.050 189.750 89.850 ;
        RECT 190.950 86.850 193.050 88.950 ;
        RECT 194.100 88.050 195.900 89.850 ;
        RECT 191.100 85.050 192.900 86.850 ;
        RECT 209.250 82.800 210.300 91.050 ;
        RECT 211.950 89.850 214.050 91.950 ;
        RECT 217.950 89.850 220.050 91.950 ;
        RECT 227.100 91.050 228.900 92.850 ;
        RECT 211.950 88.050 213.750 89.850 ;
        RECT 214.950 86.850 217.050 88.950 ;
        RECT 218.100 88.050 219.900 89.850 ;
        RECT 215.100 85.050 216.900 86.850 ;
        RECT 185.250 81.900 192.300 82.800 ;
        RECT 185.250 81.600 186.450 81.900 ;
        RECT 169.650 75.750 171.450 81.600 ;
        RECT 172.650 75.750 174.450 81.600 ;
        RECT 184.650 75.750 186.450 81.600 ;
        RECT 190.650 81.600 192.300 81.900 ;
        RECT 209.250 81.900 216.300 82.800 ;
        RECT 209.250 81.600 210.450 81.900 ;
        RECT 187.650 75.750 189.450 81.000 ;
        RECT 190.650 75.750 192.450 81.600 ;
        RECT 193.650 75.750 195.450 81.600 ;
        RECT 208.650 75.750 210.450 81.600 ;
        RECT 214.650 81.600 216.300 81.900 ;
        RECT 230.700 81.600 231.900 98.700 ;
        RECT 237.150 94.950 238.350 101.400 ;
        RECT 253.350 100.200 255.150 107.250 ;
        RECT 266.550 104.400 268.350 107.250 ;
        RECT 269.550 104.400 271.350 107.250 ;
        RECT 272.550 104.400 274.350 107.250 ;
        RECT 251.550 99.300 255.150 100.200 ;
        RECT 233.100 93.150 234.900 94.950 ;
        RECT 232.950 91.050 235.050 93.150 ;
        RECT 235.950 92.850 238.350 94.950 ;
        RECT 248.100 93.150 249.900 94.950 ;
        RECT 237.150 87.600 238.350 92.850 ;
        RECT 247.950 91.050 250.050 93.150 ;
        RECT 251.550 91.950 252.750 99.300 ;
        RECT 270.000 97.950 271.050 104.400 ;
        RECT 286.650 101.400 288.450 107.250 ;
        RECT 287.250 99.300 288.450 101.400 ;
        RECT 289.650 102.300 291.450 107.250 ;
        RECT 292.650 103.200 294.450 107.250 ;
        RECT 295.650 102.300 297.450 107.250 ;
        RECT 305.550 104.400 307.350 107.250 ;
        RECT 308.550 104.400 310.350 107.250 ;
        RECT 289.650 100.950 297.450 102.300 ;
        RECT 287.250 98.250 291.000 99.300 ;
        RECT 268.950 95.850 271.050 97.950 ;
        RECT 254.100 93.150 255.900 94.950 ;
        RECT 250.950 89.850 253.050 91.950 ;
        RECT 253.950 91.050 256.050 93.150 ;
        RECT 265.950 92.850 268.050 94.950 ;
        RECT 266.100 91.050 267.900 92.850 ;
        RECT 211.650 75.750 213.450 81.000 ;
        RECT 214.650 75.750 216.450 81.600 ;
        RECT 217.650 75.750 219.450 81.600 ;
        RECT 227.550 75.750 229.350 81.600 ;
        RECT 230.550 75.750 232.350 81.600 ;
        RECT 234.150 75.750 235.950 87.600 ;
        RECT 237.150 75.750 238.950 87.600 ;
        RECT 251.550 81.600 252.750 89.850 ;
        RECT 270.000 88.650 271.050 95.850 ;
        RECT 289.950 94.950 291.150 98.250 ;
        RECT 293.100 96.150 294.900 97.950 ;
        RECT 271.950 92.850 274.050 94.950 ;
        RECT 289.950 92.850 292.050 94.950 ;
        RECT 292.950 94.050 295.050 96.150 ;
        RECT 304.950 95.850 307.050 97.950 ;
        RECT 308.400 96.150 309.600 104.400 ;
        RECT 326.850 100.200 328.650 107.250 ;
        RECT 331.350 101.400 333.150 107.250 ;
        RECT 344.550 102.300 346.350 107.250 ;
        RECT 347.550 103.200 349.350 107.250 ;
        RECT 350.550 102.300 352.350 107.250 ;
        RECT 344.550 100.950 352.350 102.300 ;
        RECT 353.550 101.400 355.350 107.250 ;
        RECT 365.550 102.300 367.350 107.250 ;
        RECT 368.550 103.200 370.350 107.250 ;
        RECT 371.550 102.300 373.350 107.250 ;
        RECT 326.850 99.300 330.450 100.200 ;
        RECT 353.550 99.300 354.750 101.400 ;
        RECT 365.550 100.950 373.350 102.300 ;
        RECT 374.550 101.400 376.350 107.250 ;
        RECT 374.550 99.300 375.750 101.400 ;
        RECT 295.950 92.850 298.050 94.950 ;
        RECT 305.100 94.050 306.900 95.850 ;
        RECT 307.950 94.050 310.050 96.150 ;
        RECT 272.100 91.050 273.900 92.850 ;
        RECT 286.950 89.850 289.050 91.950 ;
        RECT 270.000 87.600 272.550 88.650 ;
        RECT 287.250 88.050 289.050 89.850 ;
        RECT 290.850 87.600 292.050 92.850 ;
        RECT 296.100 91.050 297.900 92.850 ;
        RECT 248.550 75.750 250.350 81.600 ;
        RECT 251.550 75.750 253.350 81.600 ;
        RECT 254.550 75.750 256.350 81.600 ;
        RECT 266.550 75.750 268.350 87.600 ;
        RECT 270.750 75.750 272.550 87.600 ;
        RECT 287.400 75.750 289.200 81.600 ;
        RECT 290.700 75.750 292.500 87.600 ;
        RECT 294.900 75.750 296.700 87.600 ;
        RECT 308.400 81.600 309.600 94.050 ;
        RECT 326.100 93.150 327.900 94.950 ;
        RECT 325.950 91.050 328.050 93.150 ;
        RECT 329.250 91.950 330.450 99.300 ;
        RECT 351.000 98.250 354.750 99.300 ;
        RECT 372.000 98.250 375.750 99.300 ;
        RECT 389.700 98.400 391.500 107.250 ;
        RECT 395.100 99.000 396.900 107.250 ;
        RECT 347.100 96.150 348.900 97.950 ;
        RECT 332.100 93.150 333.900 94.950 ;
        RECT 328.950 89.850 331.050 91.950 ;
        RECT 331.950 91.050 334.050 93.150 ;
        RECT 343.950 92.850 346.050 94.950 ;
        RECT 346.950 94.050 349.050 96.150 ;
        RECT 350.850 94.950 352.050 98.250 ;
        RECT 368.100 96.150 369.900 97.950 ;
        RECT 349.950 92.850 352.050 94.950 ;
        RECT 364.950 92.850 367.050 94.950 ;
        RECT 367.950 94.050 370.050 96.150 ;
        RECT 371.850 94.950 373.050 98.250 ;
        RECT 395.100 97.350 399.600 99.000 ;
        RECT 410.700 98.400 412.500 107.250 ;
        RECT 416.100 99.000 417.900 107.250 ;
        RECT 431.550 104.400 433.350 107.250 ;
        RECT 434.550 104.400 436.350 107.250 ;
        RECT 449.550 104.400 451.350 107.250 ;
        RECT 452.550 104.400 454.350 107.250 ;
        RECT 455.550 104.400 457.350 107.250 ;
        RECT 416.100 97.350 420.600 99.000 ;
        RECT 370.950 92.850 373.050 94.950 ;
        RECT 398.400 93.150 399.600 97.350 ;
        RECT 419.400 93.150 420.600 97.350 ;
        RECT 430.950 95.850 433.050 97.950 ;
        RECT 434.400 96.150 435.600 104.400 ;
        RECT 453.000 97.950 454.050 104.400 ;
        RECT 470.850 101.400 472.650 107.250 ;
        RECT 475.350 100.200 477.150 107.250 ;
        RECT 493.650 101.400 495.450 107.250 ;
        RECT 431.100 94.050 432.900 95.850 ;
        RECT 433.950 94.050 436.050 96.150 ;
        RECT 451.950 95.850 454.050 97.950 ;
        RECT 344.100 91.050 345.900 92.850 ;
        RECT 329.250 81.600 330.450 89.850 ;
        RECT 349.950 87.600 351.150 92.850 ;
        RECT 352.950 89.850 355.050 91.950 ;
        RECT 365.100 91.050 366.900 92.850 ;
        RECT 352.950 88.050 354.750 89.850 ;
        RECT 370.950 87.600 372.150 92.850 ;
        RECT 373.950 89.850 376.050 91.950 ;
        RECT 388.950 89.850 391.050 91.950 ;
        RECT 394.950 89.850 397.050 91.950 ;
        RECT 397.950 91.050 400.050 93.150 ;
        RECT 373.950 88.050 375.750 89.850 ;
        RECT 389.100 88.050 390.900 89.850 ;
        RECT 305.550 75.750 307.350 81.600 ;
        RECT 308.550 75.750 310.350 81.600 ;
        RECT 325.650 75.750 327.450 81.600 ;
        RECT 328.650 75.750 330.450 81.600 ;
        RECT 331.650 75.750 333.450 81.600 ;
        RECT 345.300 75.750 347.100 87.600 ;
        RECT 349.500 75.750 351.300 87.600 ;
        RECT 352.800 75.750 354.600 81.600 ;
        RECT 366.300 75.750 368.100 87.600 ;
        RECT 370.500 75.750 372.300 87.600 ;
        RECT 391.950 86.850 394.050 88.950 ;
        RECT 395.250 88.050 397.050 89.850 ;
        RECT 392.100 85.050 393.900 86.850 ;
        RECT 398.700 82.800 399.750 91.050 ;
        RECT 409.950 89.850 412.050 91.950 ;
        RECT 415.950 89.850 418.050 91.950 ;
        RECT 418.950 91.050 421.050 93.150 ;
        RECT 410.100 88.050 411.900 89.850 ;
        RECT 412.950 86.850 415.050 88.950 ;
        RECT 416.250 88.050 418.050 89.850 ;
        RECT 413.100 85.050 414.900 86.850 ;
        RECT 419.700 82.800 420.750 91.050 ;
        RECT 392.700 81.900 399.750 82.800 ;
        RECT 392.700 81.600 394.350 81.900 ;
        RECT 373.800 75.750 375.600 81.600 ;
        RECT 389.550 75.750 391.350 81.600 ;
        RECT 392.550 75.750 394.350 81.600 ;
        RECT 398.550 81.600 399.750 81.900 ;
        RECT 413.700 81.900 420.750 82.800 ;
        RECT 413.700 81.600 415.350 81.900 ;
        RECT 395.550 75.750 397.350 81.000 ;
        RECT 398.550 75.750 400.350 81.600 ;
        RECT 410.550 75.750 412.350 81.600 ;
        RECT 413.550 75.750 415.350 81.600 ;
        RECT 419.550 81.600 420.750 81.900 ;
        RECT 434.400 81.600 435.600 94.050 ;
        RECT 448.950 92.850 451.050 94.950 ;
        RECT 449.100 91.050 450.900 92.850 ;
        RECT 453.000 88.650 454.050 95.850 ;
        RECT 473.550 99.300 477.150 100.200 ;
        RECT 494.250 99.300 495.450 101.400 ;
        RECT 496.650 102.300 498.450 107.250 ;
        RECT 499.650 103.200 501.450 107.250 ;
        RECT 502.650 102.300 504.450 107.250 ;
        RECT 514.650 104.400 516.450 107.250 ;
        RECT 517.650 104.400 519.450 107.250 ;
        RECT 496.650 100.950 504.450 102.300 ;
        RECT 454.950 92.850 457.050 94.950 ;
        RECT 470.100 93.150 471.900 94.950 ;
        RECT 455.100 91.050 456.900 92.850 ;
        RECT 469.950 91.050 472.050 93.150 ;
        RECT 473.550 91.950 474.750 99.300 ;
        RECT 494.250 98.250 498.000 99.300 ;
        RECT 496.950 94.950 498.150 98.250 ;
        RECT 500.100 96.150 501.900 97.950 ;
        RECT 515.400 96.150 516.600 104.400 ;
        RECT 527.550 101.400 529.350 107.250 ;
        RECT 530.550 101.400 532.350 107.250 ;
        RECT 546.150 102.900 547.950 107.250 ;
        RECT 544.650 101.400 547.950 102.900 ;
        RECT 549.150 101.400 550.950 107.250 ;
        RECT 476.100 93.150 477.900 94.950 ;
        RECT 472.950 89.850 475.050 91.950 ;
        RECT 475.950 91.050 478.050 93.150 ;
        RECT 496.950 92.850 499.050 94.950 ;
        RECT 499.950 94.050 502.050 96.150 ;
        RECT 502.950 92.850 505.050 94.950 ;
        RECT 514.950 94.050 517.050 96.150 ;
        RECT 517.950 95.850 520.050 97.950 ;
        RECT 527.100 96.150 528.900 97.950 ;
        RECT 518.100 94.050 519.900 95.850 ;
        RECT 526.950 94.050 529.050 96.150 ;
        RECT 530.400 94.950 531.600 101.400 ;
        RECT 544.650 94.950 545.850 101.400 ;
        RECT 547.950 99.900 549.750 100.500 ;
        RECT 553.650 99.900 555.450 107.250 ;
        RECT 547.950 98.700 555.450 99.900 ;
        RECT 493.950 89.850 496.050 91.950 ;
        RECT 453.000 87.600 455.550 88.650 ;
        RECT 416.550 75.750 418.350 81.000 ;
        RECT 419.550 75.750 421.350 81.600 ;
        RECT 431.550 75.750 433.350 81.600 ;
        RECT 434.550 75.750 436.350 81.600 ;
        RECT 449.550 75.750 451.350 87.600 ;
        RECT 453.750 75.750 455.550 87.600 ;
        RECT 473.550 81.600 474.750 89.850 ;
        RECT 494.250 88.050 496.050 89.850 ;
        RECT 497.850 87.600 499.050 92.850 ;
        RECT 503.100 91.050 504.900 92.850 ;
        RECT 470.550 75.750 472.350 81.600 ;
        RECT 473.550 75.750 475.350 81.600 ;
        RECT 476.550 75.750 478.350 81.600 ;
        RECT 494.400 75.750 496.200 81.600 ;
        RECT 497.700 75.750 499.500 87.600 ;
        RECT 501.900 75.750 503.700 87.600 ;
        RECT 515.400 81.600 516.600 94.050 ;
        RECT 529.950 92.850 532.050 94.950 ;
        RECT 544.650 92.850 547.050 94.950 ;
        RECT 548.100 93.150 549.900 94.950 ;
        RECT 530.400 87.600 531.600 92.850 ;
        RECT 544.650 87.600 545.850 92.850 ;
        RECT 547.950 91.050 550.050 93.150 ;
        RECT 514.650 75.750 516.450 81.600 ;
        RECT 517.650 75.750 519.450 81.600 ;
        RECT 527.550 75.750 529.350 87.600 ;
        RECT 530.550 75.750 532.350 87.600 ;
        RECT 544.050 75.750 545.850 87.600 ;
        RECT 547.050 75.750 548.850 87.600 ;
        RECT 551.100 81.600 552.300 98.700 ;
        RECT 563.700 98.400 565.500 107.250 ;
        RECT 569.100 99.000 570.900 107.250 ;
        RECT 590.100 99.000 591.900 107.250 ;
        RECT 569.100 97.350 573.600 99.000 ;
        RECT 553.950 92.850 556.050 94.950 ;
        RECT 572.400 93.150 573.600 97.350 ;
        RECT 587.400 97.350 591.900 99.000 ;
        RECT 595.500 98.400 597.300 107.250 ;
        RECT 611.850 100.200 613.650 107.250 ;
        RECT 616.350 101.400 618.150 107.250 ;
        RECT 626.550 102.300 628.350 107.250 ;
        RECT 629.550 103.200 631.350 107.250 ;
        RECT 632.550 102.300 634.350 107.250 ;
        RECT 626.550 100.950 634.350 102.300 ;
        RECT 635.550 101.400 637.350 107.250 ;
        RECT 652.800 101.400 654.600 107.250 ;
        RECT 657.000 101.400 658.800 107.250 ;
        RECT 661.200 101.400 663.000 107.250 ;
        RECT 666.150 101.400 667.950 107.250 ;
        RECT 669.150 104.400 670.950 107.250 ;
        RECT 673.950 105.300 675.750 107.250 ;
        RECT 672.000 104.400 675.750 105.300 ;
        RECT 678.450 104.400 680.250 107.250 ;
        RECT 681.750 104.400 683.550 107.250 ;
        RECT 685.650 104.400 687.450 107.250 ;
        RECT 689.850 104.400 691.650 107.250 ;
        RECT 694.350 104.400 696.150 107.250 ;
        RECT 672.000 103.500 673.050 104.400 ;
        RECT 670.950 101.400 673.050 103.500 ;
        RECT 681.750 102.600 682.800 104.400 ;
        RECT 611.850 99.300 615.450 100.200 ;
        RECT 635.550 99.300 636.750 101.400 ;
        RECT 587.400 93.150 588.600 97.350 ;
        RECT 611.100 93.150 612.900 94.950 ;
        RECT 554.100 91.050 555.900 92.850 ;
        RECT 562.950 89.850 565.050 91.950 ;
        RECT 568.950 89.850 571.050 91.950 ;
        RECT 571.950 91.050 574.050 93.150 ;
        RECT 586.950 91.050 589.050 93.150 ;
        RECT 563.100 88.050 564.900 89.850 ;
        RECT 565.950 86.850 568.050 88.950 ;
        RECT 569.250 88.050 571.050 89.850 ;
        RECT 566.100 85.050 567.900 86.850 ;
        RECT 572.700 82.800 573.750 91.050 ;
        RECT 566.700 81.900 573.750 82.800 ;
        RECT 566.700 81.600 568.350 81.900 ;
        RECT 550.650 75.750 552.450 81.600 ;
        RECT 553.650 75.750 555.450 81.600 ;
        RECT 563.550 75.750 565.350 81.600 ;
        RECT 566.550 75.750 568.350 81.600 ;
        RECT 572.550 81.600 573.750 81.900 ;
        RECT 587.250 82.800 588.300 91.050 ;
        RECT 589.950 89.850 592.050 91.950 ;
        RECT 595.950 89.850 598.050 91.950 ;
        RECT 610.950 91.050 613.050 93.150 ;
        RECT 614.250 91.950 615.450 99.300 ;
        RECT 633.000 98.250 636.750 99.300 ;
        RECT 637.950 99.450 640.050 100.050 ;
        RECT 649.950 99.450 652.050 100.050 ;
        RECT 637.950 98.550 652.050 99.450 ;
        RECT 629.100 96.150 630.900 97.950 ;
        RECT 617.100 93.150 618.900 94.950 ;
        RECT 613.950 89.850 616.050 91.950 ;
        RECT 616.950 91.050 619.050 93.150 ;
        RECT 625.950 92.850 628.050 94.950 ;
        RECT 628.950 94.050 631.050 96.150 ;
        RECT 632.850 94.950 634.050 98.250 ;
        RECT 637.950 97.950 640.050 98.550 ;
        RECT 649.950 97.950 652.050 98.550 ;
        RECT 653.250 96.150 655.050 97.950 ;
        RECT 631.950 92.850 634.050 94.950 ;
        RECT 649.950 92.850 652.050 94.950 ;
        RECT 652.950 94.050 655.050 96.150 ;
        RECT 657.000 94.950 658.050 101.400 ;
        RECT 655.950 92.850 658.050 94.950 ;
        RECT 658.950 96.150 660.750 97.950 ;
        RECT 658.950 94.050 661.050 96.150 ;
        RECT 661.950 92.850 664.050 94.950 ;
        RECT 626.100 91.050 627.900 92.850 ;
        RECT 589.950 88.050 591.750 89.850 ;
        RECT 592.950 86.850 595.050 88.950 ;
        RECT 596.100 88.050 597.900 89.850 ;
        RECT 593.100 85.050 594.900 86.850 ;
        RECT 587.250 81.900 594.300 82.800 ;
        RECT 587.250 81.600 588.450 81.900 ;
        RECT 569.550 75.750 571.350 81.000 ;
        RECT 572.550 75.750 574.350 81.600 ;
        RECT 586.650 75.750 588.450 81.600 ;
        RECT 592.650 81.600 594.300 81.900 ;
        RECT 614.250 81.600 615.450 89.850 ;
        RECT 631.950 87.600 633.150 92.850 ;
        RECT 634.950 89.850 637.050 91.950 ;
        RECT 650.100 91.050 651.900 92.850 ;
        RECT 634.950 88.050 636.750 89.850 ;
        RECT 655.950 89.400 656.850 92.850 ;
        RECT 661.950 91.050 663.750 92.850 ;
        RECT 652.800 88.500 656.850 89.400 ;
        RECT 666.150 88.800 667.050 101.400 ;
        RECT 674.550 100.800 676.350 102.600 ;
        RECT 677.850 101.550 682.800 102.600 ;
        RECT 690.300 103.500 691.350 104.400 ;
        RECT 690.300 102.300 694.050 103.500 ;
        RECT 677.850 100.800 679.650 101.550 ;
        RECT 674.850 99.900 675.900 100.800 ;
        RECT 685.050 100.200 686.850 102.000 ;
        RECT 691.950 101.400 694.050 102.300 ;
        RECT 697.650 101.400 699.450 107.250 ;
        RECT 707.550 104.400 709.350 107.250 ;
        RECT 710.550 104.400 712.350 107.250 ;
        RECT 685.050 99.900 685.950 100.200 ;
        RECT 674.850 99.000 685.950 99.900 ;
        RECT 698.250 99.150 699.450 101.400 ;
        RECT 674.850 97.800 675.900 99.000 ;
        RECT 669.000 96.600 675.900 97.800 ;
        RECT 669.000 95.850 669.900 96.600 ;
        RECT 674.100 96.000 675.900 96.600 ;
        RECT 668.100 94.050 669.900 95.850 ;
        RECT 671.100 94.950 672.900 95.700 ;
        RECT 685.050 94.950 685.950 99.000 ;
        RECT 694.950 97.050 699.450 99.150 ;
        RECT 693.150 95.250 697.050 97.050 ;
        RECT 694.950 94.950 697.050 95.250 ;
        RECT 671.100 93.900 679.050 94.950 ;
        RECT 676.950 92.850 679.050 93.900 ;
        RECT 682.950 92.850 685.950 94.950 ;
        RECT 675.450 89.100 677.250 89.400 ;
        RECT 675.450 88.800 683.850 89.100 ;
        RECT 652.800 87.600 654.600 88.500 ;
        RECT 666.150 88.200 683.850 88.800 ;
        RECT 666.150 87.600 677.250 88.200 ;
        RECT 589.650 75.750 591.450 81.000 ;
        RECT 592.650 75.750 594.450 81.600 ;
        RECT 595.650 75.750 597.450 81.600 ;
        RECT 610.650 75.750 612.450 81.600 ;
        RECT 613.650 75.750 615.450 81.600 ;
        RECT 616.650 75.750 618.450 81.600 ;
        RECT 627.300 75.750 629.100 87.600 ;
        RECT 631.500 75.750 633.300 87.600 ;
        RECT 634.800 75.750 636.600 81.600 ;
        RECT 649.650 76.500 651.450 87.600 ;
        RECT 652.650 77.400 654.450 87.600 ;
        RECT 655.650 86.400 663.450 87.300 ;
        RECT 655.650 76.500 657.450 86.400 ;
        RECT 649.650 75.750 657.450 76.500 ;
        RECT 658.650 75.750 660.450 85.500 ;
        RECT 661.650 75.750 663.450 86.400 ;
        RECT 666.150 75.750 667.950 87.600 ;
        RECT 680.250 86.700 682.050 87.300 ;
        RECT 674.550 85.500 682.050 86.700 ;
        RECT 682.950 86.100 683.850 88.200 ;
        RECT 685.050 88.200 685.950 92.850 ;
        RECT 695.250 89.400 697.050 91.200 ;
        RECT 691.950 88.200 696.150 89.400 ;
        RECT 685.050 87.300 691.050 88.200 ;
        RECT 691.950 87.300 694.050 88.200 ;
        RECT 698.250 87.600 699.450 97.050 ;
        RECT 706.950 95.850 709.050 97.950 ;
        RECT 710.400 96.150 711.600 104.400 ;
        RECT 724.650 101.400 726.450 107.250 ;
        RECT 725.250 99.300 726.450 101.400 ;
        RECT 727.650 102.300 729.450 107.250 ;
        RECT 730.650 103.200 732.450 107.250 ;
        RECT 733.650 102.300 735.450 107.250 ;
        RECT 745.650 104.400 747.450 107.250 ;
        RECT 748.650 104.400 750.450 107.250 ;
        RECT 727.650 100.950 735.450 102.300 ;
        RECT 725.250 98.250 729.000 99.300 ;
        RECT 707.100 94.050 708.900 95.850 ;
        RECT 709.950 94.050 712.050 96.150 ;
        RECT 727.950 94.950 729.150 98.250 ;
        RECT 731.100 96.150 732.900 97.950 ;
        RECT 746.400 96.150 747.600 104.400 ;
        RECT 752.550 101.400 754.350 107.250 ;
        RECT 755.850 104.400 757.650 107.250 ;
        RECT 760.350 104.400 762.150 107.250 ;
        RECT 764.550 104.400 766.350 107.250 ;
        RECT 768.450 104.400 770.250 107.250 ;
        RECT 771.750 104.400 773.550 107.250 ;
        RECT 776.250 105.300 778.050 107.250 ;
        RECT 776.250 104.400 780.000 105.300 ;
        RECT 781.050 104.400 782.850 107.250 ;
        RECT 760.650 103.500 761.700 104.400 ;
        RECT 757.950 102.300 761.700 103.500 ;
        RECT 769.200 102.600 770.250 104.400 ;
        RECT 778.950 103.500 780.000 104.400 ;
        RECT 757.950 101.400 760.050 102.300 ;
        RECT 752.550 99.150 753.750 101.400 ;
        RECT 765.150 100.200 766.950 102.000 ;
        RECT 769.200 101.550 774.150 102.600 ;
        RECT 772.350 100.800 774.150 101.550 ;
        RECT 775.650 100.800 777.450 102.600 ;
        RECT 778.950 101.400 781.050 103.500 ;
        RECT 784.050 101.400 785.850 107.250 ;
        RECT 766.050 99.900 766.950 100.200 ;
        RECT 776.100 99.900 777.150 100.800 ;
        RECT 690.150 86.400 691.050 87.300 ;
        RECT 687.450 86.100 689.250 86.400 ;
        RECT 674.550 84.600 675.750 85.500 ;
        RECT 682.950 85.200 689.250 86.100 ;
        RECT 687.450 84.600 689.250 85.200 ;
        RECT 690.150 84.600 692.850 86.400 ;
        RECT 670.950 82.500 675.750 84.600 ;
        RECT 678.150 82.500 685.050 84.300 ;
        RECT 674.550 81.600 675.750 82.500 ;
        RECT 669.150 75.750 670.950 81.600 ;
        RECT 674.250 75.750 676.050 81.600 ;
        RECT 679.050 75.750 680.850 81.600 ;
        RECT 682.050 75.750 683.850 82.500 ;
        RECT 690.150 81.600 694.050 83.700 ;
        RECT 685.950 75.750 687.750 81.600 ;
        RECT 690.150 75.750 691.950 81.600 ;
        RECT 694.650 75.750 696.450 78.600 ;
        RECT 697.650 75.750 699.450 87.600 ;
        RECT 710.400 81.600 711.600 94.050 ;
        RECT 727.950 92.850 730.050 94.950 ;
        RECT 730.950 94.050 733.050 96.150 ;
        RECT 733.950 92.850 736.050 94.950 ;
        RECT 745.950 94.050 748.050 96.150 ;
        RECT 748.950 95.850 751.050 97.950 ;
        RECT 752.550 97.050 757.050 99.150 ;
        RECT 766.050 99.000 777.150 99.900 ;
        RECT 749.100 94.050 750.900 95.850 ;
        RECT 724.950 89.850 727.050 91.950 ;
        RECT 725.250 88.050 727.050 89.850 ;
        RECT 728.850 87.600 730.050 92.850 ;
        RECT 734.100 91.050 735.900 92.850 ;
        RECT 707.550 75.750 709.350 81.600 ;
        RECT 710.550 75.750 712.350 81.600 ;
        RECT 725.400 75.750 727.200 81.600 ;
        RECT 728.700 75.750 730.500 87.600 ;
        RECT 732.900 75.750 734.700 87.600 ;
        RECT 746.400 81.600 747.600 94.050 ;
        RECT 752.550 87.600 753.750 97.050 ;
        RECT 754.950 95.250 758.850 97.050 ;
        RECT 754.950 94.950 757.050 95.250 ;
        RECT 766.050 94.950 766.950 99.000 ;
        RECT 776.100 97.800 777.150 99.000 ;
        RECT 776.100 96.600 783.000 97.800 ;
        RECT 776.100 96.000 777.900 96.600 ;
        RECT 782.100 95.850 783.000 96.600 ;
        RECT 779.100 94.950 780.900 95.700 ;
        RECT 766.050 92.850 769.050 94.950 ;
        RECT 772.950 93.900 780.900 94.950 ;
        RECT 782.100 94.050 783.900 95.850 ;
        RECT 772.950 92.850 775.050 93.900 ;
        RECT 754.950 89.400 756.750 91.200 ;
        RECT 755.850 88.200 760.050 89.400 ;
        RECT 766.050 88.200 766.950 92.850 ;
        RECT 774.750 89.100 776.550 89.400 ;
        RECT 745.650 75.750 747.450 81.600 ;
        RECT 748.650 75.750 750.450 81.600 ;
        RECT 752.550 75.750 754.350 87.600 ;
        RECT 757.950 87.300 760.050 88.200 ;
        RECT 760.950 87.300 766.950 88.200 ;
        RECT 768.150 88.800 776.550 89.100 ;
        RECT 784.950 88.800 785.850 101.400 ;
        RECT 768.150 88.200 785.850 88.800 ;
        RECT 760.950 86.400 761.850 87.300 ;
        RECT 759.150 84.600 761.850 86.400 ;
        RECT 762.750 86.100 764.550 86.400 ;
        RECT 768.150 86.100 769.050 88.200 ;
        RECT 774.750 87.600 785.850 88.200 ;
        RECT 762.750 85.200 769.050 86.100 ;
        RECT 769.950 86.700 771.750 87.300 ;
        RECT 769.950 85.500 777.450 86.700 ;
        RECT 762.750 84.600 764.550 85.200 ;
        RECT 776.250 84.600 777.450 85.500 ;
        RECT 757.950 81.600 761.850 83.700 ;
        RECT 766.950 82.500 773.850 84.300 ;
        RECT 776.250 82.500 781.050 84.600 ;
        RECT 755.550 75.750 757.350 78.600 ;
        RECT 760.050 75.750 761.850 81.600 ;
        RECT 764.250 75.750 766.050 81.600 ;
        RECT 768.150 75.750 769.950 82.500 ;
        RECT 776.250 81.600 777.450 82.500 ;
        RECT 771.150 75.750 772.950 81.600 ;
        RECT 775.950 75.750 777.750 81.600 ;
        RECT 781.050 75.750 782.850 81.600 ;
        RECT 784.050 75.750 785.850 87.600 ;
        RECT 789.150 101.400 790.950 107.250 ;
        RECT 792.150 104.400 793.950 107.250 ;
        RECT 796.950 105.300 798.750 107.250 ;
        RECT 795.000 104.400 798.750 105.300 ;
        RECT 801.450 104.400 803.250 107.250 ;
        RECT 804.750 104.400 806.550 107.250 ;
        RECT 808.650 104.400 810.450 107.250 ;
        RECT 812.850 104.400 814.650 107.250 ;
        RECT 817.350 104.400 819.150 107.250 ;
        RECT 795.000 103.500 796.050 104.400 ;
        RECT 793.950 101.400 796.050 103.500 ;
        RECT 804.750 102.600 805.800 104.400 ;
        RECT 789.150 88.800 790.050 101.400 ;
        RECT 797.550 100.800 799.350 102.600 ;
        RECT 800.850 101.550 805.800 102.600 ;
        RECT 813.300 103.500 814.350 104.400 ;
        RECT 813.300 102.300 817.050 103.500 ;
        RECT 800.850 100.800 802.650 101.550 ;
        RECT 797.850 99.900 798.900 100.800 ;
        RECT 808.050 100.200 809.850 102.000 ;
        RECT 814.950 101.400 817.050 102.300 ;
        RECT 820.650 101.400 822.450 107.250 ;
        RECT 835.800 101.400 837.600 107.250 ;
        RECT 840.000 101.400 841.800 107.250 ;
        RECT 844.200 101.400 846.000 107.250 ;
        RECT 856.650 104.400 858.450 107.250 ;
        RECT 859.650 104.400 861.450 107.250 ;
        RECT 808.050 99.900 808.950 100.200 ;
        RECT 797.850 99.000 808.950 99.900 ;
        RECT 821.250 99.150 822.450 101.400 ;
        RECT 797.850 97.800 798.900 99.000 ;
        RECT 792.000 96.600 798.900 97.800 ;
        RECT 792.000 95.850 792.900 96.600 ;
        RECT 797.100 96.000 798.900 96.600 ;
        RECT 791.100 94.050 792.900 95.850 ;
        RECT 794.100 94.950 795.900 95.700 ;
        RECT 808.050 94.950 808.950 99.000 ;
        RECT 817.950 97.050 822.450 99.150 ;
        RECT 816.150 95.250 820.050 97.050 ;
        RECT 817.950 94.950 820.050 95.250 ;
        RECT 794.100 93.900 802.050 94.950 ;
        RECT 799.950 92.850 802.050 93.900 ;
        RECT 805.950 92.850 808.950 94.950 ;
        RECT 798.450 89.100 800.250 89.400 ;
        RECT 798.450 88.800 806.850 89.100 ;
        RECT 789.150 88.200 806.850 88.800 ;
        RECT 789.150 87.600 800.250 88.200 ;
        RECT 789.150 75.750 790.950 87.600 ;
        RECT 803.250 86.700 805.050 87.300 ;
        RECT 797.550 85.500 805.050 86.700 ;
        RECT 805.950 86.100 806.850 88.200 ;
        RECT 808.050 88.200 808.950 92.850 ;
        RECT 818.250 89.400 820.050 91.200 ;
        RECT 814.950 88.200 819.150 89.400 ;
        RECT 808.050 87.300 814.050 88.200 ;
        RECT 814.950 87.300 817.050 88.200 ;
        RECT 821.250 87.600 822.450 97.050 ;
        RECT 836.250 96.150 838.050 97.950 ;
        RECT 832.950 92.850 835.050 94.950 ;
        RECT 835.950 94.050 838.050 96.150 ;
        RECT 840.000 94.950 841.050 101.400 ;
        RECT 838.950 92.850 841.050 94.950 ;
        RECT 841.950 96.150 843.750 97.950 ;
        RECT 857.400 96.150 858.600 104.400 ;
        RECT 869.850 101.400 871.650 107.250 ;
        RECT 874.350 100.200 876.150 107.250 ;
        RECT 872.550 99.300 876.150 100.200 ;
        RECT 841.950 94.050 844.050 96.150 ;
        RECT 844.950 92.850 847.050 94.950 ;
        RECT 856.950 94.050 859.050 96.150 ;
        RECT 859.950 95.850 862.050 97.950 ;
        RECT 860.100 94.050 861.900 95.850 ;
        RECT 833.100 91.050 834.900 92.850 ;
        RECT 838.950 89.400 839.850 92.850 ;
        RECT 844.950 91.050 846.750 92.850 ;
        RECT 835.800 88.500 839.850 89.400 ;
        RECT 835.800 87.600 837.600 88.500 ;
        RECT 813.150 86.400 814.050 87.300 ;
        RECT 810.450 86.100 812.250 86.400 ;
        RECT 797.550 84.600 798.750 85.500 ;
        RECT 805.950 85.200 812.250 86.100 ;
        RECT 810.450 84.600 812.250 85.200 ;
        RECT 813.150 84.600 815.850 86.400 ;
        RECT 793.950 82.500 798.750 84.600 ;
        RECT 801.150 82.500 808.050 84.300 ;
        RECT 797.550 81.600 798.750 82.500 ;
        RECT 792.150 75.750 793.950 81.600 ;
        RECT 797.250 75.750 799.050 81.600 ;
        RECT 802.050 75.750 803.850 81.600 ;
        RECT 805.050 75.750 806.850 82.500 ;
        RECT 813.150 81.600 817.050 83.700 ;
        RECT 808.950 75.750 810.750 81.600 ;
        RECT 813.150 75.750 814.950 81.600 ;
        RECT 817.650 75.750 819.450 78.600 ;
        RECT 820.650 75.750 822.450 87.600 ;
        RECT 832.650 76.500 834.450 87.600 ;
        RECT 835.650 77.400 837.450 87.600 ;
        RECT 838.650 86.400 846.450 87.300 ;
        RECT 838.650 76.500 840.450 86.400 ;
        RECT 832.650 75.750 840.450 76.500 ;
        RECT 841.650 75.750 843.450 85.500 ;
        RECT 844.650 75.750 846.450 86.400 ;
        RECT 857.400 81.600 858.600 94.050 ;
        RECT 869.100 93.150 870.900 94.950 ;
        RECT 868.950 91.050 871.050 93.150 ;
        RECT 872.550 91.950 873.750 99.300 ;
        RECT 875.100 93.150 876.900 94.950 ;
        RECT 871.950 89.850 874.050 91.950 ;
        RECT 874.950 91.050 877.050 93.150 ;
        RECT 872.550 81.600 873.750 89.850 ;
        RECT 856.650 75.750 858.450 81.600 ;
        RECT 859.650 75.750 861.450 81.600 ;
        RECT 869.550 75.750 871.350 81.600 ;
        RECT 872.550 75.750 874.350 81.600 ;
        RECT 875.550 75.750 877.350 81.600 ;
        RECT 11.400 65.400 13.200 71.250 ;
        RECT 14.700 59.400 16.500 71.250 ;
        RECT 18.900 59.400 20.700 71.250 ;
        RECT 29.550 65.400 31.350 71.250 ;
        RECT 32.550 65.400 34.350 71.250 ;
        RECT 11.250 57.150 13.050 58.950 ;
        RECT 10.950 55.050 13.050 57.150 ;
        RECT 14.850 54.150 16.050 59.400 ;
        RECT 20.100 54.150 21.900 55.950 ;
        RECT 13.950 52.050 16.050 54.150 ;
        RECT 13.950 48.750 15.150 52.050 ;
        RECT 16.950 50.850 19.050 52.950 ;
        RECT 19.950 52.050 22.050 54.150 ;
        RECT 32.400 52.950 33.600 65.400 ;
        RECT 44.550 59.400 46.350 71.250 ;
        RECT 49.050 59.550 50.850 71.250 ;
        RECT 52.050 60.900 53.850 71.250 ;
        RECT 65.550 65.400 67.350 71.250 ;
        RECT 68.550 65.400 70.350 71.250 ;
        RECT 71.550 66.000 73.350 71.250 ;
        RECT 68.700 65.100 70.350 65.400 ;
        RECT 74.550 65.400 76.350 71.250 ;
        RECT 86.550 65.400 88.350 71.250 ;
        RECT 89.550 65.400 91.350 71.250 ;
        RECT 74.550 65.100 75.750 65.400 ;
        RECT 68.700 64.200 75.750 65.100 ;
        RECT 52.050 59.550 54.450 60.900 ;
        RECT 68.100 60.150 69.900 61.950 ;
        RECT 44.550 58.200 45.750 59.400 ;
        RECT 49.950 58.200 51.750 58.650 ;
        RECT 44.550 57.000 51.750 58.200 ;
        RECT 49.950 56.850 51.750 57.000 ;
        RECT 47.100 54.150 48.900 55.950 ;
        RECT 29.100 51.150 30.900 52.950 ;
        RECT 17.100 49.050 18.900 50.850 ;
        RECT 28.950 49.050 31.050 51.150 ;
        RECT 31.950 50.850 34.050 52.950 ;
        RECT 44.100 51.150 45.900 52.950 ;
        RECT 46.950 52.050 49.050 54.150 ;
        RECT 11.250 47.700 15.000 48.750 ;
        RECT 11.250 45.600 12.450 47.700 ;
        RECT 10.650 39.750 12.450 45.600 ;
        RECT 13.650 44.700 21.450 46.050 ;
        RECT 13.650 39.750 15.450 44.700 ;
        RECT 16.650 39.750 18.450 43.800 ;
        RECT 19.650 39.750 21.450 44.700 ;
        RECT 32.400 42.600 33.600 50.850 ;
        RECT 43.950 49.050 46.050 51.150 ;
        RECT 50.700 48.600 51.600 56.850 ;
        RECT 53.100 52.950 54.450 59.550 ;
        RECT 65.100 57.150 66.900 58.950 ;
        RECT 67.950 58.050 70.050 60.150 ;
        RECT 71.250 57.150 73.050 58.950 ;
        RECT 64.950 55.050 67.050 57.150 ;
        RECT 70.950 55.050 73.050 57.150 ;
        RECT 74.700 55.950 75.750 64.200 ;
        RECT 73.950 53.850 76.050 55.950 ;
        RECT 52.950 50.850 55.050 52.950 ;
        RECT 49.950 47.700 51.750 48.600 ;
        RECT 48.450 46.800 51.750 47.700 ;
        RECT 48.450 42.600 49.350 46.800 ;
        RECT 54.000 45.600 55.050 50.850 ;
        RECT 74.400 49.650 75.600 53.850 ;
        RECT 89.400 52.950 90.600 65.400 ;
        RECT 101.550 59.400 103.350 71.250 ;
        RECT 105.750 59.400 107.550 71.250 ;
        RECT 125.400 65.400 127.200 71.250 ;
        RECT 128.700 59.400 130.500 71.250 ;
        RECT 132.900 59.400 134.700 71.250 ;
        RECT 145.650 65.400 147.450 71.250 ;
        RECT 148.650 65.400 150.450 71.250 ;
        RECT 151.650 65.400 153.450 71.250 ;
        RECT 161.550 65.400 163.350 71.250 ;
        RECT 164.550 65.400 166.350 71.250 ;
        RECT 105.000 58.350 107.550 59.400 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 86.100 51.150 87.900 52.950 ;
        RECT 29.550 39.750 31.350 42.600 ;
        RECT 32.550 39.750 34.350 42.600 ;
        RECT 44.550 39.750 46.350 42.600 ;
        RECT 47.550 39.750 49.350 42.600 ;
        RECT 50.550 39.750 52.350 42.600 ;
        RECT 53.550 39.750 55.350 45.600 ;
        RECT 65.700 39.750 67.500 48.600 ;
        RECT 71.100 48.000 75.600 49.650 ;
        RECT 85.950 49.050 88.050 51.150 ;
        RECT 88.950 50.850 91.050 52.950 ;
        RECT 100.950 52.050 103.050 54.150 ;
        RECT 105.000 51.150 106.050 58.350 ;
        RECT 125.250 57.150 127.050 58.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 124.950 55.050 127.050 57.150 ;
        RECT 128.850 54.150 130.050 59.400 ;
        RECT 149.250 57.150 150.450 65.400 ;
        RECT 134.100 54.150 135.900 55.950 ;
        RECT 106.950 52.050 109.050 54.150 ;
        RECT 127.950 52.050 130.050 54.150 ;
        RECT 71.100 39.750 72.900 48.000 ;
        RECT 89.400 42.600 90.600 50.850 ;
        RECT 103.950 49.050 106.050 51.150 ;
        RECT 105.000 42.600 106.050 49.050 ;
        RECT 127.950 48.750 129.150 52.050 ;
        RECT 130.950 50.850 133.050 52.950 ;
        RECT 133.950 52.050 136.050 54.150 ;
        RECT 145.950 53.850 148.050 55.950 ;
        RECT 148.950 55.050 151.050 57.150 ;
        RECT 146.100 52.050 147.900 53.850 ;
        RECT 131.100 49.050 132.900 50.850 ;
        RECT 125.250 47.700 129.000 48.750 ;
        RECT 149.250 47.700 150.450 55.050 ;
        RECT 151.950 53.850 154.050 55.950 ;
        RECT 161.100 54.150 162.900 55.950 ;
        RECT 152.100 52.050 153.900 53.850 ;
        RECT 160.950 52.050 163.050 54.150 ;
        RECT 164.700 48.300 165.900 65.400 ;
        RECT 168.150 59.400 169.950 71.250 ;
        RECT 171.150 59.400 172.950 71.250 ;
        RECT 187.650 65.400 189.450 71.250 ;
        RECT 190.650 65.400 192.450 71.250 ;
        RECT 200.550 65.400 202.350 71.250 ;
        RECT 203.550 65.400 205.350 71.250 ;
        RECT 166.950 53.850 169.050 55.950 ;
        RECT 171.150 54.150 172.350 59.400 ;
        RECT 167.100 52.050 168.900 53.850 ;
        RECT 169.950 52.050 172.350 54.150 ;
        RECT 188.400 52.950 189.600 65.400 ;
        RECT 203.400 52.950 204.600 65.400 ;
        RECT 217.650 59.400 219.450 71.250 ;
        RECT 220.650 60.300 222.450 71.250 ;
        RECT 223.650 61.200 225.450 71.250 ;
        RECT 226.650 60.300 228.450 71.250 ;
        RECT 220.650 59.400 228.450 60.300 ;
        RECT 237.300 59.400 239.100 71.250 ;
        RECT 241.500 59.400 243.300 71.250 ;
        RECT 244.800 65.400 246.600 71.250 ;
        RECT 261.300 59.400 263.100 71.250 ;
        RECT 265.500 59.400 267.300 71.250 ;
        RECT 268.800 65.400 270.600 71.250 ;
        RECT 284.550 59.400 286.350 71.250 ;
        RECT 289.050 59.550 290.850 71.250 ;
        RECT 292.050 60.900 293.850 71.250 ;
        RECT 308.550 65.400 310.350 71.250 ;
        RECT 311.550 65.400 313.350 71.250 ;
        RECT 314.550 66.000 316.350 71.250 ;
        RECT 311.700 65.100 313.350 65.400 ;
        RECT 317.550 65.400 319.350 71.250 ;
        RECT 329.550 65.400 331.350 71.250 ;
        RECT 332.550 65.400 334.350 71.250 ;
        RECT 335.550 66.000 337.350 71.250 ;
        RECT 317.550 65.100 318.750 65.400 ;
        RECT 311.700 64.200 318.750 65.100 ;
        RECT 332.700 65.100 334.350 65.400 ;
        RECT 338.550 65.400 340.350 71.250 ;
        RECT 353.550 65.400 355.350 71.250 ;
        RECT 356.550 65.400 358.350 71.250 ;
        RECT 359.550 65.400 361.350 71.250 ;
        RECT 374.550 65.400 376.350 71.250 ;
        RECT 377.550 65.400 379.350 71.250 ;
        RECT 380.550 65.400 382.350 71.250 ;
        RECT 397.650 65.400 399.450 71.250 ;
        RECT 400.650 66.000 402.450 71.250 ;
        RECT 338.550 65.100 339.750 65.400 ;
        RECT 332.700 64.200 339.750 65.100 ;
        RECT 292.050 59.550 294.450 60.900 ;
        RECT 311.100 60.150 312.900 61.950 ;
        RECT 218.100 54.150 219.300 59.400 ;
        RECT 236.100 54.150 237.900 55.950 ;
        RECT 241.950 54.150 243.150 59.400 ;
        RECT 244.950 57.150 246.750 58.950 ;
        RECT 244.950 55.050 247.050 57.150 ;
        RECT 260.100 54.150 261.900 55.950 ;
        RECT 265.950 54.150 267.150 59.400 ;
        RECT 268.950 57.150 270.750 58.950 ;
        RECT 284.550 58.200 285.750 59.400 ;
        RECT 289.950 58.200 291.750 58.650 ;
        RECT 268.950 55.050 271.050 57.150 ;
        RECT 284.550 57.000 291.750 58.200 ;
        RECT 289.950 56.850 291.750 57.000 ;
        RECT 287.100 54.150 288.900 55.950 ;
        RECT 125.250 45.600 126.450 47.700 ;
        RECT 146.850 46.800 150.450 47.700 ;
        RECT 161.550 47.100 169.050 48.300 ;
        RECT 86.550 39.750 88.350 42.600 ;
        RECT 89.550 39.750 91.350 42.600 ;
        RECT 101.550 39.750 103.350 42.600 ;
        RECT 104.550 39.750 106.350 42.600 ;
        RECT 107.550 39.750 109.350 42.600 ;
        RECT 124.650 39.750 126.450 45.600 ;
        RECT 127.650 44.700 135.450 46.050 ;
        RECT 127.650 39.750 129.450 44.700 ;
        RECT 130.650 39.750 132.450 43.800 ;
        RECT 133.650 39.750 135.450 44.700 ;
        RECT 146.850 39.750 148.650 46.800 ;
        RECT 151.350 39.750 153.150 45.600 ;
        RECT 161.550 39.750 163.350 47.100 ;
        RECT 167.250 46.500 169.050 47.100 ;
        RECT 171.150 45.600 172.350 52.050 ;
        RECT 187.950 50.850 190.050 52.950 ;
        RECT 191.100 51.150 192.900 52.950 ;
        RECT 200.100 51.150 201.900 52.950 ;
        RECT 166.050 39.750 167.850 45.600 ;
        RECT 169.050 44.100 172.350 45.600 ;
        RECT 169.050 39.750 170.850 44.100 ;
        RECT 188.400 42.600 189.600 50.850 ;
        RECT 190.950 49.050 193.050 51.150 ;
        RECT 199.950 49.050 202.050 51.150 ;
        RECT 202.950 50.850 205.050 52.950 ;
        RECT 217.950 52.050 220.050 54.150 ;
        RECT 203.400 42.600 204.600 50.850 ;
        RECT 218.100 45.600 219.300 52.050 ;
        RECT 220.950 50.850 223.050 52.950 ;
        RECT 224.100 51.150 225.900 52.950 ;
        RECT 221.100 49.050 222.900 50.850 ;
        RECT 223.950 49.050 226.050 51.150 ;
        RECT 226.950 50.850 229.050 52.950 ;
        RECT 235.950 52.050 238.050 54.150 ;
        RECT 238.950 50.850 241.050 52.950 ;
        RECT 241.950 52.050 244.050 54.150 ;
        RECT 259.950 52.050 262.050 54.150 ;
        RECT 227.100 49.050 228.900 50.850 ;
        RECT 239.100 49.050 240.900 50.850 ;
        RECT 242.850 48.750 244.050 52.050 ;
        RECT 262.950 50.850 265.050 52.950 ;
        RECT 265.950 52.050 268.050 54.150 ;
        RECT 263.100 49.050 264.900 50.850 ;
        RECT 266.850 48.750 268.050 52.050 ;
        RECT 284.100 51.150 285.900 52.950 ;
        RECT 286.950 52.050 289.050 54.150 ;
        RECT 283.950 49.050 286.050 51.150 ;
        RECT 243.000 47.700 246.750 48.750 ;
        RECT 267.000 47.700 270.750 48.750 ;
        RECT 290.700 48.600 291.600 56.850 ;
        RECT 293.100 52.950 294.450 59.550 ;
        RECT 308.100 57.150 309.900 58.950 ;
        RECT 310.950 58.050 313.050 60.150 ;
        RECT 314.250 57.150 316.050 58.950 ;
        RECT 307.950 55.050 310.050 57.150 ;
        RECT 313.950 55.050 316.050 57.150 ;
        RECT 317.700 55.950 318.750 64.200 ;
        RECT 332.100 60.150 333.900 61.950 ;
        RECT 329.100 57.150 330.900 58.950 ;
        RECT 331.950 58.050 334.050 60.150 ;
        RECT 335.250 57.150 337.050 58.950 ;
        RECT 316.950 53.850 319.050 55.950 ;
        RECT 328.950 55.050 331.050 57.150 ;
        RECT 334.950 55.050 337.050 57.150 ;
        RECT 338.700 55.950 339.750 64.200 ;
        RECT 356.550 57.150 357.750 65.400 ;
        RECT 377.550 57.150 378.750 65.400 ;
        RECT 398.250 65.100 399.450 65.400 ;
        RECT 403.650 65.400 405.450 71.250 ;
        RECT 406.650 65.400 408.450 71.250 ;
        RECT 403.650 65.100 405.300 65.400 ;
        RECT 398.250 64.200 405.300 65.100 ;
        RECT 337.950 53.850 340.050 55.950 ;
        RECT 352.950 53.850 355.050 55.950 ;
        RECT 355.950 55.050 358.050 57.150 ;
        RECT 292.950 50.850 295.050 52.950 ;
        RECT 289.950 47.700 291.750 48.600 ;
        RECT 218.100 43.950 223.800 45.600 ;
        RECT 187.650 39.750 189.450 42.600 ;
        RECT 190.650 39.750 192.450 42.600 ;
        RECT 200.550 39.750 202.350 42.600 ;
        RECT 203.550 39.750 205.350 42.600 ;
        RECT 218.700 39.750 220.500 42.600 ;
        RECT 222.000 39.750 223.800 43.950 ;
        RECT 226.200 39.750 228.000 45.600 ;
        RECT 236.550 44.700 244.350 46.050 ;
        RECT 236.550 39.750 238.350 44.700 ;
        RECT 239.550 39.750 241.350 43.800 ;
        RECT 242.550 39.750 244.350 44.700 ;
        RECT 245.550 45.600 246.750 47.700 ;
        RECT 245.550 39.750 247.350 45.600 ;
        RECT 260.550 44.700 268.350 46.050 ;
        RECT 260.550 39.750 262.350 44.700 ;
        RECT 263.550 39.750 265.350 43.800 ;
        RECT 266.550 39.750 268.350 44.700 ;
        RECT 269.550 45.600 270.750 47.700 ;
        RECT 288.450 46.800 291.750 47.700 ;
        RECT 269.550 39.750 271.350 45.600 ;
        RECT 288.450 42.600 289.350 46.800 ;
        RECT 294.000 45.600 295.050 50.850 ;
        RECT 317.400 49.650 318.600 53.850 ;
        RECT 338.400 49.650 339.600 53.850 ;
        RECT 353.100 52.050 354.900 53.850 ;
        RECT 284.550 39.750 286.350 42.600 ;
        RECT 287.550 39.750 289.350 42.600 ;
        RECT 290.550 39.750 292.350 42.600 ;
        RECT 293.550 39.750 295.350 45.600 ;
        RECT 308.700 39.750 310.500 48.600 ;
        RECT 314.100 48.000 318.600 49.650 ;
        RECT 314.100 39.750 315.900 48.000 ;
        RECT 329.700 39.750 331.500 48.600 ;
        RECT 335.100 48.000 339.600 49.650 ;
        RECT 335.100 39.750 336.900 48.000 ;
        RECT 356.550 47.700 357.750 55.050 ;
        RECT 358.950 53.850 361.050 55.950 ;
        RECT 373.950 53.850 376.050 55.950 ;
        RECT 376.950 55.050 379.050 57.150 ;
        RECT 398.250 55.950 399.300 64.200 ;
        RECT 404.100 60.150 405.900 61.950 ;
        RECT 416.550 60.300 418.350 71.250 ;
        RECT 419.550 61.200 421.350 71.250 ;
        RECT 422.550 60.300 424.350 71.250 ;
        RECT 400.950 57.150 402.750 58.950 ;
        RECT 403.950 58.050 406.050 60.150 ;
        RECT 416.550 59.400 424.350 60.300 ;
        RECT 425.550 59.400 427.350 71.250 ;
        RECT 437.550 60.300 439.350 71.250 ;
        RECT 440.550 61.200 442.350 71.250 ;
        RECT 443.550 60.300 445.350 71.250 ;
        RECT 437.550 59.400 445.350 60.300 ;
        RECT 446.550 59.400 448.350 71.250 ;
        RECT 461.550 65.400 463.350 71.250 ;
        RECT 464.550 65.400 466.350 71.250 ;
        RECT 467.550 66.000 469.350 71.250 ;
        RECT 464.700 65.100 466.350 65.400 ;
        RECT 470.550 65.400 472.350 71.250 ;
        RECT 482.550 65.400 484.350 71.250 ;
        RECT 485.550 65.400 487.350 71.250 ;
        RECT 470.550 65.100 471.750 65.400 ;
        RECT 464.700 64.200 471.750 65.100 ;
        RECT 464.100 60.150 465.900 61.950 ;
        RECT 407.100 57.150 408.900 58.950 ;
        RECT 409.950 57.450 412.050 58.050 ;
        RECT 421.950 57.450 424.050 58.050 ;
        RECT 359.100 52.050 360.900 53.850 ;
        RECT 374.100 52.050 375.900 53.850 ;
        RECT 377.550 47.700 378.750 55.050 ;
        RECT 379.950 53.850 382.050 55.950 ;
        RECT 397.950 53.850 400.050 55.950 ;
        RECT 400.950 55.050 403.050 57.150 ;
        RECT 406.950 55.050 409.050 57.150 ;
        RECT 409.950 56.550 424.050 57.450 ;
        RECT 409.950 55.950 412.050 56.550 ;
        RECT 421.950 55.950 424.050 56.550 ;
        RECT 425.700 54.150 426.900 59.400 ;
        RECT 446.700 54.150 447.900 59.400 ;
        RECT 461.100 57.150 462.900 58.950 ;
        RECT 463.950 58.050 466.050 60.150 ;
        RECT 467.250 57.150 469.050 58.950 ;
        RECT 460.950 55.050 463.050 57.150 ;
        RECT 466.950 55.050 469.050 57.150 ;
        RECT 470.700 55.950 471.750 64.200 ;
        RECT 380.100 52.050 381.900 53.850 ;
        RECT 398.400 49.650 399.600 53.850 ;
        RECT 415.950 50.850 418.050 52.950 ;
        RECT 419.100 51.150 420.900 52.950 ;
        RECT 398.400 48.000 402.900 49.650 ;
        RECT 416.100 49.050 417.900 50.850 ;
        RECT 418.950 49.050 421.050 51.150 ;
        RECT 421.950 50.850 424.050 52.950 ;
        RECT 424.950 52.050 427.050 54.150 ;
        RECT 422.100 49.050 423.900 50.850 ;
        RECT 356.550 46.800 360.150 47.700 ;
        RECT 377.550 46.800 381.150 47.700 ;
        RECT 353.850 39.750 355.650 45.600 ;
        RECT 358.350 39.750 360.150 46.800 ;
        RECT 374.850 39.750 376.650 45.600 ;
        RECT 379.350 39.750 381.150 46.800 ;
        RECT 401.100 39.750 402.900 48.000 ;
        RECT 406.500 39.750 408.300 48.600 ;
        RECT 425.700 45.600 426.900 52.050 ;
        RECT 436.950 50.850 439.050 52.950 ;
        RECT 440.100 51.150 441.900 52.950 ;
        RECT 437.100 49.050 438.900 50.850 ;
        RECT 439.950 49.050 442.050 51.150 ;
        RECT 442.950 50.850 445.050 52.950 ;
        RECT 445.950 52.050 448.050 54.150 ;
        RECT 469.950 53.850 472.050 55.950 ;
        RECT 482.100 54.150 483.900 55.950 ;
        RECT 443.100 49.050 444.900 50.850 ;
        RECT 446.700 45.600 447.900 52.050 ;
        RECT 470.400 49.650 471.600 53.850 ;
        RECT 481.950 52.050 484.050 54.150 ;
        RECT 417.000 39.750 418.800 45.600 ;
        RECT 421.200 43.950 426.900 45.600 ;
        RECT 421.200 39.750 423.000 43.950 ;
        RECT 424.500 39.750 426.300 42.600 ;
        RECT 438.000 39.750 439.800 45.600 ;
        RECT 442.200 43.950 447.900 45.600 ;
        RECT 442.200 39.750 444.000 43.950 ;
        RECT 445.500 39.750 447.300 42.600 ;
        RECT 461.700 39.750 463.500 48.600 ;
        RECT 467.100 48.000 471.600 49.650 ;
        RECT 485.700 48.300 486.900 65.400 ;
        RECT 489.150 59.400 490.950 71.250 ;
        RECT 492.150 59.400 493.950 71.250 ;
        RECT 503.550 65.400 505.350 71.250 ;
        RECT 506.550 65.400 508.350 71.250 ;
        RECT 509.550 66.000 511.350 71.250 ;
        RECT 506.700 65.100 508.350 65.400 ;
        RECT 512.550 65.400 514.350 71.250 ;
        RECT 530.400 65.400 532.200 71.250 ;
        RECT 512.550 65.100 513.750 65.400 ;
        RECT 506.700 64.200 513.750 65.100 ;
        RECT 506.100 60.150 507.900 61.950 ;
        RECT 487.950 53.850 490.050 55.950 ;
        RECT 492.150 54.150 493.350 59.400 ;
        RECT 503.100 57.150 504.900 58.950 ;
        RECT 505.950 58.050 508.050 60.150 ;
        RECT 509.250 57.150 511.050 58.950 ;
        RECT 502.950 55.050 505.050 57.150 ;
        RECT 508.950 55.050 511.050 57.150 ;
        RECT 512.700 55.950 513.750 64.200 ;
        RECT 533.700 59.400 535.500 71.250 ;
        RECT 537.900 59.400 539.700 71.250 ;
        RECT 550.650 59.400 552.450 71.250 ;
        RECT 553.650 60.300 555.450 71.250 ;
        RECT 556.650 61.200 558.450 71.250 ;
        RECT 559.650 60.300 561.450 71.250 ;
        RECT 571.050 70.500 578.850 71.250 ;
        RECT 571.050 61.200 572.850 70.500 ;
        RECT 574.050 61.800 575.850 69.600 ;
        RECT 553.650 59.400 561.450 60.300 ;
        RECT 574.650 59.400 575.850 61.800 ;
        RECT 577.050 61.800 578.850 70.500 ;
        RECT 580.650 70.500 588.450 71.250 ;
        RECT 580.650 62.700 582.450 70.500 ;
        RECT 583.650 61.800 585.450 69.600 ;
        RECT 577.050 60.900 585.450 61.800 ;
        RECT 586.650 61.500 588.450 70.500 ;
        RECT 589.650 62.400 591.450 71.250 ;
        RECT 592.650 61.500 594.450 71.250 ;
        RECT 604.650 65.400 606.450 71.250 ;
        RECT 607.650 65.400 609.450 71.250 ;
        RECT 610.650 65.400 612.450 71.250 ;
        RECT 626.400 65.400 628.200 71.250 ;
        RECT 586.650 60.600 594.450 61.500 ;
        RECT 530.250 57.150 532.050 58.950 ;
        RECT 488.100 52.050 489.900 53.850 ;
        RECT 490.950 52.050 493.350 54.150 ;
        RECT 511.950 53.850 514.050 55.950 ;
        RECT 529.950 55.050 532.050 57.150 ;
        RECT 533.850 54.150 535.050 59.400 ;
        RECT 539.100 54.150 540.900 55.950 ;
        RECT 551.100 54.150 552.300 59.400 ;
        RECT 574.650 58.200 578.100 59.400 ;
        RECT 467.100 39.750 468.900 48.000 ;
        RECT 482.550 47.100 490.050 48.300 ;
        RECT 482.550 39.750 484.350 47.100 ;
        RECT 488.250 46.500 490.050 47.100 ;
        RECT 492.150 45.600 493.350 52.050 ;
        RECT 512.400 49.650 513.600 53.850 ;
        RECT 487.050 39.750 488.850 45.600 ;
        RECT 490.050 44.100 493.350 45.600 ;
        RECT 490.050 39.750 491.850 44.100 ;
        RECT 503.700 39.750 505.500 48.600 ;
        RECT 509.100 48.000 513.600 49.650 ;
        RECT 532.950 52.050 535.050 54.150 ;
        RECT 532.950 48.750 534.150 52.050 ;
        RECT 535.950 50.850 538.050 52.950 ;
        RECT 538.950 52.050 541.050 54.150 ;
        RECT 550.950 52.050 553.050 54.150 ;
        RECT 576.900 52.950 578.100 58.200 ;
        RECT 608.250 57.150 609.450 65.400 ;
        RECT 629.700 59.400 631.500 71.250 ;
        RECT 633.900 59.400 635.700 71.250 ;
        RECT 647.550 65.400 649.350 71.250 ;
        RECT 650.550 65.400 652.350 71.250 ;
        RECT 653.550 65.400 655.350 71.250 ;
        RECT 626.250 57.150 628.050 58.950 ;
        RECT 581.100 54.150 582.900 55.950 ;
        RECT 590.100 54.150 591.900 55.950 ;
        RECT 536.100 49.050 537.900 50.850 ;
        RECT 509.100 39.750 510.900 48.000 ;
        RECT 530.250 47.700 534.000 48.750 ;
        RECT 530.250 45.600 531.450 47.700 ;
        RECT 529.650 39.750 531.450 45.600 ;
        RECT 532.650 44.700 540.450 46.050 ;
        RECT 532.650 39.750 534.450 44.700 ;
        RECT 535.650 39.750 537.450 43.800 ;
        RECT 538.650 39.750 540.450 44.700 ;
        RECT 551.100 45.600 552.300 52.050 ;
        RECT 553.950 50.850 556.050 52.950 ;
        RECT 557.100 51.150 558.900 52.950 ;
        RECT 554.100 49.050 555.900 50.850 ;
        RECT 556.950 49.050 559.050 51.150 ;
        RECT 559.950 50.850 562.050 52.950 ;
        RECT 574.950 50.850 578.100 52.950 ;
        RECT 580.950 52.050 583.050 54.150 ;
        RECT 583.950 50.850 586.050 52.950 ;
        RECT 589.950 52.050 592.050 54.150 ;
        RECT 604.950 53.850 607.050 55.950 ;
        RECT 607.950 55.050 610.050 57.150 ;
        RECT 605.100 52.050 606.900 53.850 ;
        RECT 560.100 49.050 561.900 50.850 ;
        RECT 551.100 43.950 556.800 45.600 ;
        RECT 551.700 39.750 553.500 42.600 ;
        RECT 555.000 39.750 556.800 43.950 ;
        RECT 559.200 39.750 561.000 45.600 ;
        RECT 576.900 44.400 578.100 50.850 ;
        RECT 584.100 49.050 585.900 50.850 ;
        RECT 608.250 47.700 609.450 55.050 ;
        RECT 610.950 53.850 613.050 55.950 ;
        RECT 625.950 55.050 628.050 57.150 ;
        RECT 629.850 54.150 631.050 59.400 ;
        RECT 650.550 57.150 651.750 65.400 ;
        RECT 665.550 60.300 667.350 71.250 ;
        RECT 668.550 61.200 670.350 71.250 ;
        RECT 671.550 60.300 673.350 71.250 ;
        RECT 665.550 59.400 673.350 60.300 ;
        RECT 674.550 59.400 676.350 71.250 ;
        RECT 689.400 65.400 691.200 71.250 ;
        RECT 692.700 59.400 694.500 71.250 ;
        RECT 696.900 59.400 698.700 71.250 ;
        RECT 709.650 59.400 711.450 71.250 ;
        RECT 712.650 60.300 714.450 71.250 ;
        RECT 715.650 61.200 717.450 71.250 ;
        RECT 718.650 60.300 720.450 71.250 ;
        RECT 731.550 65.400 733.350 71.250 ;
        RECT 734.550 65.400 736.350 71.250 ;
        RECT 712.650 59.400 720.450 60.300 ;
        RECT 635.100 54.150 636.900 55.950 ;
        RECT 611.100 52.050 612.900 53.850 ;
        RECT 628.950 52.050 631.050 54.150 ;
        RECT 628.950 48.750 630.150 52.050 ;
        RECT 631.950 50.850 634.050 52.950 ;
        RECT 634.950 52.050 637.050 54.150 ;
        RECT 646.950 53.850 649.050 55.950 ;
        RECT 649.950 55.050 652.050 57.150 ;
        RECT 647.100 52.050 648.900 53.850 ;
        RECT 632.100 49.050 633.900 50.850 ;
        RECT 605.850 46.800 609.450 47.700 ;
        RECT 626.250 47.700 630.000 48.750 ;
        RECT 650.550 47.700 651.750 55.050 ;
        RECT 652.950 53.850 655.050 55.950 ;
        RECT 674.700 54.150 675.900 59.400 ;
        RECT 689.250 57.150 691.050 58.950 ;
        RECT 688.950 55.050 691.050 57.150 ;
        RECT 692.850 54.150 694.050 59.400 ;
        RECT 698.100 54.150 699.900 55.950 ;
        RECT 710.100 54.150 711.300 59.400 ;
        RECT 731.100 54.150 732.900 55.950 ;
        RECT 653.100 52.050 654.900 53.850 ;
        RECT 664.950 50.850 667.050 52.950 ;
        RECT 668.100 51.150 669.900 52.950 ;
        RECT 665.100 49.050 666.900 50.850 ;
        RECT 667.950 49.050 670.050 51.150 ;
        RECT 670.950 50.850 673.050 52.950 ;
        RECT 673.950 52.050 676.050 54.150 ;
        RECT 691.950 52.050 694.050 54.150 ;
        RECT 671.100 49.050 672.900 50.850 ;
        RECT 576.900 43.500 587.700 44.400 ;
        RECT 580.650 42.600 581.700 43.500 ;
        RECT 586.650 42.600 587.700 43.500 ;
        RECT 580.650 39.750 582.450 42.600 ;
        RECT 583.650 39.750 585.450 42.600 ;
        RECT 586.650 39.750 588.450 42.600 ;
        RECT 589.650 39.750 591.750 42.600 ;
        RECT 605.850 39.750 607.650 46.800 ;
        RECT 626.250 45.600 627.450 47.700 ;
        RECT 650.550 46.800 654.150 47.700 ;
        RECT 610.350 39.750 612.150 45.600 ;
        RECT 625.650 39.750 627.450 45.600 ;
        RECT 628.650 44.700 636.450 46.050 ;
        RECT 628.650 39.750 630.450 44.700 ;
        RECT 631.650 39.750 633.450 43.800 ;
        RECT 634.650 39.750 636.450 44.700 ;
        RECT 647.850 39.750 649.650 45.600 ;
        RECT 652.350 39.750 654.150 46.800 ;
        RECT 674.700 45.600 675.900 52.050 ;
        RECT 691.950 48.750 693.150 52.050 ;
        RECT 694.950 50.850 697.050 52.950 ;
        RECT 697.950 52.050 700.050 54.150 ;
        RECT 709.950 52.050 712.050 54.150 ;
        RECT 695.100 49.050 696.900 50.850 ;
        RECT 689.250 47.700 693.000 48.750 ;
        RECT 689.250 45.600 690.450 47.700 ;
        RECT 666.000 39.750 667.800 45.600 ;
        RECT 670.200 43.950 675.900 45.600 ;
        RECT 670.200 39.750 672.000 43.950 ;
        RECT 673.500 39.750 675.300 42.600 ;
        RECT 688.650 39.750 690.450 45.600 ;
        RECT 691.650 44.700 699.450 46.050 ;
        RECT 691.650 39.750 693.450 44.700 ;
        RECT 694.650 39.750 696.450 43.800 ;
        RECT 697.650 39.750 699.450 44.700 ;
        RECT 710.100 45.600 711.300 52.050 ;
        RECT 712.950 50.850 715.050 52.950 ;
        RECT 716.100 51.150 717.900 52.950 ;
        RECT 713.100 49.050 714.900 50.850 ;
        RECT 715.950 49.050 718.050 51.150 ;
        RECT 718.950 50.850 721.050 52.950 ;
        RECT 730.950 52.050 733.050 54.150 ;
        RECT 719.100 49.050 720.900 50.850 ;
        RECT 734.700 48.300 735.900 65.400 ;
        RECT 738.150 59.400 739.950 71.250 ;
        RECT 741.150 59.400 742.950 71.250 ;
        RECT 752.550 65.400 754.350 71.250 ;
        RECT 755.550 65.400 757.350 71.250 ;
        RECT 758.550 65.400 760.350 71.250 ;
        RECT 736.950 53.850 739.050 55.950 ;
        RECT 741.150 54.150 742.350 59.400 ;
        RECT 755.550 57.150 756.750 65.400 ;
        RECT 770.550 59.400 772.350 71.250 ;
        RECT 774.750 59.400 776.550 71.250 ;
        RECT 791.550 65.400 793.350 71.250 ;
        RECT 794.550 65.400 796.350 71.250 ;
        RECT 806.550 65.400 808.350 71.250 ;
        RECT 809.550 65.400 811.350 71.250 ;
        RECT 812.550 65.400 814.350 71.250 ;
        RECT 774.000 58.350 776.550 59.400 ;
        RECT 737.100 52.050 738.900 53.850 ;
        RECT 739.950 52.050 742.350 54.150 ;
        RECT 751.950 53.850 754.050 55.950 ;
        RECT 754.950 55.050 757.050 57.150 ;
        RECT 752.100 52.050 753.900 53.850 ;
        RECT 731.550 47.100 739.050 48.300 ;
        RECT 710.100 43.950 715.800 45.600 ;
        RECT 710.700 39.750 712.500 42.600 ;
        RECT 714.000 39.750 715.800 43.950 ;
        RECT 718.200 39.750 720.000 45.600 ;
        RECT 731.550 39.750 733.350 47.100 ;
        RECT 737.250 46.500 739.050 47.100 ;
        RECT 741.150 45.600 742.350 52.050 ;
        RECT 755.550 47.700 756.750 55.050 ;
        RECT 757.950 53.850 760.050 55.950 ;
        RECT 770.100 54.150 771.900 55.950 ;
        RECT 758.100 52.050 759.900 53.850 ;
        RECT 769.950 52.050 772.050 54.150 ;
        RECT 774.000 51.150 775.050 58.350 ;
        RECT 776.100 54.150 777.900 55.950 ;
        RECT 775.950 52.050 778.050 54.150 ;
        RECT 794.400 52.950 795.600 65.400 ;
        RECT 809.550 57.150 810.750 65.400 ;
        RECT 824.550 60.300 826.350 71.250 ;
        RECT 827.550 61.200 829.350 71.250 ;
        RECT 830.550 60.300 832.350 71.250 ;
        RECT 824.550 59.400 832.350 60.300 ;
        RECT 833.550 59.400 835.350 71.250 ;
        RECT 849.300 59.400 851.100 71.250 ;
        RECT 853.500 59.400 855.300 71.250 ;
        RECT 856.800 65.400 858.600 71.250 ;
        RECT 872.550 65.400 874.350 71.250 ;
        RECT 875.550 65.400 877.350 71.250 ;
        RECT 805.950 53.850 808.050 55.950 ;
        RECT 808.950 55.050 811.050 57.150 ;
        RECT 791.100 51.150 792.900 52.950 ;
        RECT 772.950 49.050 775.050 51.150 ;
        RECT 790.950 49.050 793.050 51.150 ;
        RECT 793.950 50.850 796.050 52.950 ;
        RECT 806.100 52.050 807.900 53.850 ;
        RECT 755.550 46.800 759.150 47.700 ;
        RECT 736.050 39.750 737.850 45.600 ;
        RECT 739.050 44.100 742.350 45.600 ;
        RECT 739.050 39.750 740.850 44.100 ;
        RECT 752.850 39.750 754.650 45.600 ;
        RECT 757.350 39.750 759.150 46.800 ;
        RECT 774.000 42.600 775.050 49.050 ;
        RECT 794.400 42.600 795.600 50.850 ;
        RECT 809.550 47.700 810.750 55.050 ;
        RECT 811.950 53.850 814.050 55.950 ;
        RECT 833.700 54.150 834.900 59.400 ;
        RECT 848.100 54.150 849.900 55.950 ;
        RECT 853.950 54.150 855.150 59.400 ;
        RECT 856.950 57.150 858.750 58.950 ;
        RECT 856.950 55.050 859.050 57.150 ;
        RECT 812.100 52.050 813.900 53.850 ;
        RECT 823.950 50.850 826.050 52.950 ;
        RECT 827.100 51.150 828.900 52.950 ;
        RECT 824.100 49.050 825.900 50.850 ;
        RECT 826.950 49.050 829.050 51.150 ;
        RECT 829.950 50.850 832.050 52.950 ;
        RECT 832.950 52.050 835.050 54.150 ;
        RECT 847.950 52.050 850.050 54.150 ;
        RECT 830.100 49.050 831.900 50.850 ;
        RECT 809.550 46.800 813.150 47.700 ;
        RECT 770.550 39.750 772.350 42.600 ;
        RECT 773.550 39.750 775.350 42.600 ;
        RECT 776.550 39.750 778.350 42.600 ;
        RECT 791.550 39.750 793.350 42.600 ;
        RECT 794.550 39.750 796.350 42.600 ;
        RECT 806.850 39.750 808.650 45.600 ;
        RECT 811.350 39.750 813.150 46.800 ;
        RECT 833.700 45.600 834.900 52.050 ;
        RECT 850.950 50.850 853.050 52.950 ;
        RECT 853.950 52.050 856.050 54.150 ;
        RECT 875.400 52.950 876.600 65.400 ;
        RECT 851.100 49.050 852.900 50.850 ;
        RECT 854.850 48.750 856.050 52.050 ;
        RECT 872.100 51.150 873.900 52.950 ;
        RECT 871.950 49.050 874.050 51.150 ;
        RECT 874.950 50.850 877.050 52.950 ;
        RECT 855.000 47.700 858.750 48.750 ;
        RECT 825.000 39.750 826.800 45.600 ;
        RECT 829.200 43.950 834.900 45.600 ;
        RECT 848.550 44.700 856.350 46.050 ;
        RECT 829.200 39.750 831.000 43.950 ;
        RECT 832.500 39.750 834.300 42.600 ;
        RECT 848.550 39.750 850.350 44.700 ;
        RECT 851.550 39.750 853.350 43.800 ;
        RECT 854.550 39.750 856.350 44.700 ;
        RECT 857.550 45.600 858.750 47.700 ;
        RECT 857.550 39.750 859.350 45.600 ;
        RECT 875.400 42.600 876.600 50.850 ;
        RECT 872.550 39.750 874.350 42.600 ;
        RECT 875.550 39.750 877.350 42.600 ;
        RECT 13.650 32.400 15.450 35.250 ;
        RECT 16.650 32.400 18.450 35.250 ;
        RECT 19.650 32.400 21.450 35.250 ;
        RECT 31.650 32.400 33.450 35.250 ;
        RECT 34.650 32.400 36.450 35.250 ;
        RECT 16.950 25.950 18.000 32.400 ;
        RECT 16.950 23.850 19.050 25.950 ;
        RECT 32.400 24.150 33.600 32.400 ;
        RECT 49.650 29.400 51.450 35.250 ;
        RECT 50.250 27.300 51.450 29.400 ;
        RECT 52.650 30.300 54.450 35.250 ;
        RECT 55.650 31.200 57.450 35.250 ;
        RECT 58.650 30.300 60.450 35.250 ;
        RECT 52.650 28.950 60.450 30.300 ;
        RECT 72.000 29.400 73.800 35.250 ;
        RECT 76.200 31.050 78.000 35.250 ;
        RECT 79.500 32.400 81.300 35.250 ;
        RECT 76.200 29.400 81.900 31.050 ;
        RECT 50.250 26.250 54.000 27.300 ;
        RECT 13.950 20.850 16.050 22.950 ;
        RECT 14.100 19.050 15.900 20.850 ;
        RECT 16.950 16.650 18.000 23.850 ;
        RECT 19.950 20.850 22.050 22.950 ;
        RECT 31.950 22.050 34.050 24.150 ;
        RECT 34.950 23.850 37.050 25.950 ;
        RECT 35.100 22.050 36.900 23.850 ;
        RECT 52.950 22.950 54.150 26.250 ;
        RECT 56.100 24.150 57.900 25.950 ;
        RECT 71.100 24.150 72.900 25.950 ;
        RECT 20.100 19.050 21.900 20.850 ;
        RECT 15.450 15.600 18.000 16.650 ;
        RECT 15.450 3.750 17.250 15.600 ;
        RECT 19.650 3.750 21.450 15.600 ;
        RECT 32.400 9.600 33.600 22.050 ;
        RECT 52.950 20.850 55.050 22.950 ;
        RECT 55.950 22.050 58.050 24.150 ;
        RECT 58.950 20.850 61.050 22.950 ;
        RECT 70.950 22.050 73.050 24.150 ;
        RECT 73.950 23.850 76.050 25.950 ;
        RECT 77.100 24.150 78.900 25.950 ;
        RECT 74.100 22.050 75.900 23.850 ;
        RECT 76.950 22.050 79.050 24.150 ;
        RECT 80.700 22.950 81.900 29.400 ;
        RECT 95.550 30.300 97.350 35.250 ;
        RECT 98.550 31.200 100.350 35.250 ;
        RECT 101.550 30.300 103.350 35.250 ;
        RECT 95.550 28.950 103.350 30.300 ;
        RECT 104.550 29.400 106.350 35.250 ;
        RECT 104.550 27.300 105.750 29.400 ;
        RECT 102.000 26.250 105.750 27.300 ;
        RECT 119.700 26.400 121.500 35.250 ;
        RECT 125.100 27.000 126.900 35.250 ;
        RECT 98.100 24.150 99.900 25.950 ;
        RECT 79.950 20.850 82.050 22.950 ;
        RECT 94.950 20.850 97.050 22.950 ;
        RECT 97.950 22.050 100.050 24.150 ;
        RECT 101.850 22.950 103.050 26.250 ;
        RECT 125.100 25.350 129.600 27.000 ;
        RECT 140.700 26.400 142.500 35.250 ;
        RECT 146.100 27.000 147.900 35.250 ;
        RECT 165.000 29.400 166.800 35.250 ;
        RECT 169.200 31.050 171.000 35.250 ;
        RECT 172.500 32.400 174.300 35.250 ;
        RECT 188.700 32.400 190.500 35.250 ;
        RECT 192.000 31.050 193.800 35.250 ;
        RECT 169.200 29.400 174.900 31.050 ;
        RECT 146.100 25.350 150.600 27.000 ;
        RECT 100.950 20.850 103.050 22.950 ;
        RECT 128.400 21.150 129.600 25.350 ;
        RECT 149.400 21.150 150.600 25.350 ;
        RECT 164.100 24.150 165.900 25.950 ;
        RECT 163.950 22.050 166.050 24.150 ;
        RECT 166.950 23.850 169.050 25.950 ;
        RECT 170.100 24.150 171.900 25.950 ;
        RECT 167.100 22.050 168.900 23.850 ;
        RECT 169.950 22.050 172.050 24.150 ;
        RECT 173.700 22.950 174.900 29.400 ;
        RECT 188.100 29.400 193.800 31.050 ;
        RECT 196.200 29.400 198.000 35.250 ;
        RECT 210.150 30.900 211.950 35.250 ;
        RECT 208.650 29.400 211.950 30.900 ;
        RECT 213.150 29.400 214.950 35.250 ;
        RECT 188.100 22.950 189.300 29.400 ;
        RECT 191.100 24.150 192.900 25.950 ;
        RECT 49.950 17.850 52.050 19.950 ;
        RECT 50.250 16.050 52.050 17.850 ;
        RECT 53.850 15.600 55.050 20.850 ;
        RECT 59.100 19.050 60.900 20.850 ;
        RECT 80.700 15.600 81.900 20.850 ;
        RECT 95.100 19.050 96.900 20.850 ;
        RECT 100.950 15.600 102.150 20.850 ;
        RECT 103.950 17.850 106.050 19.950 ;
        RECT 118.950 17.850 121.050 19.950 ;
        RECT 124.950 17.850 127.050 19.950 ;
        RECT 127.950 19.050 130.050 21.150 ;
        RECT 103.950 16.050 105.750 17.850 ;
        RECT 119.100 16.050 120.900 17.850 ;
        RECT 31.650 3.750 33.450 9.600 ;
        RECT 34.650 3.750 36.450 9.600 ;
        RECT 50.400 3.750 52.200 9.600 ;
        RECT 53.700 3.750 55.500 15.600 ;
        RECT 57.900 3.750 59.700 15.600 ;
        RECT 71.550 14.700 79.350 15.600 ;
        RECT 71.550 3.750 73.350 14.700 ;
        RECT 74.550 3.750 76.350 13.800 ;
        RECT 77.550 3.750 79.350 14.700 ;
        RECT 80.550 3.750 82.350 15.600 ;
        RECT 96.300 3.750 98.100 15.600 ;
        RECT 100.500 3.750 102.300 15.600 ;
        RECT 121.950 14.850 124.050 16.950 ;
        RECT 125.250 16.050 127.050 17.850 ;
        RECT 122.100 13.050 123.900 14.850 ;
        RECT 128.700 10.800 129.750 19.050 ;
        RECT 139.950 17.850 142.050 19.950 ;
        RECT 145.950 17.850 148.050 19.950 ;
        RECT 148.950 19.050 151.050 21.150 ;
        RECT 172.950 20.850 175.050 22.950 ;
        RECT 187.950 20.850 190.050 22.950 ;
        RECT 190.950 22.050 193.050 24.150 ;
        RECT 193.950 23.850 196.050 25.950 ;
        RECT 197.100 24.150 198.900 25.950 ;
        RECT 194.100 22.050 195.900 23.850 ;
        RECT 196.950 22.050 199.050 24.150 ;
        RECT 208.650 22.950 209.850 29.400 ;
        RECT 211.950 27.900 213.750 28.500 ;
        RECT 217.650 27.900 219.450 35.250 ;
        RECT 211.950 26.700 219.450 27.900 ;
        RECT 208.650 20.850 211.050 22.950 ;
        RECT 212.100 21.150 213.900 22.950 ;
        RECT 140.100 16.050 141.900 17.850 ;
        RECT 142.950 14.850 145.050 16.950 ;
        RECT 146.250 16.050 148.050 17.850 ;
        RECT 143.100 13.050 144.900 14.850 ;
        RECT 149.700 10.800 150.750 19.050 ;
        RECT 173.700 15.600 174.900 20.850 ;
        RECT 188.100 15.600 189.300 20.850 ;
        RECT 208.650 15.600 209.850 20.850 ;
        RECT 211.950 19.050 214.050 21.150 ;
        RECT 122.700 9.900 129.750 10.800 ;
        RECT 122.700 9.600 124.350 9.900 ;
        RECT 103.800 3.750 105.600 9.600 ;
        RECT 119.550 3.750 121.350 9.600 ;
        RECT 122.550 3.750 124.350 9.600 ;
        RECT 128.550 9.600 129.750 9.900 ;
        RECT 143.700 9.900 150.750 10.800 ;
        RECT 143.700 9.600 145.350 9.900 ;
        RECT 125.550 3.750 127.350 9.000 ;
        RECT 128.550 3.750 130.350 9.600 ;
        RECT 140.550 3.750 142.350 9.600 ;
        RECT 143.550 3.750 145.350 9.600 ;
        RECT 149.550 9.600 150.750 9.900 ;
        RECT 164.550 14.700 172.350 15.600 ;
        RECT 146.550 3.750 148.350 9.000 ;
        RECT 149.550 3.750 151.350 9.600 ;
        RECT 164.550 3.750 166.350 14.700 ;
        RECT 167.550 3.750 169.350 13.800 ;
        RECT 170.550 3.750 172.350 14.700 ;
        RECT 173.550 3.750 175.350 15.600 ;
        RECT 187.650 3.750 189.450 15.600 ;
        RECT 190.650 14.700 198.450 15.600 ;
        RECT 190.650 3.750 192.450 14.700 ;
        RECT 193.650 3.750 195.450 13.800 ;
        RECT 196.650 3.750 198.450 14.700 ;
        RECT 208.050 3.750 209.850 15.600 ;
        RECT 211.050 3.750 212.850 15.600 ;
        RECT 215.100 9.600 216.300 26.700 ;
        RECT 230.700 26.400 232.500 35.250 ;
        RECT 236.100 27.000 237.900 35.250 ;
        RECT 251.550 30.300 253.350 35.250 ;
        RECT 254.550 31.200 256.350 35.250 ;
        RECT 257.550 30.300 259.350 35.250 ;
        RECT 251.550 28.950 259.350 30.300 ;
        RECT 260.550 29.400 262.350 35.250 ;
        RECT 278.700 32.400 280.500 35.250 ;
        RECT 282.000 31.050 283.800 35.250 ;
        RECT 278.100 29.400 283.800 31.050 ;
        RECT 286.200 29.400 288.000 35.250 ;
        RECT 299.550 32.400 301.350 35.250 ;
        RECT 302.550 32.400 304.350 35.250 ;
        RECT 317.250 32.400 319.350 35.250 ;
        RECT 320.550 32.400 322.350 35.250 ;
        RECT 323.550 32.400 325.350 35.250 ;
        RECT 326.550 32.400 328.350 35.250 ;
        RECT 289.950 30.450 292.050 31.050 ;
        RECT 298.950 30.450 301.050 31.050 ;
        RECT 289.950 29.550 301.050 30.450 ;
        RECT 260.550 27.300 261.750 29.400 ;
        RECT 236.100 25.350 240.600 27.000 ;
        RECT 258.000 26.250 261.750 27.300 ;
        RECT 217.950 20.850 220.050 22.950 ;
        RECT 239.400 21.150 240.600 25.350 ;
        RECT 254.100 24.150 255.900 25.950 ;
        RECT 218.100 19.050 219.900 20.850 ;
        RECT 229.950 17.850 232.050 19.950 ;
        RECT 235.950 17.850 238.050 19.950 ;
        RECT 238.950 19.050 241.050 21.150 ;
        RECT 250.950 20.850 253.050 22.950 ;
        RECT 253.950 22.050 256.050 24.150 ;
        RECT 257.850 22.950 259.050 26.250 ;
        RECT 278.100 22.950 279.300 29.400 ;
        RECT 289.950 28.950 292.050 29.550 ;
        RECT 298.950 28.950 301.050 29.550 ;
        RECT 281.100 24.150 282.900 25.950 ;
        RECT 256.950 20.850 259.050 22.950 ;
        RECT 277.950 20.850 280.050 22.950 ;
        RECT 280.950 22.050 283.050 24.150 ;
        RECT 283.950 23.850 286.050 25.950 ;
        RECT 287.100 24.150 288.900 25.950 ;
        RECT 284.100 22.050 285.900 23.850 ;
        RECT 286.950 22.050 289.050 24.150 ;
        RECT 298.950 23.850 301.050 25.950 ;
        RECT 302.400 24.150 303.600 32.400 ;
        RECT 321.300 31.500 322.350 32.400 ;
        RECT 327.300 31.500 328.350 32.400 ;
        RECT 321.300 30.600 332.100 31.500 ;
        RECT 323.100 24.150 324.900 25.950 ;
        RECT 330.900 24.150 332.100 30.600 ;
        RECT 347.550 30.300 349.350 35.250 ;
        RECT 350.550 31.200 352.350 35.250 ;
        RECT 353.550 30.300 355.350 35.250 ;
        RECT 347.550 28.950 355.350 30.300 ;
        RECT 356.550 29.400 358.350 35.250 ;
        RECT 356.550 27.300 357.750 29.400 ;
        RECT 354.000 26.250 357.750 27.300 ;
        RECT 374.100 27.000 375.900 35.250 ;
        RECT 350.100 24.150 351.900 25.950 ;
        RECT 299.100 22.050 300.900 23.850 ;
        RECT 301.950 22.050 304.050 24.150 ;
        RECT 251.100 19.050 252.900 20.850 ;
        RECT 230.100 16.050 231.900 17.850 ;
        RECT 232.950 14.850 235.050 16.950 ;
        RECT 236.250 16.050 238.050 17.850 ;
        RECT 233.100 13.050 234.900 14.850 ;
        RECT 239.700 10.800 240.750 19.050 ;
        RECT 256.950 15.600 258.150 20.850 ;
        RECT 259.950 17.850 262.050 19.950 ;
        RECT 259.950 16.050 261.750 17.850 ;
        RECT 278.100 15.600 279.300 20.850 ;
        RECT 233.700 9.900 240.750 10.800 ;
        RECT 233.700 9.600 235.350 9.900 ;
        RECT 214.650 3.750 216.450 9.600 ;
        RECT 217.650 3.750 219.450 9.600 ;
        RECT 230.550 3.750 232.350 9.600 ;
        RECT 233.550 3.750 235.350 9.600 ;
        RECT 239.550 9.600 240.750 9.900 ;
        RECT 236.550 3.750 238.350 9.000 ;
        RECT 239.550 3.750 241.350 9.600 ;
        RECT 252.300 3.750 254.100 15.600 ;
        RECT 256.500 3.750 258.300 15.600 ;
        RECT 259.800 3.750 261.600 9.600 ;
        RECT 277.650 3.750 279.450 15.600 ;
        RECT 280.650 14.700 288.450 15.600 ;
        RECT 280.650 3.750 282.450 14.700 ;
        RECT 283.650 3.750 285.450 13.800 ;
        RECT 286.650 3.750 288.450 14.700 ;
        RECT 302.400 9.600 303.600 22.050 ;
        RECT 316.950 20.850 319.050 22.950 ;
        RECT 322.950 22.050 325.050 24.150 ;
        RECT 325.950 20.850 328.050 22.950 ;
        RECT 330.900 22.050 334.050 24.150 ;
        RECT 317.100 19.050 318.900 20.850 ;
        RECT 326.100 19.050 327.900 20.850 ;
        RECT 330.900 16.800 332.100 22.050 ;
        RECT 346.950 20.850 349.050 22.950 ;
        RECT 349.950 22.050 352.050 24.150 ;
        RECT 353.850 22.950 355.050 26.250 ;
        RECT 352.950 20.850 355.050 22.950 ;
        RECT 371.400 25.350 375.900 27.000 ;
        RECT 379.500 26.400 381.300 35.250 ;
        RECT 392.550 27.900 394.350 35.250 ;
        RECT 397.050 29.400 398.850 35.250 ;
        RECT 400.050 30.900 401.850 35.250 ;
        RECT 413.550 32.400 415.350 35.250 ;
        RECT 416.550 32.400 418.350 35.250 ;
        RECT 419.550 32.400 421.350 35.250 ;
        RECT 400.050 29.400 403.350 30.900 ;
        RECT 398.250 27.900 400.050 28.500 ;
        RECT 392.550 26.700 400.050 27.900 ;
        RECT 371.400 21.150 372.600 25.350 ;
        RECT 347.100 19.050 348.900 20.850 ;
        RECT 330.900 15.600 334.350 16.800 ;
        RECT 352.950 15.600 354.150 20.850 ;
        RECT 355.950 17.850 358.050 19.950 ;
        RECT 370.950 19.050 373.050 21.150 ;
        RECT 391.950 20.850 394.050 22.950 ;
        RECT 355.950 16.050 357.750 17.850 ;
        RECT 314.550 13.500 322.350 14.400 ;
        RECT 299.550 3.750 301.350 9.600 ;
        RECT 302.550 3.750 304.350 9.600 ;
        RECT 314.550 3.750 316.350 13.500 ;
        RECT 317.550 3.750 319.350 12.600 ;
        RECT 320.550 4.500 322.350 13.500 ;
        RECT 323.550 13.200 331.950 14.100 ;
        RECT 323.550 5.400 325.350 13.200 ;
        RECT 326.550 4.500 328.350 12.300 ;
        RECT 320.550 3.750 328.350 4.500 ;
        RECT 330.150 4.500 331.950 13.200 ;
        RECT 333.150 13.200 334.350 15.600 ;
        RECT 333.150 5.400 334.950 13.200 ;
        RECT 336.150 4.500 337.950 13.800 ;
        RECT 330.150 3.750 337.950 4.500 ;
        RECT 348.300 3.750 350.100 15.600 ;
        RECT 352.500 3.750 354.300 15.600 ;
        RECT 371.250 10.800 372.300 19.050 ;
        RECT 373.950 17.850 376.050 19.950 ;
        RECT 379.950 17.850 382.050 19.950 ;
        RECT 392.100 19.050 393.900 20.850 ;
        RECT 373.950 16.050 375.750 17.850 ;
        RECT 376.950 14.850 379.050 16.950 ;
        RECT 380.100 16.050 381.900 17.850 ;
        RECT 377.100 13.050 378.900 14.850 ;
        RECT 371.250 9.900 378.300 10.800 ;
        RECT 371.250 9.600 372.450 9.900 ;
        RECT 355.800 3.750 357.600 9.600 ;
        RECT 370.650 3.750 372.450 9.600 ;
        RECT 376.650 9.600 378.300 9.900 ;
        RECT 395.700 9.600 396.900 26.700 ;
        RECT 402.150 22.950 403.350 29.400 ;
        RECT 417.000 25.950 418.050 32.400 ;
        RECT 431.550 30.300 433.350 35.250 ;
        RECT 434.550 31.200 436.350 35.250 ;
        RECT 437.550 30.300 439.350 35.250 ;
        RECT 431.550 28.950 439.350 30.300 ;
        RECT 440.550 29.400 442.350 35.250 ;
        RECT 452.550 32.400 454.350 35.250 ;
        RECT 455.550 32.400 457.350 35.250 ;
        RECT 458.550 32.400 460.350 35.250 ;
        RECT 440.550 27.300 441.750 29.400 ;
        RECT 456.450 28.200 457.350 32.400 ;
        RECT 461.550 29.400 463.350 35.250 ;
        RECT 456.450 27.300 459.750 28.200 ;
        RECT 438.000 26.250 441.750 27.300 ;
        RECT 457.950 26.400 459.750 27.300 ;
        RECT 415.950 23.850 418.050 25.950 ;
        RECT 434.100 24.150 435.900 25.950 ;
        RECT 398.100 21.150 399.900 22.950 ;
        RECT 397.950 19.050 400.050 21.150 ;
        RECT 400.950 20.850 403.350 22.950 ;
        RECT 412.950 20.850 415.050 22.950 ;
        RECT 402.150 15.600 403.350 20.850 ;
        RECT 413.100 19.050 414.900 20.850 ;
        RECT 417.000 16.650 418.050 23.850 ;
        RECT 418.950 20.850 421.050 22.950 ;
        RECT 430.950 20.850 433.050 22.950 ;
        RECT 433.950 22.050 436.050 24.150 ;
        RECT 437.850 22.950 439.050 26.250 ;
        RECT 451.950 23.850 454.050 25.950 ;
        RECT 436.950 20.850 439.050 22.950 ;
        RECT 452.100 22.050 453.900 23.850 ;
        RECT 454.950 20.850 457.050 22.950 ;
        RECT 419.100 19.050 420.900 20.850 ;
        RECT 431.100 19.050 432.900 20.850 ;
        RECT 417.000 15.600 419.550 16.650 ;
        RECT 436.950 15.600 438.150 20.850 ;
        RECT 439.950 17.850 442.050 19.950 ;
        RECT 455.100 19.050 456.900 20.850 ;
        RECT 458.700 18.150 459.600 26.400 ;
        RECT 462.000 24.150 463.050 29.400 ;
        RECT 473.550 27.900 475.350 35.250 ;
        RECT 478.050 29.400 479.850 35.250 ;
        RECT 481.050 30.900 482.850 35.250 ;
        RECT 481.050 29.400 484.350 30.900 ;
        RECT 479.250 27.900 481.050 28.500 ;
        RECT 473.550 26.700 481.050 27.900 ;
        RECT 460.950 22.050 463.050 24.150 ;
        RECT 457.950 18.000 459.750 18.150 ;
        RECT 439.950 16.050 441.750 17.850 ;
        RECT 452.550 16.800 459.750 18.000 ;
        RECT 452.550 15.600 453.750 16.800 ;
        RECT 457.950 16.350 459.750 16.800 ;
        RECT 373.650 3.750 375.450 9.000 ;
        RECT 376.650 3.750 378.450 9.600 ;
        RECT 379.650 3.750 381.450 9.600 ;
        RECT 392.550 3.750 394.350 9.600 ;
        RECT 395.550 3.750 397.350 9.600 ;
        RECT 399.150 3.750 400.950 15.600 ;
        RECT 402.150 3.750 403.950 15.600 ;
        RECT 413.550 3.750 415.350 15.600 ;
        RECT 417.750 3.750 419.550 15.600 ;
        RECT 432.300 3.750 434.100 15.600 ;
        RECT 436.500 3.750 438.300 15.600 ;
        RECT 439.800 3.750 441.600 9.600 ;
        RECT 452.550 3.750 454.350 15.600 ;
        RECT 461.100 15.450 462.450 22.050 ;
        RECT 472.950 20.850 475.050 22.950 ;
        RECT 473.100 19.050 474.900 20.850 ;
        RECT 457.050 3.750 458.850 15.450 ;
        RECT 460.050 14.100 462.450 15.450 ;
        RECT 460.050 3.750 461.850 14.100 ;
        RECT 476.700 9.600 477.900 26.700 ;
        RECT 483.150 22.950 484.350 29.400 ;
        RECT 497.550 30.300 499.350 35.250 ;
        RECT 500.550 31.200 502.350 35.250 ;
        RECT 503.550 30.300 505.350 35.250 ;
        RECT 497.550 28.950 505.350 30.300 ;
        RECT 506.550 29.400 508.350 35.250 ;
        RECT 518.550 30.300 520.350 35.250 ;
        RECT 521.550 31.200 523.350 35.250 ;
        RECT 524.550 30.300 526.350 35.250 ;
        RECT 506.550 27.300 507.750 29.400 ;
        RECT 518.550 28.950 526.350 30.300 ;
        RECT 527.550 29.400 529.350 35.250 ;
        RECT 542.550 30.300 544.350 35.250 ;
        RECT 545.550 31.200 547.350 35.250 ;
        RECT 548.550 30.300 550.350 35.250 ;
        RECT 527.550 27.300 528.750 29.400 ;
        RECT 542.550 28.950 550.350 30.300 ;
        RECT 551.550 29.400 553.350 35.250 ;
        RECT 566.700 32.400 568.500 35.250 ;
        RECT 570.000 31.050 571.800 35.250 ;
        RECT 566.100 29.400 571.800 31.050 ;
        RECT 574.200 29.400 576.000 35.250 ;
        RECT 584.550 32.400 586.350 35.250 ;
        RECT 587.550 32.400 589.350 35.250 ;
        RECT 590.550 32.400 592.350 35.250 ;
        RECT 605.550 32.400 607.350 35.250 ;
        RECT 608.550 32.400 610.350 35.250 ;
        RECT 551.550 27.300 552.750 29.400 ;
        RECT 504.000 26.250 507.750 27.300 ;
        RECT 525.000 26.250 528.750 27.300 ;
        RECT 549.000 26.250 552.750 27.300 ;
        RECT 500.100 24.150 501.900 25.950 ;
        RECT 479.100 21.150 480.900 22.950 ;
        RECT 478.950 19.050 481.050 21.150 ;
        RECT 481.950 20.850 484.350 22.950 ;
        RECT 496.950 20.850 499.050 22.950 ;
        RECT 499.950 22.050 502.050 24.150 ;
        RECT 503.850 22.950 505.050 26.250 ;
        RECT 521.100 24.150 522.900 25.950 ;
        RECT 502.950 20.850 505.050 22.950 ;
        RECT 517.950 20.850 520.050 22.950 ;
        RECT 520.950 22.050 523.050 24.150 ;
        RECT 524.850 22.950 526.050 26.250 ;
        RECT 545.100 24.150 546.900 25.950 ;
        RECT 523.950 20.850 526.050 22.950 ;
        RECT 541.950 20.850 544.050 22.950 ;
        RECT 544.950 22.050 547.050 24.150 ;
        RECT 548.850 22.950 550.050 26.250 ;
        RECT 566.100 22.950 567.300 29.400 ;
        RECT 588.000 25.950 589.050 32.400 ;
        RECT 569.100 24.150 570.900 25.950 ;
        RECT 547.950 20.850 550.050 22.950 ;
        RECT 565.950 20.850 568.050 22.950 ;
        RECT 568.950 22.050 571.050 24.150 ;
        RECT 571.950 23.850 574.050 25.950 ;
        RECT 575.100 24.150 576.900 25.950 ;
        RECT 572.100 22.050 573.900 23.850 ;
        RECT 574.950 22.050 577.050 24.150 ;
        RECT 586.950 23.850 589.050 25.950 ;
        RECT 604.950 23.850 607.050 25.950 ;
        RECT 608.400 24.150 609.600 32.400 ;
        RECT 621.000 29.400 622.800 35.250 ;
        RECT 625.200 31.050 627.000 35.250 ;
        RECT 628.500 32.400 630.300 35.250 ;
        RECT 625.200 29.400 630.900 31.050 ;
        RECT 620.100 24.150 621.900 25.950 ;
        RECT 583.950 20.850 586.050 22.950 ;
        RECT 483.150 15.600 484.350 20.850 ;
        RECT 497.100 19.050 498.900 20.850 ;
        RECT 502.950 15.600 504.150 20.850 ;
        RECT 505.950 17.850 508.050 19.950 ;
        RECT 518.100 19.050 519.900 20.850 ;
        RECT 505.950 16.050 507.750 17.850 ;
        RECT 523.950 15.600 525.150 20.850 ;
        RECT 526.950 17.850 529.050 19.950 ;
        RECT 542.100 19.050 543.900 20.850 ;
        RECT 526.950 16.050 528.750 17.850 ;
        RECT 547.950 15.600 549.150 20.850 ;
        RECT 550.950 17.850 553.050 19.950 ;
        RECT 550.950 16.050 552.750 17.850 ;
        RECT 566.100 15.600 567.300 20.850 ;
        RECT 584.100 19.050 585.900 20.850 ;
        RECT 588.000 16.650 589.050 23.850 ;
        RECT 589.950 20.850 592.050 22.950 ;
        RECT 605.100 22.050 606.900 23.850 ;
        RECT 607.950 22.050 610.050 24.150 ;
        RECT 619.950 22.050 622.050 24.150 ;
        RECT 622.950 23.850 625.050 25.950 ;
        RECT 626.100 24.150 627.900 25.950 ;
        RECT 623.100 22.050 624.900 23.850 ;
        RECT 625.950 22.050 628.050 24.150 ;
        RECT 629.700 22.950 630.900 29.400 ;
        RECT 644.850 28.200 646.650 35.250 ;
        RECT 649.350 29.400 651.150 35.250 ;
        RECT 662.550 32.400 664.350 35.250 ;
        RECT 665.550 32.400 667.350 35.250 ;
        RECT 668.550 32.400 670.350 35.250 ;
        RECT 644.850 27.300 648.450 28.200 ;
        RECT 590.100 19.050 591.900 20.850 ;
        RECT 588.000 15.600 590.550 16.650 ;
        RECT 473.550 3.750 475.350 9.600 ;
        RECT 476.550 3.750 478.350 9.600 ;
        RECT 480.150 3.750 481.950 15.600 ;
        RECT 483.150 3.750 484.950 15.600 ;
        RECT 498.300 3.750 500.100 15.600 ;
        RECT 502.500 3.750 504.300 15.600 ;
        RECT 505.800 3.750 507.600 9.600 ;
        RECT 519.300 3.750 521.100 15.600 ;
        RECT 523.500 3.750 525.300 15.600 ;
        RECT 526.800 3.750 528.600 9.600 ;
        RECT 543.300 3.750 545.100 15.600 ;
        RECT 547.500 3.750 549.300 15.600 ;
        RECT 550.800 3.750 552.600 9.600 ;
        RECT 565.650 3.750 567.450 15.600 ;
        RECT 568.650 14.700 576.450 15.600 ;
        RECT 568.650 3.750 570.450 14.700 ;
        RECT 571.650 3.750 573.450 13.800 ;
        RECT 574.650 3.750 576.450 14.700 ;
        RECT 584.550 3.750 586.350 15.600 ;
        RECT 588.750 3.750 590.550 15.600 ;
        RECT 608.400 9.600 609.600 22.050 ;
        RECT 628.950 20.850 631.050 22.950 ;
        RECT 644.100 21.150 645.900 22.950 ;
        RECT 629.700 15.600 630.900 20.850 ;
        RECT 643.950 19.050 646.050 21.150 ;
        RECT 647.250 19.950 648.450 27.300 ;
        RECT 666.000 25.950 667.050 32.400 ;
        RECT 684.000 29.400 685.800 35.250 ;
        RECT 688.200 31.050 690.000 35.250 ;
        RECT 691.500 32.400 693.300 35.250 ;
        RECT 688.200 29.400 693.900 31.050 ;
        RECT 664.950 23.850 667.050 25.950 ;
        RECT 683.100 24.150 684.900 25.950 ;
        RECT 650.100 21.150 651.900 22.950 ;
        RECT 646.950 17.850 649.050 19.950 ;
        RECT 649.950 19.050 652.050 21.150 ;
        RECT 661.950 20.850 664.050 22.950 ;
        RECT 662.100 19.050 663.900 20.850 ;
        RECT 620.550 14.700 628.350 15.600 ;
        RECT 605.550 3.750 607.350 9.600 ;
        RECT 608.550 3.750 610.350 9.600 ;
        RECT 620.550 3.750 622.350 14.700 ;
        RECT 623.550 3.750 625.350 13.800 ;
        RECT 626.550 3.750 628.350 14.700 ;
        RECT 629.550 3.750 631.350 15.600 ;
        RECT 647.250 9.600 648.450 17.850 ;
        RECT 666.000 16.650 667.050 23.850 ;
        RECT 667.950 20.850 670.050 22.950 ;
        RECT 682.950 22.050 685.050 24.150 ;
        RECT 685.950 23.850 688.050 25.950 ;
        RECT 689.100 24.150 690.900 25.950 ;
        RECT 686.100 22.050 687.900 23.850 ;
        RECT 688.950 22.050 691.050 24.150 ;
        RECT 692.700 22.950 693.900 29.400 ;
        RECT 704.550 30.300 706.350 35.250 ;
        RECT 707.550 31.200 709.350 35.250 ;
        RECT 710.550 30.300 712.350 35.250 ;
        RECT 704.550 28.950 712.350 30.300 ;
        RECT 713.550 29.400 715.350 35.250 ;
        RECT 725.550 32.400 727.350 35.250 ;
        RECT 728.550 32.400 730.350 35.250 ;
        RECT 713.550 27.300 714.750 29.400 ;
        RECT 711.000 26.250 714.750 27.300 ;
        RECT 707.100 24.150 708.900 25.950 ;
        RECT 691.950 20.850 694.050 22.950 ;
        RECT 703.950 20.850 706.050 22.950 ;
        RECT 706.950 22.050 709.050 24.150 ;
        RECT 710.850 22.950 712.050 26.250 ;
        RECT 724.950 23.850 727.050 25.950 ;
        RECT 728.400 24.150 729.600 32.400 ;
        RECT 743.850 28.200 745.650 35.250 ;
        RECT 748.350 29.400 750.150 35.250 ;
        RECT 753.150 29.400 754.950 35.250 ;
        RECT 756.150 32.400 757.950 35.250 ;
        RECT 760.950 33.300 762.750 35.250 ;
        RECT 759.000 32.400 762.750 33.300 ;
        RECT 765.450 32.400 767.250 35.250 ;
        RECT 768.750 32.400 770.550 35.250 ;
        RECT 772.650 32.400 774.450 35.250 ;
        RECT 776.850 32.400 778.650 35.250 ;
        RECT 781.350 32.400 783.150 35.250 ;
        RECT 759.000 31.500 760.050 32.400 ;
        RECT 757.950 29.400 760.050 31.500 ;
        RECT 768.750 30.600 769.800 32.400 ;
        RECT 743.850 27.300 747.450 28.200 ;
        RECT 709.950 20.850 712.050 22.950 ;
        RECT 725.100 22.050 726.900 23.850 ;
        RECT 727.950 22.050 730.050 24.150 ;
        RECT 668.100 19.050 669.900 20.850 ;
        RECT 666.000 15.600 668.550 16.650 ;
        RECT 692.700 15.600 693.900 20.850 ;
        RECT 704.100 19.050 705.900 20.850 ;
        RECT 709.950 15.600 711.150 20.850 ;
        RECT 712.950 17.850 715.050 19.950 ;
        RECT 712.950 16.050 714.750 17.850 ;
        RECT 643.650 3.750 645.450 9.600 ;
        RECT 646.650 3.750 648.450 9.600 ;
        RECT 649.650 3.750 651.450 9.600 ;
        RECT 662.550 3.750 664.350 15.600 ;
        RECT 666.750 3.750 668.550 15.600 ;
        RECT 683.550 14.700 691.350 15.600 ;
        RECT 683.550 3.750 685.350 14.700 ;
        RECT 686.550 3.750 688.350 13.800 ;
        RECT 689.550 3.750 691.350 14.700 ;
        RECT 692.550 3.750 694.350 15.600 ;
        RECT 705.300 3.750 707.100 15.600 ;
        RECT 709.500 3.750 711.300 15.600 ;
        RECT 728.400 9.600 729.600 22.050 ;
        RECT 743.100 21.150 744.900 22.950 ;
        RECT 742.950 19.050 745.050 21.150 ;
        RECT 746.250 19.950 747.450 27.300 ;
        RECT 749.100 21.150 750.900 22.950 ;
        RECT 745.950 17.850 748.050 19.950 ;
        RECT 748.950 19.050 751.050 21.150 ;
        RECT 746.250 9.600 747.450 17.850 ;
        RECT 753.150 16.800 754.050 29.400 ;
        RECT 761.550 28.800 763.350 30.600 ;
        RECT 764.850 29.550 769.800 30.600 ;
        RECT 777.300 31.500 778.350 32.400 ;
        RECT 777.300 30.300 781.050 31.500 ;
        RECT 764.850 28.800 766.650 29.550 ;
        RECT 761.850 27.900 762.900 28.800 ;
        RECT 772.050 28.200 773.850 30.000 ;
        RECT 778.950 29.400 781.050 30.300 ;
        RECT 784.650 29.400 786.450 35.250 ;
        RECT 794.850 29.400 796.650 35.250 ;
        RECT 772.050 27.900 772.950 28.200 ;
        RECT 761.850 27.000 772.950 27.900 ;
        RECT 785.250 27.150 786.450 29.400 ;
        RECT 799.350 28.200 801.150 35.250 ;
        RECT 817.800 29.400 819.600 35.250 ;
        RECT 822.000 29.400 823.800 35.250 ;
        RECT 826.200 29.400 828.000 35.250 ;
        RECT 831.150 29.400 832.950 35.250 ;
        RECT 834.150 32.400 835.950 35.250 ;
        RECT 838.950 33.300 840.750 35.250 ;
        RECT 837.000 32.400 840.750 33.300 ;
        RECT 843.450 32.400 845.250 35.250 ;
        RECT 846.750 32.400 848.550 35.250 ;
        RECT 850.650 32.400 852.450 35.250 ;
        RECT 854.850 32.400 856.650 35.250 ;
        RECT 859.350 32.400 861.150 35.250 ;
        RECT 837.000 31.500 838.050 32.400 ;
        RECT 835.950 29.400 838.050 31.500 ;
        RECT 846.750 30.600 847.800 32.400 ;
        RECT 761.850 25.800 762.900 27.000 ;
        RECT 756.000 24.600 762.900 25.800 ;
        RECT 756.000 23.850 756.900 24.600 ;
        RECT 761.100 24.000 762.900 24.600 ;
        RECT 755.100 22.050 756.900 23.850 ;
        RECT 758.100 22.950 759.900 23.700 ;
        RECT 772.050 22.950 772.950 27.000 ;
        RECT 781.950 25.050 786.450 27.150 ;
        RECT 780.150 23.250 784.050 25.050 ;
        RECT 781.950 22.950 784.050 23.250 ;
        RECT 758.100 21.900 766.050 22.950 ;
        RECT 763.950 20.850 766.050 21.900 ;
        RECT 769.950 20.850 772.950 22.950 ;
        RECT 762.450 17.100 764.250 17.400 ;
        RECT 762.450 16.800 770.850 17.100 ;
        RECT 753.150 16.200 770.850 16.800 ;
        RECT 753.150 15.600 764.250 16.200 ;
        RECT 712.800 3.750 714.600 9.600 ;
        RECT 725.550 3.750 727.350 9.600 ;
        RECT 728.550 3.750 730.350 9.600 ;
        RECT 742.650 3.750 744.450 9.600 ;
        RECT 745.650 3.750 747.450 9.600 ;
        RECT 748.650 3.750 750.450 9.600 ;
        RECT 753.150 3.750 754.950 15.600 ;
        RECT 767.250 14.700 769.050 15.300 ;
        RECT 761.550 13.500 769.050 14.700 ;
        RECT 769.950 14.100 770.850 16.200 ;
        RECT 772.050 16.200 772.950 20.850 ;
        RECT 782.250 17.400 784.050 19.200 ;
        RECT 778.950 16.200 783.150 17.400 ;
        RECT 772.050 15.300 778.050 16.200 ;
        RECT 778.950 15.300 781.050 16.200 ;
        RECT 785.250 15.600 786.450 25.050 ;
        RECT 797.550 27.300 801.150 28.200 ;
        RECT 794.100 21.150 795.900 22.950 ;
        RECT 793.950 19.050 796.050 21.150 ;
        RECT 797.550 19.950 798.750 27.300 ;
        RECT 818.250 24.150 820.050 25.950 ;
        RECT 800.100 21.150 801.900 22.950 ;
        RECT 796.950 17.850 799.050 19.950 ;
        RECT 799.950 19.050 802.050 21.150 ;
        RECT 814.950 20.850 817.050 22.950 ;
        RECT 817.950 22.050 820.050 24.150 ;
        RECT 822.000 22.950 823.050 29.400 ;
        RECT 820.950 20.850 823.050 22.950 ;
        RECT 823.950 24.150 825.750 25.950 ;
        RECT 823.950 22.050 826.050 24.150 ;
        RECT 826.950 20.850 829.050 22.950 ;
        RECT 815.100 19.050 816.900 20.850 ;
        RECT 777.150 14.400 778.050 15.300 ;
        RECT 774.450 14.100 776.250 14.400 ;
        RECT 761.550 12.600 762.750 13.500 ;
        RECT 769.950 13.200 776.250 14.100 ;
        RECT 774.450 12.600 776.250 13.200 ;
        RECT 777.150 12.600 779.850 14.400 ;
        RECT 757.950 10.500 762.750 12.600 ;
        RECT 765.150 10.500 772.050 12.300 ;
        RECT 761.550 9.600 762.750 10.500 ;
        RECT 756.150 3.750 757.950 9.600 ;
        RECT 761.250 3.750 763.050 9.600 ;
        RECT 766.050 3.750 767.850 9.600 ;
        RECT 769.050 3.750 770.850 10.500 ;
        RECT 777.150 9.600 781.050 11.700 ;
        RECT 772.950 3.750 774.750 9.600 ;
        RECT 777.150 3.750 778.950 9.600 ;
        RECT 781.650 3.750 783.450 6.600 ;
        RECT 784.650 3.750 786.450 15.600 ;
        RECT 797.550 9.600 798.750 17.850 ;
        RECT 820.950 17.400 821.850 20.850 ;
        RECT 826.950 19.050 828.750 20.850 ;
        RECT 817.800 16.500 821.850 17.400 ;
        RECT 831.150 16.800 832.050 29.400 ;
        RECT 839.550 28.800 841.350 30.600 ;
        RECT 842.850 29.550 847.800 30.600 ;
        RECT 855.300 31.500 856.350 32.400 ;
        RECT 855.300 30.300 859.050 31.500 ;
        RECT 842.850 28.800 844.650 29.550 ;
        RECT 839.850 27.900 840.900 28.800 ;
        RECT 850.050 28.200 851.850 30.000 ;
        RECT 856.950 29.400 859.050 30.300 ;
        RECT 862.650 29.400 864.450 35.250 ;
        RECT 875.850 29.400 877.650 35.250 ;
        RECT 850.050 27.900 850.950 28.200 ;
        RECT 839.850 27.000 850.950 27.900 ;
        RECT 863.250 27.150 864.450 29.400 ;
        RECT 880.350 28.200 882.150 35.250 ;
        RECT 839.850 25.800 840.900 27.000 ;
        RECT 834.000 24.600 840.900 25.800 ;
        RECT 834.000 23.850 834.900 24.600 ;
        RECT 839.100 24.000 840.900 24.600 ;
        RECT 833.100 22.050 834.900 23.850 ;
        RECT 836.100 22.950 837.900 23.700 ;
        RECT 850.050 22.950 850.950 27.000 ;
        RECT 859.950 25.050 864.450 27.150 ;
        RECT 858.150 23.250 862.050 25.050 ;
        RECT 859.950 22.950 862.050 23.250 ;
        RECT 836.100 21.900 844.050 22.950 ;
        RECT 841.950 20.850 844.050 21.900 ;
        RECT 847.950 20.850 850.950 22.950 ;
        RECT 840.450 17.100 842.250 17.400 ;
        RECT 840.450 16.800 848.850 17.100 ;
        RECT 817.800 15.600 819.600 16.500 ;
        RECT 831.150 16.200 848.850 16.800 ;
        RECT 831.150 15.600 842.250 16.200 ;
        RECT 794.550 3.750 796.350 9.600 ;
        RECT 797.550 3.750 799.350 9.600 ;
        RECT 800.550 3.750 802.350 9.600 ;
        RECT 814.650 4.500 816.450 15.600 ;
        RECT 817.650 5.400 819.450 15.600 ;
        RECT 820.650 14.400 828.450 15.300 ;
        RECT 820.650 4.500 822.450 14.400 ;
        RECT 814.650 3.750 822.450 4.500 ;
        RECT 823.650 3.750 825.450 13.500 ;
        RECT 826.650 3.750 828.450 14.400 ;
        RECT 831.150 3.750 832.950 15.600 ;
        RECT 845.250 14.700 847.050 15.300 ;
        RECT 839.550 13.500 847.050 14.700 ;
        RECT 847.950 14.100 848.850 16.200 ;
        RECT 850.050 16.200 850.950 20.850 ;
        RECT 860.250 17.400 862.050 19.200 ;
        RECT 856.950 16.200 861.150 17.400 ;
        RECT 850.050 15.300 856.050 16.200 ;
        RECT 856.950 15.300 859.050 16.200 ;
        RECT 863.250 15.600 864.450 25.050 ;
        RECT 878.550 27.300 882.150 28.200 ;
        RECT 875.100 21.150 876.900 22.950 ;
        RECT 874.950 19.050 877.050 21.150 ;
        RECT 878.550 19.950 879.750 27.300 ;
        RECT 881.100 21.150 882.900 22.950 ;
        RECT 877.950 17.850 880.050 19.950 ;
        RECT 880.950 19.050 883.050 21.150 ;
        RECT 855.150 14.400 856.050 15.300 ;
        RECT 852.450 14.100 854.250 14.400 ;
        RECT 839.550 12.600 840.750 13.500 ;
        RECT 847.950 13.200 854.250 14.100 ;
        RECT 852.450 12.600 854.250 13.200 ;
        RECT 855.150 12.600 857.850 14.400 ;
        RECT 835.950 10.500 840.750 12.600 ;
        RECT 843.150 10.500 850.050 12.300 ;
        RECT 839.550 9.600 840.750 10.500 ;
        RECT 834.150 3.750 835.950 9.600 ;
        RECT 839.250 3.750 841.050 9.600 ;
        RECT 844.050 3.750 845.850 9.600 ;
        RECT 847.050 3.750 848.850 10.500 ;
        RECT 855.150 9.600 859.050 11.700 ;
        RECT 850.950 3.750 852.750 9.600 ;
        RECT 855.150 3.750 856.950 9.600 ;
        RECT 859.650 3.750 861.450 6.600 ;
        RECT 862.650 3.750 864.450 15.600 ;
        RECT 878.550 9.600 879.750 17.850 ;
        RECT 875.550 3.750 877.350 9.600 ;
        RECT 878.550 3.750 880.350 9.600 ;
        RECT 881.550 3.750 883.350 9.600 ;
      LAYER metal2 ;
        RECT 64.950 893.400 67.050 895.500 ;
        RECT 85.950 893.400 88.050 895.500 ;
        RECT 136.950 893.400 139.050 895.500 ;
        RECT 157.950 893.400 160.050 895.500 ;
        RECT 211.950 893.400 214.050 895.500 ;
        RECT 232.950 893.400 235.050 895.500 ;
        RECT 289.950 893.400 292.050 895.500 ;
        RECT 310.950 893.400 313.050 895.500 ;
        RECT 418.950 893.400 421.050 895.500 ;
        RECT 439.950 893.400 442.050 895.500 ;
        RECT 472.950 893.400 475.050 895.500 ;
        RECT 493.950 893.400 496.050 895.500 ;
        RECT 679.950 893.400 682.050 895.500 ;
        RECT 700.950 893.400 703.050 895.500 ;
        RECT 13.950 891.450 16.050 892.050 ;
        RECT 13.950 890.400 18.450 891.450 ;
        RECT 13.950 889.950 16.050 890.400 ;
        RECT 10.950 887.250 13.050 888.150 ;
        RECT 13.950 887.850 16.050 888.750 ;
        RECT 10.950 883.950 13.050 886.050 ;
        RECT 17.400 883.050 18.450 890.400 ;
        RECT 31.950 886.950 34.050 889.050 ;
        RECT 43.950 886.950 46.050 889.050 ;
        RECT 47.250 887.250 48.750 888.150 ;
        RECT 49.950 886.950 52.050 889.050 ;
        RECT 32.400 886.050 33.450 886.950 ;
        RECT 28.950 884.250 30.750 885.150 ;
        RECT 31.950 883.950 34.050 886.050 ;
        RECT 35.250 884.250 37.050 885.150 ;
        RECT 43.950 884.850 45.750 885.750 ;
        RECT 46.950 883.950 49.050 886.050 ;
        RECT 50.250 884.850 51.750 885.750 ;
        RECT 52.950 883.950 55.050 886.050 ;
        RECT 10.950 880.950 13.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 28.950 880.950 31.050 883.050 ;
        RECT 32.250 881.850 33.750 882.750 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 46.950 880.950 49.050 883.050 ;
        RECT 52.950 881.850 55.050 882.750 ;
        RECT 11.400 808.050 12.450 880.950 ;
        RECT 35.400 850.050 36.450 880.950 ;
        RECT 40.950 850.950 43.050 853.050 ;
        RECT 34.950 847.950 37.050 850.050 ;
        RECT 13.950 844.950 16.050 847.050 ;
        RECT 34.950 846.450 37.050 847.050 ;
        RECT 28.950 845.250 31.050 846.150 ;
        RECT 32.400 845.400 37.050 846.450 ;
        RECT 13.950 842.850 16.050 843.750 ;
        RECT 16.950 842.250 19.050 843.150 ;
        RECT 28.950 841.950 31.050 844.050 ;
        RECT 16.950 838.950 19.050 841.050 ;
        RECT 17.400 838.050 18.450 838.950 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 22.950 835.950 25.050 838.050 ;
        RECT 16.950 820.950 19.050 823.050 ;
        RECT 17.400 817.050 18.450 820.950 ;
        RECT 23.400 817.050 24.450 835.950 ;
        RECT 13.950 814.950 16.050 817.050 ;
        RECT 16.950 814.950 19.050 817.050 ;
        RECT 22.950 816.450 25.050 817.050 ;
        RECT 20.250 815.250 21.750 816.150 ;
        RECT 22.950 815.400 27.450 816.450 ;
        RECT 22.950 814.950 25.050 815.400 ;
        RECT 14.400 814.050 15.450 814.950 ;
        RECT 13.950 811.950 16.050 814.050 ;
        RECT 17.250 812.850 18.750 813.750 ;
        RECT 19.950 811.950 22.050 814.050 ;
        RECT 23.250 812.850 25.050 813.750 ;
        RECT 13.950 809.850 16.050 810.750 ;
        RECT 10.950 805.950 13.050 808.050 ;
        RECT 20.400 804.450 21.450 811.950 ;
        RECT 26.400 811.050 27.450 815.400 ;
        RECT 28.950 814.950 31.050 817.050 ;
        RECT 25.950 808.950 28.050 811.050 ;
        RECT 20.400 803.400 24.450 804.450 ;
        RECT 19.950 778.950 22.050 781.050 ;
        RECT 20.400 778.050 21.450 778.950 ;
        RECT 13.950 775.950 16.050 778.050 ;
        RECT 17.250 776.250 18.750 777.150 ;
        RECT 19.950 775.950 22.050 778.050 ;
        RECT 23.400 775.050 24.450 803.400 ;
        RECT 25.950 778.950 28.050 781.050 ;
        RECT 13.950 773.850 15.750 774.750 ;
        RECT 16.950 772.950 19.050 775.050 ;
        RECT 20.250 773.850 22.050 774.750 ;
        RECT 22.950 772.950 25.050 775.050 ;
        RECT 10.950 744.450 13.050 745.050 ;
        RECT 10.950 743.400 15.450 744.450 ;
        RECT 10.950 742.950 13.050 743.400 ;
        RECT 10.950 740.850 13.050 741.750 ;
        RECT 14.400 736.050 15.450 743.400 ;
        RECT 19.950 742.950 22.050 745.050 ;
        RECT 16.950 740.250 19.050 741.150 ;
        RECT 19.950 740.850 22.050 741.750 ;
        RECT 22.950 739.950 25.050 742.050 ;
        RECT 16.950 736.950 19.050 739.050 ;
        RECT 13.950 733.950 16.050 736.050 ;
        RECT 17.400 733.050 18.450 736.950 ;
        RECT 16.950 730.950 19.050 733.050 ;
        RECT 10.950 705.450 13.050 706.050 ;
        RECT 8.400 704.400 13.050 705.450 ;
        RECT 16.950 705.450 19.050 706.050 ;
        RECT 8.400 676.050 9.450 704.400 ;
        RECT 10.950 703.950 13.050 704.400 ;
        RECT 14.250 704.250 15.750 705.150 ;
        RECT 16.950 704.400 21.450 705.450 ;
        RECT 16.950 703.950 19.050 704.400 ;
        RECT 10.950 701.850 12.750 702.750 ;
        RECT 13.950 700.950 16.050 703.050 ;
        RECT 17.250 701.850 19.050 702.750 ;
        RECT 7.950 673.950 10.050 676.050 ;
        RECT 8.400 666.450 9.450 673.950 ;
        RECT 10.950 668.250 12.750 669.150 ;
        RECT 13.950 667.950 16.050 670.050 ;
        RECT 17.250 668.250 19.050 669.150 ;
        RECT 10.950 666.450 13.050 667.050 ;
        RECT 8.400 665.400 13.050 666.450 ;
        RECT 14.250 665.850 15.750 666.750 ;
        RECT 10.950 664.950 13.050 665.400 ;
        RECT 16.950 664.950 19.050 667.050 ;
        RECT 17.400 655.050 18.450 664.950 ;
        RECT 16.950 652.950 19.050 655.050 ;
        RECT 20.400 634.050 21.450 704.400 ;
        RECT 13.950 631.950 16.050 634.050 ;
        RECT 19.950 631.950 22.050 634.050 ;
        RECT 14.400 631.050 15.450 631.950 ;
        RECT 13.950 628.950 16.050 631.050 ;
        RECT 19.950 628.950 22.050 631.050 ;
        RECT 13.950 626.850 16.050 627.750 ;
        RECT 16.950 626.250 19.050 627.150 ;
        RECT 16.950 622.950 19.050 625.050 ;
        RECT 13.950 603.450 16.050 604.050 ;
        RECT 13.950 602.400 18.450 603.450 ;
        RECT 13.950 601.950 16.050 602.400 ;
        RECT 10.950 599.250 13.050 600.150 ;
        RECT 13.950 599.850 16.050 600.750 ;
        RECT 10.950 595.950 13.050 598.050 ;
        RECT 13.950 557.250 16.050 558.150 ;
        RECT 13.950 555.450 16.050 556.050 ;
        RECT 17.400 555.450 18.450 602.400 ;
        RECT 20.400 588.450 21.450 628.950 ;
        RECT 23.400 592.050 24.450 739.950 ;
        RECT 26.400 739.050 27.450 778.950 ;
        RECT 29.400 778.050 30.450 814.950 ;
        RECT 32.400 814.050 33.450 845.400 ;
        RECT 34.950 844.950 37.050 845.400 ;
        RECT 38.250 845.250 40.050 846.150 ;
        RECT 34.950 842.850 36.750 843.750 ;
        RECT 37.950 841.950 40.050 844.050 ;
        RECT 38.400 820.050 39.450 841.950 ;
        RECT 37.950 817.950 40.050 820.050 ;
        RECT 41.400 817.050 42.450 850.950 ;
        RECT 43.950 844.950 46.050 847.050 ;
        RECT 43.950 842.850 46.050 843.750 ;
        RECT 47.400 817.050 48.450 880.950 ;
        RECT 65.400 876.600 66.600 893.400 ;
        RECT 70.950 886.950 73.050 889.050 ;
        RECT 76.950 886.950 79.050 889.050 ;
        RECT 70.950 884.850 73.050 885.750 ;
        RECT 76.950 884.850 79.050 885.750 ;
        RECT 86.250 881.400 87.450 893.400 ;
        RECT 88.950 890.250 91.050 891.150 ;
        RECT 88.950 886.950 91.050 889.050 ;
        RECT 89.400 883.050 90.450 886.950 ;
        RECT 100.950 884.250 102.750 885.150 ;
        RECT 103.950 883.950 106.050 886.050 ;
        RECT 107.250 884.250 109.050 885.150 ;
        RECT 121.950 884.250 123.750 885.150 ;
        RECT 124.950 883.950 127.050 886.050 ;
        RECT 128.250 884.250 130.050 885.150 ;
        RECT 85.950 879.300 88.050 881.400 ;
        RECT 88.950 880.950 91.050 883.050 ;
        RECT 100.950 880.950 103.050 883.050 ;
        RECT 104.250 881.850 105.750 882.750 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 125.250 881.850 126.750 882.750 ;
        RECT 127.950 880.950 130.050 883.050 ;
        RECT 101.400 880.050 102.450 880.950 ;
        RECT 64.950 874.500 67.050 876.600 ;
        RECT 86.250 875.700 87.450 879.300 ;
        RECT 100.950 877.950 103.050 880.050 ;
        RECT 85.950 873.600 88.050 875.700 ;
        RECT 107.400 871.050 108.450 880.950 ;
        RECT 106.950 868.950 109.050 871.050 ;
        RECT 128.400 868.050 129.450 880.950 ;
        RECT 137.400 876.600 138.600 893.400 ;
        RECT 142.950 888.450 145.050 889.050 ;
        RECT 148.950 888.450 151.050 889.050 ;
        RECT 142.950 887.400 147.450 888.450 ;
        RECT 142.950 886.950 145.050 887.400 ;
        RECT 142.950 884.850 145.050 885.750 ;
        RECT 146.400 882.450 147.450 887.400 ;
        RECT 148.950 887.400 153.450 888.450 ;
        RECT 148.950 886.950 151.050 887.400 ;
        RECT 148.950 884.850 151.050 885.750 ;
        RECT 146.400 881.400 150.450 882.450 ;
        RECT 136.950 874.500 139.050 876.600 ;
        RECT 127.950 865.950 130.050 868.050 ;
        RECT 133.950 854.400 136.050 856.500 ;
        RECT 61.950 850.950 64.050 853.050 ;
        RECT 91.950 850.950 94.050 853.050 ;
        RECT 124.950 850.950 127.050 853.050 ;
        RECT 62.400 847.050 63.450 850.950 ;
        RECT 67.950 848.250 70.050 849.150 ;
        RECT 82.950 847.950 85.050 850.050 ;
        RECT 83.400 847.050 84.450 847.950 ;
        RECT 58.950 845.250 60.750 846.150 ;
        RECT 61.950 844.950 64.050 847.050 ;
        RECT 65.250 845.250 66.750 846.150 ;
        RECT 67.950 844.950 70.050 847.050 ;
        RECT 82.950 844.950 85.050 847.050 ;
        RECT 58.950 841.950 61.050 844.050 ;
        RECT 62.250 842.850 63.750 843.750 ;
        RECT 64.950 841.950 67.050 844.050 ;
        RECT 58.950 817.950 61.050 820.050 ;
        RECT 64.950 817.950 67.050 820.050 ;
        RECT 34.950 814.950 37.050 817.050 ;
        RECT 38.250 815.250 39.750 816.150 ;
        RECT 40.950 814.950 43.050 817.050 ;
        RECT 46.950 816.450 49.050 817.050 ;
        RECT 44.250 815.250 45.750 816.150 ;
        RECT 46.950 815.400 51.450 816.450 ;
        RECT 58.950 815.850 61.050 816.750 ;
        RECT 46.950 814.950 49.050 815.400 ;
        RECT 50.400 814.050 51.450 815.400 ;
        RECT 61.950 815.250 64.050 816.150 ;
        RECT 31.950 811.950 34.050 814.050 ;
        RECT 34.950 812.850 36.750 813.750 ;
        RECT 37.950 811.950 40.050 814.050 ;
        RECT 41.250 812.850 42.750 813.750 ;
        RECT 43.950 811.950 46.050 814.050 ;
        RECT 47.250 812.850 49.050 813.750 ;
        RECT 49.950 811.950 52.050 814.050 ;
        RECT 61.950 811.950 64.050 814.050 ;
        RECT 31.950 805.950 34.050 808.050 ;
        RECT 28.950 775.950 31.050 778.050 ;
        RECT 29.400 742.050 30.450 775.950 ;
        RECT 32.400 775.050 33.450 805.950 ;
        RECT 38.400 781.050 39.450 811.950 ;
        RECT 44.400 811.050 45.450 811.950 ;
        RECT 43.950 808.950 46.050 811.050 ;
        RECT 37.950 778.950 40.050 781.050 ;
        RECT 31.950 772.950 34.050 775.050 ;
        RECT 37.950 773.250 40.050 774.150 ;
        RECT 31.950 770.850 34.050 771.750 ;
        RECT 37.950 769.950 40.050 772.050 ;
        RECT 41.250 770.250 43.050 771.150 ;
        RECT 38.400 769.050 39.450 769.950 ;
        RECT 37.950 766.950 40.050 769.050 ;
        RECT 40.950 766.950 43.050 769.050 ;
        RECT 38.400 745.050 39.450 766.950 ;
        RECT 41.400 763.050 42.450 766.950 ;
        RECT 40.950 760.950 43.050 763.050 ;
        RECT 37.950 742.950 40.050 745.050 ;
        RECT 38.400 742.050 39.450 742.950 ;
        RECT 28.950 739.950 31.050 742.050 ;
        RECT 31.950 739.950 34.050 742.050 ;
        RECT 37.950 739.950 40.050 742.050 ;
        RECT 41.250 740.250 43.050 741.150 ;
        RECT 25.950 736.950 28.050 739.050 ;
        RECT 31.950 737.850 33.750 738.750 ;
        RECT 34.950 736.950 37.050 739.050 ;
        RECT 38.250 737.850 39.750 738.750 ;
        RECT 40.950 736.950 43.050 739.050 ;
        RECT 26.400 631.050 27.450 736.950 ;
        RECT 44.400 736.050 45.450 808.950 ;
        RECT 55.950 772.950 58.050 775.050 ;
        RECT 65.400 772.050 66.450 817.950 ;
        RECT 68.400 811.050 69.450 844.950 ;
        RECT 79.950 842.250 82.050 843.150 ;
        RECT 82.950 842.850 85.050 843.750 ;
        RECT 79.950 838.950 82.050 841.050 ;
        RECT 80.400 814.050 81.450 838.950 ;
        RECT 88.950 820.950 91.050 823.050 ;
        RECT 82.950 817.950 85.050 820.050 ;
        RECT 83.400 817.050 84.450 817.950 ;
        RECT 89.400 817.050 90.450 820.950 ;
        RECT 92.400 820.050 93.450 850.950 ;
        RECT 125.400 850.050 126.450 850.950 ;
        RECT 97.950 847.950 100.050 850.050 ;
        RECT 103.950 849.450 106.050 850.050 ;
        RECT 101.250 848.250 102.750 849.150 ;
        RECT 103.950 848.400 108.450 849.450 ;
        RECT 103.950 847.950 106.050 848.400 ;
        RECT 97.950 845.850 99.750 846.750 ;
        RECT 100.950 844.950 103.050 847.050 ;
        RECT 104.250 845.850 106.050 846.750 ;
        RECT 107.400 841.050 108.450 848.400 ;
        RECT 118.950 847.950 121.050 850.050 ;
        RECT 122.250 848.250 123.750 849.150 ;
        RECT 124.950 847.950 127.050 850.050 ;
        RECT 118.950 845.850 120.750 846.750 ;
        RECT 121.950 844.950 124.050 847.050 ;
        RECT 125.250 845.850 127.050 846.750 ;
        RECT 100.950 838.950 103.050 841.050 ;
        RECT 106.950 838.950 109.050 841.050 ;
        RECT 97.950 820.950 100.050 823.050 ;
        RECT 91.950 817.950 94.050 820.050 ;
        RECT 82.950 814.950 85.050 817.050 ;
        RECT 86.250 815.250 87.750 816.150 ;
        RECT 88.950 814.950 91.050 817.050 ;
        RECT 79.950 813.450 82.050 814.050 ;
        RECT 77.400 812.400 82.050 813.450 ;
        RECT 83.250 812.850 84.750 813.750 ;
        RECT 67.950 808.950 70.050 811.050 ;
        RECT 77.400 808.050 78.450 812.400 ;
        RECT 79.950 811.950 82.050 812.400 ;
        RECT 85.950 811.950 88.050 814.050 ;
        RECT 89.250 812.850 91.050 813.750 ;
        RECT 79.950 809.850 82.050 810.750 ;
        RECT 67.950 805.950 70.050 808.050 ;
        RECT 76.950 805.950 79.050 808.050 ;
        RECT 52.950 770.250 55.050 771.150 ;
        RECT 55.950 770.850 58.050 771.750 ;
        RECT 64.950 769.950 67.050 772.050 ;
        RECT 52.950 766.950 55.050 769.050 ;
        RECT 68.400 768.450 69.450 805.950 ;
        RECT 70.950 773.250 72.750 774.150 ;
        RECT 73.950 772.950 76.050 775.050 ;
        RECT 79.950 774.450 82.050 775.050 ;
        RECT 79.950 773.400 84.450 774.450 ;
        RECT 79.950 772.950 82.050 773.400 ;
        RECT 70.950 769.950 73.050 772.050 ;
        RECT 74.250 770.850 76.050 771.750 ;
        RECT 76.950 770.250 79.050 771.150 ;
        RECT 79.950 770.850 82.050 771.750 ;
        RECT 68.400 767.400 72.450 768.450 ;
        RECT 58.950 760.950 61.050 763.050 ;
        RECT 67.950 760.950 70.050 763.050 ;
        RECT 59.400 742.050 60.450 760.950 ;
        RECT 64.950 745.950 67.050 748.050 ;
        RECT 52.950 739.950 55.050 742.050 ;
        RECT 55.950 740.250 57.750 741.150 ;
        RECT 58.950 739.950 61.050 742.050 ;
        RECT 62.250 740.250 64.050 741.150 ;
        RECT 53.400 738.450 54.450 739.950 ;
        RECT 55.950 738.450 58.050 739.050 ;
        RECT 53.400 737.400 58.050 738.450 ;
        RECT 59.250 737.850 60.750 738.750 ;
        RECT 61.950 738.450 64.050 739.050 ;
        RECT 65.400 738.450 66.450 745.950 ;
        RECT 68.400 742.050 69.450 760.950 ;
        RECT 67.950 739.950 70.050 742.050 ;
        RECT 55.950 736.950 58.050 737.400 ;
        RECT 61.950 737.400 66.450 738.450 ;
        RECT 71.400 738.450 72.450 767.400 ;
        RECT 76.950 766.950 79.050 769.050 ;
        RECT 77.400 763.050 78.450 766.950 ;
        RECT 76.950 760.950 79.050 763.050 ;
        RECT 83.400 748.050 84.450 773.400 ;
        RECT 76.950 745.950 79.050 748.050 ;
        RECT 82.950 745.950 85.050 748.050 ;
        RECT 73.950 743.250 76.050 744.150 ;
        RECT 76.950 743.850 79.050 744.750 ;
        RECT 82.950 744.450 85.050 745.050 ;
        RECT 86.400 744.450 87.450 811.950 ;
        RECT 92.400 775.050 93.450 817.950 ;
        RECT 98.400 817.050 99.450 820.950 ;
        RECT 101.400 820.050 102.450 838.950 ;
        RECT 134.400 837.600 135.600 854.400 ;
        RECT 142.950 850.950 145.050 853.050 ;
        RECT 136.950 847.950 139.050 850.050 ;
        RECT 133.950 835.500 136.050 837.600 ;
        RECT 100.950 817.950 103.050 820.050 ;
        RECT 97.950 814.950 100.050 817.050 ;
        RECT 101.250 815.850 102.750 816.750 ;
        RECT 103.950 814.950 106.050 817.050 ;
        RECT 133.950 814.950 136.050 817.050 ;
        RECT 97.950 812.850 100.050 813.750 ;
        RECT 103.950 812.850 106.050 813.750 ;
        RECT 121.950 812.250 123.750 813.150 ;
        RECT 124.950 811.950 127.050 814.050 ;
        RECT 128.250 812.250 130.050 813.150 ;
        RECT 121.950 810.450 124.050 811.050 ;
        RECT 119.400 809.400 124.050 810.450 ;
        RECT 125.250 809.850 126.750 810.750 ;
        RECT 100.950 781.950 103.050 784.050 ;
        RECT 94.950 775.950 97.050 778.050 ;
        RECT 95.400 775.050 96.450 775.950 ;
        RECT 88.950 774.450 91.050 775.050 ;
        RECT 91.950 774.450 94.050 775.050 ;
        RECT 88.950 773.400 94.050 774.450 ;
        RECT 88.950 772.950 91.050 773.400 ;
        RECT 91.950 772.950 94.050 773.400 ;
        RECT 94.950 772.950 97.050 775.050 ;
        RECT 98.250 773.250 100.050 774.150 ;
        RECT 88.950 770.850 91.050 771.750 ;
        RECT 91.950 770.250 94.050 771.150 ;
        RECT 94.950 770.850 96.750 771.750 ;
        RECT 97.950 771.450 100.050 772.050 ;
        RECT 101.400 771.450 102.450 781.950 ;
        RECT 112.950 779.250 115.050 780.150 ;
        RECT 119.400 778.050 120.450 809.400 ;
        RECT 121.950 808.950 124.050 809.400 ;
        RECT 127.950 808.950 130.050 811.050 ;
        RECT 106.950 775.950 109.050 778.050 ;
        RECT 109.950 776.250 111.750 777.150 ;
        RECT 112.950 775.950 115.050 778.050 ;
        RECT 116.250 776.250 117.750 777.150 ;
        RECT 118.950 775.950 121.050 778.050 ;
        RECT 97.950 770.400 102.450 771.450 ;
        RECT 97.950 769.950 100.050 770.400 ;
        RECT 91.950 766.950 94.050 769.050 ;
        RECT 79.950 743.250 81.750 744.150 ;
        RECT 82.950 743.400 87.450 744.450 ;
        RECT 82.950 742.950 85.050 743.400 ;
        RECT 73.950 739.950 76.050 742.050 ;
        RECT 79.950 739.950 82.050 742.050 ;
        RECT 83.250 740.850 85.050 741.750 ;
        RECT 80.400 739.050 81.450 739.950 ;
        RECT 71.400 737.400 75.450 738.450 ;
        RECT 61.950 736.950 64.050 737.400 ;
        RECT 31.950 733.950 34.050 736.050 ;
        RECT 34.950 734.850 37.050 735.750 ;
        RECT 43.950 733.950 46.050 736.050 ;
        RECT 28.950 730.950 31.050 733.050 ;
        RECT 29.400 673.050 30.450 730.950 ;
        RECT 32.400 706.050 33.450 733.950 ;
        RECT 37.950 707.250 40.050 708.150 ;
        RECT 31.950 703.950 34.050 706.050 ;
        RECT 35.250 704.250 36.750 705.150 ;
        RECT 37.950 703.950 40.050 706.050 ;
        RECT 41.250 704.250 43.050 705.150 ;
        RECT 64.950 703.950 67.050 706.050 ;
        RECT 70.950 703.950 73.050 706.050 ;
        RECT 31.950 701.850 33.750 702.750 ;
        RECT 34.950 700.950 37.050 703.050 ;
        RECT 38.400 673.050 39.450 703.950 ;
        RECT 40.950 700.950 43.050 703.050 ;
        RECT 52.950 700.950 55.050 703.050 ;
        RECT 41.400 673.050 42.450 700.950 ;
        RECT 52.950 698.850 55.050 699.750 ;
        RECT 55.950 698.250 58.050 699.150 ;
        RECT 55.950 694.950 58.050 697.050 ;
        RECT 52.950 673.950 55.050 676.050 ;
        RECT 53.400 673.050 54.450 673.950 ;
        RECT 28.950 670.950 31.050 673.050 ;
        RECT 37.950 670.950 40.050 673.050 ;
        RECT 40.950 670.950 43.050 673.050 ;
        RECT 52.950 670.950 55.050 673.050 ;
        RECT 58.950 672.450 61.050 673.050 ;
        RECT 56.250 671.250 57.750 672.150 ;
        RECT 58.950 671.400 63.450 672.450 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 28.950 668.250 30.750 669.150 ;
        RECT 31.950 667.950 34.050 670.050 ;
        RECT 37.950 669.450 40.050 670.050 ;
        RECT 49.950 669.450 52.050 670.050 ;
        RECT 37.950 668.400 42.450 669.450 ;
        RECT 37.950 667.950 40.050 668.400 ;
        RECT 28.950 664.950 31.050 667.050 ;
        RECT 32.250 665.850 33.750 666.750 ;
        RECT 34.950 664.950 37.050 667.050 ;
        RECT 38.250 665.850 40.050 666.750 ;
        RECT 41.400 664.050 42.450 668.400 ;
        RECT 47.400 668.400 52.050 669.450 ;
        RECT 53.250 668.850 54.750 669.750 ;
        RECT 43.950 664.950 46.050 667.050 ;
        RECT 28.950 661.950 31.050 664.050 ;
        RECT 34.950 662.850 37.050 663.750 ;
        RECT 40.950 661.950 43.050 664.050 ;
        RECT 25.950 628.950 28.050 631.050 ;
        RECT 29.400 628.050 30.450 661.950 ;
        RECT 44.400 661.050 45.450 664.950 ;
        RECT 31.950 658.950 34.050 661.050 ;
        RECT 43.950 658.950 46.050 661.050 ;
        RECT 32.400 634.050 33.450 658.950 ;
        RECT 43.950 652.950 46.050 655.050 ;
        RECT 37.950 635.250 40.050 636.150 ;
        RECT 44.400 634.050 45.450 652.950 ;
        RECT 31.950 631.950 34.050 634.050 ;
        RECT 35.250 632.250 36.750 633.150 ;
        RECT 37.950 631.950 40.050 634.050 ;
        RECT 41.250 632.250 43.050 633.150 ;
        RECT 43.950 631.950 46.050 634.050 ;
        RECT 31.950 629.850 33.750 630.750 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 37.950 628.950 40.050 631.050 ;
        RECT 40.950 628.950 43.050 631.050 ;
        RECT 28.950 625.950 31.050 628.050 ;
        RECT 34.950 625.950 37.050 628.050 ;
        RECT 28.950 601.950 31.050 604.050 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 25.950 599.250 28.050 600.150 ;
        RECT 28.950 599.850 31.050 600.750 ;
        RECT 25.950 595.950 28.050 598.050 ;
        RECT 22.950 589.950 25.050 592.050 ;
        RECT 20.400 587.400 24.450 588.450 ;
        RECT 19.950 556.950 22.050 559.050 ;
        RECT 10.950 554.250 12.750 555.150 ;
        RECT 13.950 554.400 18.450 555.450 ;
        RECT 19.950 554.850 22.050 555.750 ;
        RECT 13.950 553.950 16.050 554.400 ;
        RECT 10.950 550.950 13.050 553.050 ;
        RECT 14.400 541.050 15.450 553.950 ;
        RECT 13.950 538.950 16.050 541.050 ;
        RECT 7.950 533.400 10.050 535.500 ;
        RECT 8.400 516.600 9.600 533.400 ;
        RECT 13.950 526.950 16.050 529.050 ;
        RECT 19.950 528.450 22.050 529.050 ;
        RECT 17.400 527.400 22.050 528.450 ;
        RECT 13.950 524.850 16.050 525.750 ;
        RECT 7.950 514.500 10.050 516.600 ;
        RECT 17.400 498.450 18.450 527.400 ;
        RECT 19.950 526.950 22.050 527.400 ;
        RECT 19.950 524.850 22.050 525.750 ;
        RECT 17.400 497.400 21.450 498.450 ;
        RECT 10.950 485.250 13.050 486.150 ;
        RECT 16.950 485.250 19.050 486.150 ;
        RECT 10.950 481.950 13.050 484.050 ;
        RECT 14.250 482.250 15.750 483.150 ;
        RECT 16.950 481.950 19.050 484.050 ;
        RECT 11.400 472.050 12.450 481.950 ;
        RECT 13.950 478.950 16.050 481.050 ;
        RECT 10.950 469.950 13.050 472.050 ;
        RECT 14.400 463.050 15.450 478.950 ;
        RECT 17.400 475.050 18.450 481.950 ;
        RECT 16.950 472.950 19.050 475.050 ;
        RECT 20.400 469.050 21.450 497.400 ;
        RECT 19.950 466.950 22.050 469.050 ;
        RECT 7.950 460.950 10.050 463.050 ;
        RECT 13.950 460.950 16.050 463.050 ;
        RECT 8.400 457.050 9.450 460.950 ;
        RECT 23.400 460.050 24.450 587.400 ;
        RECT 26.400 532.050 27.450 595.950 ;
        RECT 32.400 538.050 33.450 601.950 ;
        RECT 35.400 598.050 36.450 625.950 ;
        RECT 38.400 604.050 39.450 628.950 ;
        RECT 41.400 619.050 42.450 628.950 ;
        RECT 44.400 625.050 45.450 631.950 ;
        RECT 43.950 622.950 46.050 625.050 ;
        RECT 40.950 616.950 43.050 619.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 37.950 599.850 39.750 600.750 ;
        RECT 40.950 600.450 43.050 601.050 ;
        RECT 44.400 600.450 45.450 622.950 ;
        RECT 47.400 619.050 48.450 668.400 ;
        RECT 49.950 667.950 52.050 668.400 ;
        RECT 55.950 667.950 58.050 670.050 ;
        RECT 59.250 668.850 61.050 669.750 ;
        RECT 49.950 665.850 52.050 666.750 ;
        RECT 52.950 664.950 55.050 667.050 ;
        RECT 53.400 634.050 54.450 664.950 ;
        RECT 56.400 649.050 57.450 667.950 ;
        RECT 62.400 667.050 63.450 671.400 ;
        RECT 61.950 664.950 64.050 667.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 635.250 61.050 636.150 ;
        RECT 52.950 631.950 55.050 634.050 ;
        RECT 56.250 632.250 57.750 633.150 ;
        RECT 58.950 631.950 61.050 634.050 ;
        RECT 62.250 632.250 64.050 633.150 ;
        RECT 52.950 629.850 54.750 630.750 ;
        RECT 55.950 628.950 58.050 631.050 ;
        RECT 56.400 625.050 57.450 628.950 ;
        RECT 59.400 628.050 60.450 631.950 ;
        RECT 61.950 628.950 64.050 631.050 ;
        RECT 58.950 625.950 61.050 628.050 ;
        RECT 55.950 622.950 58.050 625.050 ;
        RECT 62.400 619.050 63.450 628.950 ;
        RECT 65.400 622.050 66.450 703.950 ;
        RECT 67.950 701.250 70.050 702.150 ;
        RECT 70.950 701.850 73.050 702.750 ;
        RECT 74.400 700.050 75.450 737.400 ;
        RECT 79.950 736.950 82.050 739.050 ;
        RECT 92.400 736.050 93.450 766.950 ;
        RECT 100.950 760.950 103.050 763.050 ;
        RECT 101.400 745.050 102.450 760.950 ;
        RECT 100.950 742.950 103.050 745.050 ;
        RECT 100.950 740.850 103.050 741.750 ;
        RECT 103.950 740.250 106.050 741.150 ;
        RECT 103.950 736.950 106.050 739.050 ;
        RECT 104.400 736.050 105.450 736.950 ;
        RECT 79.950 733.950 82.050 736.050 ;
        RECT 91.950 733.950 94.050 736.050 ;
        RECT 103.950 733.950 106.050 736.050 ;
        RECT 76.950 701.250 79.050 702.150 ;
        RECT 67.950 697.950 70.050 700.050 ;
        RECT 73.950 697.950 76.050 700.050 ;
        RECT 76.950 699.450 79.050 700.050 ;
        RECT 80.400 699.450 81.450 733.950 ;
        RECT 94.950 704.250 97.050 705.150 ;
        RECT 85.950 701.250 87.750 702.150 ;
        RECT 88.950 700.950 91.050 703.050 ;
        RECT 92.250 701.250 93.750 702.150 ;
        RECT 94.950 700.950 97.050 703.050 ;
        RECT 76.950 698.400 81.450 699.450 ;
        RECT 76.950 697.950 79.050 698.400 ;
        RECT 85.950 697.950 88.050 700.050 ;
        RECT 89.250 698.850 90.750 699.750 ;
        RECT 91.950 697.950 94.050 700.050 ;
        RECT 67.950 673.950 70.050 676.050 ;
        RECT 73.950 673.950 76.050 676.050 ;
        RECT 67.950 671.850 70.050 672.750 ;
        RECT 70.950 671.250 73.050 672.150 ;
        RECT 70.950 667.950 73.050 670.050 ;
        RECT 71.400 667.050 72.450 667.950 ;
        RECT 70.950 664.950 73.050 667.050 ;
        RECT 74.400 634.050 75.450 673.950 ;
        RECT 77.400 643.050 78.450 697.950 ;
        RECT 79.950 694.950 82.050 697.050 ;
        RECT 80.400 664.050 81.450 694.950 ;
        RECT 86.400 694.050 87.450 697.950 ;
        RECT 85.950 691.950 88.050 694.050 ;
        RECT 82.950 670.950 85.050 673.050 ;
        RECT 95.400 672.450 96.450 700.950 ;
        RECT 104.400 700.050 105.450 733.950 ;
        RECT 103.950 697.950 106.050 700.050 ;
        RECT 107.400 697.050 108.450 775.950 ;
        RECT 109.950 772.950 112.050 775.050 ;
        RECT 115.950 772.950 118.050 775.050 ;
        RECT 119.250 773.850 121.050 774.750 ;
        RECT 110.400 769.050 111.450 772.950 ;
        RECT 115.950 769.950 118.050 772.050 ;
        RECT 109.950 766.950 112.050 769.050 ;
        RECT 109.950 742.950 112.050 745.050 ;
        RECT 109.950 740.850 112.050 741.750 ;
        RECT 116.400 738.450 117.450 769.950 ;
        RECT 121.950 742.950 124.050 745.050 ;
        RECT 122.400 742.050 123.450 742.950 ;
        RECT 118.950 740.250 120.750 741.150 ;
        RECT 121.950 739.950 124.050 742.050 ;
        RECT 125.250 740.250 127.050 741.150 ;
        RECT 118.950 738.450 121.050 739.050 ;
        RECT 116.400 737.400 121.050 738.450 ;
        RECT 122.250 737.850 123.750 738.750 ;
        RECT 112.950 703.950 115.050 706.050 ;
        RECT 113.400 703.050 114.450 703.950 ;
        RECT 116.400 703.050 117.450 737.400 ;
        RECT 118.950 736.950 121.050 737.400 ;
        RECT 124.950 736.950 127.050 739.050 ;
        RECT 109.950 701.250 111.750 702.150 ;
        RECT 112.950 700.950 115.050 703.050 ;
        RECT 115.950 700.950 118.050 703.050 ;
        RECT 118.950 702.450 121.050 703.050 ;
        RECT 118.950 701.400 123.450 702.450 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 122.400 700.050 123.450 701.400 ;
        RECT 109.950 697.950 112.050 700.050 ;
        RECT 113.250 698.850 115.050 699.750 ;
        RECT 115.950 698.250 118.050 699.150 ;
        RECT 118.950 698.850 121.050 699.750 ;
        RECT 121.950 697.950 124.050 700.050 ;
        RECT 106.950 694.950 109.050 697.050 ;
        RECT 112.950 694.950 115.050 697.050 ;
        RECT 115.950 694.950 118.050 697.050 ;
        RECT 125.400 696.450 126.450 736.950 ;
        RECT 128.400 718.050 129.450 808.950 ;
        RECT 134.400 784.050 135.450 814.950 ;
        RECT 137.400 811.050 138.450 847.950 ;
        RECT 143.400 847.050 144.450 850.950 ;
        RECT 139.950 845.250 142.050 846.150 ;
        RECT 142.950 844.950 145.050 847.050 ;
        RECT 145.950 845.250 148.050 846.150 ;
        RECT 149.400 844.050 150.450 881.400 ;
        RECT 139.950 841.950 142.050 844.050 ;
        RECT 145.950 841.950 148.050 844.050 ;
        RECT 148.950 841.950 151.050 844.050 ;
        RECT 140.400 838.050 141.450 841.950 ;
        RECT 146.400 841.050 147.450 841.950 ;
        RECT 152.400 841.050 153.450 887.400 ;
        RECT 158.250 881.400 159.450 893.400 ;
        RECT 160.950 890.250 163.050 891.150 ;
        RECT 175.950 889.950 178.050 892.050 ;
        RECT 160.950 886.950 163.050 889.050 ;
        RECT 175.950 887.850 178.050 888.750 ;
        RECT 178.950 887.250 181.050 888.150 ;
        RECT 178.950 883.950 181.050 886.050 ;
        RECT 196.950 884.250 198.750 885.150 ;
        RECT 199.950 883.950 202.050 886.050 ;
        RECT 203.250 884.250 205.050 885.150 ;
        RECT 179.400 883.050 180.450 883.950 ;
        RECT 157.950 879.300 160.050 881.400 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 187.950 880.950 190.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 200.250 881.850 201.750 882.750 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 158.250 875.700 159.450 879.300 ;
        RECT 157.950 873.600 160.050 875.700 ;
        RECT 178.950 865.950 181.050 868.050 ;
        RECT 154.950 855.300 157.050 857.400 ;
        RECT 155.250 851.700 156.450 855.300 ;
        RECT 154.950 849.600 157.050 851.700 ;
        RECT 145.950 838.950 148.050 841.050 ;
        RECT 151.950 838.950 154.050 841.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 155.250 837.600 156.450 849.600 ;
        RECT 172.950 848.250 175.050 849.150 ;
        RECT 179.400 847.050 180.450 865.950 ;
        RECT 172.950 844.950 175.050 847.050 ;
        RECT 176.250 845.250 177.750 846.150 ;
        RECT 178.950 844.950 181.050 847.050 ;
        RECT 182.250 845.250 184.050 846.150 ;
        RECT 184.950 844.950 187.050 847.050 ;
        RECT 157.950 843.450 160.050 844.050 ;
        RECT 157.950 842.400 162.450 843.450 ;
        RECT 157.950 841.950 160.050 842.400 ;
        RECT 157.950 839.850 160.050 840.750 ;
        RECT 146.400 817.050 147.450 835.950 ;
        RECT 154.950 835.500 157.050 837.600 ;
        RECT 161.400 820.050 162.450 842.400 ;
        RECT 172.950 841.950 175.050 844.050 ;
        RECT 175.950 841.950 178.050 844.050 ;
        RECT 179.250 842.850 180.750 843.750 ;
        RECT 181.950 841.950 184.050 844.050 ;
        RECT 160.950 817.950 163.050 820.050 ;
        RECT 173.400 817.050 174.450 841.950 ;
        RECT 178.950 835.950 181.050 838.050 ;
        RECT 179.400 817.050 180.450 835.950 ;
        RECT 139.950 814.950 142.050 817.050 ;
        RECT 143.250 815.250 144.750 816.150 ;
        RECT 145.950 814.950 148.050 817.050 ;
        RECT 151.950 816.450 154.050 817.050 ;
        RECT 149.250 815.250 150.750 816.150 ;
        RECT 151.950 815.400 156.450 816.450 ;
        RECT 151.950 814.950 154.050 815.400 ;
        RECT 139.950 812.850 141.750 813.750 ;
        RECT 142.950 811.950 145.050 814.050 ;
        RECT 146.250 812.850 147.750 813.750 ;
        RECT 148.950 811.950 151.050 814.050 ;
        RECT 152.250 812.850 154.050 813.750 ;
        RECT 136.950 808.950 139.050 811.050 ;
        RECT 133.950 781.950 136.050 784.050 ;
        RECT 149.400 778.050 150.450 811.950 ;
        RECT 155.400 811.050 156.450 815.400 ;
        RECT 157.950 814.950 160.050 817.050 ;
        RECT 166.950 814.950 169.050 817.050 ;
        RECT 170.250 815.250 171.750 816.150 ;
        RECT 172.950 814.950 175.050 817.050 ;
        RECT 176.250 815.250 177.750 816.150 ;
        RECT 178.950 814.950 181.050 817.050 ;
        RECT 154.950 808.950 157.050 811.050 ;
        RECT 148.950 775.950 151.050 778.050 ;
        RECT 158.400 775.050 159.450 814.950 ;
        RECT 182.400 814.050 183.450 841.950 ;
        RECT 166.950 812.850 168.750 813.750 ;
        RECT 169.950 811.950 172.050 814.050 ;
        RECT 173.250 812.850 174.750 813.750 ;
        RECT 175.950 811.950 178.050 814.050 ;
        RECT 179.250 812.850 181.050 813.750 ;
        RECT 181.950 811.950 184.050 814.050 ;
        RECT 170.400 799.050 171.450 811.950 ;
        RECT 176.400 808.050 177.450 811.950 ;
        RECT 175.950 805.950 178.050 808.050 ;
        RECT 169.950 796.950 172.050 799.050 ;
        RECT 181.950 796.950 184.050 799.050 ;
        RECT 130.950 773.250 133.050 774.150 ;
        RECT 136.950 773.250 139.050 774.150 ;
        RECT 151.950 773.250 154.050 774.150 ;
        RECT 157.950 772.950 160.050 775.050 ;
        RECT 169.950 774.450 172.050 775.050 ;
        RECT 167.400 773.400 172.050 774.450 ;
        RECT 130.950 769.950 133.050 772.050 ;
        RECT 134.250 770.250 135.750 771.150 ;
        RECT 136.950 769.950 139.050 772.050 ;
        RECT 148.950 770.250 150.750 771.150 ;
        RECT 151.950 769.950 154.050 772.050 ;
        RECT 157.950 770.850 160.050 771.750 ;
        RECT 133.950 766.950 136.050 769.050 ;
        RECT 137.400 766.050 138.450 769.950 ;
        RECT 148.950 766.950 151.050 769.050 ;
        RECT 136.950 763.950 139.050 766.050 ;
        RECT 152.400 765.450 153.450 769.950 ;
        RECT 167.400 769.050 168.450 773.400 ;
        RECT 169.950 772.950 172.050 773.400 ;
        RECT 175.950 772.950 178.050 775.050 ;
        RECT 179.250 773.250 181.050 774.150 ;
        RECT 169.950 770.850 172.050 771.750 ;
        RECT 172.950 770.250 175.050 771.150 ;
        RECT 175.950 770.850 177.750 771.750 ;
        RECT 178.950 771.450 181.050 772.050 ;
        RECT 182.400 771.450 183.450 796.950 ;
        RECT 185.400 778.050 186.450 844.950 ;
        RECT 188.400 838.050 189.450 880.950 ;
        RECT 197.400 880.050 198.450 880.950 ;
        RECT 196.950 877.950 199.050 880.050 ;
        RECT 203.400 871.050 204.450 880.950 ;
        RECT 212.400 876.600 213.600 893.400 ;
        RECT 217.950 888.450 220.050 889.050 ;
        RECT 223.950 888.450 226.050 889.050 ;
        RECT 217.950 887.400 222.450 888.450 ;
        RECT 217.950 886.950 220.050 887.400 ;
        RECT 221.400 886.050 222.450 887.400 ;
        RECT 223.950 887.400 228.450 888.450 ;
        RECT 223.950 886.950 226.050 887.400 ;
        RECT 214.950 883.950 217.050 886.050 ;
        RECT 217.950 884.850 220.050 885.750 ;
        RECT 220.950 883.950 223.050 886.050 ;
        RECT 223.950 884.850 226.050 885.750 ;
        RECT 211.950 874.500 214.050 876.600 ;
        RECT 199.950 868.950 202.050 871.050 ;
        RECT 202.950 868.950 205.050 871.050 ;
        RECT 208.950 868.950 211.050 871.050 ;
        RECT 190.950 854.400 193.050 856.500 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 191.400 837.600 192.600 854.400 ;
        RECT 200.400 847.050 201.450 868.950 ;
        RECT 196.950 845.250 199.050 846.150 ;
        RECT 199.950 844.950 202.050 847.050 ;
        RECT 202.950 845.250 205.050 846.150 ;
        RECT 196.950 841.950 199.050 844.050 ;
        RECT 190.950 835.500 193.050 837.600 ;
        RECT 190.950 817.950 193.050 820.050 ;
        RECT 190.950 815.850 193.050 816.750 ;
        RECT 193.950 815.250 196.050 816.150 ;
        RECT 193.950 811.950 196.050 814.050 ;
        RECT 194.400 811.050 195.450 811.950 ;
        RECT 193.950 808.950 196.050 811.050 ;
        RECT 200.400 808.050 201.450 844.950 ;
        RECT 202.950 841.950 205.050 844.050 ;
        RECT 203.400 841.050 204.450 841.950 ;
        RECT 202.950 838.950 205.050 841.050 ;
        RECT 209.400 835.050 210.450 868.950 ;
        RECT 211.950 855.300 214.050 857.400 ;
        RECT 215.400 856.050 216.450 883.950 ;
        RECT 227.400 880.050 228.450 887.400 ;
        RECT 233.250 881.400 234.450 893.400 ;
        RECT 235.950 890.250 238.050 891.150 ;
        RECT 250.950 889.950 253.050 892.050 ;
        RECT 235.950 886.950 238.050 889.050 ;
        RECT 250.950 887.850 253.050 888.750 ;
        RECT 253.950 887.250 256.050 888.150 ;
        RECT 274.950 886.950 277.050 889.050 ;
        RECT 280.950 888.450 283.050 889.050 ;
        RECT 278.250 887.250 279.750 888.150 ;
        RECT 280.950 887.400 285.450 888.450 ;
        RECT 280.950 886.950 283.050 887.400 ;
        RECT 247.950 883.950 250.050 886.050 ;
        RECT 253.950 883.950 256.050 886.050 ;
        RECT 271.950 885.450 274.050 886.050 ;
        RECT 269.400 884.400 274.050 885.450 ;
        RECT 275.250 884.850 276.750 885.750 ;
        RECT 226.950 877.950 229.050 880.050 ;
        RECT 232.950 879.300 235.050 881.400 ;
        RECT 233.250 875.700 234.450 879.300 ;
        RECT 232.950 873.600 235.050 875.700 ;
        RECT 212.250 851.700 213.450 855.300 ;
        RECT 214.950 853.950 217.050 856.050 ;
        RECT 211.950 849.600 214.050 851.700 ;
        RECT 226.950 850.950 229.050 853.050 ;
        RECT 238.950 850.950 241.050 853.050 ;
        RECT 212.250 837.600 213.450 849.600 ;
        RECT 214.950 841.950 217.050 844.050 ;
        RECT 220.950 841.950 223.050 844.050 ;
        RECT 227.400 843.450 228.450 850.950 ;
        RECT 232.950 847.950 235.050 850.050 ;
        RECT 233.400 847.050 234.450 847.950 ;
        RECT 239.400 847.050 240.450 850.950 ;
        RECT 229.950 845.250 231.750 846.150 ;
        RECT 232.950 844.950 235.050 847.050 ;
        RECT 236.250 845.250 237.750 846.150 ;
        RECT 238.950 844.950 241.050 847.050 ;
        RECT 242.250 845.250 244.050 846.150 ;
        RECT 244.950 844.950 247.050 847.050 ;
        RECT 229.950 843.450 232.050 844.050 ;
        RECT 227.400 842.400 232.050 843.450 ;
        RECT 233.250 842.850 234.750 843.750 ;
        RECT 229.950 841.950 232.050 842.400 ;
        RECT 235.950 841.950 238.050 844.050 ;
        RECT 239.250 842.850 240.750 843.750 ;
        RECT 241.950 843.450 244.050 844.050 ;
        RECT 245.400 843.450 246.450 844.950 ;
        RECT 241.950 842.400 246.450 843.450 ;
        RECT 241.950 841.950 244.050 842.400 ;
        RECT 214.950 839.850 217.050 840.750 ;
        RECT 211.950 835.500 214.050 837.600 ;
        RECT 208.950 832.950 211.050 835.050 ;
        RECT 221.400 820.050 222.450 841.950 ;
        RECT 232.950 832.950 235.050 835.050 ;
        RECT 211.950 817.950 214.050 820.050 ;
        RECT 220.950 817.950 223.050 820.050 ;
        RECT 208.950 815.250 211.050 816.150 ;
        RECT 211.950 815.850 214.050 816.750 ;
        RECT 208.950 811.950 211.050 814.050 ;
        RECT 221.400 810.450 222.450 817.950 ;
        RECT 223.950 812.250 225.750 813.150 ;
        RECT 226.950 811.950 229.050 814.050 ;
        RECT 230.250 812.250 232.050 813.150 ;
        RECT 223.950 810.450 226.050 811.050 ;
        RECT 221.400 809.400 226.050 810.450 ;
        RECT 227.250 809.850 228.750 810.750 ;
        RECT 229.950 810.450 232.050 811.050 ;
        RECT 233.400 810.450 234.450 832.950 ;
        RECT 248.400 817.050 249.450 883.950 ;
        RECT 250.950 854.400 253.050 856.500 ;
        RECT 251.400 837.600 252.600 854.400 ;
        RECT 250.950 835.500 253.050 837.600 ;
        RECT 254.400 826.050 255.450 883.950 ;
        RECT 269.400 883.050 270.450 884.400 ;
        RECT 271.950 883.950 274.050 884.400 ;
        RECT 277.950 883.950 280.050 886.050 ;
        RECT 281.250 884.850 283.050 885.750 ;
        RECT 284.400 883.050 285.450 887.400 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 881.850 274.050 882.750 ;
        RECT 283.950 880.950 286.050 883.050 ;
        RECT 290.400 876.600 291.600 893.400 ;
        RECT 295.950 886.950 298.050 889.050 ;
        RECT 301.950 888.450 304.050 889.050 ;
        RECT 301.950 887.400 306.450 888.450 ;
        RECT 301.950 886.950 304.050 887.400 ;
        RECT 295.950 884.850 298.050 885.750 ;
        RECT 301.950 884.850 304.050 885.750 ;
        RECT 305.400 880.050 306.450 887.400 ;
        RECT 311.250 881.400 312.450 893.400 ;
        RECT 313.950 890.250 316.050 891.150 ;
        RECT 325.950 889.950 328.050 892.050 ;
        RECT 340.950 889.950 343.050 892.050 ;
        RECT 382.950 889.950 385.050 892.050 ;
        RECT 397.950 889.950 400.050 892.050 ;
        RECT 341.400 889.050 342.450 889.950 ;
        RECT 398.400 889.050 399.450 889.950 ;
        RECT 313.950 886.950 316.050 889.050 ;
        RECT 325.950 887.850 328.050 888.750 ;
        RECT 328.950 887.250 331.050 888.150 ;
        RECT 340.950 886.950 343.050 889.050 ;
        RECT 379.950 888.450 382.050 889.050 ;
        RECT 377.400 887.400 382.050 888.450 ;
        RECT 383.250 887.850 384.750 888.750 ;
        RECT 385.950 888.450 388.050 889.050 ;
        RECT 328.950 883.950 331.050 886.050 ;
        RECT 340.950 884.850 343.050 885.750 ;
        RECT 346.950 884.850 349.050 885.750 ;
        RECT 364.950 884.250 366.750 885.150 ;
        RECT 367.950 883.950 370.050 886.050 ;
        RECT 371.250 884.250 373.050 885.150 ;
        RECT 304.950 877.950 307.050 880.050 ;
        RECT 310.950 879.300 313.050 881.400 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 364.950 880.950 367.050 883.050 ;
        RECT 368.250 881.850 369.750 882.750 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 289.950 874.500 292.050 876.600 ;
        RECT 271.950 855.300 274.050 857.400 ;
        RECT 272.250 851.700 273.450 855.300 ;
        RECT 298.950 853.950 301.050 856.050 ;
        RECT 271.950 849.600 274.050 851.700 ;
        RECT 256.950 845.250 259.050 846.150 ;
        RECT 262.950 845.250 265.050 846.150 ;
        RECT 256.950 841.950 259.050 844.050 ;
        RECT 262.950 843.450 265.050 844.050 ;
        RECT 260.400 842.400 265.050 843.450 ;
        RECT 260.400 841.050 261.450 842.400 ;
        RECT 262.950 841.950 265.050 842.400 ;
        RECT 259.950 838.950 262.050 841.050 ;
        RECT 253.950 823.950 256.050 826.050 ;
        RECT 254.400 817.050 255.450 823.950 ;
        RECT 247.950 814.950 250.050 817.050 ;
        RECT 251.250 815.250 252.750 816.150 ;
        RECT 253.950 814.950 256.050 817.050 ;
        RECT 244.950 813.450 247.050 814.050 ;
        RECT 223.950 808.950 226.050 809.400 ;
        RECT 229.950 809.400 234.450 810.450 ;
        RECT 242.400 812.400 247.050 813.450 ;
        RECT 248.250 812.850 249.750 813.750 ;
        RECT 229.950 808.950 232.050 809.400 ;
        RECT 199.950 805.950 202.050 808.050 ;
        RECT 242.400 807.450 243.450 812.400 ;
        RECT 244.950 811.950 247.050 812.400 ;
        RECT 250.950 811.950 253.050 814.050 ;
        RECT 254.250 812.850 256.050 813.750 ;
        RECT 244.950 809.850 247.050 810.750 ;
        RECT 242.400 806.400 246.450 807.450 ;
        RECT 184.950 775.950 187.050 778.050 ;
        RECT 235.950 777.450 238.050 778.050 ;
        RECT 220.950 776.250 223.050 777.150 ;
        RECT 233.400 776.400 238.050 777.450 ;
        RECT 184.950 772.950 187.050 775.050 ;
        RECT 193.950 773.250 196.050 774.150 ;
        RECT 199.950 773.250 202.050 774.150 ;
        RECT 211.950 773.250 213.750 774.150 ;
        RECT 214.950 772.950 217.050 775.050 ;
        RECT 218.250 773.250 219.750 774.150 ;
        RECT 220.950 772.950 223.050 775.050 ;
        RECT 178.950 770.400 183.450 771.450 ;
        RECT 178.950 769.950 181.050 770.400 ;
        RECT 166.950 766.950 169.050 769.050 ;
        RECT 172.950 766.950 175.050 769.050 ;
        RECT 175.950 766.950 178.050 769.050 ;
        RECT 149.400 764.400 153.450 765.450 ;
        RECT 149.400 745.050 150.450 764.400 ;
        RECT 152.400 763.050 153.450 764.400 ;
        RECT 173.400 763.050 174.450 766.950 ;
        RECT 151.950 760.950 154.050 763.050 ;
        RECT 172.950 760.950 175.050 763.050 ;
        RECT 160.950 745.950 163.050 748.050 ;
        RECT 139.950 744.450 142.050 745.050 ;
        RECT 137.400 743.400 142.050 744.450 ;
        RECT 137.400 736.050 138.450 743.400 ;
        RECT 139.950 742.950 142.050 743.400 ;
        RECT 148.950 742.950 151.050 745.050 ;
        RECT 139.950 740.850 142.050 741.750 ;
        RECT 145.950 740.250 148.050 741.150 ;
        RECT 148.950 740.850 151.050 741.750 ;
        RECT 145.950 736.950 148.050 739.050 ;
        RECT 161.400 738.450 162.450 745.950 ;
        RECT 166.950 742.950 169.050 745.050 ;
        RECT 169.950 742.950 172.050 745.050 ;
        RECT 167.400 742.050 168.450 742.950 ;
        RECT 163.950 740.250 165.750 741.150 ;
        RECT 166.950 739.950 169.050 742.050 ;
        RECT 170.400 739.050 171.450 742.950 ;
        RECT 172.950 739.950 175.050 742.050 ;
        RECT 163.950 738.450 166.050 739.050 ;
        RECT 161.400 737.400 166.050 738.450 ;
        RECT 167.250 737.850 168.750 738.750 ;
        RECT 163.950 736.950 166.050 737.400 ;
        RECT 169.950 736.950 172.050 739.050 ;
        RECT 173.250 737.850 175.050 738.750 ;
        RECT 136.950 733.950 139.050 736.050 ;
        RECT 169.950 734.850 172.050 735.750 ;
        RECT 127.950 715.950 130.050 718.050 ;
        RECT 154.950 715.950 157.050 718.050 ;
        RECT 133.950 707.250 136.050 708.150 ;
        RECT 130.950 704.250 132.750 705.150 ;
        RECT 133.950 703.950 136.050 706.050 ;
        RECT 137.250 704.250 138.750 705.150 ;
        RECT 139.950 703.950 142.050 706.050 ;
        RECT 130.950 700.950 133.050 703.050 ;
        RECT 134.400 697.050 135.450 703.950 ;
        RECT 136.950 700.950 139.050 703.050 ;
        RECT 140.250 701.850 142.050 702.750 ;
        RECT 137.400 700.050 138.450 700.950 ;
        RECT 136.950 697.950 139.050 700.050 ;
        RECT 155.400 699.450 156.450 715.950 ;
        RECT 176.400 709.050 177.450 766.950 ;
        RECT 185.400 766.050 186.450 772.950 ;
        RECT 193.950 771.450 196.050 772.050 ;
        RECT 191.400 770.400 196.050 771.450 ;
        RECT 184.950 763.950 187.050 766.050 ;
        RECT 185.400 745.050 186.450 763.950 ;
        RECT 184.950 742.950 187.050 745.050 ;
        RECT 184.950 740.850 187.050 741.750 ;
        RECT 187.950 740.250 190.050 741.150 ;
        RECT 191.400 739.050 192.450 770.400 ;
        RECT 193.950 769.950 196.050 770.400 ;
        RECT 197.250 770.250 198.750 771.150 ;
        RECT 199.950 769.950 202.050 772.050 ;
        RECT 211.950 769.950 214.050 772.050 ;
        RECT 215.250 770.850 216.750 771.750 ;
        RECT 217.950 769.950 220.050 772.050 ;
        RECT 196.950 766.950 199.050 769.050 ;
        RECT 200.400 745.050 201.450 769.950 ;
        RECT 212.400 769.050 213.450 769.950 ;
        RECT 211.950 766.950 214.050 769.050 ;
        RECT 221.400 751.050 222.450 772.950 ;
        RECT 233.400 772.050 234.450 776.400 ;
        RECT 235.950 775.950 238.050 776.400 ;
        RECT 239.250 776.250 240.750 777.150 ;
        RECT 241.950 775.950 244.050 778.050 ;
        RECT 245.400 775.050 246.450 806.400 ;
        RECT 251.400 778.050 252.450 811.950 ;
        RECT 250.950 775.950 253.050 778.050 ;
        RECT 235.950 773.850 237.750 774.750 ;
        RECT 238.950 772.950 241.050 775.050 ;
        RECT 242.250 773.850 244.050 774.750 ;
        RECT 244.950 772.950 247.050 775.050 ;
        RECT 256.950 772.950 259.050 775.050 ;
        RECT 232.950 769.950 235.050 772.050 ;
        RECT 253.950 770.250 256.050 771.150 ;
        RECT 256.950 770.850 259.050 771.750 ;
        RECT 253.950 768.450 256.050 769.050 ;
        RECT 251.400 767.400 256.050 768.450 ;
        RECT 220.950 748.950 223.050 751.050 ;
        RECT 244.950 745.950 247.050 748.050 ;
        RECT 193.950 742.950 196.050 745.050 ;
        RECT 199.950 742.950 202.050 745.050 ;
        RECT 211.950 742.950 214.050 745.050 ;
        RECT 217.950 744.450 220.050 745.050 ;
        RECT 215.250 743.250 216.750 744.150 ;
        RECT 217.950 743.400 222.450 744.450 ;
        RECT 217.950 742.950 220.050 743.400 ;
        RECT 193.950 740.850 196.050 741.750 ;
        RECT 208.950 739.950 211.050 742.050 ;
        RECT 212.250 740.850 213.750 741.750 ;
        RECT 214.950 739.950 217.050 742.050 ;
        RECT 218.250 740.850 220.050 741.750 ;
        RECT 215.400 739.050 216.450 739.950 ;
        RECT 187.950 736.950 190.050 739.050 ;
        RECT 190.950 736.950 193.050 739.050 ;
        RECT 208.950 737.850 211.050 738.750 ;
        RECT 211.950 736.950 214.050 739.050 ;
        RECT 214.950 736.950 217.050 739.050 ;
        RECT 160.950 706.950 163.050 709.050 ;
        RECT 175.950 706.950 178.050 709.050 ;
        RECT 161.400 703.050 162.450 706.950 ;
        RECT 175.950 703.950 178.050 706.050 ;
        RECT 157.950 701.250 159.750 702.150 ;
        RECT 160.950 700.950 163.050 703.050 ;
        RECT 163.950 700.950 166.050 703.050 ;
        RECT 172.950 701.250 175.050 702.150 ;
        RECT 175.950 701.850 178.050 702.750 ;
        RECT 181.950 701.250 184.050 702.150 ;
        RECT 157.950 699.450 160.050 700.050 ;
        RECT 155.400 698.400 160.050 699.450 ;
        RECT 161.250 698.850 163.050 699.750 ;
        RECT 157.950 697.950 160.050 698.400 ;
        RECT 122.400 695.400 126.450 696.450 ;
        RECT 95.400 671.400 99.450 672.450 ;
        RECT 79.950 661.950 82.050 664.050 ;
        RECT 76.950 640.950 79.050 643.050 ;
        RECT 73.950 631.950 76.050 634.050 ;
        RECT 79.950 632.250 82.050 633.150 ;
        RECT 70.950 629.250 72.750 630.150 ;
        RECT 73.950 628.950 76.050 631.050 ;
        RECT 77.250 629.250 78.750 630.150 ;
        RECT 79.950 628.950 82.050 631.050 ;
        RECT 70.950 625.950 73.050 628.050 ;
        RECT 74.250 626.850 75.750 627.750 ;
        RECT 76.950 625.950 79.050 628.050 ;
        RECT 64.950 619.950 67.050 622.050 ;
        RECT 73.950 619.950 76.050 622.050 ;
        RECT 46.950 616.950 49.050 619.050 ;
        RECT 61.950 616.950 64.050 619.050 ;
        RECT 40.950 599.400 45.450 600.450 ;
        RECT 40.950 598.950 43.050 599.400 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 40.950 596.850 43.050 597.750 ;
        RECT 44.400 592.050 45.450 599.400 ;
        RECT 46.950 599.250 49.050 600.150 ;
        RECT 61.950 598.950 64.050 601.050 ;
        RECT 65.250 599.250 66.750 600.150 ;
        RECT 67.950 598.950 70.050 601.050 ;
        RECT 70.950 598.950 73.050 601.050 ;
        RECT 71.400 598.050 72.450 598.950 ;
        RECT 46.950 595.950 49.050 598.050 ;
        RECT 61.950 596.850 63.750 597.750 ;
        RECT 64.950 595.950 67.050 598.050 ;
        RECT 68.250 596.850 69.750 597.750 ;
        RECT 70.950 595.950 73.050 598.050 ;
        RECT 70.950 593.850 73.050 594.750 ;
        RECT 34.950 589.950 37.050 592.050 ;
        RECT 43.950 589.950 46.050 592.050 ;
        RECT 64.950 589.950 67.050 592.050 ;
        RECT 74.400 591.450 75.450 619.950 ;
        RECT 71.400 590.400 75.450 591.450 ;
        RECT 35.400 562.050 36.450 589.950 ;
        RECT 40.950 563.250 43.050 564.150 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 38.250 560.250 39.750 561.150 ;
        RECT 40.950 559.950 43.050 562.050 ;
        RECT 44.250 560.250 46.050 561.150 ;
        RECT 46.950 559.950 49.050 562.050 ;
        RECT 52.950 559.950 55.050 562.050 ;
        RECT 56.250 560.250 57.750 561.150 ;
        RECT 58.950 559.950 61.050 562.050 ;
        RECT 61.950 559.950 64.050 562.050 ;
        RECT 41.400 559.050 42.450 559.950 ;
        RECT 34.950 557.850 36.750 558.750 ;
        RECT 37.950 556.950 40.050 559.050 ;
        RECT 40.950 556.950 43.050 559.050 ;
        RECT 43.950 556.950 46.050 559.050 ;
        RECT 34.950 538.950 37.050 541.050 ;
        RECT 31.950 535.950 34.050 538.050 ;
        RECT 28.950 533.400 31.050 535.500 ;
        RECT 25.950 529.950 28.050 532.050 ;
        RECT 29.250 521.400 30.450 533.400 ;
        RECT 31.950 530.250 34.050 531.150 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 32.400 526.050 33.450 526.950 ;
        RECT 31.950 523.950 34.050 526.050 ;
        RECT 28.950 519.300 31.050 521.400 ;
        RECT 29.250 515.700 30.450 519.300 ;
        RECT 28.950 513.600 31.050 515.700 ;
        RECT 25.950 494.400 28.050 496.500 ;
        RECT 26.400 477.600 27.600 494.400 ;
        RECT 35.400 490.050 36.450 538.950 ;
        RECT 37.950 535.950 40.050 538.050 ;
        RECT 38.400 526.050 39.450 535.950 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 38.400 496.050 39.450 523.950 ;
        RECT 37.950 493.950 40.050 496.050 ;
        RECT 34.950 487.950 37.050 490.050 ;
        RECT 31.950 485.250 34.050 486.150 ;
        RECT 25.950 475.500 28.050 477.600 ;
        RECT 35.400 475.050 36.450 487.950 ;
        RECT 37.950 485.250 40.050 486.150 ;
        RECT 37.950 481.950 40.050 484.050 ;
        RECT 34.950 472.950 37.050 475.050 ;
        RECT 31.950 469.950 34.050 472.050 ;
        RECT 32.400 463.050 33.450 469.950 ;
        RECT 31.950 460.950 34.050 463.050 ;
        RECT 13.950 457.950 16.050 460.050 ;
        RECT 22.950 457.950 25.050 460.050 ;
        RECT 14.400 457.050 15.450 457.950 ;
        RECT 32.400 457.050 33.450 460.950 ;
        RECT 7.950 454.950 10.050 457.050 ;
        RECT 11.250 455.250 12.750 456.150 ;
        RECT 13.950 454.950 16.050 457.050 ;
        RECT 31.950 454.950 34.050 457.050 ;
        RECT 7.950 452.850 9.750 453.750 ;
        RECT 10.950 451.950 13.050 454.050 ;
        RECT 14.250 452.850 15.750 453.750 ;
        RECT 16.950 451.950 19.050 454.050 ;
        RECT 22.950 451.950 25.050 454.050 ;
        RECT 31.950 452.850 34.050 453.750 ;
        RECT 16.950 449.850 19.050 450.750 ;
        RECT 10.950 416.250 13.050 417.150 ;
        RECT 7.950 412.950 10.050 415.050 ;
        RECT 10.950 412.950 13.050 415.050 ;
        RECT 14.250 413.250 15.750 414.150 ;
        RECT 16.950 412.950 19.050 415.050 ;
        RECT 20.250 413.250 22.050 414.150 ;
        RECT 8.400 378.450 9.450 412.950 ;
        RECT 11.400 408.450 12.450 412.950 ;
        RECT 13.950 409.950 16.050 412.050 ;
        RECT 17.250 410.850 18.750 411.750 ;
        RECT 19.950 411.450 22.050 412.050 ;
        RECT 23.400 411.450 24.450 451.950 ;
        RECT 35.400 450.450 36.450 472.950 ;
        RECT 38.400 469.050 39.450 481.950 ;
        RECT 44.400 475.050 45.450 556.950 ;
        RECT 47.400 541.050 48.450 559.950 ;
        RECT 52.950 557.850 54.750 558.750 ;
        RECT 55.950 556.950 58.050 559.050 ;
        RECT 59.250 557.850 61.050 558.750 ;
        RECT 62.400 553.050 63.450 559.950 ;
        RECT 61.950 550.950 64.050 553.050 ;
        RECT 46.950 538.950 49.050 541.050 ;
        RECT 46.950 529.950 49.050 532.050 ;
        RECT 47.400 529.050 48.450 529.950 ;
        RECT 46.950 526.950 49.050 529.050 ;
        RECT 50.250 527.250 51.750 528.150 ;
        RECT 52.950 526.950 55.050 529.050 ;
        RECT 46.950 524.850 48.750 525.750 ;
        RECT 49.950 523.950 52.050 526.050 ;
        RECT 53.250 524.850 54.750 525.750 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 50.400 522.450 51.450 523.950 ;
        RECT 50.400 521.400 54.450 522.450 ;
        RECT 55.950 521.850 58.050 522.750 ;
        RECT 53.400 517.050 54.450 521.400 ;
        RECT 52.950 514.950 55.050 517.050 ;
        RECT 46.950 495.300 49.050 497.400 ;
        RECT 49.950 496.950 52.050 499.050 ;
        RECT 47.250 491.700 48.450 495.300 ;
        RECT 46.950 489.600 49.050 491.700 ;
        RECT 47.250 477.600 48.450 489.600 ;
        RECT 50.400 484.050 51.450 496.950 ;
        RECT 49.950 481.950 52.050 484.050 ;
        RECT 49.950 479.850 52.050 480.750 ;
        RECT 46.950 475.500 49.050 477.600 ;
        RECT 43.950 472.950 46.050 475.050 ;
        RECT 43.950 469.950 46.050 472.050 ;
        RECT 37.950 466.950 40.050 469.050 ;
        RECT 40.950 454.950 43.050 457.050 ;
        RECT 37.950 452.250 40.050 453.150 ;
        RECT 40.950 452.850 43.050 453.750 ;
        RECT 37.950 450.450 40.050 451.050 ;
        RECT 35.400 449.400 40.050 450.450 ;
        RECT 37.950 448.950 40.050 449.400 ;
        RECT 28.950 422.400 31.050 424.500 ;
        RECT 19.950 410.400 24.450 411.450 ;
        RECT 19.950 409.950 22.050 410.400 ;
        RECT 11.400 407.400 15.450 408.450 ;
        RECT 14.400 382.050 15.450 407.400 ;
        RECT 22.950 406.950 25.050 409.050 ;
        RECT 10.950 380.250 12.750 381.150 ;
        RECT 13.950 379.950 16.050 382.050 ;
        RECT 17.250 380.250 19.050 381.150 ;
        RECT 10.950 378.450 13.050 379.050 ;
        RECT 8.400 377.400 13.050 378.450 ;
        RECT 14.250 377.850 15.750 378.750 ;
        RECT 10.950 376.950 13.050 377.400 ;
        RECT 11.400 298.050 12.450 376.950 ;
        RECT 13.950 370.950 16.050 373.050 ;
        RECT 14.400 343.050 15.450 370.950 ;
        RECT 13.950 340.950 16.050 343.050 ;
        RECT 19.950 340.950 22.050 343.050 ;
        RECT 13.950 338.850 16.050 339.750 ;
        RECT 16.950 338.250 19.050 339.150 ;
        RECT 16.950 336.450 19.050 337.050 ;
        RECT 20.400 336.450 21.450 340.950 ;
        RECT 16.950 335.400 21.450 336.450 ;
        RECT 16.950 334.950 19.050 335.400 ;
        RECT 13.950 308.250 15.750 309.150 ;
        RECT 16.950 307.950 19.050 310.050 ;
        RECT 20.250 308.250 22.050 309.150 ;
        RECT 13.950 304.950 16.050 307.050 ;
        RECT 17.250 305.850 18.750 306.750 ;
        RECT 19.950 304.950 22.050 307.050 ;
        RECT 14.400 304.050 15.450 304.950 ;
        RECT 20.400 304.050 21.450 304.950 ;
        RECT 13.950 301.950 16.050 304.050 ;
        RECT 19.950 301.950 22.050 304.050 ;
        RECT 10.950 295.950 13.050 298.050 ;
        RECT 7.950 278.400 10.050 280.500 ;
        RECT 8.400 261.600 9.600 278.400 ;
        RECT 13.950 269.250 16.050 270.150 ;
        RECT 19.950 269.250 22.050 270.150 ;
        RECT 13.950 265.950 16.050 268.050 ;
        RECT 19.950 267.450 22.050 268.050 ;
        RECT 23.400 267.450 24.450 406.950 ;
        RECT 29.400 405.600 30.600 422.400 ;
        RECT 34.950 413.250 37.050 414.150 ;
        RECT 34.950 409.950 37.050 412.050 ;
        RECT 28.950 403.500 31.050 405.600 ;
        RECT 34.950 385.950 37.050 388.050 ;
        RECT 31.950 383.250 34.050 384.150 ;
        RECT 34.950 383.850 37.050 384.750 ;
        RECT 31.950 379.950 34.050 382.050 ;
        RECT 32.400 379.050 33.450 379.950 ;
        RECT 31.950 376.950 34.050 379.050 ;
        RECT 38.400 370.050 39.450 448.950 ;
        RECT 40.950 413.250 43.050 414.150 ;
        RECT 40.950 409.950 43.050 412.050 ;
        RECT 41.400 409.050 42.450 409.950 ;
        RECT 40.950 406.950 43.050 409.050 ;
        RECT 28.950 367.950 31.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 29.400 339.450 30.450 367.950 ;
        RECT 40.950 343.950 43.050 346.050 ;
        RECT 41.400 343.050 42.450 343.950 ;
        RECT 31.950 341.250 33.750 342.150 ;
        RECT 34.950 340.950 37.050 343.050 ;
        RECT 40.950 340.950 43.050 343.050 ;
        RECT 31.950 339.450 34.050 340.050 ;
        RECT 29.400 338.400 34.050 339.450 ;
        RECT 35.250 338.850 37.050 339.750 ;
        RECT 31.950 337.950 34.050 338.400 ;
        RECT 37.950 338.250 40.050 339.150 ;
        RECT 40.950 338.850 43.050 339.750 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 34.950 316.950 37.050 319.050 ;
        RECT 35.400 310.050 36.450 316.950 ;
        RECT 38.400 316.050 39.450 334.950 ;
        RECT 44.400 319.050 45.450 469.950 ;
        RECT 46.950 466.950 49.050 469.050 ;
        RECT 47.400 460.050 48.450 466.950 ;
        RECT 46.950 457.950 49.050 460.050 ;
        RECT 47.400 409.050 48.450 457.950 ;
        RECT 49.950 423.300 52.050 425.400 ;
        RECT 50.250 419.700 51.450 423.300 ;
        RECT 49.950 417.600 52.050 419.700 ;
        RECT 46.950 406.950 49.050 409.050 ;
        RECT 50.250 405.600 51.450 417.600 ;
        RECT 53.400 415.050 54.450 514.950 ;
        RECT 62.400 487.050 63.450 550.950 ;
        RECT 61.950 484.950 64.050 487.050 ;
        RECT 58.950 472.950 61.050 475.050 ;
        RECT 59.400 460.050 60.450 472.950 ;
        RECT 62.400 463.050 63.450 484.950 ;
        RECT 65.400 481.050 66.450 589.950 ;
        RECT 67.950 568.950 70.050 571.050 ;
        RECT 68.400 517.050 69.450 568.950 ;
        RECT 71.400 556.050 72.450 590.400 ;
        RECT 77.400 562.050 78.450 625.950 ;
        RECT 80.400 619.050 81.450 628.950 ;
        RECT 79.950 616.950 82.050 619.050 ;
        RECT 80.400 601.050 81.450 616.950 ;
        RECT 83.400 604.050 84.450 670.950 ;
        RECT 88.950 668.250 90.750 669.150 ;
        RECT 91.950 667.950 94.050 670.050 ;
        RECT 95.250 668.250 97.050 669.150 ;
        RECT 88.950 664.950 91.050 667.050 ;
        RECT 92.250 665.850 93.750 666.750 ;
        RECT 94.950 664.950 97.050 667.050 ;
        RECT 89.400 649.050 90.450 664.950 ;
        RECT 95.400 660.450 96.450 664.950 ;
        RECT 92.400 659.400 96.450 660.450 ;
        RECT 88.950 646.950 91.050 649.050 ;
        RECT 92.400 631.050 93.450 659.400 ;
        RECT 98.400 640.050 99.450 671.400 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 107.400 670.050 108.450 670.950 ;
        RECT 103.950 668.250 105.750 669.150 ;
        RECT 106.950 667.950 109.050 670.050 ;
        RECT 110.250 668.250 112.050 669.150 ;
        RECT 103.950 664.950 106.050 667.050 ;
        RECT 107.250 665.850 108.750 666.750 ;
        RECT 109.950 664.950 112.050 667.050 ;
        RECT 103.950 661.950 106.050 664.050 ;
        RECT 97.950 637.950 100.050 640.050 ;
        RECT 97.950 635.250 100.050 636.150 ;
        RECT 104.400 634.050 105.450 661.950 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 94.950 632.250 96.750 633.150 ;
        RECT 97.950 631.950 100.050 634.050 ;
        RECT 101.250 632.250 102.750 633.150 ;
        RECT 103.950 631.950 106.050 634.050 ;
        RECT 91.950 628.950 94.050 631.050 ;
        RECT 94.950 628.950 97.050 631.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 79.950 598.950 82.050 601.050 ;
        RECT 85.950 598.950 88.050 601.050 ;
        RECT 91.950 598.950 94.050 601.050 ;
        RECT 85.950 596.850 88.050 597.750 ;
        RECT 88.950 595.950 91.050 598.050 ;
        RECT 91.950 596.850 94.050 597.750 ;
        RECT 73.950 560.250 76.050 561.150 ;
        RECT 76.950 559.950 79.050 562.050 ;
        RECT 73.950 556.950 76.050 559.050 ;
        RECT 77.250 557.250 78.750 558.150 ;
        RECT 79.950 556.950 82.050 559.050 ;
        RECT 83.250 557.250 85.050 558.150 ;
        RECT 70.950 553.950 73.050 556.050 ;
        RECT 74.400 550.050 75.450 556.950 ;
        RECT 89.400 556.050 90.450 595.950 ;
        RECT 98.400 595.050 99.450 631.950 ;
        RECT 107.400 631.050 108.450 646.950 ;
        RECT 109.950 640.950 112.050 643.050 ;
        RECT 100.950 628.950 103.050 631.050 ;
        RECT 104.250 629.850 106.050 630.750 ;
        RECT 106.950 628.950 109.050 631.050 ;
        RECT 103.950 599.250 106.050 600.150 ;
        RECT 106.950 598.950 109.050 601.050 ;
        RECT 91.950 592.950 94.050 595.050 ;
        RECT 97.950 592.950 100.050 595.050 ;
        RECT 76.950 553.950 79.050 556.050 ;
        RECT 80.250 554.850 81.750 555.750 ;
        RECT 82.950 555.450 85.050 556.050 ;
        RECT 82.950 554.400 87.450 555.450 ;
        RECT 82.950 553.950 85.050 554.400 ;
        RECT 73.950 547.950 76.050 550.050 ;
        RECT 82.950 547.950 85.050 550.050 ;
        RECT 70.950 524.250 72.750 525.150 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 77.250 524.250 79.050 525.150 ;
        RECT 70.950 520.950 73.050 523.050 ;
        RECT 74.250 521.850 75.750 522.750 ;
        RECT 71.400 517.050 72.450 520.950 ;
        RECT 67.950 514.950 70.050 517.050 ;
        RECT 70.950 514.950 73.050 517.050 ;
        RECT 67.950 488.250 70.050 489.150 ;
        RECT 73.950 487.950 76.050 490.050 ;
        RECT 74.400 487.050 75.450 487.950 ;
        RECT 67.950 484.950 70.050 487.050 ;
        RECT 71.250 485.250 72.750 486.150 ;
        RECT 73.950 484.950 76.050 487.050 ;
        RECT 77.250 485.250 79.050 486.150 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 74.250 482.850 75.750 483.750 ;
        RECT 76.950 481.950 79.050 484.050 ;
        RECT 64.950 478.950 67.050 481.050 ;
        RECT 83.400 466.050 84.450 547.950 ;
        RECT 86.400 538.050 87.450 554.400 ;
        RECT 88.950 553.950 91.050 556.050 ;
        RECT 92.400 550.050 93.450 592.950 ;
        RECT 94.950 557.250 97.050 558.150 ;
        RECT 100.950 557.250 103.050 558.150 ;
        RECT 94.950 553.950 97.050 556.050 ;
        RECT 98.250 554.250 99.750 555.150 ;
        RECT 100.950 553.950 103.050 556.050 ;
        RECT 91.950 547.950 94.050 550.050 ;
        RECT 85.950 535.950 88.050 538.050 ;
        RECT 91.950 529.950 94.050 532.050 ;
        RECT 95.400 529.050 96.450 553.950 ;
        RECT 97.950 550.950 100.050 553.050 ;
        RECT 97.950 547.950 100.050 550.050 ;
        RECT 88.950 528.450 91.050 529.050 ;
        RECT 86.400 527.400 91.050 528.450 ;
        RECT 92.250 527.850 93.750 528.750 ;
        RECT 86.400 522.450 87.450 527.400 ;
        RECT 88.950 526.950 91.050 527.400 ;
        RECT 94.950 526.950 97.050 529.050 ;
        RECT 88.950 524.850 91.050 525.750 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 94.950 524.850 97.050 525.750 ;
        RECT 86.400 521.400 90.450 522.450 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 82.950 463.950 85.050 466.050 ;
        RECT 61.950 460.950 64.050 463.050 ;
        RECT 67.950 461.400 70.050 463.500 ;
        RECT 58.950 459.450 61.050 460.050 ;
        RECT 58.950 458.400 63.450 459.450 ;
        RECT 58.950 457.950 61.050 458.400 ;
        RECT 55.950 455.250 58.050 456.150 ;
        RECT 58.950 455.850 61.050 456.750 ;
        RECT 55.950 451.950 58.050 454.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 62.400 412.050 63.450 458.400 ;
        RECT 64.950 458.250 67.050 459.150 ;
        RECT 64.950 454.950 67.050 457.050 ;
        RECT 65.400 451.050 66.450 454.950 ;
        RECT 64.950 448.950 67.050 451.050 ;
        RECT 68.550 449.400 69.750 461.400 ;
        RECT 76.950 457.950 79.050 460.050 ;
        RECT 77.400 457.050 78.450 457.950 ;
        RECT 76.950 454.950 79.050 457.050 ;
        RECT 82.950 454.950 85.050 457.050 ;
        RECT 70.950 451.950 73.050 454.050 ;
        RECT 76.950 452.850 79.050 453.750 ;
        RECT 82.950 452.850 85.050 453.750 ;
        RECT 52.950 409.950 55.050 412.050 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 52.950 407.850 55.050 408.750 ;
        RECT 49.950 403.500 52.050 405.600 ;
        RECT 55.950 403.950 58.050 406.050 ;
        RECT 46.950 380.250 48.750 381.150 ;
        RECT 49.950 379.950 52.050 382.050 ;
        RECT 53.250 380.250 55.050 381.150 ;
        RECT 46.950 376.950 49.050 379.050 ;
        RECT 50.250 377.850 51.750 378.750 ;
        RECT 52.950 378.450 55.050 379.050 ;
        RECT 56.400 378.450 57.450 403.950 ;
        RECT 65.400 388.050 66.450 448.950 ;
        RECT 67.950 447.300 70.050 449.400 ;
        RECT 68.550 443.700 69.750 447.300 ;
        RECT 67.950 441.600 70.050 443.700 ;
        RECT 71.400 415.050 72.450 451.950 ;
        RECT 86.400 451.050 87.450 490.950 ;
        RECT 89.400 490.050 90.450 521.400 ;
        RECT 88.950 487.950 91.050 490.050 ;
        RECT 92.400 487.050 93.450 523.950 ;
        RECT 88.950 484.950 91.050 487.050 ;
        RECT 91.950 484.950 94.050 487.050 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 88.950 482.850 91.050 483.750 ;
        RECT 91.950 482.250 94.050 483.150 ;
        RECT 95.400 481.050 96.450 484.950 ;
        RECT 91.950 478.950 94.050 481.050 ;
        RECT 94.950 478.950 97.050 481.050 ;
        RECT 92.400 478.050 93.450 478.950 ;
        RECT 91.950 475.950 94.050 478.050 ;
        RECT 91.950 472.950 94.050 475.050 ;
        RECT 88.950 461.400 91.050 463.500 ;
        RECT 85.950 448.950 88.050 451.050 ;
        RECT 79.950 442.950 82.050 445.050 ;
        RECT 89.400 444.600 90.600 461.400 ;
        RECT 92.400 445.050 93.450 472.950 ;
        RECT 94.950 448.950 97.050 451.050 ;
        RECT 76.950 416.250 79.050 417.150 ;
        RECT 67.950 413.250 69.750 414.150 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 74.250 413.250 75.750 414.150 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 71.250 410.850 72.750 411.750 ;
        RECT 73.950 409.950 76.050 412.050 ;
        RECT 68.400 406.050 69.450 409.950 ;
        RECT 67.950 403.950 70.050 406.050 ;
        RECT 70.950 391.950 73.050 394.050 ;
        RECT 64.950 385.950 67.050 388.050 ;
        RECT 71.400 385.050 72.450 391.950 ;
        RECT 74.400 391.050 75.450 409.950 ;
        RECT 73.950 388.950 76.050 391.050 ;
        RECT 76.950 385.950 79.050 388.050 ;
        RECT 77.400 385.050 78.450 385.950 ;
        RECT 70.950 382.950 73.050 385.050 ;
        RECT 74.250 383.250 75.750 384.150 ;
        RECT 76.950 382.950 79.050 385.050 ;
        RECT 67.950 379.950 70.050 382.050 ;
        RECT 71.250 380.850 72.750 381.750 ;
        RECT 73.950 379.950 76.050 382.050 ;
        RECT 77.250 380.850 79.050 381.750 ;
        RECT 52.950 377.400 57.450 378.450 ;
        RECT 67.950 377.850 70.050 378.750 ;
        RECT 52.950 376.950 55.050 377.400 ;
        RECT 46.950 373.950 49.050 376.050 ;
        RECT 47.400 319.050 48.450 373.950 ;
        RECT 56.400 349.050 57.450 377.400 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 80.400 378.450 81.450 442.950 ;
        RECT 88.950 442.500 91.050 444.600 ;
        RECT 91.950 442.950 94.050 445.050 ;
        RECT 95.400 418.050 96.450 448.950 ;
        RECT 88.950 417.450 91.050 418.050 ;
        RECT 86.400 416.400 91.050 417.450 ;
        RECT 82.950 406.950 85.050 409.050 ;
        RECT 83.400 379.050 84.450 406.950 ;
        RECT 86.400 406.050 87.450 416.400 ;
        RECT 88.950 415.950 91.050 416.400 ;
        RECT 92.250 416.250 93.750 417.150 ;
        RECT 94.950 415.950 97.050 418.050 ;
        RECT 88.950 413.850 90.750 414.750 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 95.250 413.850 97.050 414.750 ;
        RECT 88.950 409.950 91.050 412.050 ;
        RECT 85.950 403.950 88.050 406.050 ;
        RECT 85.950 400.950 88.050 403.050 ;
        RECT 77.400 377.400 81.450 378.450 ;
        RECT 55.950 346.950 58.050 349.050 ;
        RECT 67.950 346.950 70.050 349.050 ;
        RECT 49.950 340.950 52.050 343.050 ;
        RECT 52.950 341.250 54.750 342.150 ;
        RECT 55.950 340.950 58.050 343.050 ;
        RECT 61.950 342.450 64.050 343.050 ;
        RECT 61.950 341.400 66.450 342.450 ;
        RECT 61.950 340.950 64.050 341.400 ;
        RECT 40.950 316.950 43.050 319.050 ;
        RECT 43.950 316.950 46.050 319.050 ;
        RECT 46.950 316.950 49.050 319.050 ;
        RECT 37.950 313.950 40.050 316.050 ;
        RECT 31.950 308.250 33.750 309.150 ;
        RECT 34.950 307.950 37.050 310.050 ;
        RECT 38.250 308.250 40.050 309.150 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 35.250 305.850 36.750 306.750 ;
        RECT 37.950 304.950 40.050 307.050 ;
        RECT 31.950 301.950 34.050 304.050 ;
        RECT 38.400 303.450 39.450 304.950 ;
        RECT 35.400 302.400 39.450 303.450 ;
        RECT 28.950 279.300 31.050 281.400 ;
        RECT 29.250 275.700 30.450 279.300 ;
        RECT 28.950 273.600 31.050 275.700 ;
        RECT 19.950 266.400 24.450 267.450 ;
        RECT 19.950 265.950 22.050 266.400 ;
        RECT 7.950 259.500 10.050 261.600 ;
        RECT 14.400 241.050 15.450 265.950 ;
        RECT 13.950 238.950 16.050 241.050 ;
        RECT 17.250 239.250 18.750 240.150 ;
        RECT 19.950 238.950 22.050 241.050 ;
        RECT 4.950 235.950 7.050 238.050 ;
        RECT 10.950 235.950 13.050 238.050 ;
        RECT 14.250 236.850 15.750 237.750 ;
        RECT 16.950 235.950 19.050 238.050 ;
        RECT 20.250 236.850 22.050 237.750 ;
        RECT 5.400 199.050 6.450 235.950 ;
        RECT 10.950 233.850 13.050 234.750 ;
        RECT 17.400 234.450 18.450 235.950 ;
        RECT 14.400 233.400 18.450 234.450 ;
        RECT 14.400 204.450 15.450 233.400 ;
        RECT 11.400 203.400 15.450 204.450 ;
        RECT 11.400 202.050 12.450 203.400 ;
        RECT 10.950 201.450 13.050 202.050 ;
        RECT 8.400 200.400 13.050 201.450 ;
        RECT 4.950 196.950 7.050 199.050 ;
        RECT 8.400 166.050 9.450 200.400 ;
        RECT 10.950 199.950 13.050 200.400 ;
        RECT 14.250 200.250 15.750 201.150 ;
        RECT 23.400 199.050 24.450 266.400 ;
        RECT 29.250 261.600 30.450 273.600 ;
        RECT 32.400 268.050 33.450 301.950 ;
        RECT 31.950 265.950 34.050 268.050 ;
        RECT 31.950 263.850 34.050 264.750 ;
        RECT 28.950 259.500 31.050 261.600 ;
        RECT 28.950 238.950 31.050 241.050 ;
        RECT 29.400 234.450 30.450 238.950 ;
        RECT 35.400 238.050 36.450 302.400 ;
        RECT 41.400 238.050 42.450 316.950 ;
        RECT 50.400 316.050 51.450 340.950 ;
        RECT 52.950 337.950 55.050 340.050 ;
        RECT 56.250 338.850 58.050 339.750 ;
        RECT 58.950 338.250 61.050 339.150 ;
        RECT 61.950 338.850 64.050 339.750 ;
        RECT 53.400 331.050 54.450 337.950 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 59.400 334.050 60.450 334.950 ;
        RECT 58.950 331.950 61.050 334.050 ;
        RECT 52.950 328.950 55.050 331.050 ;
        RECT 59.400 316.050 60.450 331.950 ;
        RECT 65.400 328.050 66.450 341.400 ;
        RECT 64.950 325.950 67.050 328.050 ;
        RECT 64.950 316.950 67.050 319.050 ;
        RECT 65.400 316.050 66.450 316.950 ;
        RECT 68.400 316.050 69.450 346.950 ;
        RECT 46.950 313.950 49.050 316.050 ;
        RECT 49.950 313.950 52.050 316.050 ;
        RECT 58.950 313.950 61.050 316.050 ;
        RECT 64.950 313.950 67.050 316.050 ;
        RECT 67.950 313.950 70.050 316.050 ;
        RECT 47.400 313.050 48.450 313.950 ;
        RECT 46.950 310.950 49.050 313.050 ;
        RECT 50.250 311.850 51.750 312.750 ;
        RECT 52.950 312.450 55.050 313.050 ;
        RECT 55.950 312.450 58.050 313.050 ;
        RECT 52.950 311.400 58.050 312.450 ;
        RECT 52.950 310.950 55.050 311.400 ;
        RECT 55.950 310.950 58.050 311.400 ;
        RECT 46.950 308.850 49.050 309.750 ;
        RECT 52.950 308.850 55.050 309.750 ;
        RECT 56.400 304.050 57.450 310.950 ;
        RECT 55.950 301.950 58.050 304.050 ;
        RECT 43.950 295.950 46.050 298.050 ;
        RECT 31.950 236.250 33.750 237.150 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 38.250 236.250 40.050 237.150 ;
        RECT 40.950 235.950 43.050 238.050 ;
        RECT 31.950 234.450 34.050 235.050 ;
        RECT 29.400 233.400 34.050 234.450 ;
        RECT 35.250 233.850 36.750 234.750 ;
        RECT 31.950 232.950 34.050 233.400 ;
        RECT 37.950 232.950 40.050 235.050 ;
        RECT 25.950 226.950 28.050 229.050 ;
        RECT 10.950 197.850 12.750 198.750 ;
        RECT 13.950 196.950 16.050 199.050 ;
        RECT 17.250 197.850 19.050 198.750 ;
        RECT 22.950 196.950 25.050 199.050 ;
        RECT 26.400 172.050 27.450 226.950 ;
        RECT 28.950 196.950 31.050 199.050 ;
        RECT 28.950 194.850 31.050 195.750 ;
        RECT 10.950 169.950 13.050 172.050 ;
        RECT 25.950 169.950 28.050 172.050 ;
        RECT 11.400 169.050 12.450 169.950 ;
        RECT 10.950 166.950 13.050 169.050 ;
        RECT 14.250 167.250 15.750 168.150 ;
        RECT 16.950 166.950 19.050 169.050 ;
        RECT 22.950 166.950 25.050 169.050 ;
        RECT 7.950 163.950 10.050 166.050 ;
        RECT 10.950 164.850 12.750 165.750 ;
        RECT 13.950 163.950 16.050 166.050 ;
        RECT 17.250 164.850 18.750 165.750 ;
        RECT 19.950 163.950 22.050 166.050 ;
        RECT 14.400 163.050 15.450 163.950 ;
        RECT 13.950 160.950 16.050 163.050 ;
        RECT 19.950 161.850 22.050 162.750 ;
        RECT 7.950 135.300 10.050 137.400 ;
        RECT 8.550 131.700 9.750 135.300 ;
        RECT 7.950 129.600 10.050 131.700 ;
        RECT 4.950 121.950 7.050 124.050 ;
        RECT 4.950 119.850 7.050 120.750 ;
        RECT 8.550 117.600 9.750 129.600 ;
        RECT 23.400 129.450 24.450 166.950 ;
        RECT 20.400 128.400 24.450 129.450 ;
        RECT 16.950 125.250 19.050 126.150 ;
        RECT 10.950 121.950 13.050 124.050 ;
        RECT 13.950 121.950 16.050 124.050 ;
        RECT 16.950 121.950 19.050 124.050 ;
        RECT 20.400 123.450 21.450 128.400 ;
        RECT 22.950 125.250 25.050 126.150 ;
        RECT 26.400 124.050 27.450 169.950 ;
        RECT 34.950 164.250 36.750 165.150 ;
        RECT 37.950 163.950 40.050 166.050 ;
        RECT 41.250 164.250 43.050 165.150 ;
        RECT 34.950 160.950 37.050 163.050 ;
        RECT 38.250 161.850 39.750 162.750 ;
        RECT 44.400 154.050 45.450 295.950 ;
        RECT 49.950 270.450 52.050 271.050 ;
        RECT 49.950 269.400 54.450 270.450 ;
        RECT 49.950 268.950 52.050 269.400 ;
        RECT 46.950 266.250 49.050 267.150 ;
        RECT 49.950 266.850 52.050 267.750 ;
        RECT 46.950 262.950 49.050 265.050 ;
        RECT 53.400 247.050 54.450 269.400 ;
        RECT 52.950 244.950 55.050 247.050 ;
        RECT 53.400 241.050 54.450 244.950 ;
        RECT 56.400 244.050 57.450 301.950 ;
        RECT 59.400 250.050 60.450 313.950 ;
        RECT 64.950 311.850 67.050 312.750 ;
        RECT 67.950 311.250 70.050 312.150 ;
        RECT 67.950 307.950 70.050 310.050 ;
        RECT 68.400 280.050 69.450 307.950 ;
        RECT 67.950 277.950 70.050 280.050 ;
        RECT 71.400 277.050 72.450 376.950 ;
        RECT 73.950 343.950 76.050 346.050 ;
        RECT 74.400 343.050 75.450 343.950 ;
        RECT 73.950 340.950 76.050 343.050 ;
        RECT 73.950 338.850 76.050 339.750 ;
        RECT 73.950 313.950 76.050 316.050 ;
        RECT 70.950 274.950 73.050 277.050 ;
        RECT 74.400 274.050 75.450 313.950 ;
        RECT 77.400 310.050 78.450 377.400 ;
        RECT 82.950 376.950 85.050 379.050 ;
        RECT 79.950 341.250 82.050 342.150 ;
        RECT 79.950 337.950 82.050 340.050 ;
        RECT 83.250 338.250 85.050 339.150 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 86.400 331.050 87.450 400.950 ;
        RECT 89.400 385.050 90.450 409.950 ;
        RECT 98.400 403.050 99.450 547.950 ;
        RECT 107.400 547.050 108.450 598.950 ;
        RECT 106.950 544.950 109.050 547.050 ;
        RECT 100.950 532.950 103.050 535.050 ;
        RECT 101.400 484.050 102.450 532.950 ;
        RECT 110.400 529.050 111.450 640.950 ;
        RECT 113.400 621.450 114.450 694.950 ;
        RECT 116.400 661.050 117.450 694.950 ;
        RECT 122.400 666.450 123.450 695.400 ;
        RECT 133.950 694.950 136.050 697.050 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 128.400 670.050 129.450 670.950 ;
        RECT 124.950 668.250 126.750 669.150 ;
        RECT 127.950 667.950 130.050 670.050 ;
        RECT 133.950 667.950 136.050 670.050 ;
        RECT 137.400 667.050 138.450 697.950 ;
        RECT 148.950 691.950 151.050 694.050 ;
        RECT 149.400 673.050 150.450 691.950 ;
        RECT 154.950 676.950 157.050 679.050 ;
        RECT 155.400 676.050 156.450 676.950 ;
        RECT 154.950 673.950 157.050 676.050 ;
        RECT 148.950 670.950 151.050 673.050 ;
        RECT 152.250 671.250 154.050 672.150 ;
        RECT 154.950 671.850 157.050 672.750 ;
        RECT 157.950 671.250 160.050 672.150 ;
        RECT 148.950 668.850 150.750 669.750 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 157.950 667.950 160.050 670.050 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 124.950 666.450 127.050 667.050 ;
        RECT 122.400 665.400 127.050 666.450 ;
        RECT 128.250 665.850 129.750 666.750 ;
        RECT 124.950 664.950 127.050 665.400 ;
        RECT 130.950 664.950 133.050 667.050 ;
        RECT 134.250 665.850 136.050 666.750 ;
        RECT 136.950 664.950 139.050 667.050 ;
        RECT 130.950 662.850 133.050 663.750 ;
        RECT 115.950 658.950 118.050 661.050 ;
        RECT 130.950 637.950 133.050 640.050 ;
        RECT 124.950 635.250 127.050 636.150 ;
        RECT 118.950 633.450 121.050 634.050 ;
        RECT 116.400 632.400 121.050 633.450 ;
        RECT 116.400 625.050 117.450 632.400 ;
        RECT 118.950 631.950 121.050 632.400 ;
        RECT 122.250 632.250 123.750 633.150 ;
        RECT 124.950 631.950 127.050 634.050 ;
        RECT 128.250 632.250 130.050 633.150 ;
        RECT 118.950 629.850 120.750 630.750 ;
        RECT 121.950 628.950 124.050 631.050 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 122.400 625.050 123.450 628.950 ;
        RECT 115.950 622.950 118.050 625.050 ;
        RECT 121.950 622.950 124.050 625.050 ;
        RECT 113.400 620.400 117.450 621.450 ;
        RECT 116.400 559.050 117.450 620.400 ;
        RECT 124.950 599.250 127.050 600.150 ;
        RECT 124.950 595.950 127.050 598.050 ;
        RECT 112.950 557.250 115.050 558.150 ;
        RECT 115.950 556.950 118.050 559.050 ;
        RECT 118.950 557.250 121.050 558.150 ;
        RECT 112.950 553.950 115.050 556.050 ;
        RECT 116.250 554.250 117.750 555.150 ;
        RECT 118.950 553.950 121.050 556.050 ;
        RECT 113.400 553.050 114.450 553.950 ;
        RECT 112.950 550.950 115.050 553.050 ;
        RECT 115.950 550.950 118.050 553.050 ;
        RECT 121.950 550.950 124.050 553.050 ;
        RECT 116.400 531.450 117.450 550.950 ;
        RECT 116.400 530.400 120.450 531.450 ;
        RECT 109.950 526.950 112.050 529.050 ;
        RECT 113.250 527.250 114.750 528.150 ;
        RECT 115.950 526.950 118.050 529.050 ;
        RECT 119.400 526.050 120.450 530.400 ;
        RECT 122.400 528.450 123.450 550.950 ;
        RECT 125.400 550.050 126.450 595.950 ;
        RECT 131.400 568.050 132.450 637.950 ;
        RECT 152.400 634.050 153.450 667.950 ;
        RECT 158.400 649.050 159.450 667.950 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 151.950 631.950 154.050 634.050 ;
        RECT 139.950 628.950 142.050 631.050 ;
        RECT 154.950 628.950 157.050 631.050 ;
        RECT 136.950 626.250 139.050 627.150 ;
        RECT 139.950 626.850 142.050 627.750 ;
        RECT 154.950 626.850 157.050 627.750 ;
        RECT 157.950 626.250 160.050 627.150 ;
        RECT 136.950 622.950 139.050 625.050 ;
        RECT 154.950 624.450 157.050 625.050 ;
        RECT 157.950 624.450 160.050 625.050 ;
        RECT 154.950 623.400 160.050 624.450 ;
        RECT 154.950 622.950 157.050 623.400 ;
        RECT 157.950 622.950 160.050 623.400 ;
        RECT 137.400 598.050 138.450 622.950 ;
        RECT 145.950 619.950 148.050 622.050 ;
        RECT 146.400 601.050 147.450 619.950 ;
        RECT 145.950 598.950 148.050 601.050 ;
        RECT 149.250 599.250 150.750 600.150 ;
        RECT 151.950 598.950 154.050 601.050 ;
        RECT 155.400 598.050 156.450 622.950 ;
        RECT 157.950 610.950 160.050 613.050 ;
        RECT 158.400 601.050 159.450 610.950 ;
        RECT 157.950 598.950 160.050 601.050 ;
        RECT 133.950 595.950 136.050 598.050 ;
        RECT 136.950 595.950 139.050 598.050 ;
        RECT 142.950 595.950 145.050 598.050 ;
        RECT 146.250 596.850 147.750 597.750 ;
        RECT 148.950 595.950 151.050 598.050 ;
        RECT 152.250 596.850 154.050 597.750 ;
        RECT 154.950 595.950 157.050 598.050 ;
        RECT 130.950 565.950 133.050 568.050 ;
        RECT 130.950 559.950 133.050 562.050 ;
        RECT 124.950 547.950 127.050 550.050 ;
        RECT 127.950 535.950 130.050 538.050 ;
        RECT 128.400 532.050 129.450 535.950 ;
        RECT 131.400 532.050 132.450 559.950 ;
        RECT 134.400 537.450 135.450 595.950 ;
        RECT 142.950 593.850 145.050 594.750 ;
        RECT 136.950 562.950 139.050 565.050 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 137.400 562.050 138.450 562.950 ;
        RECT 136.950 559.950 139.050 562.050 ;
        RECT 140.250 560.250 141.750 561.150 ;
        RECT 142.950 559.950 145.050 562.050 ;
        RECT 136.950 557.850 138.750 558.750 ;
        RECT 139.950 556.950 142.050 559.050 ;
        RECT 143.250 557.850 145.050 558.750 ;
        RECT 139.950 550.950 142.050 553.050 ;
        RECT 134.400 536.400 138.450 537.450 ;
        RECT 127.950 529.950 130.050 532.050 ;
        RECT 130.950 529.950 133.050 532.050 ;
        RECT 124.950 528.450 127.050 529.050 ;
        RECT 122.400 527.400 127.050 528.450 ;
        RECT 128.250 527.850 129.750 528.750 ;
        RECT 130.950 528.450 133.050 529.050 ;
        RECT 106.950 525.450 109.050 526.050 ;
        RECT 104.400 524.400 109.050 525.450 ;
        RECT 110.250 524.850 111.750 525.750 ;
        RECT 104.400 493.050 105.450 524.400 ;
        RECT 106.950 523.950 109.050 524.400 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 116.250 524.850 118.050 525.750 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 122.400 523.050 123.450 527.400 ;
        RECT 124.950 526.950 127.050 527.400 ;
        RECT 130.950 527.400 135.450 528.450 ;
        RECT 130.950 526.950 133.050 527.400 ;
        RECT 124.950 524.850 127.050 525.750 ;
        RECT 130.950 524.850 133.050 525.750 ;
        RECT 106.950 521.850 109.050 522.750 ;
        RECT 115.950 520.950 118.050 523.050 ;
        RECT 121.950 520.950 124.050 523.050 ;
        RECT 130.950 520.950 133.050 523.050 ;
        RECT 112.950 517.950 115.050 520.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 103.950 485.250 106.050 486.150 ;
        RECT 109.950 485.250 112.050 486.150 ;
        RECT 100.950 481.950 103.050 484.050 ;
        RECT 103.950 481.950 106.050 484.050 ;
        RECT 107.250 482.250 108.750 483.150 ;
        RECT 109.950 481.950 112.050 484.050 ;
        RECT 104.400 481.050 105.450 481.950 ;
        RECT 100.950 478.950 103.050 481.050 ;
        RECT 103.950 478.950 106.050 481.050 ;
        RECT 106.950 478.950 109.050 481.050 ;
        RECT 101.400 412.050 102.450 478.950 ;
        RECT 113.400 475.050 114.450 517.950 ;
        RECT 116.400 478.050 117.450 520.950 ;
        RECT 121.950 487.950 124.050 490.050 ;
        RECT 127.950 488.250 130.050 489.150 ;
        RECT 122.400 487.050 123.450 487.950 ;
        RECT 118.950 485.250 120.750 486.150 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 125.250 485.250 126.750 486.150 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 118.950 481.950 121.050 484.050 ;
        RECT 122.250 482.850 123.750 483.750 ;
        RECT 124.950 481.950 127.050 484.050 ;
        RECT 119.400 481.050 120.450 481.950 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 115.950 475.950 118.050 478.050 ;
        RECT 121.950 475.950 124.050 478.050 ;
        RECT 112.950 472.950 115.050 475.050 ;
        RECT 103.950 463.950 106.050 466.050 ;
        RECT 104.400 456.450 105.450 463.950 ;
        RECT 106.950 456.450 109.050 457.050 ;
        RECT 104.400 455.400 109.050 456.450 ;
        RECT 100.950 409.950 103.050 412.050 ;
        RECT 104.400 409.050 105.450 455.400 ;
        RECT 106.950 454.950 109.050 455.400 ;
        RECT 110.250 455.250 111.750 456.150 ;
        RECT 112.950 454.950 115.050 457.050 ;
        RECT 106.950 452.850 108.750 453.750 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 113.250 452.850 114.750 453.750 ;
        RECT 115.950 451.950 118.050 454.050 ;
        RECT 110.400 451.050 111.450 451.950 ;
        RECT 109.950 448.950 112.050 451.050 ;
        RECT 115.950 449.850 118.050 450.750 ;
        RECT 109.950 416.250 112.050 417.150 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 113.250 413.250 114.750 414.150 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 119.250 413.250 121.050 414.150 ;
        RECT 103.950 406.950 106.050 409.050 ;
        RECT 110.400 408.450 111.450 412.950 ;
        RECT 112.950 409.950 115.050 412.050 ;
        RECT 116.250 410.850 117.750 411.750 ;
        RECT 118.950 409.950 121.050 412.050 ;
        RECT 110.400 407.400 114.450 408.450 ;
        RECT 97.950 400.950 100.050 403.050 ;
        RECT 109.950 391.950 112.050 394.050 ;
        RECT 106.950 388.950 109.050 391.050 ;
        RECT 103.950 385.950 106.050 388.050 ;
        RECT 88.950 382.950 91.050 385.050 ;
        RECT 92.250 383.250 94.050 384.150 ;
        RECT 97.950 382.950 100.050 385.050 ;
        RECT 101.250 383.250 103.050 384.150 ;
        RECT 88.950 380.850 90.750 381.750 ;
        RECT 91.950 379.950 94.050 382.050 ;
        RECT 97.950 380.850 99.750 381.750 ;
        RECT 100.950 379.950 103.050 382.050 ;
        RECT 92.400 349.050 93.450 379.950 ;
        RECT 101.400 379.050 102.450 379.950 ;
        RECT 104.400 379.050 105.450 385.950 ;
        RECT 100.950 376.950 103.050 379.050 ;
        RECT 103.950 376.950 106.050 379.050 ;
        RECT 103.950 349.950 106.050 352.050 ;
        RECT 91.950 346.950 94.050 349.050 ;
        RECT 100.950 344.250 103.050 345.150 ;
        RECT 91.950 341.250 93.750 342.150 ;
        RECT 94.950 340.950 97.050 343.050 ;
        RECT 100.950 342.450 103.050 343.050 ;
        RECT 104.400 342.450 105.450 349.950 ;
        RECT 98.250 341.250 99.750 342.150 ;
        RECT 100.950 341.400 105.450 342.450 ;
        RECT 100.950 340.950 103.050 341.400 ;
        RECT 88.950 339.450 91.050 340.050 ;
        RECT 91.950 339.450 94.050 340.050 ;
        RECT 88.950 338.400 94.050 339.450 ;
        RECT 95.250 338.850 96.750 339.750 ;
        RECT 88.950 337.950 91.050 338.400 ;
        RECT 91.950 337.950 94.050 338.400 ;
        RECT 97.950 337.950 100.050 340.050 ;
        RECT 85.950 328.950 88.050 331.050 ;
        RECT 89.400 316.050 90.450 337.950 ;
        RECT 107.400 319.050 108.450 388.950 ;
        RECT 110.400 382.050 111.450 391.950 ;
        RECT 109.950 379.950 112.050 382.050 ;
        RECT 113.400 381.450 114.450 407.400 ;
        RECT 119.400 394.050 120.450 409.950 ;
        RECT 118.950 391.950 121.050 394.050 ;
        RECT 122.400 390.450 123.450 475.950 ;
        RECT 128.400 472.050 129.450 484.950 ;
        RECT 131.400 484.050 132.450 520.950 ;
        RECT 134.400 490.050 135.450 527.400 ;
        RECT 133.950 487.950 136.050 490.050 ;
        RECT 130.950 481.950 133.050 484.050 ;
        RECT 127.950 469.950 130.050 472.050 ;
        RECT 127.950 452.250 129.750 453.150 ;
        RECT 130.950 451.950 133.050 454.050 ;
        RECT 134.250 452.250 136.050 453.150 ;
        RECT 131.250 449.850 132.750 450.750 ;
        RECT 133.950 448.950 136.050 451.050 ;
        RECT 137.400 445.050 138.450 536.400 ;
        RECT 140.400 451.050 141.450 550.950 ;
        RECT 142.950 535.950 145.050 538.050 ;
        RECT 143.400 526.050 144.450 535.950 ;
        RECT 152.400 529.050 153.450 562.950 ;
        RECT 154.950 557.250 157.050 558.150 ;
        RECT 154.950 553.950 157.050 556.050 ;
        RECT 158.400 535.050 159.450 598.950 ;
        RECT 161.400 562.050 162.450 667.950 ;
        RECT 160.950 559.950 163.050 562.050 ;
        RECT 164.400 559.050 165.450 700.950 ;
        RECT 188.400 700.050 189.450 736.950 ;
        RECT 190.950 703.950 193.050 706.050 ;
        RECT 172.950 697.950 175.050 700.050 ;
        RECT 181.950 697.950 184.050 700.050 ;
        RECT 187.950 697.950 190.050 700.050 ;
        RECT 191.400 699.450 192.450 703.950 ;
        RECT 193.950 701.250 195.750 702.150 ;
        RECT 196.950 700.950 199.050 703.050 ;
        RECT 202.950 700.950 205.050 703.050 ;
        RECT 208.950 700.950 211.050 703.050 ;
        RECT 193.950 699.450 196.050 700.050 ;
        RECT 191.400 698.400 196.050 699.450 ;
        RECT 197.250 698.850 199.050 699.750 ;
        RECT 193.950 697.950 196.050 698.400 ;
        RECT 199.950 698.250 202.050 699.150 ;
        RECT 202.950 698.850 205.050 699.750 ;
        RECT 182.400 697.050 183.450 697.950 ;
        RECT 181.950 694.950 184.050 697.050 ;
        RECT 190.950 694.950 193.050 697.050 ;
        RECT 199.950 694.950 202.050 697.050 ;
        RECT 202.950 694.950 205.050 697.050 ;
        RECT 191.400 670.050 192.450 694.950 ;
        RECT 166.950 668.250 168.750 669.150 ;
        RECT 169.950 667.950 172.050 670.050 ;
        RECT 173.250 668.250 175.050 669.150 ;
        RECT 187.950 668.250 189.750 669.150 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 194.250 668.250 196.050 669.150 ;
        RECT 200.400 667.050 201.450 694.950 ;
        RECT 203.400 682.050 204.450 694.950 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 203.400 670.050 204.450 679.950 ;
        RECT 209.400 670.050 210.450 700.950 ;
        RECT 212.400 699.450 213.450 736.950 ;
        RECT 221.400 733.050 222.450 743.400 ;
        RECT 245.400 742.050 246.450 745.950 ;
        RECT 251.400 742.050 252.450 767.400 ;
        RECT 253.950 766.950 256.050 767.400 ;
        RECT 260.400 742.050 261.450 838.950 ;
        RECT 272.250 837.600 273.450 849.600 ;
        RECT 295.950 848.250 298.050 849.150 ;
        RECT 280.950 844.950 283.050 847.050 ;
        RECT 286.950 845.250 288.750 846.150 ;
        RECT 289.950 844.950 292.050 847.050 ;
        RECT 295.950 846.450 298.050 847.050 ;
        RECT 299.400 846.450 300.450 853.950 ;
        RECT 293.250 845.250 294.750 846.150 ;
        RECT 295.950 845.400 300.450 846.450 ;
        RECT 295.950 844.950 298.050 845.400 ;
        RECT 274.950 841.950 277.050 844.050 ;
        RECT 274.950 839.850 277.050 840.750 ;
        RECT 271.950 835.500 274.050 837.600 ;
        RECT 262.950 832.950 265.050 835.050 ;
        RECT 263.400 817.050 264.450 832.950 ;
        RECT 262.950 814.950 265.050 817.050 ;
        RECT 266.250 815.250 267.750 816.150 ;
        RECT 268.950 814.950 271.050 817.050 ;
        RECT 281.400 814.050 282.450 844.950 ;
        RECT 283.950 841.950 286.050 844.050 ;
        RECT 286.950 841.950 289.050 844.050 ;
        RECT 290.250 842.850 291.750 843.750 ;
        RECT 292.950 841.950 295.050 844.050 ;
        RECT 284.400 820.050 285.450 841.950 ;
        RECT 287.400 835.050 288.450 841.950 ;
        RECT 286.950 832.950 289.050 835.050 ;
        RECT 293.400 829.050 294.450 841.950 ;
        RECT 305.400 841.050 306.450 877.950 ;
        RECT 311.250 875.700 312.450 879.300 ;
        RECT 310.950 873.600 313.050 875.700 ;
        RECT 307.950 854.400 310.050 856.500 ;
        RECT 328.950 855.300 331.050 857.400 ;
        RECT 304.950 838.950 307.050 841.050 ;
        RECT 308.400 837.600 309.600 854.400 ;
        RECT 329.250 851.700 330.450 855.300 ;
        RECT 328.950 849.600 331.050 851.700 ;
        RECT 313.950 845.250 316.050 846.150 ;
        RECT 319.950 845.250 322.050 846.150 ;
        RECT 313.950 843.450 316.050 844.050 ;
        RECT 311.400 842.400 316.050 843.450 ;
        RECT 307.950 835.500 310.050 837.600 ;
        RECT 292.950 826.950 295.050 829.050 ;
        RECT 283.950 817.950 286.050 820.050 ;
        RECT 311.400 817.050 312.450 842.400 ;
        RECT 313.950 841.950 316.050 842.400 ;
        RECT 319.950 841.950 322.050 844.050 ;
        RECT 320.400 841.050 321.450 841.950 ;
        RECT 319.950 838.950 322.050 841.050 ;
        RECT 283.950 815.850 286.050 816.750 ;
        RECT 286.950 815.250 289.050 816.150 ;
        RECT 298.950 814.950 301.050 817.050 ;
        RECT 304.950 816.450 307.050 817.050 ;
        RECT 302.400 815.400 307.050 816.450 ;
        RECT 262.950 812.850 264.750 813.750 ;
        RECT 265.950 811.950 268.050 814.050 ;
        RECT 269.250 812.850 270.750 813.750 ;
        RECT 271.950 811.950 274.050 814.050 ;
        RECT 280.950 811.950 283.050 814.050 ;
        RECT 286.950 811.950 289.050 814.050 ;
        RECT 266.400 811.050 267.450 811.950 ;
        RECT 265.950 808.950 268.050 811.050 ;
        RECT 271.950 809.850 274.050 810.750 ;
        RECT 299.400 802.050 300.450 814.950 ;
        RECT 298.950 799.950 301.050 802.050 ;
        RECT 295.950 777.450 298.050 778.050 ;
        RECT 271.950 776.250 274.050 777.150 ;
        RECT 293.400 776.400 298.050 777.450 ;
        RECT 271.950 772.950 274.050 775.050 ;
        RECT 275.250 773.250 276.750 774.150 ;
        RECT 277.950 772.950 280.050 775.050 ;
        RECT 281.250 773.250 283.050 774.150 ;
        RECT 286.950 772.950 289.050 775.050 ;
        RECT 289.950 773.250 292.050 774.150 ;
        RECT 265.950 745.950 268.050 748.050 ;
        RECT 265.950 743.850 268.050 744.750 ;
        RECT 268.950 743.250 271.050 744.150 ;
        RECT 229.950 740.250 231.750 741.150 ;
        RECT 232.950 739.950 235.050 742.050 ;
        RECT 238.950 741.450 241.050 742.050 ;
        RECT 238.950 740.400 243.450 741.450 ;
        RECT 238.950 739.950 241.050 740.400 ;
        RECT 242.400 739.050 243.450 740.400 ;
        RECT 244.950 739.950 247.050 742.050 ;
        RECT 247.950 740.250 249.750 741.150 ;
        RECT 250.950 739.950 253.050 742.050 ;
        RECT 254.250 740.250 256.050 741.150 ;
        RECT 259.950 739.950 262.050 742.050 ;
        RECT 265.950 739.950 268.050 742.050 ;
        RECT 268.950 739.950 271.050 742.050 ;
        RECT 229.950 736.950 232.050 739.050 ;
        RECT 233.250 737.850 234.750 738.750 ;
        RECT 235.950 736.950 238.050 739.050 ;
        RECT 239.250 737.850 241.050 738.750 ;
        RECT 241.950 736.950 244.050 739.050 ;
        RECT 235.950 734.850 238.050 735.750 ;
        RECT 220.950 730.950 223.050 733.050 ;
        RECT 217.950 703.950 220.050 706.050 ;
        RECT 218.400 703.050 219.450 703.950 ;
        RECT 214.950 701.250 216.750 702.150 ;
        RECT 217.950 700.950 220.050 703.050 ;
        RECT 223.950 700.950 226.050 703.050 ;
        RECT 238.950 700.950 241.050 703.050 ;
        RECT 214.950 699.450 217.050 700.050 ;
        RECT 212.400 698.400 217.050 699.450 ;
        RECT 218.250 698.850 220.050 699.750 ;
        RECT 214.950 697.950 217.050 698.400 ;
        RECT 220.950 698.250 223.050 699.150 ;
        RECT 223.950 698.850 226.050 699.750 ;
        RECT 238.950 698.850 241.050 699.750 ;
        RECT 241.950 698.250 244.050 699.150 ;
        RECT 220.950 696.450 223.050 697.050 ;
        RECT 218.400 695.400 223.050 696.450 ;
        RECT 202.950 667.950 205.050 670.050 ;
        RECT 208.950 667.950 211.050 670.050 ;
        RECT 212.250 668.250 214.050 669.150 ;
        RECT 218.400 667.050 219.450 695.400 ;
        RECT 220.950 694.950 223.050 695.400 ;
        RECT 241.950 694.950 244.050 697.050 ;
        RECT 221.400 694.050 222.450 694.950 ;
        RECT 220.950 691.950 223.050 694.050 ;
        RECT 245.400 688.050 246.450 739.950 ;
        RECT 247.950 736.950 250.050 739.050 ;
        RECT 251.250 737.850 252.750 738.750 ;
        RECT 253.950 736.950 256.050 739.050 ;
        RECT 259.950 736.950 262.050 739.050 ;
        RECT 244.950 685.950 247.050 688.050 ;
        RECT 248.400 685.050 249.450 736.950 ;
        RECT 254.400 736.050 255.450 736.950 ;
        RECT 253.950 733.950 256.050 736.050 ;
        RECT 250.950 710.400 253.050 712.500 ;
        RECT 251.400 693.600 252.600 710.400 ;
        RECT 254.400 694.050 255.450 733.950 ;
        RECT 256.950 701.250 259.050 702.150 ;
        RECT 256.950 697.950 259.050 700.050 ;
        RECT 257.400 694.050 258.450 697.950 ;
        RECT 260.400 697.050 261.450 736.950 ;
        RECT 262.950 701.250 265.050 702.150 ;
        RECT 266.400 700.050 267.450 739.950 ;
        RECT 272.400 718.050 273.450 772.950 ;
        RECT 274.950 769.950 277.050 772.050 ;
        RECT 278.250 770.850 279.750 771.750 ;
        RECT 280.950 769.950 283.050 772.050 ;
        RECT 287.400 771.450 288.450 772.950 ;
        RECT 293.400 772.050 294.450 776.400 ;
        RECT 295.950 775.950 298.050 776.400 ;
        RECT 295.950 773.850 298.050 774.750 ;
        RECT 298.950 773.250 301.050 774.150 ;
        RECT 289.950 771.450 292.050 772.050 ;
        RECT 287.400 770.400 292.050 771.450 ;
        RECT 275.400 769.050 276.450 769.950 ;
        RECT 274.950 766.950 277.050 769.050 ;
        RECT 287.400 745.050 288.450 770.400 ;
        RECT 289.950 769.950 292.050 770.400 ;
        RECT 292.950 769.950 295.050 772.050 ;
        RECT 298.950 769.950 301.050 772.050 ;
        RECT 302.400 769.050 303.450 815.400 ;
        RECT 304.950 814.950 307.050 815.400 ;
        RECT 308.250 815.250 309.750 816.150 ;
        RECT 310.950 814.950 313.050 817.050 ;
        RECT 314.250 815.250 315.750 816.150 ;
        RECT 316.950 814.950 319.050 817.050 ;
        RECT 304.950 812.850 306.750 813.750 ;
        RECT 307.950 811.950 310.050 814.050 ;
        RECT 311.250 812.850 312.750 813.750 ;
        RECT 313.950 811.950 316.050 814.050 ;
        RECT 317.250 812.850 319.050 813.750 ;
        RECT 308.400 772.050 309.450 811.950 ;
        RECT 320.400 811.050 321.450 838.950 ;
        RECT 329.250 837.600 330.450 849.600 ;
        RECT 331.950 843.450 334.050 844.050 ;
        RECT 331.950 842.400 336.450 843.450 ;
        RECT 331.950 841.950 334.050 842.400 ;
        RECT 331.950 839.850 334.050 840.750 ;
        RECT 328.950 835.500 331.050 837.600 ;
        RECT 335.400 822.450 336.450 842.400 ;
        RECT 337.950 841.950 340.050 844.050 ;
        RECT 332.400 821.400 336.450 822.450 ;
        RECT 332.400 820.050 333.450 821.400 ;
        RECT 331.950 817.950 334.050 820.050 ;
        RECT 325.950 814.950 328.050 817.050 ;
        RECT 328.950 815.250 331.050 816.150 ;
        RECT 331.950 815.850 334.050 816.750 ;
        RECT 326.400 813.450 327.450 814.950 ;
        RECT 328.950 813.450 331.050 814.050 ;
        RECT 326.400 812.400 331.050 813.450 ;
        RECT 328.950 811.950 331.050 812.400 ;
        RECT 329.400 811.050 330.450 811.950 ;
        RECT 313.950 808.950 316.050 811.050 ;
        RECT 319.950 808.950 322.050 811.050 ;
        RECT 328.950 808.950 331.050 811.050 ;
        RECT 314.400 775.050 315.450 808.950 ;
        RECT 338.400 805.050 339.450 841.950 ;
        RECT 341.400 814.050 342.450 880.950 ;
        RECT 358.950 850.950 361.050 853.050 ;
        RECT 352.950 847.950 355.050 850.050 ;
        RECT 353.400 847.050 354.450 847.950 ;
        RECT 359.400 847.050 360.450 850.950 ;
        RECT 365.400 847.050 366.450 880.950 ;
        RECT 377.400 880.050 378.450 887.400 ;
        RECT 379.950 886.950 382.050 887.400 ;
        RECT 385.950 887.400 390.450 888.450 ;
        RECT 385.950 886.950 388.050 887.400 ;
        RECT 379.950 884.850 382.050 885.750 ;
        RECT 385.950 884.850 388.050 885.750 ;
        RECT 389.400 882.450 390.450 887.400 ;
        RECT 397.950 886.950 400.050 889.050 ;
        RECT 401.250 887.250 402.750 888.150 ;
        RECT 403.950 886.950 406.050 889.050 ;
        RECT 397.950 884.850 399.750 885.750 ;
        RECT 400.950 883.950 403.050 886.050 ;
        RECT 404.250 884.850 405.750 885.750 ;
        RECT 406.950 883.950 409.050 886.050 ;
        RECT 386.400 881.400 390.450 882.450 ;
        RECT 406.950 881.850 409.050 882.750 ;
        RECT 370.950 877.950 373.050 880.050 ;
        RECT 376.950 877.950 379.050 880.050 ;
        RECT 371.400 850.050 372.450 877.950 ;
        RECT 386.400 850.050 387.450 881.400 ;
        RECT 419.400 876.600 420.600 893.400 ;
        RECT 424.950 886.950 427.050 889.050 ;
        RECT 430.950 888.450 433.050 889.050 ;
        RECT 433.950 888.450 436.050 889.050 ;
        RECT 430.950 887.400 436.050 888.450 ;
        RECT 430.950 886.950 433.050 887.400 ;
        RECT 433.950 886.950 436.050 887.400 ;
        RECT 424.950 884.850 427.050 885.750 ;
        RECT 430.950 884.850 433.050 885.750 ;
        RECT 418.950 874.500 421.050 876.600 ;
        RECT 388.950 854.400 391.050 856.500 ;
        RECT 409.950 855.300 412.050 857.400 ;
        RECT 370.950 849.450 373.050 850.050 ;
        RECT 368.400 848.400 373.050 849.450 ;
        RECT 349.950 845.250 351.750 846.150 ;
        RECT 352.950 844.950 355.050 847.050 ;
        RECT 356.250 845.250 357.750 846.150 ;
        RECT 358.950 844.950 361.050 847.050 ;
        RECT 362.250 845.250 364.050 846.150 ;
        RECT 364.950 844.950 367.050 847.050 ;
        RECT 349.950 841.950 352.050 844.050 ;
        RECT 353.250 842.850 354.750 843.750 ;
        RECT 355.950 841.950 358.050 844.050 ;
        RECT 359.250 842.850 360.750 843.750 ;
        RECT 361.950 841.950 364.050 844.050 ;
        RECT 368.400 843.450 369.450 848.400 ;
        RECT 370.950 847.950 373.050 848.400 ;
        RECT 374.250 848.250 375.750 849.150 ;
        RECT 376.950 847.950 379.050 850.050 ;
        RECT 385.950 847.950 388.050 850.050 ;
        RECT 370.950 845.850 372.750 846.750 ;
        RECT 373.950 844.950 376.050 847.050 ;
        RECT 377.250 845.850 379.050 846.750 ;
        RECT 382.950 844.950 385.050 847.050 ;
        RECT 365.400 842.400 369.450 843.450 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 344.400 817.050 345.450 835.950 ;
        RECT 355.950 820.950 358.050 823.050 ;
        RECT 356.400 817.050 357.450 820.950 ;
        RECT 362.400 820.050 363.450 841.950 ;
        RECT 361.950 817.950 364.050 820.050 ;
        RECT 343.950 814.950 346.050 817.050 ;
        RECT 347.250 815.250 348.750 816.150 ;
        RECT 349.950 814.950 352.050 817.050 ;
        RECT 353.250 815.250 354.750 816.150 ;
        RECT 355.950 814.950 358.050 817.050 ;
        RECT 361.950 814.950 364.050 817.050 ;
        RECT 340.950 811.950 343.050 814.050 ;
        RECT 343.950 812.850 345.750 813.750 ;
        RECT 346.950 811.950 349.050 814.050 ;
        RECT 350.250 812.850 351.750 813.750 ;
        RECT 352.950 811.950 355.050 814.050 ;
        RECT 356.250 812.850 358.050 813.750 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 313.950 772.950 316.050 775.050 ;
        RECT 307.950 769.950 310.050 772.050 ;
        RECT 313.950 770.850 316.050 771.750 ;
        RECT 334.950 770.850 337.050 771.750 ;
        RECT 301.950 766.950 304.050 769.050 ;
        RECT 322.950 747.450 325.050 748.050 ;
        RECT 320.400 746.400 325.050 747.450 ;
        RECT 280.950 742.950 283.050 745.050 ;
        RECT 284.250 743.250 285.750 744.150 ;
        RECT 286.950 742.950 289.050 745.050 ;
        RECT 316.950 742.950 319.050 745.050 ;
        RECT 280.950 740.850 282.750 741.750 ;
        RECT 283.950 739.950 286.050 742.050 ;
        RECT 287.250 740.850 288.750 741.750 ;
        RECT 289.950 739.950 292.050 742.050 ;
        RECT 307.950 740.250 309.750 741.150 ;
        RECT 310.950 739.950 313.050 742.050 ;
        RECT 314.250 740.250 316.050 741.150 ;
        RECT 284.400 739.050 285.450 739.950 ;
        RECT 283.950 736.950 286.050 739.050 ;
        RECT 289.950 737.850 292.050 738.750 ;
        RECT 307.950 736.950 310.050 739.050 ;
        RECT 311.250 737.850 312.750 738.750 ;
        RECT 313.950 738.450 316.050 739.050 ;
        RECT 317.400 738.450 318.450 742.950 ;
        RECT 320.400 739.050 321.450 746.400 ;
        RECT 322.950 745.950 325.050 746.400 ;
        RECT 341.400 745.050 342.450 811.950 ;
        RECT 347.400 808.050 348.450 811.950 ;
        RECT 353.400 811.050 354.450 811.950 ;
        RECT 352.950 808.950 355.050 811.050 ;
        RECT 346.950 805.950 349.050 808.050 ;
        RECT 362.400 805.050 363.450 814.950 ;
        RECT 365.400 811.050 366.450 842.400 ;
        RECT 367.950 823.950 370.050 826.050 ;
        RECT 368.400 817.050 369.450 823.950 ;
        RECT 379.950 820.950 382.050 823.050 ;
        RECT 380.400 817.050 381.450 820.950 ;
        RECT 383.400 820.050 384.450 844.950 ;
        RECT 382.950 817.950 385.050 820.050 ;
        RECT 367.950 814.950 370.050 817.050 ;
        RECT 371.250 815.250 372.750 816.150 ;
        RECT 373.950 814.950 376.050 817.050 ;
        RECT 377.250 815.250 378.750 816.150 ;
        RECT 379.950 814.950 382.050 817.050 ;
        RECT 383.400 814.050 384.450 817.950 ;
        RECT 367.950 812.850 369.750 813.750 ;
        RECT 370.950 811.950 373.050 814.050 ;
        RECT 374.250 812.850 375.750 813.750 ;
        RECT 376.950 811.950 379.050 814.050 ;
        RECT 380.250 812.850 382.050 813.750 ;
        RECT 382.950 811.950 385.050 814.050 ;
        RECT 364.950 808.950 367.050 811.050 ;
        RECT 371.400 808.050 372.450 811.950 ;
        RECT 373.950 808.950 376.050 811.050 ;
        RECT 370.950 805.950 373.050 808.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 361.950 802.950 364.050 805.050 ;
        RECT 322.950 743.850 324.750 744.750 ;
        RECT 325.950 742.950 328.050 745.050 ;
        RECT 331.950 743.250 334.050 744.150 ;
        RECT 340.950 742.950 343.050 745.050 ;
        RECT 347.400 742.050 348.450 802.950 ;
        RECT 349.950 775.950 352.050 778.050 ;
        RECT 350.400 771.450 351.450 775.950 ;
        RECT 374.400 775.050 375.450 808.950 ;
        RECT 352.950 773.250 355.050 774.150 ;
        RECT 358.950 773.250 361.050 774.150 ;
        RECT 373.950 772.950 376.050 775.050 ;
        RECT 386.400 772.050 387.450 847.950 ;
        RECT 389.400 837.600 390.600 854.400 ;
        RECT 410.250 851.700 411.450 855.300 ;
        RECT 409.950 849.600 412.050 851.700 ;
        RECT 394.950 845.250 397.050 846.150 ;
        RECT 400.950 845.250 403.050 846.150 ;
        RECT 394.950 841.950 397.050 844.050 ;
        RECT 400.950 841.950 403.050 844.050 ;
        RECT 401.400 841.050 402.450 841.950 ;
        RECT 400.950 838.950 403.050 841.050 ;
        RECT 410.250 837.600 411.450 849.600 ;
        RECT 427.950 844.950 430.050 847.050 ;
        RECT 412.950 841.950 415.050 844.050 ;
        RECT 421.950 841.950 424.050 844.050 ;
        RECT 424.950 842.250 427.050 843.150 ;
        RECT 427.950 842.850 430.050 843.750 ;
        RECT 412.950 839.850 415.050 840.750 ;
        RECT 422.400 840.450 423.450 841.950 ;
        RECT 434.400 841.050 435.450 886.950 ;
        RECT 440.250 881.400 441.450 893.400 ;
        RECT 442.950 890.250 445.050 891.150 ;
        RECT 442.950 886.950 445.050 889.050 ;
        RECT 443.400 883.050 444.450 886.950 ;
        RECT 454.950 884.250 456.750 885.150 ;
        RECT 457.950 883.950 460.050 886.050 ;
        RECT 461.250 884.250 463.050 885.150 ;
        RECT 439.950 879.300 442.050 881.400 ;
        RECT 442.950 880.950 445.050 883.050 ;
        RECT 454.950 880.950 457.050 883.050 ;
        RECT 458.250 881.850 459.750 882.750 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 440.250 875.700 441.450 879.300 ;
        RECT 439.950 873.600 442.050 875.700 ;
        RECT 439.950 854.400 442.050 856.500 ;
        RECT 455.400 856.050 456.450 880.950 ;
        RECT 473.400 876.600 474.600 893.400 ;
        RECT 478.950 888.450 481.050 889.050 ;
        RECT 478.950 887.400 483.450 888.450 ;
        RECT 478.950 886.950 481.050 887.400 ;
        RECT 482.400 886.050 483.450 887.400 ;
        RECT 484.950 886.950 487.050 889.050 ;
        RECT 478.950 884.850 481.050 885.750 ;
        RECT 481.950 883.950 484.050 886.050 ;
        RECT 484.950 884.850 487.050 885.750 ;
        RECT 481.950 880.950 484.050 883.050 ;
        RECT 494.250 881.400 495.450 893.400 ;
        RECT 508.950 891.450 511.050 892.050 ;
        RECT 523.950 891.450 526.050 892.050 ;
        RECT 496.950 890.250 499.050 891.150 ;
        RECT 506.400 890.400 511.050 891.450 ;
        RECT 506.400 889.050 507.450 890.400 ;
        RECT 508.950 889.950 511.050 890.400 ;
        RECT 521.400 890.400 526.050 891.450 ;
        RECT 496.950 886.950 499.050 889.050 ;
        RECT 505.950 886.950 508.050 889.050 ;
        RECT 508.950 887.850 511.050 888.750 ;
        RECT 511.950 887.250 514.050 888.150 ;
        RECT 502.950 883.950 505.050 886.050 ;
        RECT 511.950 883.950 514.050 886.050 ;
        RECT 472.950 874.500 475.050 876.600 ;
        RECT 424.950 840.450 427.050 841.050 ;
        RECT 422.400 839.400 427.050 840.450 ;
        RECT 424.950 838.950 427.050 839.400 ;
        RECT 433.950 838.950 436.050 841.050 ;
        RECT 440.400 837.600 441.600 854.400 ;
        RECT 454.950 853.950 457.050 856.050 ;
        RECT 460.950 855.300 463.050 857.400 ;
        RECT 461.250 851.700 462.450 855.300 ;
        RECT 482.400 853.050 483.450 880.950 ;
        RECT 493.950 879.300 496.050 881.400 ;
        RECT 494.250 875.700 495.450 879.300 ;
        RECT 493.950 873.600 496.050 875.700 ;
        RECT 460.950 849.600 463.050 851.700 ;
        RECT 481.950 850.950 484.050 853.050 ;
        RECT 445.950 845.250 448.050 846.150 ;
        RECT 451.950 845.250 454.050 846.150 ;
        RECT 442.950 841.950 445.050 844.050 ;
        RECT 445.950 841.950 448.050 844.050 ;
        RECT 451.950 841.950 454.050 844.050 ;
        RECT 388.950 835.500 391.050 837.600 ;
        RECT 409.950 835.500 412.050 837.600 ;
        RECT 439.950 835.500 442.050 837.600 ;
        RECT 394.950 829.950 397.050 832.050 ;
        RECT 391.950 817.950 394.050 820.050 ;
        RECT 392.400 802.050 393.450 817.950 ;
        RECT 395.400 817.050 396.450 829.950 ;
        RECT 418.950 826.950 421.050 829.050 ;
        RECT 419.400 820.050 420.450 826.950 ;
        RECT 427.950 823.950 430.050 826.050 ;
        RECT 400.950 817.950 403.050 820.050 ;
        RECT 406.950 817.950 409.050 820.050 ;
        RECT 418.950 817.950 421.050 820.050 ;
        RECT 394.950 814.950 397.050 817.050 ;
        RECT 398.250 815.250 400.050 816.150 ;
        RECT 400.950 815.850 403.050 816.750 ;
        RECT 403.950 815.250 406.050 816.150 ;
        RECT 394.950 812.850 396.750 813.750 ;
        RECT 397.950 811.950 400.050 814.050 ;
        RECT 403.950 811.950 406.050 814.050 ;
        RECT 398.400 805.050 399.450 811.950 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 391.950 799.950 394.050 802.050 ;
        RECT 404.400 799.050 405.450 811.950 ;
        RECT 407.400 808.050 408.450 817.950 ;
        RECT 415.950 815.250 418.050 816.150 ;
        RECT 418.950 815.850 421.050 816.750 ;
        RECT 421.950 815.250 423.750 816.150 ;
        RECT 424.950 814.950 427.050 817.050 ;
        RECT 415.950 811.950 418.050 814.050 ;
        RECT 421.950 811.950 424.050 814.050 ;
        RECT 425.250 812.850 427.050 813.750 ;
        RECT 406.950 805.950 409.050 808.050 ;
        RECT 416.400 799.050 417.450 811.950 ;
        RECT 403.950 796.950 406.050 799.050 ;
        RECT 415.950 796.950 418.050 799.050 ;
        RECT 391.950 776.250 394.050 777.150 ;
        RECT 397.950 775.950 400.050 778.050 ;
        RECT 406.950 775.950 409.050 778.050 ;
        RECT 398.400 775.050 399.450 775.950 ;
        RECT 391.950 772.950 394.050 775.050 ;
        RECT 395.250 773.250 396.750 774.150 ;
        RECT 397.950 772.950 400.050 775.050 ;
        RECT 401.250 773.250 403.050 774.150 ;
        RECT 403.950 772.950 406.050 775.050 ;
        RECT 352.950 771.450 355.050 772.050 ;
        RECT 350.400 770.400 355.050 771.450 ;
        RECT 352.950 769.950 355.050 770.400 ;
        RECT 358.950 769.950 361.050 772.050 ;
        RECT 370.950 770.250 373.050 771.150 ;
        RECT 373.950 770.850 376.050 771.750 ;
        RECT 385.950 769.950 388.050 772.050 ;
        RECT 394.950 769.950 397.050 772.050 ;
        RECT 398.250 770.850 399.750 771.750 ;
        RECT 400.950 769.950 403.050 772.050 ;
        RECT 359.400 760.050 360.450 769.950 ;
        RECT 370.950 768.450 373.050 769.050 ;
        RECT 373.950 768.450 376.050 769.050 ;
        RECT 370.950 767.400 376.050 768.450 ;
        RECT 370.950 766.950 373.050 767.400 ;
        RECT 373.950 766.950 376.050 767.400 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 362.400 745.050 363.450 757.950 ;
        RECT 358.950 742.950 361.050 745.050 ;
        RECT 361.950 742.950 364.050 745.050 ;
        RECT 367.950 742.950 370.050 745.050 ;
        RECT 325.950 740.850 328.050 741.750 ;
        RECT 331.950 739.950 334.050 742.050 ;
        RECT 340.950 739.950 343.050 742.050 ;
        RECT 343.950 740.250 345.750 741.150 ;
        RECT 346.950 739.950 349.050 742.050 ;
        RECT 350.250 740.250 352.050 741.150 ;
        RECT 332.400 739.050 333.450 739.950 ;
        RECT 313.950 737.400 318.450 738.450 ;
        RECT 313.950 736.950 316.050 737.400 ;
        RECT 319.950 736.950 322.050 739.050 ;
        RECT 331.950 736.950 334.050 739.050 ;
        RECT 341.400 738.450 342.450 739.950 ;
        RECT 343.950 738.450 346.050 739.050 ;
        RECT 341.400 737.400 346.050 738.450 ;
        RECT 347.250 737.850 348.750 738.750 ;
        RECT 343.950 736.950 346.050 737.400 ;
        RECT 349.950 736.950 352.050 739.050 ;
        RECT 284.400 733.050 285.450 736.950 ;
        RECT 283.950 730.950 286.050 733.050 ;
        RECT 271.950 715.950 274.050 718.050 ;
        RECT 271.950 711.300 274.050 713.400 ;
        RECT 272.250 707.700 273.450 711.300 ;
        RECT 271.950 705.600 274.050 707.700 ;
        RECT 262.950 697.950 265.050 700.050 ;
        RECT 265.950 697.950 268.050 700.050 ;
        RECT 259.950 694.950 262.050 697.050 ;
        RECT 250.950 691.500 253.050 693.600 ;
        RECT 253.950 691.950 256.050 694.050 ;
        RECT 256.950 691.950 259.050 694.050 ;
        RECT 250.950 685.950 253.050 688.050 ;
        RECT 247.950 682.950 250.050 685.050 ;
        RECT 235.950 676.950 238.050 679.050 ;
        RECT 229.950 670.950 232.050 673.050 ;
        RECT 230.400 670.050 231.450 670.950 ;
        RECT 236.400 670.050 237.450 676.950 ;
        RECT 251.400 673.050 252.450 685.950 ;
        RECT 260.400 673.050 261.450 694.950 ;
        RECT 272.250 693.600 273.450 705.600 ;
        RECT 274.950 703.950 277.050 706.050 ;
        RECT 275.400 700.050 276.450 703.950 ;
        RECT 280.950 700.950 283.050 703.050 ;
        RECT 274.950 697.950 277.050 700.050 ;
        RECT 274.950 695.850 277.050 696.750 ;
        RECT 271.950 691.500 274.050 693.600 ;
        RECT 274.950 691.950 277.050 694.050 ;
        RECT 275.400 673.050 276.450 691.950 ;
        RECT 281.400 673.050 282.450 700.950 ;
        RECT 241.950 670.950 244.050 673.050 ;
        RECT 250.950 670.950 253.050 673.050 ;
        RECT 259.950 670.950 262.050 673.050 ;
        RECT 268.950 670.950 271.050 673.050 ;
        RECT 274.950 670.950 277.050 673.050 ;
        RECT 278.250 671.250 279.750 672.150 ;
        RECT 280.950 670.950 283.050 673.050 ;
        RECT 226.950 668.250 228.750 669.150 ;
        RECT 229.950 667.950 232.050 670.050 ;
        RECT 235.950 667.950 238.050 670.050 ;
        RECT 166.950 664.950 169.050 667.050 ;
        RECT 170.250 665.850 171.750 666.750 ;
        RECT 172.950 664.950 175.050 667.050 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 191.250 665.850 192.750 666.750 ;
        RECT 193.950 664.950 196.050 667.050 ;
        RECT 199.950 664.950 202.050 667.050 ;
        RECT 202.950 665.850 204.750 666.750 ;
        RECT 205.950 664.950 208.050 667.050 ;
        RECT 209.250 665.850 210.750 666.750 ;
        RECT 211.950 664.950 214.050 667.050 ;
        RECT 217.950 664.950 220.050 667.050 ;
        RECT 226.950 664.950 229.050 667.050 ;
        RECT 230.250 665.850 231.750 666.750 ;
        RECT 232.950 664.950 235.050 667.050 ;
        RECT 236.250 665.850 238.050 666.750 ;
        RECT 167.400 661.050 168.450 664.950 ;
        RECT 173.400 663.450 174.450 664.950 ;
        RECT 170.400 662.400 174.450 663.450 ;
        RECT 166.950 658.950 169.050 661.050 ;
        RECT 167.400 622.050 168.450 658.950 ;
        RECT 170.400 634.050 171.450 662.400 ;
        RECT 194.400 652.050 195.450 664.950 ;
        RECT 205.950 662.850 208.050 663.750 ;
        RECT 208.950 661.950 211.050 664.050 ;
        RECT 229.950 661.950 232.050 664.050 ;
        RECT 232.950 662.850 235.050 663.750 ;
        RECT 193.950 649.950 196.050 652.050 ;
        RECT 205.950 649.950 208.050 652.050 ;
        RECT 193.950 646.950 196.050 649.050 ;
        RECT 175.950 635.250 178.050 636.150 ;
        RECT 194.400 634.050 195.450 646.950 ;
        RECT 199.950 635.250 202.050 636.150 ;
        RECT 169.950 631.950 172.050 634.050 ;
        RECT 173.250 632.250 174.750 633.150 ;
        RECT 175.950 631.950 178.050 634.050 ;
        RECT 179.250 632.250 181.050 633.150 ;
        RECT 193.950 631.950 196.050 634.050 ;
        RECT 197.250 632.250 198.750 633.150 ;
        RECT 199.950 631.950 202.050 634.050 ;
        RECT 203.250 632.250 205.050 633.150 ;
        RECT 169.950 629.850 171.750 630.750 ;
        RECT 172.950 628.950 175.050 631.050 ;
        RECT 176.400 628.050 177.450 631.950 ;
        RECT 178.950 628.950 181.050 631.050 ;
        RECT 193.950 629.850 195.750 630.750 ;
        RECT 196.950 628.950 199.050 631.050 ;
        RECT 175.950 625.950 178.050 628.050 ;
        RECT 179.400 625.050 180.450 628.950 ;
        RECT 178.950 622.950 181.050 625.050 ;
        RECT 166.950 619.950 169.050 622.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 173.400 601.050 174.450 601.950 ;
        RECT 166.950 599.250 169.050 600.150 ;
        RECT 172.950 598.950 175.050 601.050 ;
        RECT 176.250 599.250 178.050 600.150 ;
        RECT 166.950 595.950 169.050 598.050 ;
        RECT 172.950 596.850 174.750 597.750 ;
        RECT 175.950 595.950 178.050 598.050 ;
        RECT 176.400 595.050 177.450 595.950 ;
        RECT 175.950 592.950 178.050 595.050 ;
        RECT 179.400 588.450 180.450 622.950 ;
        RECT 197.400 619.050 198.450 628.950 ;
        RECT 200.400 628.050 201.450 631.950 ;
        RECT 202.950 628.950 205.050 631.050 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 196.950 616.950 199.050 619.050 ;
        RECT 197.400 604.050 198.450 616.950 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 200.400 601.050 201.450 601.950 ;
        RECT 181.950 598.950 184.050 601.050 ;
        RECT 193.950 598.950 196.050 601.050 ;
        RECT 197.250 599.850 198.750 600.750 ;
        RECT 199.950 598.950 202.050 601.050 ;
        RECT 203.400 598.050 204.450 628.950 ;
        RECT 181.950 596.850 184.050 597.750 ;
        RECT 193.950 596.850 196.050 597.750 ;
        RECT 199.950 596.850 202.050 597.750 ;
        RECT 202.950 595.950 205.050 598.050 ;
        RECT 199.950 592.950 202.050 595.050 ;
        RECT 179.400 587.400 183.450 588.450 ;
        RECT 166.950 565.950 169.050 568.050 ;
        RECT 169.950 567.300 172.050 569.400 ;
        RECT 160.950 557.250 163.050 558.150 ;
        RECT 163.950 556.950 166.050 559.050 ;
        RECT 167.400 556.050 168.450 565.950 ;
        RECT 170.550 563.700 171.750 567.300 ;
        RECT 169.950 561.600 172.050 563.700 ;
        RECT 160.950 553.950 163.050 556.050 ;
        RECT 166.950 555.450 169.050 556.050 ;
        RECT 164.400 554.400 169.050 555.450 ;
        RECT 161.400 547.050 162.450 553.950 ;
        RECT 160.950 544.950 163.050 547.050 ;
        RECT 157.950 532.950 160.050 535.050 ;
        RECT 158.400 529.050 159.450 532.950 ;
        RECT 164.400 531.450 165.450 554.400 ;
        RECT 166.950 553.950 169.050 554.400 ;
        RECT 166.950 551.850 169.050 552.750 ;
        RECT 170.550 549.600 171.750 561.600 ;
        RECT 172.950 559.950 175.050 562.050 ;
        RECT 169.950 547.500 172.050 549.600 ;
        RECT 166.950 531.450 169.050 532.050 ;
        RECT 164.400 530.400 169.050 531.450 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 155.250 527.250 156.750 528.150 ;
        RECT 157.950 526.950 160.050 529.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 148.950 525.450 151.050 526.050 ;
        RECT 146.400 524.400 151.050 525.450 ;
        RECT 152.250 524.850 153.750 525.750 ;
        RECT 146.400 520.050 147.450 524.400 ;
        RECT 148.950 523.950 151.050 524.400 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 158.250 524.850 160.050 525.750 ;
        RECT 148.950 521.850 151.050 522.750 ;
        RECT 145.950 517.950 148.050 520.050 ;
        RECT 142.950 493.950 145.050 496.050 ;
        RECT 145.950 493.950 148.050 496.050 ;
        RECT 139.950 448.950 142.050 451.050 ;
        RECT 127.950 442.950 130.050 445.050 ;
        RECT 136.950 442.950 139.050 445.050 ;
        RECT 124.950 391.950 127.050 394.050 ;
        RECT 119.400 389.400 123.450 390.450 ;
        RECT 119.400 385.050 120.450 389.400 ;
        RECT 125.400 385.050 126.450 391.950 ;
        RECT 118.950 382.950 121.050 385.050 ;
        RECT 122.250 383.250 123.750 384.150 ;
        RECT 124.950 382.950 127.050 385.050 ;
        RECT 115.950 381.450 118.050 382.050 ;
        RECT 113.400 380.400 118.050 381.450 ;
        RECT 119.250 380.850 120.750 381.750 ;
        RECT 113.400 373.050 114.450 380.400 ;
        RECT 115.950 379.950 118.050 380.400 ;
        RECT 121.950 379.950 124.050 382.050 ;
        RECT 125.250 380.850 127.050 381.750 ;
        RECT 115.950 377.850 118.050 378.750 ;
        RECT 122.400 378.450 123.450 379.950 ;
        RECT 119.400 377.400 123.450 378.450 ;
        RECT 112.950 370.950 115.050 373.050 ;
        RECT 109.950 343.950 112.050 346.050 ;
        RECT 110.400 340.050 111.450 343.950 ;
        RECT 119.400 343.050 120.450 377.400 ;
        RECT 124.950 344.250 127.050 345.150 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 115.950 341.250 117.750 342.150 ;
        RECT 118.950 340.950 121.050 343.050 ;
        RECT 122.250 341.250 123.750 342.150 ;
        RECT 124.950 340.950 127.050 343.050 ;
        RECT 109.950 337.950 112.050 340.050 ;
        RECT 106.950 316.950 109.050 319.050 ;
        RECT 88.950 313.950 91.050 316.050 ;
        RECT 100.950 313.950 103.050 316.050 ;
        RECT 106.950 313.950 109.050 316.050 ;
        RECT 85.950 310.950 88.050 313.050 ;
        RECT 89.250 311.850 90.750 312.750 ;
        RECT 91.950 310.950 94.050 313.050 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 85.950 308.850 88.050 309.750 ;
        RECT 91.950 308.850 94.050 309.750 ;
        RECT 101.400 307.050 102.450 313.950 ;
        RECT 113.400 313.050 114.450 340.950 ;
        RECT 128.400 340.050 129.450 442.950 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 130.950 410.850 133.050 411.750 ;
        RECT 133.950 410.250 136.050 411.150 ;
        RECT 133.950 406.950 136.050 409.050 ;
        RECT 134.400 403.050 135.450 406.950 ;
        RECT 133.950 400.950 136.050 403.050 ;
        RECT 136.950 385.950 139.050 388.050 ;
        RECT 137.400 385.050 138.450 385.950 ;
        RECT 133.950 383.250 135.750 384.150 ;
        RECT 136.950 382.950 139.050 385.050 ;
        RECT 133.950 379.950 136.050 382.050 ;
        RECT 137.250 380.850 139.050 381.750 ;
        RECT 134.400 379.050 135.450 379.950 ;
        RECT 133.950 376.950 136.050 379.050 ;
        RECT 140.400 376.050 141.450 448.950 ;
        RECT 143.400 387.450 144.450 493.950 ;
        RECT 146.400 490.050 147.450 493.950 ;
        RECT 164.400 492.450 165.450 530.400 ;
        RECT 166.950 529.950 169.050 530.400 ;
        RECT 173.400 529.050 174.450 559.950 ;
        RECT 178.950 557.250 181.050 558.150 ;
        RECT 182.400 556.050 183.450 587.400 ;
        RECT 190.950 566.400 193.050 568.500 ;
        RECT 184.950 557.250 187.050 558.150 ;
        RECT 178.950 553.950 181.050 556.050 ;
        RECT 181.950 553.950 184.050 556.050 ;
        RECT 184.950 555.450 187.050 556.050 ;
        RECT 184.950 554.400 189.450 555.450 ;
        RECT 184.950 553.950 187.050 554.400 ;
        RECT 179.400 550.050 180.450 553.950 ;
        RECT 178.950 547.950 181.050 550.050 ;
        RECT 179.400 538.050 180.450 547.950 ;
        RECT 178.950 535.950 181.050 538.050 ;
        RECT 188.400 529.050 189.450 554.400 ;
        RECT 191.400 549.600 192.600 566.400 ;
        RECT 193.950 556.950 196.050 559.050 ;
        RECT 190.950 547.500 193.050 549.600 ;
        RECT 166.950 527.850 169.050 528.750 ;
        RECT 169.950 527.250 172.050 528.150 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 185.250 527.250 186.750 528.150 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 169.950 525.450 172.050 526.050 ;
        RECT 173.400 525.450 174.450 526.950 ;
        RECT 169.950 524.400 174.450 525.450 ;
        RECT 181.950 524.850 183.750 525.750 ;
        RECT 169.950 523.950 172.050 524.400 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 188.250 524.850 189.750 525.750 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 161.400 491.400 165.450 492.450 ;
        RECT 145.950 487.950 148.050 490.050 ;
        RECT 151.950 489.450 154.050 490.050 ;
        RECT 149.250 488.250 150.750 489.150 ;
        RECT 151.950 488.400 156.450 489.450 ;
        RECT 151.950 487.950 154.050 488.400 ;
        RECT 145.950 485.850 147.750 486.750 ;
        RECT 148.950 484.950 151.050 487.050 ;
        RECT 152.250 485.850 154.050 486.750 ;
        RECT 155.400 478.050 156.450 488.400 ;
        RECT 151.950 475.950 154.050 478.050 ;
        RECT 154.950 475.950 157.050 478.050 ;
        RECT 152.400 457.050 153.450 475.950 ;
        RECT 161.400 457.050 162.450 491.400 ;
        RECT 163.950 488.250 166.050 489.150 ;
        RECT 170.400 487.050 171.450 523.950 ;
        RECT 185.400 517.050 186.450 523.950 ;
        RECT 190.950 521.850 193.050 522.750 ;
        RECT 184.950 514.950 187.050 517.050 ;
        RECT 178.950 499.950 181.050 502.050 ;
        RECT 187.950 499.950 190.050 502.050 ;
        RECT 163.950 484.950 166.050 487.050 ;
        RECT 167.250 485.250 168.750 486.150 ;
        RECT 169.950 484.950 172.050 487.050 ;
        RECT 173.250 485.250 175.050 486.150 ;
        RECT 179.400 484.050 180.450 499.950 ;
        RECT 181.950 495.300 184.050 497.400 ;
        RECT 182.550 491.700 183.750 495.300 ;
        RECT 181.950 489.600 184.050 491.700 ;
        RECT 166.950 481.950 169.050 484.050 ;
        RECT 170.250 482.850 171.750 483.750 ;
        RECT 172.950 481.950 175.050 484.050 ;
        RECT 178.950 481.950 181.050 484.050 ;
        RECT 163.950 478.950 166.050 481.050 ;
        RECT 164.400 460.050 165.450 478.950 ;
        RECT 167.400 463.050 168.450 481.950 ;
        RECT 173.400 478.050 174.450 481.950 ;
        RECT 178.950 479.850 181.050 480.750 ;
        RECT 172.950 475.950 175.050 478.050 ;
        RECT 182.550 477.600 183.750 489.600 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 185.400 478.050 186.450 484.950 ;
        RECT 181.950 475.500 184.050 477.600 ;
        RECT 184.950 475.950 187.050 478.050 ;
        RECT 166.950 460.950 169.050 463.050 ;
        RECT 163.950 457.950 166.050 460.050 ;
        RECT 151.950 454.950 154.050 457.050 ;
        RECT 160.950 454.950 163.050 457.050 ;
        RECT 166.950 454.950 169.050 457.050 ;
        RECT 169.950 454.950 172.050 457.050 ;
        RECT 173.250 455.250 175.050 456.150 ;
        RECT 178.950 454.950 181.050 457.050 ;
        RECT 182.250 455.250 184.050 456.150 ;
        RECT 151.950 452.850 154.050 453.750 ;
        RECT 157.950 452.850 160.050 453.750 ;
        RECT 167.400 418.050 168.450 454.950 ;
        RECT 169.950 452.850 171.750 453.750 ;
        RECT 172.950 451.950 175.050 454.050 ;
        RECT 178.950 452.850 180.750 453.750 ;
        RECT 181.950 453.450 184.050 454.050 ;
        RECT 185.400 453.450 186.450 475.950 ;
        RECT 188.400 459.450 189.450 499.950 ;
        RECT 190.950 485.250 193.050 486.150 ;
        RECT 190.950 481.950 193.050 484.050 ;
        RECT 191.400 481.050 192.450 481.950 ;
        RECT 190.950 478.950 193.050 481.050 ;
        RECT 194.400 460.050 195.450 556.950 ;
        RECT 196.950 485.250 199.050 486.150 ;
        RECT 196.950 481.950 199.050 484.050 ;
        RECT 197.400 478.050 198.450 481.950 ;
        RECT 196.950 475.950 199.050 478.050 ;
        RECT 190.950 459.450 193.050 460.050 ;
        RECT 188.400 458.400 193.050 459.450 ;
        RECT 188.400 457.050 189.450 458.400 ;
        RECT 190.950 457.950 193.050 458.400 ;
        RECT 193.950 457.950 196.050 460.050 ;
        RECT 196.950 457.950 199.050 460.050 ;
        RECT 187.950 454.950 190.050 457.050 ;
        RECT 190.950 455.850 193.050 456.750 ;
        RECT 193.950 455.250 196.050 456.150 ;
        RECT 181.950 452.400 186.450 453.450 ;
        RECT 193.950 453.450 196.050 454.050 ;
        RECT 197.400 453.450 198.450 457.950 ;
        RECT 193.950 452.400 198.450 453.450 ;
        RECT 181.950 451.950 184.050 452.400 ;
        RECT 193.950 451.950 196.050 452.400 ;
        RECT 173.400 451.050 174.450 451.950 ;
        RECT 172.950 448.950 175.050 451.050 ;
        RECT 178.950 448.950 181.050 451.050 ;
        RECT 172.950 421.950 175.050 424.050 ;
        RECT 173.400 418.050 174.450 421.950 ;
        RECT 166.950 417.450 169.050 418.050 ;
        RECT 164.400 416.400 169.050 417.450 ;
        RECT 145.950 413.250 148.050 414.150 ;
        RECT 151.950 413.250 154.050 414.150 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 146.400 406.050 147.450 409.950 ;
        RECT 148.950 406.950 151.050 409.050 ;
        RECT 145.950 403.950 148.050 406.050 ;
        RECT 143.400 386.400 147.450 387.450 ;
        RECT 146.400 385.050 147.450 386.400 ;
        RECT 142.950 383.250 144.750 384.150 ;
        RECT 145.950 382.950 148.050 385.050 ;
        RECT 142.950 379.950 145.050 382.050 ;
        RECT 146.250 380.850 148.050 381.750 ;
        RECT 139.950 373.950 142.050 376.050 ;
        RECT 143.400 370.050 144.450 379.950 ;
        RECT 149.400 379.050 150.450 406.950 ;
        RECT 151.950 400.950 154.050 403.050 ;
        RECT 148.950 376.950 151.050 379.050 ;
        RECT 148.950 370.950 151.050 373.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 133.950 346.950 136.050 349.050 ;
        RECT 136.950 346.950 139.050 349.050 ;
        RECT 115.950 337.950 118.050 340.050 ;
        RECT 119.250 338.850 120.750 339.750 ;
        RECT 121.950 337.950 124.050 340.050 ;
        RECT 127.950 337.950 130.050 340.050 ;
        RECT 116.400 334.050 117.450 337.950 ;
        RECT 115.950 331.950 118.050 334.050 ;
        RECT 124.950 316.950 127.050 319.050 ;
        RECT 103.950 311.250 106.050 312.150 ;
        RECT 106.950 311.850 109.050 312.750 ;
        RECT 109.950 311.250 111.750 312.150 ;
        RECT 112.950 310.950 115.050 313.050 ;
        RECT 103.950 307.950 106.050 310.050 ;
        RECT 109.950 307.950 112.050 310.050 ;
        RECT 113.250 308.850 115.050 309.750 ;
        RECT 100.950 304.950 103.050 307.050 ;
        RECT 82.950 277.950 85.050 280.050 ;
        RECT 67.950 273.450 70.050 274.050 ;
        RECT 65.400 272.400 70.050 273.450 ;
        RECT 65.400 265.050 66.450 272.400 ;
        RECT 67.950 271.950 70.050 272.400 ;
        RECT 71.250 272.250 72.750 273.150 ;
        RECT 73.950 271.950 76.050 274.050 ;
        RECT 79.950 271.950 82.050 274.050 ;
        RECT 67.950 269.850 69.750 270.750 ;
        RECT 70.950 268.950 73.050 271.050 ;
        RECT 74.250 269.850 76.050 270.750 ;
        RECT 80.400 268.050 81.450 271.950 ;
        RECT 79.950 265.950 82.050 268.050 ;
        RECT 64.950 262.950 67.050 265.050 ;
        RECT 73.950 262.950 76.050 265.050 ;
        RECT 58.950 247.950 61.050 250.050 ;
        RECT 55.950 241.950 58.050 244.050 ;
        RECT 64.950 241.950 67.050 244.050 ;
        RECT 52.950 238.950 55.050 241.050 ;
        RECT 61.950 238.950 64.050 241.050 ;
        RECT 52.950 236.250 54.750 237.150 ;
        RECT 55.950 235.950 58.050 238.050 ;
        RECT 59.250 236.250 61.050 237.150 ;
        RECT 52.950 232.950 55.050 235.050 ;
        RECT 56.250 233.850 57.750 234.750 ;
        RECT 58.950 234.450 61.050 235.050 ;
        RECT 62.400 234.450 63.450 238.950 ;
        RECT 58.950 233.400 63.450 234.450 ;
        RECT 58.950 232.950 61.050 233.400 ;
        RECT 65.400 199.050 66.450 241.950 ;
        RECT 74.400 241.050 75.450 262.950 ;
        RECT 80.400 241.050 81.450 265.950 ;
        RECT 73.950 238.950 76.050 241.050 ;
        RECT 77.250 239.250 78.750 240.150 ;
        RECT 79.950 238.950 82.050 241.050 ;
        RECT 70.950 235.950 73.050 238.050 ;
        RECT 74.250 236.850 75.750 237.750 ;
        RECT 76.950 235.950 79.050 238.050 ;
        RECT 80.250 236.850 82.050 237.750 ;
        RECT 70.950 233.850 73.050 234.750 ;
        RECT 73.950 232.950 76.050 235.050 ;
        RECT 52.950 196.950 55.050 199.050 ;
        RECT 64.950 196.950 67.050 199.050 ;
        RECT 49.950 194.850 52.050 195.750 ;
        RECT 53.400 174.450 54.450 196.950 ;
        RECT 74.400 196.050 75.450 232.950 ;
        RECT 77.400 229.050 78.450 235.950 ;
        RECT 76.950 226.950 79.050 229.050 ;
        RECT 76.950 207.300 79.050 209.400 ;
        RECT 77.550 203.700 78.750 207.300 ;
        RECT 76.950 201.600 79.050 203.700 ;
        RECT 64.950 194.850 67.050 195.750 ;
        RECT 73.950 195.450 76.050 196.050 ;
        RECT 67.950 194.250 70.050 195.150 ;
        RECT 71.400 194.400 76.050 195.450 ;
        RECT 67.950 192.450 70.050 193.050 ;
        RECT 71.400 192.450 72.450 194.400 ;
        RECT 73.950 193.950 76.050 194.400 ;
        RECT 67.950 191.400 72.450 192.450 ;
        RECT 73.950 191.850 76.050 192.750 ;
        RECT 67.950 190.950 70.050 191.400 ;
        RECT 55.950 187.950 58.050 190.050 ;
        RECT 77.550 189.600 78.750 201.600 ;
        RECT 50.400 173.400 54.450 174.450 ;
        RECT 50.400 169.050 51.450 173.400 ;
        RECT 56.400 169.050 57.450 187.950 ;
        RECT 76.950 187.500 79.050 189.600 ;
        RECT 49.950 166.950 52.050 169.050 ;
        RECT 53.250 167.250 54.750 168.150 ;
        RECT 55.950 166.950 58.050 169.050 ;
        RECT 61.950 166.950 64.050 169.050 ;
        RECT 49.950 164.850 51.750 165.750 ;
        RECT 52.950 163.950 55.050 166.050 ;
        RECT 56.250 164.850 57.750 165.750 ;
        RECT 58.950 163.950 61.050 166.050 ;
        RECT 53.400 163.050 54.450 163.950 ;
        RECT 52.950 160.950 55.050 163.050 ;
        RECT 58.950 161.850 61.050 162.750 ;
        RECT 43.950 151.950 46.050 154.050 ;
        RECT 28.950 134.400 31.050 136.500 ;
        RECT 22.950 123.450 25.050 124.050 ;
        RECT 20.400 122.400 25.050 123.450 ;
        RECT 22.950 121.950 25.050 122.400 ;
        RECT 25.950 121.950 28.050 124.050 ;
        RECT 7.950 115.500 10.050 117.600 ;
        RECT 11.400 111.450 12.450 121.950 ;
        RECT 8.400 110.400 12.450 111.450 ;
        RECT 8.400 100.050 9.450 110.400 ;
        RECT 7.950 99.450 10.050 100.050 ;
        RECT 5.400 98.400 10.050 99.450 ;
        RECT 5.400 55.050 6.450 98.400 ;
        RECT 7.950 97.950 10.050 98.400 ;
        RECT 7.950 95.850 10.050 96.750 ;
        RECT 10.950 95.250 13.050 96.150 ;
        RECT 10.950 93.450 13.050 94.050 ;
        RECT 14.400 93.450 15.450 121.950 ;
        RECT 17.400 121.050 18.450 121.950 ;
        RECT 16.950 118.950 19.050 121.050 ;
        RECT 29.400 117.600 30.600 134.400 ;
        RECT 58.950 127.950 61.050 130.050 ;
        RECT 46.950 124.950 49.050 127.050 ;
        RECT 52.950 125.250 55.050 126.150 ;
        RECT 46.950 122.850 49.050 123.750 ;
        RECT 52.950 121.950 55.050 124.050 ;
        RECT 56.250 122.250 58.050 123.150 ;
        RECT 55.950 120.450 58.050 121.050 ;
        RECT 59.400 120.450 60.450 127.950 ;
        RECT 53.400 119.400 60.450 120.450 ;
        RECT 28.950 115.500 31.050 117.600 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 35.400 100.050 36.450 100.950 ;
        RECT 34.950 97.950 37.050 100.050 ;
        RECT 53.400 97.050 54.450 119.400 ;
        RECT 55.950 118.950 58.050 119.400 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 28.950 96.450 31.050 97.050 ;
        RECT 10.950 92.400 15.450 93.450 ;
        RECT 26.400 95.400 31.050 96.450 ;
        RECT 10.950 91.950 13.050 92.400 ;
        RECT 11.400 61.050 12.450 91.950 ;
        RECT 10.950 58.950 13.050 61.050 ;
        RECT 10.950 56.250 13.050 57.150 ;
        RECT 4.950 52.950 7.050 55.050 ;
        RECT 10.950 52.950 13.050 55.050 ;
        RECT 14.250 53.250 15.750 54.150 ;
        RECT 16.950 52.950 19.050 55.050 ;
        RECT 20.250 53.250 22.050 54.150 ;
        RECT 26.400 52.050 27.450 95.400 ;
        RECT 28.950 94.950 31.050 95.400 ;
        RECT 32.250 95.250 34.050 96.150 ;
        RECT 34.950 95.850 37.050 96.750 ;
        RECT 37.950 95.250 40.050 96.150 ;
        RECT 46.950 94.950 49.050 97.050 ;
        RECT 50.250 95.250 51.750 96.150 ;
        RECT 52.950 94.950 55.050 97.050 ;
        RECT 56.400 94.050 57.450 100.950 ;
        RECT 62.400 97.050 63.450 166.950 ;
        RECT 73.950 164.250 75.750 165.150 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 80.250 164.250 82.050 165.150 ;
        RECT 73.950 160.950 76.050 163.050 ;
        RECT 77.250 161.850 78.750 162.750 ;
        RECT 83.400 130.050 84.450 277.950 ;
        RECT 91.950 274.950 94.050 277.050 ;
        RECT 85.950 272.250 88.050 273.150 ;
        RECT 92.400 271.050 93.450 274.950 ;
        RECT 85.950 268.950 88.050 271.050 ;
        RECT 89.250 269.250 90.750 270.150 ;
        RECT 91.950 268.950 94.050 271.050 ;
        RECT 95.250 269.250 97.050 270.150 ;
        RECT 88.950 265.950 91.050 268.050 ;
        RECT 92.250 266.850 93.750 267.750 ;
        RECT 94.950 265.950 97.050 268.050 ;
        RECT 89.400 262.050 90.450 265.950 ;
        RECT 101.400 265.050 102.450 304.950 ;
        RECT 104.400 274.050 105.450 307.950 ;
        RECT 103.950 271.950 106.050 274.050 ;
        RECT 118.950 271.950 121.050 274.050 ;
        RECT 109.950 269.250 112.050 270.150 ;
        RECT 115.950 269.250 118.050 270.150 ;
        RECT 109.950 265.950 112.050 268.050 ;
        RECT 115.950 267.450 118.050 268.050 ;
        RECT 119.400 267.450 120.450 271.950 ;
        RECT 121.950 268.950 124.050 271.050 ;
        RECT 113.250 266.250 114.750 267.150 ;
        RECT 115.950 266.400 120.450 267.450 ;
        RECT 115.950 265.950 118.050 266.400 ;
        RECT 100.950 262.950 103.050 265.050 ;
        RECT 88.950 259.950 91.050 262.050 ;
        RECT 89.400 235.050 90.450 259.950 ;
        RECT 97.950 247.950 100.050 250.050 ;
        RECT 91.950 244.950 94.050 247.050 ;
        RECT 92.400 241.050 93.450 244.950 ;
        RECT 94.950 241.950 97.050 244.050 ;
        RECT 98.400 241.050 99.450 247.950 ;
        RECT 110.400 247.050 111.450 265.950 ;
        RECT 122.400 265.050 123.450 268.950 ;
        RECT 125.400 265.050 126.450 316.950 ;
        RECT 134.400 316.050 135.450 346.950 ;
        RECT 137.400 343.050 138.450 346.950 ;
        RECT 136.950 340.950 139.050 343.050 ;
        RECT 139.950 341.250 142.050 342.150 ;
        RECT 145.950 341.250 148.050 342.150 ;
        RECT 139.950 339.450 142.050 340.050 ;
        RECT 137.400 338.400 142.050 339.450 ;
        RECT 145.950 339.450 148.050 340.050 ;
        RECT 149.400 339.450 150.450 370.950 ;
        RECT 133.950 313.950 136.050 316.050 ;
        RECT 130.950 310.950 133.050 313.050 ;
        RECT 131.400 310.050 132.450 310.950 ;
        RECT 137.400 310.050 138.450 338.400 ;
        RECT 139.950 337.950 142.050 338.400 ;
        RECT 143.250 338.250 144.750 339.150 ;
        RECT 145.950 338.400 150.450 339.450 ;
        RECT 145.950 337.950 148.050 338.400 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 152.400 334.050 153.450 400.950 ;
        RECT 164.400 388.050 165.450 416.400 ;
        RECT 166.950 415.950 169.050 416.400 ;
        RECT 170.250 416.250 171.750 417.150 ;
        RECT 172.950 415.950 175.050 418.050 ;
        RECT 166.950 413.850 168.750 414.750 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 173.250 413.850 175.050 414.750 ;
        RECT 175.950 391.950 178.050 394.050 ;
        RECT 163.950 385.950 166.050 388.050 ;
        RECT 163.950 384.450 166.050 385.050 ;
        RECT 169.950 384.450 172.050 385.050 ;
        RECT 163.950 383.400 168.450 384.450 ;
        RECT 163.950 382.950 166.050 383.400 ;
        RECT 163.950 380.850 166.050 381.750 ;
        RECT 167.400 373.050 168.450 383.400 ;
        RECT 169.950 383.400 174.450 384.450 ;
        RECT 169.950 382.950 172.050 383.400 ;
        RECT 169.950 380.850 172.050 381.750 ;
        RECT 166.950 370.950 169.050 373.050 ;
        RECT 169.950 349.950 172.050 352.050 ;
        RECT 170.400 346.050 171.450 349.950 ;
        RECT 154.950 343.950 157.050 346.050 ;
        RECT 157.950 344.250 160.050 345.150 ;
        RECT 169.950 343.950 172.050 346.050 ;
        RECT 155.400 342.450 156.450 343.950 ;
        RECT 157.950 342.450 160.050 343.050 ;
        RECT 155.400 341.400 160.050 342.450 ;
        RECT 157.950 340.950 160.050 341.400 ;
        RECT 161.250 341.250 162.750 342.150 ;
        RECT 163.950 340.950 166.050 343.050 ;
        RECT 167.250 341.250 169.050 342.150 ;
        RECT 160.950 337.950 163.050 340.050 ;
        RECT 164.250 338.850 165.750 339.750 ;
        RECT 166.950 339.450 169.050 340.050 ;
        RECT 170.400 339.450 171.450 343.950 ;
        RECT 166.950 338.400 171.450 339.450 ;
        RECT 173.400 339.450 174.450 383.400 ;
        RECT 176.400 346.050 177.450 391.950 ;
        RECT 175.950 343.950 178.050 346.050 ;
        RECT 175.950 341.250 178.050 342.150 ;
        RECT 175.950 339.450 178.050 340.050 ;
        RECT 173.400 338.400 178.050 339.450 ;
        RECT 166.950 337.950 169.050 338.400 ;
        RECT 175.950 337.950 178.050 338.400 ;
        RECT 151.950 331.950 154.050 334.050 ;
        RECT 172.950 331.950 175.050 334.050 ;
        RECT 148.950 325.950 151.050 328.050 ;
        RECT 149.400 319.050 150.450 325.950 ;
        RECT 148.950 316.950 151.050 319.050 ;
        RECT 149.400 313.050 150.450 316.950 ;
        RECT 166.950 313.950 169.050 316.050 ;
        RECT 142.950 312.450 145.050 313.050 ;
        RECT 140.400 311.400 145.050 312.450 ;
        RECT 127.950 308.250 129.750 309.150 ;
        RECT 130.950 307.950 133.050 310.050 ;
        RECT 134.250 308.250 136.050 309.150 ;
        RECT 136.950 307.950 139.050 310.050 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 131.250 305.850 132.750 306.750 ;
        RECT 133.950 304.950 136.050 307.050 ;
        RECT 134.400 304.050 135.450 304.950 ;
        RECT 133.950 301.950 136.050 304.050 ;
        RECT 134.400 277.050 135.450 301.950 ;
        RECT 140.400 301.050 141.450 311.400 ;
        RECT 142.950 310.950 145.050 311.400 ;
        RECT 146.250 311.250 147.750 312.150 ;
        RECT 148.950 310.950 151.050 313.050 ;
        RECT 142.950 308.850 144.750 309.750 ;
        RECT 145.950 307.950 148.050 310.050 ;
        RECT 149.250 308.850 150.750 309.750 ;
        RECT 151.950 307.950 154.050 310.050 ;
        RECT 139.950 298.950 142.050 301.050 ;
        RECT 133.950 274.950 136.050 277.050 ;
        RECT 139.950 274.950 142.050 277.050 ;
        RECT 127.950 271.950 130.050 274.050 ;
        RECT 128.400 271.050 129.450 271.950 ;
        RECT 127.950 268.950 130.050 271.050 ;
        RECT 133.950 268.950 136.050 271.050 ;
        RECT 137.250 269.250 139.050 270.150 ;
        RECT 127.950 266.850 130.050 267.750 ;
        RECT 130.950 266.250 133.050 267.150 ;
        RECT 133.950 266.850 135.750 267.750 ;
        RECT 136.950 265.950 139.050 268.050 ;
        RECT 112.950 262.950 115.050 265.050 ;
        RECT 121.950 262.950 124.050 265.050 ;
        RECT 124.950 262.950 127.050 265.050 ;
        RECT 130.950 262.950 133.050 265.050 ;
        RECT 131.400 262.050 132.450 262.950 ;
        RECT 130.950 259.950 133.050 262.050 ;
        RECT 137.400 247.050 138.450 265.950 ;
        RECT 109.950 244.950 112.050 247.050 ;
        RECT 112.950 244.950 115.050 247.050 ;
        RECT 136.950 244.950 139.050 247.050 ;
        RECT 106.950 241.950 109.050 244.050 ;
        RECT 91.950 238.950 94.050 241.050 ;
        RECT 95.250 239.850 96.750 240.750 ;
        RECT 97.950 238.950 100.050 241.050 ;
        RECT 91.950 236.850 94.050 237.750 ;
        RECT 97.950 236.850 100.050 237.750 ;
        RECT 88.950 232.950 91.050 235.050 ;
        RECT 107.400 232.050 108.450 241.950 ;
        RECT 113.400 240.450 114.450 244.950 ;
        RECT 140.400 244.050 141.450 274.950 ;
        RECT 121.950 241.950 124.050 244.050 ;
        RECT 139.950 241.950 142.050 244.050 ;
        RECT 110.400 239.400 114.450 240.450 ;
        RECT 106.950 229.950 109.050 232.050 ;
        RECT 97.950 206.400 100.050 208.500 ;
        RECT 85.950 197.250 88.050 198.150 ;
        RECT 91.950 197.250 94.050 198.150 ;
        RECT 85.950 193.950 88.050 196.050 ;
        RECT 91.950 193.950 94.050 196.050 ;
        RECT 86.400 175.050 87.450 193.950 ;
        RECT 92.400 190.050 93.450 193.950 ;
        RECT 91.950 187.950 94.050 190.050 ;
        RECT 98.400 189.600 99.600 206.400 ;
        RECT 97.950 187.500 100.050 189.600 ;
        RECT 103.950 187.950 106.050 190.050 ;
        RECT 94.950 175.950 97.050 178.050 ;
        RECT 85.950 172.950 88.050 175.050 ;
        RECT 88.950 172.950 91.050 175.050 ;
        RECT 85.950 134.400 88.050 136.500 ;
        RECT 70.950 127.950 73.050 130.050 ;
        RECT 74.250 128.250 75.750 129.150 ;
        RECT 76.950 127.950 79.050 130.050 ;
        RECT 82.950 127.950 85.050 130.050 ;
        RECT 67.950 124.950 70.050 127.050 ;
        RECT 70.950 125.850 72.750 126.750 ;
        RECT 73.950 124.950 76.050 127.050 ;
        RECT 77.250 125.850 79.050 126.750 ;
        RECT 61.950 94.950 64.050 97.050 ;
        RECT 28.950 92.850 30.750 93.750 ;
        RECT 31.950 91.950 34.050 94.050 ;
        RECT 34.950 91.950 37.050 94.050 ;
        RECT 37.950 91.950 40.050 94.050 ;
        RECT 46.950 92.850 48.750 93.750 ;
        RECT 49.950 91.950 52.050 94.050 ;
        RECT 53.250 92.850 54.750 93.750 ;
        RECT 55.950 91.950 58.050 94.050 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 13.950 49.950 16.050 52.050 ;
        RECT 17.250 50.850 18.750 51.750 ;
        RECT 19.950 49.950 22.050 52.050 ;
        RECT 25.950 49.950 28.050 52.050 ;
        RECT 28.950 50.250 31.050 51.150 ;
        RECT 31.950 50.850 34.050 51.750 ;
        RECT 14.400 46.050 15.450 49.950 ;
        RECT 16.950 46.950 19.050 49.050 ;
        RECT 26.400 48.450 27.450 49.950 ;
        RECT 28.950 48.450 31.050 49.050 ;
        RECT 26.400 47.400 31.050 48.450 ;
        RECT 28.950 46.950 31.050 47.400 ;
        RECT 13.950 43.950 16.050 46.050 ;
        RECT 13.950 34.950 16.050 37.050 ;
        RECT 14.400 25.050 15.450 34.950 ;
        RECT 17.400 28.050 18.450 46.950 ;
        RECT 35.400 28.050 36.450 91.950 ;
        RECT 38.400 85.050 39.450 91.950 ;
        RECT 50.400 85.050 51.450 91.950 ;
        RECT 55.950 89.850 58.050 90.750 ;
        RECT 68.400 90.450 69.450 124.950 ;
        RECT 74.400 97.050 75.450 124.950 ;
        RECT 83.400 124.050 84.450 127.950 ;
        RECT 82.950 121.950 85.050 124.050 ;
        RECT 86.400 117.600 87.600 134.400 ;
        RECT 89.400 124.050 90.450 172.950 ;
        RECT 95.400 166.050 96.450 175.950 ;
        RECT 104.400 169.050 105.450 187.950 ;
        RECT 106.950 169.950 109.050 172.050 ;
        RECT 97.950 166.950 100.050 169.050 ;
        RECT 101.250 167.250 102.750 168.150 ;
        RECT 103.950 166.950 106.050 169.050 ;
        RECT 94.950 163.950 97.050 166.050 ;
        RECT 98.250 164.850 99.750 165.750 ;
        RECT 100.950 163.950 103.050 166.050 ;
        RECT 104.250 164.850 106.050 165.750 ;
        RECT 94.950 161.850 97.050 162.750 ;
        RECT 107.400 141.450 108.450 169.950 ;
        RECT 110.400 166.050 111.450 239.400 ;
        RECT 112.950 236.250 114.750 237.150 ;
        RECT 115.950 235.950 118.050 238.050 ;
        RECT 119.250 236.250 121.050 237.150 ;
        RECT 112.950 232.950 115.050 235.050 ;
        RECT 116.250 233.850 117.750 234.750 ;
        RECT 118.950 234.450 121.050 235.050 ;
        RECT 122.400 234.450 123.450 241.950 ;
        RECT 140.400 241.050 141.450 241.950 ;
        RECT 124.950 238.950 127.050 241.050 ;
        RECT 133.950 238.950 136.050 241.050 ;
        RECT 137.250 239.250 138.750 240.150 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 118.950 233.400 123.450 234.450 ;
        RECT 118.950 232.950 121.050 233.400 ;
        RECT 118.950 226.950 121.050 229.050 ;
        RECT 119.400 202.050 120.450 226.950 ;
        RECT 125.400 202.050 126.450 238.950 ;
        RECT 130.950 235.950 133.050 238.050 ;
        RECT 134.250 236.850 135.750 237.750 ;
        RECT 136.950 235.950 139.050 238.050 ;
        RECT 140.250 236.850 142.050 237.750 ;
        RECT 130.950 233.850 133.050 234.750 ;
        RECT 146.400 202.050 147.450 307.950 ;
        RECT 151.950 305.850 154.050 306.750 ;
        RECT 148.950 298.950 151.050 301.050 ;
        RECT 149.400 274.050 150.450 298.950 ;
        RECT 148.950 271.950 151.050 274.050 ;
        RECT 149.400 271.050 150.450 271.950 ;
        RECT 148.950 268.950 151.050 271.050 ;
        RECT 154.950 268.950 157.050 271.050 ;
        RECT 158.250 269.250 160.050 270.150 ;
        RECT 167.400 268.050 168.450 313.950 ;
        RECT 173.400 313.050 174.450 331.950 ;
        RECT 176.400 322.050 177.450 337.950 ;
        RECT 179.400 334.050 180.450 448.950 ;
        RECT 182.400 424.050 183.450 451.950 ;
        RECT 181.950 421.950 184.050 424.050 ;
        RECT 182.400 409.050 183.450 421.950 ;
        RECT 194.400 417.450 195.450 451.950 ;
        RECT 200.400 450.450 201.450 592.950 ;
        RECT 206.400 564.450 207.450 649.950 ;
        RECT 209.400 622.050 210.450 661.950 ;
        RECT 223.950 632.250 226.050 633.150 ;
        RECT 214.950 629.250 216.750 630.150 ;
        RECT 217.950 628.950 220.050 631.050 ;
        RECT 221.250 629.250 222.750 630.150 ;
        RECT 223.950 628.950 226.050 631.050 ;
        RECT 224.400 628.050 225.450 628.950 ;
        RECT 211.950 625.950 214.050 628.050 ;
        RECT 214.950 625.950 217.050 628.050 ;
        RECT 218.250 626.850 219.750 627.750 ;
        RECT 220.950 625.950 223.050 628.050 ;
        RECT 223.950 625.950 226.050 628.050 ;
        RECT 208.950 619.950 211.050 622.050 ;
        RECT 212.400 604.050 213.450 625.950 ;
        RECT 215.400 613.050 216.450 625.950 ;
        RECT 221.400 622.050 222.450 625.950 ;
        RECT 220.950 619.950 223.050 622.050 ;
        RECT 226.950 616.950 229.050 619.050 ;
        RECT 214.950 610.950 217.050 613.050 ;
        RECT 223.950 610.950 226.050 613.050 ;
        RECT 211.950 603.450 214.050 604.050 ;
        RECT 209.400 602.400 214.050 603.450 ;
        RECT 209.400 595.050 210.450 602.400 ;
        RECT 211.950 601.950 214.050 602.400 ;
        RECT 211.950 599.850 214.050 600.750 ;
        RECT 214.950 599.250 217.050 600.150 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 214.950 595.950 217.050 598.050 ;
        RECT 208.950 592.950 211.050 595.050 ;
        RECT 203.400 563.400 207.450 564.450 ;
        RECT 203.400 502.050 204.450 563.400 ;
        RECT 208.950 561.450 211.050 562.050 ;
        RECT 206.400 560.400 211.050 561.450 ;
        RECT 206.400 553.050 207.450 560.400 ;
        RECT 208.950 559.950 211.050 560.400 ;
        RECT 212.250 560.250 213.750 561.150 ;
        RECT 208.950 557.850 210.750 558.750 ;
        RECT 211.950 556.950 214.050 559.050 ;
        RECT 215.250 557.850 217.050 558.750 ;
        RECT 205.950 550.950 208.050 553.050 ;
        RECT 218.400 532.050 219.450 598.950 ;
        RECT 224.400 538.050 225.450 610.950 ;
        RECT 227.400 598.050 228.450 616.950 ;
        RECT 230.400 601.050 231.450 661.950 ;
        RECT 242.400 634.050 243.450 670.950 ;
        RECT 244.950 667.950 247.050 670.050 ;
        RECT 250.950 668.850 253.050 669.750 ;
        RECT 253.950 668.250 256.050 669.150 ;
        RECT 259.950 668.850 262.050 669.750 ;
        RECT 241.950 631.950 244.050 634.050 ;
        RECT 242.400 631.050 243.450 631.950 ;
        RECT 241.950 628.950 244.050 631.050 ;
        RECT 235.950 625.950 238.050 628.050 ;
        RECT 238.950 626.250 241.050 627.150 ;
        RECT 241.950 626.850 244.050 627.750 ;
        RECT 236.400 601.050 237.450 625.950 ;
        RECT 245.400 625.050 246.450 667.950 ;
        RECT 253.950 666.450 256.050 667.050 ;
        RECT 251.400 665.400 256.050 666.450 ;
        RECT 238.950 622.950 241.050 625.050 ;
        RECT 244.950 622.950 247.050 625.050 ;
        RECT 239.400 619.050 240.450 622.950 ;
        RECT 238.950 616.950 241.050 619.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 229.950 598.950 232.050 601.050 ;
        RECT 232.950 598.950 235.050 601.050 ;
        RECT 235.950 598.950 238.050 601.050 ;
        RECT 239.250 599.250 240.750 600.150 ;
        RECT 241.950 598.950 244.050 601.050 ;
        RECT 233.400 598.050 234.450 598.950 ;
        RECT 226.950 595.950 229.050 598.050 ;
        RECT 232.950 595.950 235.050 598.050 ;
        RECT 236.250 596.850 237.750 597.750 ;
        RECT 238.950 595.950 241.050 598.050 ;
        RECT 242.250 596.850 244.050 597.750 ;
        RECT 232.950 593.850 235.050 594.750 ;
        RECT 232.950 571.950 235.050 574.050 ;
        RECT 233.400 562.050 234.450 571.950 ;
        RECT 245.400 568.050 246.450 601.950 ;
        RECT 251.400 592.050 252.450 665.400 ;
        RECT 253.950 664.950 256.050 665.400 ;
        RECT 259.950 635.250 262.050 636.150 ;
        RECT 256.950 632.250 258.750 633.150 ;
        RECT 259.950 631.950 262.050 634.050 ;
        RECT 263.250 632.250 264.750 633.150 ;
        RECT 265.950 631.950 268.050 634.050 ;
        RECT 260.400 631.050 261.450 631.950 ;
        RECT 256.950 628.950 259.050 631.050 ;
        RECT 259.950 628.950 262.050 631.050 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 266.250 629.850 268.050 630.750 ;
        RECT 257.400 625.050 258.450 628.950 ;
        RECT 256.950 622.950 259.050 625.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 253.950 600.450 256.050 601.050 ;
        RECT 253.950 599.400 258.450 600.450 ;
        RECT 253.950 598.950 256.050 599.400 ;
        RECT 253.950 596.850 256.050 597.750 ;
        RECT 250.950 589.950 253.050 592.050 ;
        RECT 257.400 589.050 258.450 599.400 ;
        RECT 259.950 598.950 262.050 601.050 ;
        RECT 259.950 596.850 262.050 597.750 ;
        RECT 256.950 586.950 259.050 589.050 ;
        RECT 259.950 580.950 262.050 583.050 ;
        RECT 244.950 565.950 247.050 568.050 ;
        RECT 226.950 560.250 229.050 561.150 ;
        RECT 232.950 559.950 235.050 562.050 ;
        RECT 233.400 559.050 234.450 559.950 ;
        RECT 245.400 559.050 246.450 565.950 ;
        RECT 226.950 556.950 229.050 559.050 ;
        RECT 230.250 557.250 231.750 558.150 ;
        RECT 232.950 556.950 235.050 559.050 ;
        RECT 236.250 557.250 238.050 558.150 ;
        RECT 244.950 556.950 247.050 559.050 ;
        RECT 250.950 556.950 253.050 559.050 ;
        RECT 254.250 557.250 256.050 558.150 ;
        RECT 229.950 553.950 232.050 556.050 ;
        RECT 233.250 554.850 234.750 555.750 ;
        RECT 235.950 553.950 238.050 556.050 ;
        RECT 244.950 554.850 247.050 555.750 ;
        RECT 247.950 554.250 250.050 555.150 ;
        RECT 250.950 554.850 252.750 555.750 ;
        RECT 253.950 553.950 256.050 556.050 ;
        RECT 223.950 535.950 226.050 538.050 ;
        RECT 220.950 533.400 223.050 535.500 ;
        RECT 217.950 529.950 220.050 532.050 ;
        RECT 205.950 524.250 207.750 525.150 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 212.250 524.250 214.050 525.150 ;
        RECT 205.950 520.950 208.050 523.050 ;
        RECT 209.250 521.850 210.750 522.750 ;
        RECT 206.400 517.050 207.450 520.950 ;
        RECT 205.950 514.950 208.050 517.050 ;
        RECT 221.400 516.600 222.600 533.400 ;
        RECT 226.950 528.450 229.050 529.050 ;
        RECT 230.400 528.450 231.450 553.950 ;
        RECT 236.400 553.050 237.450 553.950 ;
        RECT 235.950 550.950 238.050 553.050 ;
        RECT 247.950 550.950 250.050 553.050 ;
        RECT 247.950 541.950 250.050 544.050 ;
        RECT 232.950 535.950 235.050 538.050 ;
        RECT 233.400 529.050 234.450 535.950 ;
        RECT 238.950 532.950 241.050 535.050 ;
        RECT 241.950 533.400 244.050 535.500 ;
        RECT 226.950 527.400 231.450 528.450 ;
        RECT 226.950 526.950 229.050 527.400 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 226.950 524.850 229.050 525.750 ;
        RECT 232.950 524.850 235.050 525.750 ;
        RECT 202.950 499.950 205.050 502.050 ;
        RECT 202.950 494.400 205.050 496.500 ;
        RECT 203.400 477.600 204.600 494.400 ;
        RECT 202.950 475.500 205.050 477.600 ;
        RECT 202.950 460.950 205.050 463.050 ;
        RECT 184.950 416.250 187.050 417.150 ;
        RECT 191.400 416.400 195.450 417.450 ;
        RECT 197.400 449.400 201.450 450.450 ;
        RECT 191.400 415.050 192.450 416.400 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 188.250 413.250 189.750 414.150 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 194.250 413.250 196.050 414.150 ;
        RECT 187.950 409.950 190.050 412.050 ;
        RECT 191.250 410.850 192.750 411.750 ;
        RECT 193.950 409.950 196.050 412.050 ;
        RECT 194.400 409.050 195.450 409.950 ;
        RECT 181.950 406.950 184.050 409.050 ;
        RECT 193.950 406.950 196.050 409.050 ;
        RECT 184.950 384.450 187.050 385.050 ;
        RECT 182.400 383.400 187.050 384.450 ;
        RECT 182.400 364.050 183.450 383.400 ;
        RECT 184.950 382.950 187.050 383.400 ;
        RECT 188.250 383.250 189.750 384.150 ;
        RECT 190.950 382.950 193.050 385.050 ;
        RECT 184.950 380.850 186.750 381.750 ;
        RECT 187.950 379.950 190.050 382.050 ;
        RECT 191.250 380.850 192.750 381.750 ;
        RECT 193.950 379.950 196.050 382.050 ;
        RECT 193.950 377.850 196.050 378.750 ;
        RECT 181.950 361.950 184.050 364.050 ;
        RECT 181.950 341.250 184.050 342.150 ;
        RECT 184.950 340.950 187.050 343.050 ;
        RECT 181.950 339.450 184.050 340.050 ;
        RECT 185.400 339.450 186.450 340.950 ;
        RECT 197.400 340.050 198.450 449.400 ;
        RECT 199.950 415.950 202.050 418.050 ;
        RECT 200.400 403.050 201.450 415.950 ;
        RECT 199.950 400.950 202.050 403.050 ;
        RECT 203.400 379.050 204.450 460.950 ;
        RECT 206.400 454.050 207.450 514.950 ;
        RECT 220.950 514.500 223.050 516.600 ;
        RECT 226.950 499.950 229.050 502.050 ;
        RECT 227.400 490.050 228.450 499.950 ;
        RECT 220.950 489.450 223.050 490.050 ;
        RECT 218.400 488.400 223.050 489.450 ;
        RECT 218.400 487.050 219.450 488.400 ;
        RECT 220.950 487.950 223.050 488.400 ;
        RECT 224.250 488.250 225.750 489.150 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 217.950 484.950 220.050 487.050 ;
        RECT 220.950 485.850 222.750 486.750 ;
        RECT 223.950 484.950 226.050 487.050 ;
        RECT 227.250 485.850 229.050 486.750 ;
        RECT 239.400 483.450 240.450 532.950 ;
        RECT 242.250 521.400 243.450 533.400 ;
        RECT 244.950 530.250 247.050 531.150 ;
        RECT 244.950 528.450 247.050 529.050 ;
        RECT 248.400 528.450 249.450 541.950 ;
        RECT 250.950 529.950 253.050 532.050 ;
        RECT 244.950 527.400 249.450 528.450 ;
        RECT 244.950 526.950 247.050 527.400 ;
        RECT 241.950 519.300 244.050 521.400 ;
        RECT 242.250 515.700 243.450 519.300 ;
        RECT 241.950 513.600 244.050 515.700 ;
        RECT 241.950 485.250 244.050 486.150 ;
        RECT 241.950 483.450 244.050 484.050 ;
        RECT 239.400 482.400 244.050 483.450 ;
        RECT 245.400 483.450 246.450 526.950 ;
        RECT 247.950 485.250 250.050 486.150 ;
        RECT 247.950 483.450 250.050 484.050 ;
        RECT 245.400 482.400 250.050 483.450 ;
        RECT 241.950 481.950 244.050 482.400 ;
        RECT 247.950 481.950 250.050 482.400 ;
        RECT 214.950 475.950 217.050 478.050 ;
        RECT 208.950 457.950 211.050 460.050 ;
        RECT 209.400 457.050 210.450 457.950 ;
        RECT 215.400 457.050 216.450 475.950 ;
        RECT 238.950 457.950 241.050 460.050 ;
        RECT 208.950 454.950 211.050 457.050 ;
        RECT 212.250 455.250 213.750 456.150 ;
        RECT 214.950 454.950 217.050 457.050 ;
        RECT 205.950 451.950 208.050 454.050 ;
        RECT 208.950 452.850 210.750 453.750 ;
        RECT 211.950 451.950 214.050 454.050 ;
        RECT 215.250 452.850 216.750 453.750 ;
        RECT 217.950 451.950 220.050 454.050 ;
        RECT 229.950 452.250 231.750 453.150 ;
        RECT 232.950 451.950 235.050 454.050 ;
        RECT 236.250 452.250 238.050 453.150 ;
        RECT 212.400 451.050 213.450 451.950 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 217.950 449.850 220.050 450.750 ;
        RECT 233.250 449.850 234.750 450.750 ;
        RECT 235.950 448.950 238.050 451.050 ;
        RECT 205.950 415.950 208.050 418.050 ;
        RECT 211.950 417.450 214.050 418.050 ;
        RECT 209.250 416.250 210.750 417.150 ;
        RECT 211.950 416.400 216.450 417.450 ;
        RECT 211.950 415.950 214.050 416.400 ;
        RECT 205.950 413.850 207.750 414.750 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 212.250 413.850 214.050 414.750 ;
        RECT 215.400 409.050 216.450 416.400 ;
        RECT 217.950 415.950 220.050 418.050 ;
        RECT 226.950 417.450 229.050 418.050 ;
        RECT 224.400 416.400 229.050 417.450 ;
        RECT 214.950 406.950 217.050 409.050 ;
        RECT 215.400 394.050 216.450 406.950 ;
        RECT 214.950 391.950 217.050 394.050 ;
        RECT 205.950 380.250 207.750 381.150 ;
        RECT 208.950 379.950 211.050 382.050 ;
        RECT 212.250 380.250 214.050 381.150 ;
        RECT 202.950 376.950 205.050 379.050 ;
        RECT 205.950 376.950 208.050 379.050 ;
        RECT 209.250 377.850 210.750 378.750 ;
        RECT 211.950 376.950 214.050 379.050 ;
        RECT 202.950 370.950 205.050 373.050 ;
        RECT 199.950 341.250 202.050 342.150 ;
        RECT 181.950 338.400 186.450 339.450 ;
        RECT 181.950 337.950 184.050 338.400 ;
        RECT 196.950 337.950 199.050 340.050 ;
        RECT 199.950 339.450 202.050 340.050 ;
        RECT 203.400 339.450 204.450 370.950 ;
        RECT 206.400 364.050 207.450 376.950 ;
        RECT 218.400 373.050 219.450 415.950 ;
        RECT 224.400 412.050 225.450 416.400 ;
        RECT 226.950 415.950 229.050 416.400 ;
        RECT 230.250 416.250 231.750 417.150 ;
        RECT 232.950 415.950 235.050 418.050 ;
        RECT 226.950 413.850 228.750 414.750 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 233.250 413.850 235.050 414.750 ;
        RECT 223.950 409.950 226.050 412.050 ;
        RECT 224.400 385.050 225.450 409.950 ;
        RECT 230.400 403.050 231.450 412.950 ;
        RECT 229.950 400.950 232.050 403.050 ;
        RECT 239.400 385.050 240.450 457.950 ;
        RECT 244.950 448.950 247.050 451.050 ;
        RECT 220.950 382.950 223.050 385.050 ;
        RECT 223.950 382.950 226.050 385.050 ;
        RECT 226.950 383.250 228.750 384.150 ;
        RECT 229.950 382.950 232.050 385.050 ;
        RECT 235.950 383.250 237.750 384.150 ;
        RECT 238.950 382.950 241.050 385.050 ;
        RECT 217.950 370.950 220.050 373.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 205.950 361.950 208.050 364.050 ;
        RECT 205.950 341.250 208.050 342.150 ;
        RECT 199.950 338.400 204.450 339.450 ;
        RECT 199.950 337.950 202.050 338.400 ;
        RECT 178.950 331.950 181.050 334.050 ;
        RECT 196.950 328.950 199.050 331.050 ;
        RECT 197.400 322.050 198.450 328.950 ;
        RECT 175.950 319.950 178.050 322.050 ;
        RECT 196.950 319.950 199.050 322.050 ;
        RECT 197.400 313.050 198.450 319.950 ;
        RECT 212.400 313.050 213.450 367.950 ;
        RECT 214.950 361.950 217.050 364.050 ;
        RECT 215.400 343.050 216.450 361.950 ;
        RECT 214.950 340.950 217.050 343.050 ;
        RECT 218.250 341.250 220.050 342.150 ;
        RECT 214.950 338.850 216.750 339.750 ;
        RECT 217.950 337.950 220.050 340.050 ;
        RECT 218.400 334.050 219.450 337.950 ;
        RECT 217.950 331.950 220.050 334.050 ;
        RECT 169.950 310.950 172.050 313.050 ;
        RECT 172.950 310.950 175.050 313.050 ;
        RECT 176.250 311.250 177.750 312.150 ;
        RECT 178.950 310.950 181.050 313.050 ;
        RECT 187.950 310.950 190.050 313.050 ;
        RECT 190.950 312.450 193.050 313.050 ;
        RECT 190.950 311.400 195.450 312.450 ;
        RECT 190.950 310.950 193.050 311.400 ;
        RECT 170.400 310.050 171.450 310.950 ;
        RECT 169.950 307.950 172.050 310.050 ;
        RECT 173.250 308.850 174.750 309.750 ;
        RECT 175.950 307.950 178.050 310.050 ;
        RECT 179.250 308.850 181.050 309.750 ;
        RECT 169.950 305.850 172.050 306.750 ;
        RECT 176.400 292.050 177.450 307.950 ;
        RECT 188.400 304.050 189.450 310.950 ;
        RECT 190.950 308.850 193.050 309.750 ;
        RECT 194.400 307.050 195.450 311.400 ;
        RECT 196.950 310.950 199.050 313.050 ;
        RECT 211.950 310.950 214.050 313.050 ;
        RECT 196.950 308.850 199.050 309.750 ;
        RECT 208.950 308.250 210.750 309.150 ;
        RECT 211.950 307.950 214.050 310.050 ;
        RECT 215.250 308.250 217.050 309.150 ;
        RECT 193.950 304.950 196.050 307.050 ;
        RECT 208.950 304.950 211.050 307.050 ;
        RECT 212.250 305.850 213.750 306.750 ;
        RECT 214.950 304.950 217.050 307.050 ;
        RECT 187.950 301.950 190.050 304.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 172.950 274.950 175.050 277.050 ;
        RECT 148.950 266.850 151.050 267.750 ;
        RECT 151.950 266.250 154.050 267.150 ;
        RECT 154.950 266.850 156.750 267.750 ;
        RECT 157.950 265.950 160.050 268.050 ;
        RECT 166.950 265.950 169.050 268.050 ;
        RECT 151.950 262.950 154.050 265.050 ;
        RECT 158.400 244.050 159.450 265.950 ;
        RECT 173.400 265.050 174.450 274.950 ;
        RECT 188.400 271.050 189.450 301.950 ;
        RECT 194.400 274.050 195.450 304.950 ;
        RECT 193.950 271.950 196.050 274.050 ;
        RECT 196.950 271.950 199.050 274.050 ;
        RECT 178.950 270.450 181.050 271.050 ;
        RECT 175.950 269.250 177.750 270.150 ;
        RECT 178.950 269.400 183.450 270.450 ;
        RECT 178.950 268.950 181.050 269.400 ;
        RECT 175.950 265.950 178.050 268.050 ;
        RECT 179.250 266.850 181.050 267.750 ;
        RECT 172.950 262.950 175.050 265.050 ;
        RECT 148.950 241.950 151.050 244.050 ;
        RECT 157.950 241.950 160.050 244.050 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 166.950 241.950 169.050 244.050 ;
        RECT 149.400 241.050 150.450 241.950 ;
        RECT 148.950 238.950 151.050 241.050 ;
        RECT 154.950 238.950 157.050 241.050 ;
        RECT 149.400 234.450 150.450 238.950 ;
        RECT 155.400 238.050 156.450 238.950 ;
        RECT 151.950 236.250 153.750 237.150 ;
        RECT 154.950 235.950 157.050 238.050 ;
        RECT 158.250 236.250 160.050 237.150 ;
        RECT 151.950 234.450 154.050 235.050 ;
        RECT 149.400 233.400 154.050 234.450 ;
        RECT 155.250 233.850 156.750 234.750 ;
        RECT 151.950 232.950 154.050 233.400 ;
        RECT 157.950 232.950 160.050 235.050 ;
        RECT 158.400 222.450 159.450 232.950 ;
        RECT 155.400 221.400 159.450 222.450 ;
        RECT 112.950 199.950 115.050 202.050 ;
        RECT 118.950 199.950 121.050 202.050 ;
        RECT 124.950 201.450 127.050 202.050 ;
        RECT 122.250 200.250 123.750 201.150 ;
        RECT 124.950 200.400 129.450 201.450 ;
        RECT 124.950 199.950 127.050 200.400 ;
        RECT 113.400 172.050 114.450 199.950 ;
        RECT 118.950 197.850 120.750 198.750 ;
        RECT 121.950 196.950 124.050 199.050 ;
        RECT 125.250 197.850 127.050 198.750 ;
        RECT 128.400 193.050 129.450 200.400 ;
        RECT 136.950 200.250 139.050 201.150 ;
        RECT 142.950 199.950 145.050 202.050 ;
        RECT 145.950 199.950 148.050 202.050 ;
        RECT 143.400 199.050 144.450 199.950 ;
        RECT 136.950 196.950 139.050 199.050 ;
        RECT 140.250 197.250 141.750 198.150 ;
        RECT 142.950 196.950 145.050 199.050 ;
        RECT 146.250 197.250 148.050 198.150 ;
        RECT 139.950 193.950 142.050 196.050 ;
        RECT 143.250 194.850 144.750 195.750 ;
        RECT 145.950 193.950 148.050 196.050 ;
        RECT 146.400 193.050 147.450 193.950 ;
        RECT 127.950 190.950 130.050 193.050 ;
        RECT 145.950 190.950 148.050 193.050 ;
        RECT 155.400 190.050 156.450 221.400 ;
        RECT 164.400 211.050 165.450 241.950 ;
        RECT 166.950 239.850 169.050 240.750 ;
        RECT 169.950 239.250 172.050 240.150 ;
        RECT 176.400 238.050 177.450 265.950 ;
        RECT 182.400 253.050 183.450 269.400 ;
        RECT 184.950 269.250 186.750 270.150 ;
        RECT 187.950 268.950 190.050 271.050 ;
        RECT 184.950 265.950 187.050 268.050 ;
        RECT 188.250 266.850 190.050 267.750 ;
        RECT 185.400 265.050 186.450 265.950 ;
        RECT 184.950 262.950 187.050 265.050 ;
        RECT 181.950 250.950 184.050 253.050 ;
        RECT 190.950 247.950 193.050 250.050 ;
        RECT 191.400 244.050 192.450 247.950 ;
        RECT 190.950 241.950 193.050 244.050 ;
        RECT 184.950 240.450 187.050 241.050 ;
        RECT 182.400 239.400 187.050 240.450 ;
        RECT 169.950 235.950 172.050 238.050 ;
        RECT 175.950 235.950 178.050 238.050 ;
        RECT 163.950 208.950 166.050 211.050 ;
        RECT 157.950 200.250 160.050 201.150 ;
        RECT 164.400 199.050 165.450 208.950 ;
        RECT 170.400 199.050 171.450 235.950 ;
        RECT 182.400 202.050 183.450 239.400 ;
        RECT 184.950 238.950 187.050 239.400 ;
        RECT 188.250 239.250 190.050 240.150 ;
        RECT 190.950 239.850 193.050 240.750 ;
        RECT 193.950 239.250 196.050 240.150 ;
        RECT 184.950 236.850 186.750 237.750 ;
        RECT 187.950 235.950 190.050 238.050 ;
        RECT 193.950 237.450 196.050 238.050 ;
        RECT 197.400 237.450 198.450 271.950 ;
        RECT 202.950 269.250 205.050 270.150 ;
        RECT 208.950 269.250 211.050 270.150 ;
        RECT 202.950 265.950 205.050 268.050 ;
        RECT 215.400 259.050 216.450 304.950 ;
        RECT 218.400 265.050 219.450 331.950 ;
        RECT 221.400 274.050 222.450 382.950 ;
        RECT 226.950 379.950 229.050 382.050 ;
        RECT 230.250 380.850 232.050 381.750 ;
        RECT 235.950 379.950 238.050 382.050 ;
        RECT 239.250 380.850 241.050 381.750 ;
        RECT 227.400 364.050 228.450 379.950 ;
        RECT 226.950 361.950 229.050 364.050 ;
        RECT 236.400 358.050 237.450 379.950 ;
        RECT 235.950 355.950 238.050 358.050 ;
        RECT 223.950 349.950 226.050 352.050 ;
        RECT 224.400 343.050 225.450 349.950 ;
        RECT 229.950 346.950 232.050 349.050 ;
        RECT 230.400 343.050 231.450 346.950 ;
        RECT 223.950 340.950 226.050 343.050 ;
        RECT 227.250 341.250 229.050 342.150 ;
        RECT 229.950 340.950 232.050 343.050 ;
        RECT 223.950 338.850 225.750 339.750 ;
        RECT 226.950 337.950 229.050 340.050 ;
        RECT 236.400 330.450 237.450 355.950 ;
        RECT 241.950 341.250 244.050 342.150 ;
        RECT 241.950 337.950 244.050 340.050 ;
        RECT 236.400 329.400 240.450 330.450 ;
        RECT 226.950 310.950 229.050 313.050 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 220.950 271.950 223.050 274.050 ;
        RECT 224.400 271.050 225.450 307.950 ;
        RECT 227.400 306.450 228.450 310.950 ;
        RECT 229.950 308.250 231.750 309.150 ;
        RECT 232.950 307.950 235.050 310.050 ;
        RECT 236.250 308.250 238.050 309.150 ;
        RECT 229.950 306.450 232.050 307.050 ;
        RECT 227.400 305.400 232.050 306.450 ;
        RECT 233.250 305.850 234.750 306.750 ;
        RECT 229.950 304.950 232.050 305.400 ;
        RECT 235.950 304.950 238.050 307.050 ;
        RECT 232.950 301.950 235.050 304.050 ;
        RECT 220.950 269.250 223.050 270.150 ;
        RECT 223.950 268.950 226.050 271.050 ;
        RECT 226.950 269.250 229.050 270.150 ;
        RECT 233.400 268.050 234.450 301.950 ;
        RECT 236.400 301.050 237.450 304.950 ;
        RECT 239.400 304.050 240.450 329.400 ;
        RECT 238.950 301.950 241.050 304.050 ;
        RECT 235.950 298.950 238.050 301.050 ;
        RECT 242.400 298.050 243.450 337.950 ;
        RECT 245.400 322.050 246.450 448.950 ;
        RECT 251.400 418.050 252.450 529.950 ;
        RECT 254.400 529.050 255.450 553.950 ;
        RECT 260.400 547.050 261.450 580.950 ;
        RECT 259.950 544.950 262.050 547.050 ;
        RECT 263.400 534.450 264.450 601.950 ;
        RECT 269.400 583.050 270.450 670.950 ;
        RECT 271.950 667.950 274.050 670.050 ;
        RECT 275.250 668.850 276.750 669.750 ;
        RECT 277.950 667.950 280.050 670.050 ;
        RECT 281.250 668.850 283.050 669.750 ;
        RECT 278.400 667.050 279.450 667.950 ;
        RECT 271.950 665.850 274.050 666.750 ;
        RECT 277.950 664.950 280.050 667.050 ;
        RECT 284.400 649.050 285.450 730.950 ;
        RECT 340.950 706.950 343.050 709.050 ;
        RECT 343.950 706.950 346.050 709.050 ;
        RECT 295.950 703.950 298.050 706.050 ;
        RECT 310.950 703.950 313.050 706.050 ;
        RECT 328.950 703.950 331.050 706.050 ;
        RECT 289.950 700.950 292.050 703.050 ;
        RECT 289.950 698.850 292.050 699.750 ;
        RECT 292.950 698.250 295.050 699.150 ;
        RECT 292.950 696.450 295.050 697.050 ;
        RECT 296.400 696.450 297.450 703.950 ;
        RECT 329.400 703.050 330.450 703.950 ;
        RECT 307.950 701.250 310.050 702.150 ;
        RECT 310.950 701.850 313.050 702.750 ;
        RECT 316.950 701.250 319.050 702.150 ;
        RECT 328.950 700.950 331.050 703.050 ;
        RECT 307.950 697.950 310.050 700.050 ;
        RECT 316.950 697.950 319.050 700.050 ;
        RECT 319.950 697.950 322.050 700.050 ;
        RECT 325.950 698.250 328.050 699.150 ;
        RECT 328.950 698.850 331.050 699.750 ;
        RECT 292.950 695.400 297.450 696.450 ;
        RECT 292.950 694.950 295.050 695.400 ;
        RECT 308.400 694.050 309.450 697.950 ;
        RECT 317.400 697.050 318.450 697.950 ;
        RECT 316.950 694.950 319.050 697.050 ;
        RECT 307.950 691.950 310.050 694.050 ;
        RECT 286.950 682.950 289.050 685.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 280.950 635.250 283.050 636.150 ;
        RECT 287.400 634.050 288.450 682.950 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 292.950 668.250 294.750 669.150 ;
        RECT 295.950 667.950 298.050 670.050 ;
        RECT 299.250 668.250 301.050 669.150 ;
        RECT 296.250 665.850 297.750 666.750 ;
        RECT 298.950 664.950 301.050 667.050 ;
        RECT 299.400 664.050 300.450 664.950 ;
        RECT 298.950 661.950 301.050 664.050 ;
        RECT 299.400 660.450 300.450 661.950 ;
        RECT 296.400 659.400 300.450 660.450 ;
        RECT 277.950 632.250 279.750 633.150 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 284.250 632.250 285.750 633.150 ;
        RECT 286.950 631.950 289.050 634.050 ;
        RECT 277.950 628.950 280.050 631.050 ;
        RECT 278.400 625.050 279.450 628.950 ;
        RECT 281.400 628.050 282.450 631.950 ;
        RECT 283.950 628.950 286.050 631.050 ;
        RECT 287.250 629.850 289.050 630.750 ;
        RECT 280.950 625.950 283.050 628.050 ;
        RECT 277.950 622.950 280.050 625.050 ;
        RECT 292.950 622.950 295.050 625.050 ;
        RECT 277.950 598.950 280.050 601.050 ;
        RECT 268.950 580.950 271.050 583.050 ;
        RECT 268.950 563.250 271.050 564.150 ;
        RECT 265.950 560.250 267.750 561.150 ;
        RECT 268.950 559.950 271.050 562.050 ;
        RECT 272.250 560.250 273.750 561.150 ;
        RECT 274.950 559.950 277.050 562.050 ;
        RECT 269.400 559.050 270.450 559.950 ;
        RECT 265.950 556.950 268.050 559.050 ;
        RECT 268.950 556.950 271.050 559.050 ;
        RECT 271.950 556.950 274.050 559.050 ;
        RECT 275.250 557.850 277.050 558.750 ;
        RECT 266.400 553.050 267.450 556.950 ;
        RECT 265.950 550.950 268.050 553.050 ;
        RECT 263.400 533.400 267.450 534.450 ;
        RECT 262.950 529.950 265.050 532.050 ;
        RECT 253.950 526.950 256.050 529.050 ;
        RECT 259.950 527.250 262.050 528.150 ;
        RECT 262.950 527.850 265.050 528.750 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 266.400 523.050 267.450 533.400 ;
        RECT 269.400 526.050 270.450 556.950 ;
        RECT 278.400 550.050 279.450 598.950 ;
        RECT 280.950 596.250 282.750 597.150 ;
        RECT 283.950 595.950 286.050 598.050 ;
        RECT 287.250 596.250 289.050 597.150 ;
        RECT 280.950 592.950 283.050 595.050 ;
        RECT 284.250 593.850 285.750 594.750 ;
        RECT 280.950 565.950 283.050 568.050 ;
        RECT 281.400 559.050 282.450 565.950 ;
        RECT 293.400 565.050 294.450 622.950 ;
        RECT 296.400 595.050 297.450 659.400 ;
        RECT 302.400 631.050 303.450 679.950 ;
        RECT 310.950 677.400 313.050 679.500 ;
        RECT 311.400 660.600 312.600 677.400 ;
        RECT 316.950 670.950 319.050 673.050 ;
        RECT 320.400 672.450 321.450 697.950 ;
        RECT 325.950 694.950 328.050 697.050 ;
        RECT 326.400 694.050 327.450 694.950 ;
        RECT 325.950 691.950 328.050 694.050 ;
        RECT 331.950 677.400 334.050 679.500 ;
        RECT 322.950 672.450 325.050 673.050 ;
        RECT 320.400 671.400 325.050 672.450 ;
        RECT 316.950 668.850 319.050 669.750 ;
        RECT 310.950 658.500 313.050 660.600 ;
        RECT 313.950 639.300 316.050 641.400 ;
        RECT 314.550 635.700 315.750 639.300 ;
        RECT 313.950 633.600 316.050 635.700 ;
        RECT 301.950 630.450 304.050 631.050 ;
        RECT 299.400 629.400 304.050 630.450 ;
        RECT 299.400 604.050 300.450 629.400 ;
        RECT 301.950 628.950 304.050 629.400 ;
        RECT 301.950 626.850 304.050 627.750 ;
        RECT 310.950 627.450 313.050 628.050 ;
        RECT 304.950 626.250 307.050 627.150 ;
        RECT 308.400 626.400 313.050 627.450 ;
        RECT 308.400 625.050 309.450 626.400 ;
        RECT 310.950 625.950 313.050 626.400 ;
        RECT 304.950 622.950 307.050 625.050 ;
        RECT 307.950 622.950 310.050 625.050 ;
        RECT 310.950 623.850 313.050 624.750 ;
        RECT 314.550 621.600 315.750 633.600 ;
        RECT 320.400 627.450 321.450 671.400 ;
        RECT 322.950 670.950 325.050 671.400 ;
        RECT 322.950 668.850 325.050 669.750 ;
        RECT 332.250 665.400 333.450 677.400 ;
        RECT 334.950 674.250 337.050 675.150 ;
        RECT 337.950 673.950 340.050 676.050 ;
        RECT 334.950 672.450 337.050 673.050 ;
        RECT 338.400 672.450 339.450 673.950 ;
        RECT 334.950 671.400 339.450 672.450 ;
        RECT 334.950 670.950 337.050 671.400 ;
        RECT 331.950 663.300 334.050 665.400 ;
        RECT 332.250 659.700 333.450 663.300 ;
        RECT 331.950 657.600 334.050 659.700 ;
        RECT 334.950 638.400 337.050 640.500 ;
        RECT 322.950 629.250 325.050 630.150 ;
        RECT 328.950 629.250 331.050 630.150 ;
        RECT 322.950 627.450 325.050 628.050 ;
        RECT 320.400 626.400 325.050 627.450 ;
        RECT 322.950 625.950 325.050 626.400 ;
        RECT 328.950 625.950 331.050 628.050 ;
        RECT 313.950 619.500 316.050 621.600 ;
        RECT 323.400 613.050 324.450 625.950 ;
        RECT 322.950 610.950 325.050 613.050 ;
        RECT 329.400 610.050 330.450 625.950 ;
        RECT 335.400 621.600 336.600 638.400 ;
        RECT 341.400 625.050 342.450 706.950 ;
        RECT 344.400 700.050 345.450 706.950 ;
        RECT 346.950 704.250 349.050 705.150 ;
        RECT 346.950 700.950 349.050 703.050 ;
        RECT 350.250 701.250 351.750 702.150 ;
        RECT 352.950 700.950 355.050 703.050 ;
        RECT 356.250 701.250 358.050 702.150 ;
        RECT 343.950 697.950 346.050 700.050 ;
        RECT 349.950 697.950 352.050 700.050 ;
        RECT 353.250 698.850 354.750 699.750 ;
        RECT 355.950 697.950 358.050 700.050 ;
        RECT 352.950 694.950 355.050 697.050 ;
        RECT 346.950 691.950 349.050 694.050 ;
        RECT 340.950 622.950 343.050 625.050 ;
        RECT 334.950 619.500 337.050 621.600 ;
        RECT 301.950 607.950 304.050 610.050 ;
        RECT 328.950 607.950 331.050 610.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 299.400 601.050 300.450 601.950 ;
        RECT 302.400 601.050 303.450 607.950 ;
        RECT 322.950 603.450 325.050 604.050 ;
        RECT 322.950 602.400 327.450 603.450 ;
        RECT 322.950 601.950 325.050 602.400 ;
        RECT 298.950 598.950 301.050 601.050 ;
        RECT 301.950 598.950 304.050 601.050 ;
        RECT 305.250 599.250 306.750 600.150 ;
        RECT 307.950 598.950 310.050 601.050 ;
        RECT 319.950 599.250 322.050 600.150 ;
        RECT 322.950 599.850 325.050 600.750 ;
        RECT 298.950 595.950 301.050 598.050 ;
        RECT 302.250 596.850 303.750 597.750 ;
        RECT 304.950 595.950 307.050 598.050 ;
        RECT 308.250 596.850 310.050 597.750 ;
        RECT 319.950 595.950 322.050 598.050 ;
        RECT 305.400 595.050 306.450 595.950 ;
        RECT 295.950 592.950 298.050 595.050 ;
        RECT 298.950 593.850 301.050 594.750 ;
        RECT 304.950 592.950 307.050 595.050 ;
        RECT 322.950 592.950 325.050 595.050 ;
        RECT 295.950 589.950 298.050 592.050 ;
        RECT 289.950 563.250 292.050 564.150 ;
        RECT 292.950 562.950 295.050 565.050 ;
        RECT 296.400 562.050 297.450 589.950 ;
        RECT 304.950 562.950 307.050 565.050 ;
        RECT 286.950 560.250 288.750 561.150 ;
        RECT 289.950 559.950 292.050 562.050 ;
        RECT 293.250 560.250 294.750 561.150 ;
        RECT 295.950 559.950 298.050 562.050 ;
        RECT 301.950 559.950 304.050 562.050 ;
        RECT 280.950 556.950 283.050 559.050 ;
        RECT 286.950 556.950 289.050 559.050 ;
        RECT 277.950 547.950 280.050 550.050 ;
        RECT 277.950 544.950 280.050 547.050 ;
        RECT 278.400 529.050 279.450 544.950 ;
        RECT 271.950 526.950 274.050 529.050 ;
        RECT 275.250 527.250 276.750 528.150 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 280.950 526.950 283.050 529.050 ;
        RECT 281.400 526.050 282.450 526.950 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 271.950 524.850 273.750 525.750 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 278.250 524.850 279.750 525.750 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 265.950 520.950 268.050 523.050 ;
        RECT 280.950 521.850 283.050 522.750 ;
        RECT 253.950 499.950 256.050 502.050 ;
        RECT 254.400 457.050 255.450 499.950 ;
        RECT 259.950 488.250 262.050 489.150 ;
        RECT 266.400 487.050 267.450 520.950 ;
        RECT 287.400 514.050 288.450 556.950 ;
        RECT 290.400 535.050 291.450 559.950 ;
        RECT 292.950 556.950 295.050 559.050 ;
        RECT 296.250 557.850 298.050 558.750 ;
        RECT 292.950 547.950 295.050 550.050 ;
        RECT 289.950 532.950 292.050 535.050 ;
        RECT 286.950 511.950 289.050 514.050 ;
        RECT 287.400 493.050 288.450 511.950 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 281.400 487.050 282.450 490.950 ;
        RECT 286.950 488.250 289.050 489.150 ;
        RECT 259.950 484.950 262.050 487.050 ;
        RECT 263.250 485.250 264.750 486.150 ;
        RECT 265.950 484.950 268.050 487.050 ;
        RECT 269.250 485.250 271.050 486.150 ;
        RECT 277.950 485.250 279.750 486.150 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 284.250 485.250 285.750 486.150 ;
        RECT 286.950 484.950 289.050 487.050 ;
        RECT 262.950 481.950 265.050 484.050 ;
        RECT 266.250 482.850 267.750 483.750 ;
        RECT 268.950 481.950 271.050 484.050 ;
        RECT 277.950 481.950 280.050 484.050 ;
        RECT 281.250 482.850 282.750 483.750 ;
        RECT 283.950 481.950 286.050 484.050 ;
        RECT 263.400 481.050 264.450 481.950 ;
        RECT 262.950 478.950 265.050 481.050 ;
        RECT 262.950 460.950 265.050 463.050 ;
        RECT 263.400 457.050 264.450 460.950 ;
        RECT 253.950 454.950 256.050 457.050 ;
        RECT 257.250 455.250 259.050 456.150 ;
        RECT 262.950 454.950 265.050 457.050 ;
        RECT 266.250 455.250 268.050 456.150 ;
        RECT 253.950 452.850 255.750 453.750 ;
        RECT 256.950 453.450 259.050 454.050 ;
        RECT 256.950 452.400 261.450 453.450 ;
        RECT 262.950 452.850 264.750 453.750 ;
        RECT 265.950 453.450 268.050 454.050 ;
        RECT 269.400 453.450 270.450 481.950 ;
        RECT 271.950 478.950 274.050 481.050 ;
        RECT 278.400 480.450 279.450 481.950 ;
        RECT 278.400 479.400 282.450 480.450 ;
        RECT 256.950 451.950 259.050 452.400 ;
        RECT 253.950 421.950 256.050 424.050 ;
        RECT 247.950 416.250 250.050 417.150 ;
        RECT 250.950 415.950 253.050 418.050 ;
        RECT 254.400 415.050 255.450 421.950 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 251.250 413.250 252.750 414.150 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 257.250 413.250 259.050 414.150 ;
        RECT 250.950 409.950 253.050 412.050 ;
        RECT 254.250 410.850 255.750 411.750 ;
        RECT 256.950 409.950 259.050 412.050 ;
        RECT 257.400 409.050 258.450 409.950 ;
        RECT 256.950 406.950 259.050 409.050 ;
        RECT 253.950 385.950 256.050 388.050 ;
        RECT 254.400 382.050 255.450 385.950 ;
        RECT 250.950 380.250 252.750 381.150 ;
        RECT 253.950 379.950 256.050 382.050 ;
        RECT 257.250 380.250 259.050 381.150 ;
        RECT 250.950 376.950 253.050 379.050 ;
        RECT 254.250 377.850 255.750 378.750 ;
        RECT 256.950 376.950 259.050 379.050 ;
        RECT 251.400 373.050 252.450 376.950 ;
        RECT 260.400 375.450 261.450 452.400 ;
        RECT 265.950 452.400 270.450 453.450 ;
        RECT 265.950 451.950 268.050 452.400 ;
        RECT 272.400 421.050 273.450 478.950 ;
        RECT 281.400 457.050 282.450 479.400 ;
        RECT 284.400 460.050 285.450 481.950 ;
        RECT 283.950 457.950 286.050 460.050 ;
        RECT 280.950 454.950 283.050 457.050 ;
        RECT 283.950 454.950 286.050 457.050 ;
        RECT 274.950 452.850 277.050 453.750 ;
        RECT 280.950 452.850 283.050 453.750 ;
        RECT 280.950 442.950 283.050 445.050 ;
        RECT 268.950 419.250 271.050 420.150 ;
        RECT 271.950 418.950 274.050 421.050 ;
        RECT 262.950 415.950 265.050 418.050 ;
        RECT 265.950 416.250 267.750 417.150 ;
        RECT 268.950 415.950 271.050 418.050 ;
        RECT 272.250 416.250 273.750 417.150 ;
        RECT 274.950 415.950 277.050 418.050 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 263.400 409.050 264.450 415.950 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 275.250 413.850 277.050 414.750 ;
        RECT 266.400 412.050 267.450 412.950 ;
        RECT 265.950 409.950 268.050 412.050 ;
        RECT 262.950 406.950 265.050 409.050 ;
        RECT 262.950 382.950 265.050 385.050 ;
        RECT 263.400 379.050 264.450 382.950 ;
        RECT 266.400 379.050 267.450 409.950 ;
        RECT 269.400 406.050 270.450 412.950 ;
        RECT 268.950 403.950 271.050 406.050 ;
        RECT 272.400 403.050 273.450 412.950 ;
        RECT 278.400 409.050 279.450 415.950 ;
        RECT 281.400 412.050 282.450 442.950 ;
        RECT 280.950 409.950 283.050 412.050 ;
        RECT 277.950 406.950 280.050 409.050 ;
        RECT 271.950 400.950 274.050 403.050 ;
        RECT 274.950 388.950 277.050 391.050 ;
        RECT 268.950 383.250 270.750 384.150 ;
        RECT 271.950 382.950 274.050 385.050 ;
        RECT 268.950 379.950 271.050 382.050 ;
        RECT 272.250 380.850 274.050 381.750 ;
        RECT 275.400 381.450 276.450 388.950 ;
        RECT 277.950 383.250 279.750 384.150 ;
        RECT 280.950 382.950 283.050 385.050 ;
        RECT 277.950 381.450 280.050 382.050 ;
        RECT 275.400 380.400 280.050 381.450 ;
        RECT 281.250 380.850 283.050 381.750 ;
        RECT 277.950 379.950 280.050 380.400 ;
        RECT 262.950 376.950 265.050 379.050 ;
        RECT 265.950 376.950 268.050 379.050 ;
        RECT 257.400 374.400 261.450 375.450 ;
        RECT 250.950 370.950 253.050 373.050 ;
        RECT 250.950 343.950 253.050 346.050 ;
        RECT 247.950 341.250 250.050 342.150 ;
        RECT 247.950 339.450 250.050 340.050 ;
        RECT 251.400 339.450 252.450 343.950 ;
        RECT 247.950 338.400 252.450 339.450 ;
        RECT 247.950 337.950 250.050 338.400 ;
        RECT 257.400 325.050 258.450 374.400 ;
        RECT 269.400 364.050 270.450 379.950 ;
        RECT 277.950 376.950 280.050 379.050 ;
        RECT 268.950 361.950 271.050 364.050 ;
        RECT 259.950 346.950 262.050 349.050 ;
        RECT 260.400 346.050 261.450 346.950 ;
        RECT 259.950 343.950 262.050 346.050 ;
        RECT 265.950 345.450 268.050 346.050 ;
        RECT 263.250 344.250 264.750 345.150 ;
        RECT 265.950 344.400 270.450 345.450 ;
        RECT 265.950 343.950 268.050 344.400 ;
        RECT 259.950 341.850 261.750 342.750 ;
        RECT 262.950 340.950 265.050 343.050 ;
        RECT 266.250 341.850 268.050 342.750 ;
        RECT 269.400 334.050 270.450 344.400 ;
        RECT 278.400 339.450 279.450 376.950 ;
        RECT 280.950 341.250 283.050 342.150 ;
        RECT 280.950 339.450 283.050 340.050 ;
        RECT 278.400 338.400 283.050 339.450 ;
        RECT 280.950 337.950 283.050 338.400 ;
        RECT 268.950 331.950 271.050 334.050 ;
        RECT 277.950 331.950 280.050 334.050 ;
        RECT 256.950 322.950 259.050 325.050 ;
        RECT 244.950 319.950 247.050 322.050 ;
        RECT 257.400 313.050 258.450 322.950 ;
        RECT 265.950 319.950 268.050 322.050 ;
        RECT 262.950 313.950 265.050 316.050 ;
        RECT 244.950 311.250 246.750 312.150 ;
        RECT 247.950 310.950 250.050 313.050 ;
        RECT 253.950 311.250 255.750 312.150 ;
        RECT 256.950 310.950 259.050 313.050 ;
        RECT 244.950 307.950 247.050 310.050 ;
        RECT 248.250 308.850 250.050 309.750 ;
        RECT 253.950 307.950 256.050 310.050 ;
        RECT 257.250 308.850 259.050 309.750 ;
        RECT 245.400 301.050 246.450 307.950 ;
        RECT 244.950 298.950 247.050 301.050 ;
        RECT 250.950 298.950 253.050 301.050 ;
        RECT 235.950 295.950 238.050 298.050 ;
        RECT 241.950 295.950 244.050 298.050 ;
        RECT 236.400 268.050 237.450 295.950 ;
        RECT 244.950 274.950 247.050 277.050 ;
        RECT 238.950 272.250 241.050 273.150 ;
        RECT 245.400 271.050 246.450 274.950 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 242.250 269.250 243.750 270.150 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 248.250 269.250 250.050 270.150 ;
        RECT 220.950 265.950 223.050 268.050 ;
        RECT 226.950 265.950 229.050 268.050 ;
        RECT 232.950 265.950 235.050 268.050 ;
        RECT 235.950 265.950 238.050 268.050 ;
        RECT 238.950 265.950 241.050 268.050 ;
        RECT 241.950 265.950 244.050 268.050 ;
        RECT 245.250 266.850 246.750 267.750 ;
        RECT 247.950 267.450 250.050 268.050 ;
        RECT 251.400 267.450 252.450 298.950 ;
        RECT 247.950 266.400 252.450 267.450 ;
        RECT 247.950 265.950 250.050 266.400 ;
        RECT 217.950 262.950 220.050 265.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 202.950 253.950 205.050 256.050 ;
        RECT 203.400 253.050 204.450 253.950 ;
        RECT 202.950 250.950 205.050 253.050 ;
        RECT 193.950 236.400 198.450 237.450 ;
        RECT 193.950 235.950 196.050 236.400 ;
        RECT 188.400 232.050 189.450 235.950 ;
        RECT 197.400 235.050 198.450 236.400 ;
        RECT 196.950 232.950 199.050 235.050 ;
        RECT 203.400 234.450 204.450 250.950 ;
        RECT 217.950 244.950 220.050 247.050 ;
        RECT 205.950 236.250 207.750 237.150 ;
        RECT 208.950 235.950 211.050 238.050 ;
        RECT 212.250 236.250 214.050 237.150 ;
        RECT 214.950 235.950 217.050 238.050 ;
        RECT 205.950 234.450 208.050 235.050 ;
        RECT 203.400 233.400 208.050 234.450 ;
        RECT 209.250 233.850 210.750 234.750 ;
        RECT 205.950 232.950 208.050 233.400 ;
        RECT 211.950 232.950 214.050 235.050 ;
        RECT 187.950 229.950 190.050 232.050 ;
        RECT 196.950 229.950 199.050 232.050 ;
        RECT 181.950 199.950 184.050 202.050 ;
        RECT 184.950 200.250 187.050 201.150 ;
        RECT 187.950 199.950 190.050 202.050 ;
        RECT 157.950 196.950 160.050 199.050 ;
        RECT 161.250 197.250 162.750 198.150 ;
        RECT 163.950 196.950 166.050 199.050 ;
        RECT 167.250 197.250 169.050 198.150 ;
        RECT 169.950 196.950 172.050 199.050 ;
        RECT 175.950 197.250 177.750 198.150 ;
        RECT 178.950 196.950 181.050 199.050 ;
        RECT 182.250 197.250 183.750 198.150 ;
        RECT 184.950 196.950 187.050 199.050 ;
        RECT 158.400 196.050 159.450 196.950 ;
        RECT 185.400 196.050 186.450 196.950 ;
        RECT 157.950 193.950 160.050 196.050 ;
        RECT 160.950 193.950 163.050 196.050 ;
        RECT 164.250 194.850 165.750 195.750 ;
        RECT 166.950 193.950 169.050 196.050 ;
        RECT 175.950 193.950 178.050 196.050 ;
        RECT 179.250 194.850 180.750 195.750 ;
        RECT 181.950 193.950 184.050 196.050 ;
        RECT 184.950 193.950 187.050 196.050 ;
        RECT 154.950 187.950 157.050 190.050 ;
        RECT 158.400 178.050 159.450 193.950 ;
        RECT 157.950 175.950 160.050 178.050 ;
        RECT 127.950 173.400 130.050 175.500 ;
        RECT 112.950 169.950 115.050 172.050 ;
        RECT 112.950 167.850 115.050 168.750 ;
        RECT 115.950 167.250 118.050 168.150 ;
        RECT 109.950 163.950 112.050 166.050 ;
        RECT 115.950 163.950 118.050 166.050 ;
        RECT 116.400 163.050 117.450 163.950 ;
        RECT 115.950 160.950 118.050 163.050 ;
        RECT 107.400 140.400 111.450 141.450 ;
        RECT 106.950 135.300 109.050 137.400 ;
        RECT 107.250 131.700 108.450 135.300 ;
        RECT 106.950 129.600 109.050 131.700 ;
        RECT 91.950 125.250 94.050 126.150 ;
        RECT 94.950 124.950 97.050 127.050 ;
        RECT 97.950 125.250 100.050 126.150 ;
        RECT 88.950 121.950 91.050 124.050 ;
        RECT 91.950 123.450 94.050 124.050 ;
        RECT 95.400 123.450 96.450 124.950 ;
        RECT 91.950 122.400 96.450 123.450 ;
        RECT 91.950 121.950 94.050 122.400 ;
        RECT 97.950 121.950 100.050 124.050 ;
        RECT 89.400 121.050 90.450 121.950 ;
        RECT 88.950 118.950 91.050 121.050 ;
        RECT 107.250 117.600 108.450 129.600 ;
        RECT 110.400 124.050 111.450 140.400 ;
        RECT 116.400 126.450 117.450 160.950 ;
        RECT 128.400 156.600 129.600 173.400 ;
        RECT 139.950 172.950 142.050 175.050 ;
        RECT 148.950 173.400 151.050 175.500 ;
        RECT 140.400 169.050 141.450 172.950 ;
        RECT 133.950 166.950 136.050 169.050 ;
        RECT 139.950 166.950 142.050 169.050 ;
        RECT 133.950 164.850 136.050 165.750 ;
        RECT 139.950 164.850 142.050 165.750 ;
        RECT 149.250 161.400 150.450 173.400 ;
        RECT 151.950 170.250 154.050 171.150 ;
        RECT 151.950 166.950 154.050 169.050 ;
        RECT 161.400 168.450 162.450 193.950 ;
        RECT 167.400 190.050 168.450 193.950 ;
        RECT 176.400 190.050 177.450 193.950 ;
        RECT 166.950 187.950 169.050 190.050 ;
        RECT 175.950 187.950 178.050 190.050 ;
        RECT 158.400 167.400 162.450 168.450 ;
        RECT 148.950 159.300 151.050 161.400 ;
        RECT 152.400 160.050 153.450 166.950 ;
        RECT 127.950 154.500 130.050 156.600 ;
        RECT 149.250 155.700 150.450 159.300 ;
        RECT 151.950 157.950 154.050 160.050 ;
        RECT 124.950 151.950 127.050 154.050 ;
        RECT 148.950 153.600 151.050 155.700 ;
        RECT 125.400 130.050 126.450 151.950 ;
        RECT 124.950 127.950 127.050 130.050 ;
        RECT 130.950 128.250 133.050 129.150 ;
        RECT 149.250 128.250 150.750 129.150 ;
        RECT 151.950 127.950 154.050 130.050 ;
        RECT 125.400 127.050 126.450 127.950 ;
        RECT 116.400 125.400 120.450 126.450 ;
        RECT 109.950 121.950 112.050 124.050 ;
        RECT 115.950 121.950 118.050 124.050 ;
        RECT 119.400 123.450 120.450 125.400 ;
        RECT 121.950 125.250 123.750 126.150 ;
        RECT 124.950 124.950 127.050 127.050 ;
        RECT 128.250 125.250 129.750 126.150 ;
        RECT 130.950 124.950 133.050 127.050 ;
        RECT 145.950 125.850 147.750 126.750 ;
        RECT 148.950 124.950 151.050 127.050 ;
        RECT 152.250 125.850 154.050 126.750 ;
        RECT 121.950 123.450 124.050 124.050 ;
        RECT 119.400 122.400 124.050 123.450 ;
        RECT 125.250 122.850 126.750 123.750 ;
        RECT 121.950 121.950 124.050 122.400 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 109.950 119.850 112.050 120.750 ;
        RECT 85.950 115.500 88.050 117.600 ;
        RECT 106.950 115.500 109.050 117.600 ;
        RECT 97.950 103.950 100.050 106.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 92.400 97.050 93.450 100.950 ;
        RECT 98.400 97.050 99.450 103.950 ;
        RECT 73.950 94.950 76.050 97.050 ;
        RECT 91.950 94.950 94.050 97.050 ;
        RECT 97.950 94.950 100.050 97.050 ;
        RECT 70.950 92.250 72.750 93.150 ;
        RECT 73.950 91.950 76.050 94.050 ;
        RECT 77.250 92.250 79.050 93.150 ;
        RECT 79.950 91.950 82.050 94.050 ;
        RECT 91.950 92.850 94.050 93.750 ;
        RECT 97.950 92.850 100.050 93.750 ;
        RECT 106.950 92.250 108.750 93.150 ;
        RECT 109.950 91.950 112.050 94.050 ;
        RECT 113.250 92.250 115.050 93.150 ;
        RECT 70.950 90.450 73.050 91.050 ;
        RECT 68.400 89.400 73.050 90.450 ;
        RECT 74.250 89.850 75.750 90.750 ;
        RECT 70.950 88.950 73.050 89.400 ;
        RECT 76.950 88.950 79.050 91.050 ;
        RECT 80.400 85.050 81.450 91.950 ;
        RECT 106.950 88.950 109.050 91.050 ;
        RECT 110.250 89.850 111.750 90.750 ;
        RECT 112.950 88.950 115.050 91.050 ;
        RECT 37.950 82.950 40.050 85.050 ;
        RECT 49.950 82.950 52.050 85.050 ;
        RECT 79.950 82.950 82.050 85.050 ;
        RECT 61.950 58.950 64.050 61.050 ;
        RECT 67.950 59.250 70.050 60.150 ;
        RECT 46.950 53.250 49.050 54.150 ;
        RECT 52.950 52.950 55.050 55.050 ;
        RECT 62.400 54.450 63.450 58.950 ;
        RECT 107.400 58.050 108.450 88.950 ;
        RECT 109.950 61.950 112.050 64.050 ;
        RECT 64.950 56.250 66.750 57.150 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 73.950 57.450 76.050 58.050 ;
        RECT 71.250 56.250 72.750 57.150 ;
        RECT 73.950 56.400 78.450 57.450 ;
        RECT 73.950 55.950 76.050 56.400 ;
        RECT 68.400 55.050 69.450 55.950 ;
        RECT 64.950 54.450 67.050 55.050 ;
        RECT 62.400 53.400 67.050 54.450 ;
        RECT 64.950 52.950 67.050 53.400 ;
        RECT 67.950 52.950 70.050 55.050 ;
        RECT 70.950 52.950 73.050 55.050 ;
        RECT 74.250 53.850 76.050 54.750 ;
        RECT 71.400 52.050 72.450 52.950 ;
        RECT 43.950 50.250 45.750 51.150 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 52.950 50.850 55.050 51.750 ;
        RECT 70.950 49.950 73.050 52.050 ;
        RECT 43.950 46.950 46.050 49.050 ;
        RECT 44.400 37.050 45.450 46.950 ;
        RECT 43.950 34.950 46.050 37.050 ;
        RECT 16.950 25.950 19.050 28.050 ;
        RECT 34.950 25.950 37.050 28.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 17.250 23.850 18.750 24.750 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 31.950 23.250 34.050 24.150 ;
        RECT 34.950 23.850 37.050 24.750 ;
        RECT 47.400 22.050 48.450 49.950 ;
        RECT 77.400 49.050 78.450 56.400 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 88.950 52.950 91.050 55.050 ;
        RECT 100.950 53.250 103.050 54.150 ;
        RECT 106.950 53.250 109.050 54.150 ;
        RECT 85.950 50.250 88.050 51.150 ;
        RECT 88.950 50.850 91.050 51.750 ;
        RECT 100.950 49.950 103.050 52.050 ;
        RECT 106.950 51.450 109.050 52.050 ;
        RECT 110.400 51.450 111.450 61.950 ;
        RECT 104.250 50.250 105.750 51.150 ;
        RECT 106.950 50.400 111.450 51.450 ;
        RECT 106.950 49.950 109.050 50.400 ;
        RECT 76.950 46.950 79.050 49.050 ;
        RECT 85.950 46.950 88.050 49.050 ;
        RECT 103.950 46.950 106.050 49.050 ;
        RECT 86.400 37.050 87.450 46.950 ;
        RECT 52.950 34.950 55.050 37.050 ;
        RECT 58.950 34.950 61.050 37.050 ;
        RECT 85.950 34.950 88.050 37.050 ;
        RECT 49.950 31.950 52.050 34.050 ;
        RECT 50.400 22.050 51.450 31.950 ;
        RECT 53.400 25.050 54.450 34.950 ;
        RECT 59.400 25.050 60.450 34.950 ;
        RECT 73.950 31.950 76.050 34.050 ;
        RECT 67.950 28.950 70.050 31.050 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 56.250 23.250 57.750 24.150 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 68.400 22.050 69.450 28.950 ;
        RECT 74.400 28.050 75.450 31.950 ;
        RECT 73.950 25.950 76.050 28.050 ;
        RECT 70.950 23.250 73.050 24.150 ;
        RECT 73.950 23.850 76.050 24.750 ;
        RECT 76.950 23.250 78.750 24.150 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 86.400 22.050 87.450 34.950 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 98.250 23.250 99.750 24.150 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 104.400 24.450 105.450 46.950 ;
        RECT 104.400 23.400 108.450 24.450 ;
        RECT 13.950 20.850 16.050 21.750 ;
        RECT 19.950 20.850 22.050 21.750 ;
        RECT 31.950 19.950 34.050 22.050 ;
        RECT 46.950 19.950 49.050 22.050 ;
        RECT 49.950 19.950 52.050 22.050 ;
        RECT 53.250 20.850 54.750 21.750 ;
        RECT 55.950 19.950 58.050 22.050 ;
        RECT 59.250 20.850 61.050 21.750 ;
        RECT 67.950 21.450 70.050 22.050 ;
        RECT 70.950 21.450 73.050 22.050 ;
        RECT 67.950 20.400 73.050 21.450 ;
        RECT 67.950 19.950 70.050 20.400 ;
        RECT 70.950 19.950 73.050 20.400 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 80.250 20.850 82.050 21.750 ;
        RECT 85.950 19.950 88.050 22.050 ;
        RECT 94.950 20.850 96.750 21.750 ;
        RECT 97.950 19.950 100.050 22.050 ;
        RECT 101.250 20.850 102.750 21.750 ;
        RECT 103.950 19.950 106.050 22.050 ;
        RECT 98.400 19.050 99.450 19.950 ;
        RECT 107.400 19.050 108.450 23.400 ;
        RECT 116.400 22.050 117.450 121.950 ;
        RECT 122.400 109.050 123.450 121.950 ;
        RECT 154.950 112.950 157.050 115.050 ;
        RECT 127.950 109.950 130.050 112.050 ;
        RECT 121.950 106.950 124.050 109.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 119.400 64.050 120.450 100.950 ;
        RECT 121.950 97.950 124.050 100.050 ;
        RECT 122.400 91.050 123.450 97.950 ;
        RECT 128.400 97.050 129.450 109.950 ;
        RECT 142.950 106.950 145.050 109.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 131.400 97.050 132.450 100.950 ;
        RECT 124.950 94.950 127.050 97.050 ;
        RECT 127.950 94.950 130.050 97.050 ;
        RECT 130.950 94.950 133.050 97.050 ;
        RECT 134.250 95.250 135.750 96.150 ;
        RECT 136.950 94.950 139.050 97.050 ;
        RECT 121.950 88.950 124.050 91.050 ;
        RECT 118.950 61.950 121.050 64.050 ;
        RECT 125.400 61.050 126.450 94.950 ;
        RECT 128.400 94.050 129.450 94.950 ;
        RECT 127.950 91.950 130.050 94.050 ;
        RECT 131.250 92.850 132.750 93.750 ;
        RECT 133.950 91.950 136.050 94.050 ;
        RECT 137.250 92.850 139.050 93.750 ;
        RECT 127.950 89.850 130.050 90.750 ;
        RECT 130.950 88.950 133.050 91.050 ;
        RECT 118.950 58.950 121.050 61.050 ;
        RECT 124.950 58.950 127.050 61.050 ;
        RECT 119.400 34.050 120.450 58.950 ;
        RECT 124.950 56.250 127.050 57.150 ;
        RECT 131.400 55.050 132.450 88.950 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 124.950 52.950 127.050 55.050 ;
        RECT 128.250 53.250 129.750 54.150 ;
        RECT 130.950 52.950 133.050 55.050 ;
        RECT 134.250 53.250 136.050 54.150 ;
        RECT 127.950 49.950 130.050 52.050 ;
        RECT 131.250 50.850 132.750 51.750 ;
        RECT 133.950 49.950 136.050 52.050 ;
        RECT 121.950 34.950 124.050 37.050 ;
        RECT 118.950 31.950 121.050 34.050 ;
        RECT 119.400 22.050 120.450 31.950 ;
        RECT 115.950 19.950 118.050 22.050 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 122.400 19.050 123.450 34.950 ;
        RECT 128.400 34.050 129.450 49.950 ;
        RECT 140.400 49.050 141.450 55.950 ;
        RECT 139.950 46.950 142.050 49.050 ;
        RECT 127.950 31.950 130.050 34.050 ;
        RECT 124.950 28.950 127.050 31.050 ;
        RECT 125.400 22.050 126.450 28.950 ;
        RECT 136.950 25.950 139.050 28.050 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 128.250 20.250 130.050 21.150 ;
        RECT 137.400 19.050 138.450 25.950 ;
        RECT 143.400 25.050 144.450 106.950 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 149.400 97.050 150.450 100.950 ;
        RECT 151.950 97.950 154.050 100.050 ;
        RECT 155.400 97.050 156.450 112.950 ;
        RECT 148.950 94.950 151.050 97.050 ;
        RECT 152.250 95.850 153.750 96.750 ;
        RECT 154.950 94.950 157.050 97.050 ;
        RECT 148.950 92.850 151.050 93.750 ;
        RECT 154.950 92.850 157.050 93.750 ;
        RECT 158.400 78.450 159.450 167.400 ;
        RECT 169.950 166.950 172.050 169.050 ;
        RECT 175.950 168.450 178.050 169.050 ;
        RECT 173.250 167.250 174.750 168.150 ;
        RECT 175.950 167.400 180.450 168.450 ;
        RECT 175.950 166.950 178.050 167.400 ;
        RECT 160.950 163.950 163.050 166.050 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 170.250 164.850 171.750 165.750 ;
        RECT 172.950 163.950 175.050 166.050 ;
        RECT 176.250 164.850 178.050 165.750 ;
        RECT 161.400 127.050 162.450 163.950 ;
        RECT 166.950 161.850 169.050 162.750 ;
        RECT 173.400 154.050 174.450 163.950 ;
        RECT 169.950 151.950 172.050 154.050 ;
        RECT 172.950 151.950 175.050 154.050 ;
        RECT 170.400 130.050 171.450 151.950 ;
        RECT 179.400 133.050 180.450 167.400 ;
        RECT 178.950 130.950 181.050 133.050 ;
        RECT 167.250 128.250 168.750 129.150 ;
        RECT 169.950 127.950 172.050 130.050 ;
        RECT 179.400 127.050 180.450 130.950 ;
        RECT 160.950 124.950 163.050 127.050 ;
        RECT 163.950 125.850 165.750 126.750 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 170.250 125.850 172.050 126.750 ;
        RECT 178.950 124.950 181.050 127.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 173.400 100.050 174.450 100.950 ;
        RECT 182.400 100.050 183.450 193.950 ;
        RECT 188.400 130.050 189.450 199.950 ;
        RECT 197.400 192.450 198.450 229.950 ;
        RECT 212.400 229.050 213.450 232.950 ;
        RECT 211.950 226.950 214.050 229.050 ;
        RECT 211.950 223.950 214.050 226.050 ;
        RECT 202.950 196.950 205.050 199.050 ;
        RECT 199.950 194.250 202.050 195.150 ;
        RECT 202.950 194.850 205.050 195.750 ;
        RECT 199.950 192.450 202.050 193.050 ;
        RECT 197.400 191.400 202.050 192.450 ;
        RECT 199.950 190.950 202.050 191.400 ;
        RECT 212.400 169.050 213.450 223.950 ;
        RECT 215.400 202.050 216.450 235.950 ;
        RECT 214.950 199.950 217.050 202.050 ;
        RECT 218.400 199.050 219.450 244.950 ;
        RECT 221.400 244.050 222.450 265.950 ;
        RECT 220.950 241.950 223.050 244.050 ;
        RECT 235.950 241.950 238.050 244.050 ;
        RECT 236.400 241.050 237.450 241.950 ;
        RECT 223.950 238.950 226.050 241.050 ;
        RECT 229.950 238.950 232.050 241.050 ;
        RECT 233.250 239.250 234.750 240.150 ;
        RECT 235.950 238.950 238.050 241.050 ;
        RECT 224.400 208.050 225.450 238.950 ;
        RECT 239.400 238.050 240.450 265.950 ;
        RECT 242.400 238.050 243.450 265.950 ;
        RECT 254.400 265.050 255.450 307.950 ;
        RECT 256.950 304.950 259.050 307.050 ;
        RECT 257.400 292.050 258.450 304.950 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 253.950 262.950 256.050 265.050 ;
        RECT 244.950 244.950 247.050 247.050 ;
        RECT 245.400 241.050 246.450 244.950 ;
        RECT 244.950 238.950 247.050 241.050 ;
        RECT 248.250 239.250 249.750 240.150 ;
        RECT 250.950 238.950 253.050 241.050 ;
        RECT 226.950 235.950 229.050 238.050 ;
        RECT 230.250 236.850 231.750 237.750 ;
        RECT 232.950 235.950 235.050 238.050 ;
        RECT 236.250 236.850 238.050 237.750 ;
        RECT 238.950 235.950 241.050 238.050 ;
        RECT 241.950 235.950 244.050 238.050 ;
        RECT 244.950 236.850 246.750 237.750 ;
        RECT 247.950 235.950 250.050 238.050 ;
        RECT 251.250 236.850 252.750 237.750 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 226.950 233.850 229.050 234.750 ;
        RECT 253.950 233.850 256.050 234.750 ;
        RECT 235.950 226.950 238.050 229.050 ;
        RECT 223.950 205.950 226.050 208.050 ;
        RECT 223.950 200.250 226.050 201.150 ;
        RECT 214.950 197.250 216.750 198.150 ;
        RECT 217.950 196.950 220.050 199.050 ;
        RECT 221.250 197.250 222.750 198.150 ;
        RECT 223.950 196.950 226.050 199.050 ;
        RECT 214.950 193.950 217.050 196.050 ;
        RECT 218.250 194.850 219.750 195.750 ;
        RECT 220.950 193.950 223.050 196.050 ;
        RECT 236.400 195.450 237.450 226.950 ;
        RECT 257.400 226.050 258.450 289.950 ;
        RECT 259.950 269.250 262.050 270.150 ;
        RECT 259.950 265.950 262.050 268.050 ;
        RECT 260.400 247.050 261.450 265.950 ;
        RECT 263.400 259.050 264.450 313.950 ;
        RECT 266.400 277.050 267.450 319.950 ;
        RECT 278.400 313.050 279.450 331.950 ;
        RECT 271.950 310.950 274.050 313.050 ;
        RECT 275.250 311.250 276.750 312.150 ;
        RECT 277.950 310.950 280.050 313.050 ;
        RECT 271.950 308.850 273.750 309.750 ;
        RECT 274.950 307.950 277.050 310.050 ;
        RECT 278.250 308.850 279.750 309.750 ;
        RECT 280.950 307.950 283.050 310.050 ;
        RECT 275.400 307.050 276.450 307.950 ;
        RECT 274.950 304.950 277.050 307.050 ;
        RECT 277.950 304.950 280.050 307.050 ;
        RECT 280.950 305.850 283.050 306.750 ;
        RECT 265.950 274.950 268.050 277.050 ;
        RECT 278.400 274.050 279.450 304.950 ;
        RECT 277.950 271.950 280.050 274.050 ;
        RECT 274.950 270.450 277.050 271.050 ;
        RECT 265.950 269.250 268.050 270.150 ;
        RECT 274.950 269.400 279.450 270.450 ;
        RECT 274.950 268.950 277.050 269.400 ;
        RECT 265.950 265.950 268.050 268.050 ;
        RECT 274.950 266.850 277.050 267.750 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 266.400 262.050 267.450 262.950 ;
        RECT 265.950 259.950 268.050 262.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 259.950 244.950 262.050 247.050 ;
        RECT 260.400 229.050 261.450 244.950 ;
        RECT 259.950 226.950 262.050 229.050 ;
        RECT 256.950 223.950 259.050 226.050 ;
        RECT 241.950 208.950 244.050 211.050 ;
        RECT 242.400 199.050 243.450 208.950 ;
        RECT 260.400 202.050 261.450 226.950 ;
        RECT 266.400 202.050 267.450 259.950 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 271.950 244.950 274.050 247.050 ;
        RECT 272.400 244.050 273.450 244.950 ;
        RECT 271.950 241.950 274.050 244.050 ;
        RECT 268.950 239.250 271.050 240.150 ;
        RECT 271.950 239.850 274.050 240.750 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 247.950 200.250 250.050 201.150 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 263.250 200.250 264.750 201.150 ;
        RECT 265.950 199.950 268.050 202.050 ;
        RECT 238.950 197.250 240.750 198.150 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 245.250 197.250 246.750 198.150 ;
        RECT 247.950 196.950 250.050 199.050 ;
        RECT 259.950 197.850 261.750 198.750 ;
        RECT 262.950 196.950 265.050 199.050 ;
        RECT 266.250 197.850 268.050 198.750 ;
        RECT 238.950 195.450 241.050 196.050 ;
        RECT 236.400 194.400 241.050 195.450 ;
        RECT 242.250 194.850 243.750 195.750 ;
        RECT 215.400 193.050 216.450 193.950 ;
        RECT 214.950 190.950 217.050 193.050 ;
        RECT 199.950 166.950 202.050 169.050 ;
        RECT 211.950 166.950 214.050 169.050 ;
        RECT 215.250 167.250 216.750 168.150 ;
        RECT 217.950 166.950 220.050 169.050 ;
        RECT 190.950 164.250 192.750 165.150 ;
        RECT 193.950 163.950 196.050 166.050 ;
        RECT 197.250 164.250 199.050 165.150 ;
        RECT 190.950 160.950 193.050 163.050 ;
        RECT 194.250 161.850 195.750 162.750 ;
        RECT 196.950 162.450 199.050 163.050 ;
        RECT 200.400 162.450 201.450 166.950 ;
        RECT 208.950 163.950 211.050 166.050 ;
        RECT 212.250 164.850 213.750 165.750 ;
        RECT 214.950 163.950 217.050 166.050 ;
        RECT 218.250 164.850 220.050 165.750 ;
        RECT 215.400 163.050 216.450 163.950 ;
        RECT 196.950 161.400 201.450 162.450 ;
        RECT 208.950 161.850 211.050 162.750 ;
        RECT 196.950 160.950 199.050 161.400 ;
        RECT 214.950 160.950 217.050 163.050 ;
        RECT 217.950 160.950 220.050 163.050 ;
        RECT 215.400 160.050 216.450 160.950 ;
        RECT 214.950 157.950 217.050 160.050 ;
        RECT 187.950 127.950 190.050 130.050 ;
        RECT 193.950 127.950 196.050 130.050 ;
        RECT 187.950 124.950 190.050 127.050 ;
        RECT 190.950 124.950 193.050 127.050 ;
        RECT 184.950 122.250 187.050 123.150 ;
        RECT 187.950 122.850 190.050 123.750 ;
        RECT 184.950 118.950 187.050 121.050 ;
        RECT 185.400 118.050 186.450 118.950 ;
        RECT 184.950 115.950 187.050 118.050 ;
        RECT 191.400 109.050 192.450 124.950 ;
        RECT 190.950 106.950 193.050 109.050 ;
        RECT 172.950 97.950 175.050 100.050 ;
        RECT 181.950 97.950 184.050 100.050 ;
        RECT 169.950 95.250 172.050 96.150 ;
        RECT 172.950 95.850 175.050 96.750 ;
        RECT 187.950 94.950 190.050 97.050 ;
        RECT 188.400 94.050 189.450 94.950 ;
        RECT 169.950 91.950 172.050 94.050 ;
        RECT 184.950 92.250 186.750 93.150 ;
        RECT 187.950 91.950 190.050 94.050 ;
        RECT 170.400 91.050 171.450 91.950 ;
        RECT 191.400 91.050 192.450 106.950 ;
        RECT 194.400 94.050 195.450 127.950 ;
        RECT 199.950 126.450 202.050 127.050 ;
        RECT 197.400 125.400 202.050 126.450 ;
        RECT 197.400 115.050 198.450 125.400 ;
        RECT 199.950 124.950 202.050 125.400 ;
        RECT 205.950 124.950 208.050 127.050 ;
        RECT 209.250 125.250 211.050 126.150 ;
        RECT 199.950 122.850 202.050 123.750 ;
        RECT 202.950 122.250 205.050 123.150 ;
        RECT 205.950 122.850 207.750 123.750 ;
        RECT 208.950 121.950 211.050 124.050 ;
        RECT 202.950 118.950 205.050 121.050 ;
        RECT 214.950 118.950 217.050 121.050 ;
        RECT 196.950 112.950 199.050 115.050 ;
        RECT 203.400 112.050 204.450 118.950 ;
        RECT 202.950 109.950 205.050 112.050 ;
        RECT 193.950 91.950 196.050 94.050 ;
        RECT 208.950 92.250 210.750 93.150 ;
        RECT 211.950 91.950 214.050 94.050 ;
        RECT 215.400 91.050 216.450 118.950 ;
        RECT 218.400 118.050 219.450 160.950 ;
        RECT 217.950 115.950 220.050 118.050 ;
        RECT 218.400 94.050 219.450 115.950 ;
        RECT 221.400 100.050 222.450 193.950 ;
        RECT 236.400 193.050 237.450 194.400 ;
        RECT 238.950 193.950 241.050 194.400 ;
        RECT 244.950 193.950 247.050 196.050 ;
        RECT 235.950 190.950 238.050 193.050 ;
        RECT 245.400 175.050 246.450 193.950 ;
        RECT 244.950 172.950 247.050 175.050 ;
        RECT 275.400 169.050 276.450 256.950 ;
        RECT 278.400 244.050 279.450 269.400 ;
        RECT 280.950 268.950 283.050 271.050 ;
        RECT 280.950 266.850 283.050 267.750 ;
        RECT 284.400 253.050 285.450 454.950 ;
        RECT 290.400 451.050 291.450 490.950 ;
        RECT 293.400 457.050 294.450 547.950 ;
        RECT 295.950 532.950 298.050 535.050 ;
        RECT 296.400 532.050 297.450 532.950 ;
        RECT 302.400 532.050 303.450 559.950 ;
        RECT 295.950 529.950 298.050 532.050 ;
        RECT 301.950 529.950 304.050 532.050 ;
        RECT 295.950 527.850 298.050 528.750 ;
        RECT 298.950 527.250 301.050 528.150 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 299.400 490.050 300.450 490.950 ;
        RECT 305.400 490.050 306.450 562.950 ;
        RECT 307.950 559.950 310.050 562.050 ;
        RECT 313.950 561.450 316.050 562.050 ;
        RECT 311.250 560.250 312.750 561.150 ;
        RECT 313.950 560.400 318.450 561.450 ;
        RECT 313.950 559.950 316.050 560.400 ;
        RECT 307.950 557.850 309.750 558.750 ;
        RECT 310.950 556.950 313.050 559.050 ;
        RECT 314.250 557.850 316.050 558.750 ;
        RECT 317.400 556.050 318.450 560.400 ;
        RECT 316.950 553.950 319.050 556.050 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 313.950 524.250 315.750 525.150 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 320.250 524.250 322.050 525.150 ;
        RECT 298.950 489.450 301.050 490.050 ;
        RECT 296.400 488.400 301.050 489.450 ;
        RECT 296.400 484.050 297.450 488.400 ;
        RECT 298.950 487.950 301.050 488.400 ;
        RECT 302.250 488.250 303.750 489.150 ;
        RECT 304.950 487.950 307.050 490.050 ;
        RECT 298.950 485.850 300.750 486.750 ;
        RECT 301.950 484.950 304.050 487.050 ;
        RECT 305.250 485.850 307.050 486.750 ;
        RECT 295.950 481.950 298.050 484.050 ;
        RECT 307.950 457.950 310.050 460.050 ;
        RECT 292.950 454.950 295.050 457.050 ;
        RECT 292.950 451.950 295.050 454.050 ;
        RECT 298.950 452.250 300.750 453.150 ;
        RECT 301.950 451.950 304.050 454.050 ;
        RECT 305.250 452.250 307.050 453.150 ;
        RECT 289.950 448.950 292.050 451.050 ;
        RECT 293.400 421.050 294.450 451.950 ;
        RECT 298.950 448.950 301.050 451.050 ;
        RECT 302.250 449.850 303.750 450.750 ;
        RECT 304.950 450.450 307.050 451.050 ;
        RECT 308.400 450.450 309.450 457.950 ;
        RECT 304.950 449.400 309.450 450.450 ;
        RECT 304.950 448.950 307.050 449.400 ;
        RECT 304.950 427.950 307.050 430.050 ;
        RECT 305.400 424.050 306.450 427.950 ;
        RECT 304.950 421.950 307.050 424.050 ;
        RECT 292.950 418.950 295.050 421.050 ;
        RECT 295.950 419.250 298.050 420.150 ;
        RECT 286.950 417.450 289.050 418.050 ;
        RECT 289.950 417.450 292.050 418.050 ;
        RECT 286.950 416.400 292.050 417.450 ;
        RECT 286.950 415.950 289.050 416.400 ;
        RECT 289.950 415.950 292.050 416.400 ;
        RECT 293.250 416.250 294.750 417.150 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 299.250 416.250 301.050 417.150 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 289.950 413.850 291.750 414.750 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 287.400 385.050 288.450 412.950 ;
        RECT 289.950 409.950 292.050 412.050 ;
        RECT 286.950 382.950 289.050 385.050 ;
        RECT 287.400 379.050 288.450 382.950 ;
        RECT 286.950 376.950 289.050 379.050 ;
        RECT 290.400 343.050 291.450 409.950 ;
        RECT 299.400 409.050 300.450 412.950 ;
        RECT 298.950 406.950 301.050 409.050 ;
        RECT 302.400 406.050 303.450 412.950 ;
        RECT 301.950 403.950 304.050 406.050 ;
        RECT 295.950 380.250 297.750 381.150 ;
        RECT 298.950 379.950 301.050 382.050 ;
        RECT 302.250 380.250 304.050 381.150 ;
        RECT 295.950 376.950 298.050 379.050 ;
        RECT 299.250 377.850 300.750 378.750 ;
        RECT 301.950 376.950 304.050 379.050 ;
        RECT 296.400 364.050 297.450 376.950 ;
        RECT 295.950 361.950 298.050 364.050 ;
        RECT 305.400 361.050 306.450 421.950 ;
        RECT 311.400 421.050 312.450 523.950 ;
        RECT 313.950 520.950 316.050 523.050 ;
        RECT 317.250 521.850 318.750 522.750 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 320.400 520.050 321.450 520.950 ;
        RECT 319.950 517.950 322.050 520.050 ;
        RECT 320.400 493.050 321.450 517.950 ;
        RECT 323.400 508.050 324.450 592.950 ;
        RECT 326.400 565.050 327.450 602.400 ;
        RECT 334.950 600.450 337.050 601.050 ;
        RECT 332.400 599.400 337.050 600.450 ;
        RECT 332.400 589.050 333.450 599.400 ;
        RECT 334.950 598.950 337.050 599.400 ;
        RECT 338.250 599.250 339.750 600.150 ;
        RECT 340.950 598.950 343.050 601.050 ;
        RECT 334.950 596.850 336.750 597.750 ;
        RECT 337.950 595.950 340.050 598.050 ;
        RECT 341.250 596.850 342.750 597.750 ;
        RECT 343.950 595.950 346.050 598.050 ;
        RECT 343.950 593.850 346.050 594.750 ;
        RECT 331.950 586.950 334.050 589.050 ;
        RECT 347.400 574.050 348.450 691.950 ;
        RECT 349.950 676.950 352.050 679.050 ;
        RECT 350.400 673.050 351.450 676.950 ;
        RECT 353.400 676.050 354.450 694.950 ;
        RECT 356.400 682.050 357.450 697.950 ;
        RECT 355.950 679.950 358.050 682.050 ;
        RECT 352.950 673.950 355.050 676.050 ;
        RECT 356.400 673.050 357.450 679.950 ;
        RECT 349.950 670.950 352.050 673.050 ;
        RECT 353.250 671.850 354.750 672.750 ;
        RECT 355.950 670.950 358.050 673.050 ;
        RECT 349.950 668.850 352.050 669.750 ;
        RECT 355.950 668.850 358.050 669.750 ;
        RECT 359.400 636.450 360.450 742.950 ;
        RECT 361.950 740.850 364.050 741.750 ;
        RECT 367.950 740.850 370.050 741.750 ;
        RECT 364.950 706.950 367.050 709.050 ;
        RECT 365.400 706.050 366.450 706.950 ;
        RECT 364.950 703.950 367.050 706.050 ;
        RECT 368.250 704.250 369.750 705.150 ;
        RECT 370.950 703.950 373.050 706.050 ;
        RECT 374.400 703.050 375.450 766.950 ;
        RECT 388.950 745.950 391.050 748.050 ;
        RECT 397.950 745.950 400.050 748.050 ;
        RECT 389.400 745.050 390.450 745.950 ;
        RECT 385.950 742.950 388.050 745.050 ;
        RECT 388.950 742.950 391.050 745.050 ;
        RECT 392.250 743.250 393.750 744.150 ;
        RECT 394.950 742.950 397.050 745.050 ;
        RECT 386.400 742.050 387.450 742.950 ;
        RECT 385.950 739.950 388.050 742.050 ;
        RECT 389.250 740.850 390.750 741.750 ;
        RECT 391.950 739.950 394.050 742.050 ;
        RECT 395.250 740.850 397.050 741.750 ;
        RECT 385.950 737.850 388.050 738.750 ;
        RECT 392.400 730.050 393.450 739.950 ;
        RECT 398.400 733.050 399.450 745.950 ;
        RECT 401.400 745.050 402.450 769.950 ;
        RECT 400.950 742.950 403.050 745.050 ;
        RECT 404.400 739.050 405.450 772.950 ;
        RECT 403.950 736.950 406.050 739.050 ;
        RECT 397.950 730.950 400.050 733.050 ;
        RECT 391.950 727.950 394.050 730.050 ;
        RECT 394.950 704.250 397.050 705.150 ;
        RECT 361.950 700.950 364.050 703.050 ;
        RECT 364.950 701.850 366.750 702.750 ;
        RECT 367.950 700.950 370.050 703.050 ;
        RECT 371.250 701.850 373.050 702.750 ;
        RECT 373.950 700.950 376.050 703.050 ;
        RECT 385.950 701.250 387.750 702.150 ;
        RECT 388.950 700.950 391.050 703.050 ;
        RECT 392.250 701.250 393.750 702.150 ;
        RECT 394.950 700.950 397.050 703.050 ;
        RECT 362.400 679.050 363.450 700.950 ;
        RECT 385.950 697.950 388.050 700.050 ;
        RECT 389.250 698.850 390.750 699.750 ;
        RECT 391.950 697.950 394.050 700.050 ;
        RECT 386.400 685.050 387.450 697.950 ;
        RECT 404.400 685.050 405.450 736.950 ;
        RECT 407.400 730.050 408.450 775.950 ;
        RECT 409.950 773.250 412.050 774.150 ;
        RECT 415.950 773.250 418.050 774.150 ;
        RECT 428.400 772.050 429.450 823.950 ;
        RECT 443.400 820.050 444.450 841.950 ;
        RECT 446.400 826.050 447.450 841.950 ;
        RECT 452.400 841.050 453.450 841.950 ;
        RECT 451.950 838.950 454.050 841.050 ;
        RECT 445.950 823.950 448.050 826.050 ;
        RECT 442.950 819.450 445.050 820.050 ;
        RECT 442.950 818.400 447.450 819.450 ;
        RECT 442.950 817.950 445.050 818.400 ;
        RECT 439.950 815.250 442.050 816.150 ;
        RECT 442.950 815.850 445.050 816.750 ;
        RECT 439.950 811.950 442.050 814.050 ;
        RECT 440.400 808.050 441.450 811.950 ;
        RECT 446.400 811.050 447.450 818.400 ;
        RECT 445.950 808.950 448.050 811.050 ;
        RECT 439.950 805.950 442.050 808.050 ;
        RECT 445.950 805.950 448.050 808.050 ;
        RECT 433.950 777.450 436.050 778.050 ;
        RECT 431.400 776.400 436.050 777.450 ;
        RECT 439.950 777.450 442.050 778.050 ;
        RECT 409.950 769.950 412.050 772.050 ;
        RECT 413.250 770.250 414.750 771.150 ;
        RECT 415.950 769.950 418.050 772.050 ;
        RECT 427.950 769.950 430.050 772.050 ;
        RECT 410.400 745.050 411.450 769.950 ;
        RECT 416.400 769.050 417.450 769.950 ;
        RECT 412.950 766.950 415.050 769.050 ;
        RECT 415.950 766.950 418.050 769.050 ;
        RECT 413.400 766.050 414.450 766.950 ;
        RECT 431.400 766.050 432.450 776.400 ;
        RECT 433.950 775.950 436.050 776.400 ;
        RECT 437.250 776.250 438.750 777.150 ;
        RECT 439.950 776.400 444.450 777.450 ;
        RECT 439.950 775.950 442.050 776.400 ;
        RECT 433.950 773.850 435.750 774.750 ;
        RECT 436.950 772.950 439.050 775.050 ;
        RECT 440.250 773.850 442.050 774.750 ;
        RECT 439.950 769.950 442.050 772.050 ;
        RECT 412.950 763.950 415.050 766.050 ;
        RECT 430.950 763.950 433.050 766.050 ;
        RECT 418.950 748.950 421.050 751.050 ;
        RECT 409.950 742.950 412.050 745.050 ;
        RECT 412.950 742.950 415.050 745.050 ;
        RECT 413.400 742.050 414.450 742.950 ;
        RECT 409.950 740.250 411.750 741.150 ;
        RECT 412.950 739.950 415.050 742.050 ;
        RECT 416.250 740.250 418.050 741.150 ;
        RECT 409.950 736.950 412.050 739.050 ;
        RECT 413.250 737.850 414.750 738.750 ;
        RECT 415.950 736.950 418.050 739.050 ;
        RECT 406.950 727.950 409.050 730.050 ;
        RECT 409.950 718.950 412.050 721.050 ;
        RECT 410.400 706.050 411.450 718.950 ;
        RECT 409.950 705.450 412.050 706.050 ;
        RECT 407.400 704.400 412.050 705.450 ;
        RECT 407.400 694.050 408.450 704.400 ;
        RECT 409.950 703.950 412.050 704.400 ;
        RECT 413.250 704.250 414.750 705.150 ;
        RECT 409.950 701.850 411.750 702.750 ;
        RECT 412.950 700.950 415.050 703.050 ;
        RECT 416.250 701.850 418.050 702.750 ;
        RECT 406.950 691.950 409.050 694.050 ;
        RECT 385.950 682.950 388.050 685.050 ;
        RECT 403.950 682.950 406.050 685.050 ;
        RECT 382.950 679.950 385.050 682.050 ;
        RECT 361.950 676.950 364.050 679.050 ;
        RECT 370.950 670.950 373.050 673.050 ;
        RECT 376.950 672.450 379.050 673.050 ;
        RECT 374.250 671.250 375.750 672.150 ;
        RECT 376.950 671.400 381.450 672.450 ;
        RECT 376.950 670.950 379.050 671.400 ;
        RECT 380.400 670.050 381.450 671.400 ;
        RECT 367.950 669.450 370.050 670.050 ;
        RECT 365.400 668.400 370.050 669.450 ;
        RECT 371.250 668.850 372.750 669.750 ;
        RECT 359.400 635.400 363.450 636.450 ;
        RECT 358.950 632.250 361.050 633.150 ;
        RECT 349.950 629.250 351.750 630.150 ;
        RECT 352.950 628.950 355.050 631.050 ;
        RECT 358.950 630.450 361.050 631.050 ;
        RECT 362.400 630.450 363.450 635.400 ;
        RECT 365.400 631.050 366.450 668.400 ;
        RECT 367.950 667.950 370.050 668.400 ;
        RECT 373.950 667.950 376.050 670.050 ;
        RECT 377.250 668.850 379.050 669.750 ;
        RECT 379.950 667.950 382.050 670.050 ;
        RECT 367.950 665.850 370.050 666.750 ;
        RECT 374.400 664.050 375.450 667.950 ;
        RECT 373.950 661.950 376.050 664.050 ;
        RECT 376.950 661.950 379.050 664.050 ;
        RECT 377.400 634.050 378.450 661.950 ;
        RECT 374.250 632.250 375.750 633.150 ;
        RECT 376.950 631.950 379.050 634.050 ;
        RECT 356.250 629.250 357.750 630.150 ;
        RECT 358.950 629.400 363.450 630.450 ;
        RECT 358.950 628.950 361.050 629.400 ;
        RECT 364.950 628.950 367.050 631.050 ;
        RECT 370.950 629.850 372.750 630.750 ;
        RECT 373.950 628.950 376.050 631.050 ;
        RECT 377.250 629.850 379.050 630.750 ;
        RECT 349.950 625.950 352.050 628.050 ;
        RECT 353.250 626.850 354.750 627.750 ;
        RECT 355.950 625.950 358.050 628.050 ;
        RECT 358.950 625.950 361.050 628.050 ;
        RECT 346.950 571.950 349.050 574.050 ;
        RECT 325.950 562.950 328.050 565.050 ;
        RECT 337.950 562.950 340.050 565.050 ;
        RECT 331.950 560.250 334.050 561.150 ;
        RECT 338.400 559.050 339.450 562.950 ;
        RECT 343.950 559.950 346.050 562.050 ;
        RECT 331.950 556.950 334.050 559.050 ;
        RECT 335.250 557.250 336.750 558.150 ;
        RECT 337.950 556.950 340.050 559.050 ;
        RECT 341.250 557.250 343.050 558.150 ;
        RECT 344.400 556.050 345.450 559.950 ;
        RECT 334.950 553.950 337.050 556.050 ;
        RECT 338.250 554.850 339.750 555.750 ;
        RECT 340.950 553.950 343.050 556.050 ;
        RECT 343.950 553.950 346.050 556.050 ;
        RECT 350.400 553.050 351.450 625.950 ;
        RECT 356.400 625.050 357.450 625.950 ;
        RECT 355.950 622.950 358.050 625.050 ;
        RECT 352.950 595.950 355.050 598.050 ;
        RECT 353.400 559.050 354.450 595.950 ;
        RECT 355.950 562.950 358.050 565.050 ;
        RECT 356.400 559.050 357.450 562.950 ;
        RECT 352.950 556.950 355.050 559.050 ;
        RECT 355.950 556.950 358.050 559.050 ;
        RECT 352.950 554.850 355.050 555.750 ;
        RECT 355.950 554.250 358.050 555.150 ;
        RECT 343.950 550.950 346.050 553.050 ;
        RECT 349.950 550.950 352.050 553.050 ;
        RECT 355.950 550.950 358.050 553.050 ;
        RECT 328.950 529.950 331.050 532.050 ;
        RECT 331.950 529.950 334.050 532.050 ;
        RECT 340.950 529.950 343.050 532.050 ;
        RECT 322.950 505.950 325.050 508.050 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 313.950 487.950 316.050 490.050 ;
        RECT 314.400 463.050 315.450 487.950 ;
        RECT 313.950 460.950 316.050 463.050 ;
        RECT 314.400 457.050 315.450 460.950 ;
        RECT 313.950 454.950 316.050 457.050 ;
        RECT 317.400 454.050 318.450 490.950 ;
        RECT 323.400 487.050 324.450 490.950 ;
        RECT 319.950 485.250 321.750 486.150 ;
        RECT 322.950 484.950 325.050 487.050 ;
        RECT 319.950 481.950 322.050 484.050 ;
        RECT 323.250 482.850 325.050 483.750 ;
        RECT 320.400 460.050 321.450 481.950 ;
        RECT 319.950 457.950 322.050 460.050 ;
        RECT 329.400 457.050 330.450 529.950 ;
        RECT 331.950 527.850 334.050 528.750 ;
        RECT 334.950 527.250 337.050 528.150 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 335.400 514.050 336.450 523.950 ;
        RECT 341.400 523.050 342.450 529.950 ;
        RECT 340.950 520.950 343.050 523.050 ;
        RECT 344.400 520.050 345.450 550.950 ;
        RECT 359.400 529.050 360.450 625.950 ;
        RECT 383.400 625.050 384.450 679.950 ;
        RECT 385.950 673.950 388.050 676.050 ;
        RECT 397.950 673.950 400.050 676.050 ;
        RECT 385.950 671.850 388.050 672.750 ;
        RECT 388.950 671.250 391.050 672.150 ;
        RECT 388.950 667.950 391.050 670.050 ;
        RECT 398.400 666.450 399.450 673.950 ;
        RECT 404.400 670.050 405.450 682.950 ;
        RECT 409.950 673.950 412.050 676.050 ;
        RECT 400.950 668.250 402.750 669.150 ;
        RECT 403.950 667.950 406.050 670.050 ;
        RECT 407.250 668.250 409.050 669.150 ;
        RECT 400.950 666.450 403.050 667.050 ;
        RECT 398.400 665.400 403.050 666.450 ;
        RECT 404.250 665.850 405.750 666.750 ;
        RECT 406.950 666.450 409.050 667.050 ;
        RECT 410.400 666.450 411.450 673.950 ;
        RECT 400.950 664.950 403.050 665.400 ;
        RECT 406.950 665.400 411.450 666.450 ;
        RECT 406.950 664.950 409.050 665.400 ;
        RECT 400.950 661.950 403.050 664.050 ;
        RECT 388.950 629.250 391.050 630.150 ;
        RECT 394.950 629.250 397.050 630.150 ;
        RECT 388.950 625.950 391.050 628.050 ;
        RECT 392.250 626.250 393.750 627.150 ;
        RECT 394.950 625.950 397.050 628.050 ;
        RECT 382.950 622.950 385.050 625.050 ;
        RECT 389.400 622.050 390.450 625.950 ;
        RECT 391.950 622.950 394.050 625.050 ;
        RECT 388.950 619.950 391.050 622.050 ;
        RECT 388.950 616.950 391.050 619.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 365.400 601.050 366.450 601.950 ;
        RECT 364.950 598.950 367.050 601.050 ;
        RECT 365.400 598.050 366.450 598.950 ;
        RECT 374.400 598.050 375.450 601.950 ;
        RECT 361.950 596.250 363.750 597.150 ;
        RECT 364.950 595.950 367.050 598.050 ;
        RECT 370.950 595.950 373.050 598.050 ;
        RECT 373.950 595.950 376.050 598.050 ;
        RECT 361.950 592.950 364.050 595.050 ;
        RECT 365.250 593.850 366.750 594.750 ;
        RECT 367.950 592.950 370.050 595.050 ;
        RECT 371.250 593.850 373.050 594.750 ;
        RECT 377.400 592.050 378.450 601.950 ;
        RECT 389.400 601.050 390.450 616.950 ;
        RECT 379.950 599.250 382.050 600.150 ;
        RECT 382.950 599.850 385.050 600.750 ;
        RECT 385.950 599.250 387.750 600.150 ;
        RECT 388.950 598.950 391.050 601.050 ;
        RECT 379.950 595.950 382.050 598.050 ;
        RECT 385.950 595.950 388.050 598.050 ;
        RECT 389.250 596.850 391.050 597.750 ;
        RECT 386.400 595.050 387.450 595.950 ;
        RECT 395.400 595.050 396.450 625.950 ;
        RECT 385.950 592.950 388.050 595.050 ;
        RECT 388.950 592.950 391.050 595.050 ;
        RECT 394.950 592.950 397.050 595.050 ;
        RECT 367.950 590.850 370.050 591.750 ;
        RECT 370.950 589.950 373.050 592.050 ;
        RECT 376.950 589.950 379.050 592.050 ;
        RECT 371.400 562.050 372.450 589.950 ;
        RECT 376.950 563.250 379.050 564.150 ;
        RECT 370.950 559.950 373.050 562.050 ;
        RECT 374.250 560.250 375.750 561.150 ;
        RECT 376.950 559.950 379.050 562.050 ;
        RECT 380.250 560.250 382.050 561.150 ;
        RECT 382.950 559.950 385.050 562.050 ;
        RECT 370.950 557.850 372.750 558.750 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 379.950 556.950 382.050 559.050 ;
        RECT 380.400 556.050 381.450 556.950 ;
        RECT 379.950 553.950 382.050 556.050 ;
        RECT 383.400 553.050 384.450 559.950 ;
        RECT 382.950 550.950 385.050 553.050 ;
        RECT 376.950 532.950 379.050 535.050 ;
        RECT 373.950 529.950 376.050 532.050 ;
        RECT 358.950 526.950 361.050 529.050 ;
        RECT 364.950 526.950 367.050 529.050 ;
        RECT 370.950 527.250 373.050 528.150 ;
        RECT 373.950 527.850 376.050 528.750 ;
        RECT 346.950 524.250 348.750 525.150 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 353.250 524.250 355.050 525.150 ;
        RECT 355.950 523.950 358.050 526.050 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 346.950 520.950 349.050 523.050 ;
        RECT 350.250 521.850 351.750 522.750 ;
        RECT 352.950 520.950 355.050 523.050 ;
        RECT 347.400 520.050 348.450 520.950 ;
        RECT 343.950 517.950 346.050 520.050 ;
        RECT 346.950 517.950 349.050 520.050 ;
        RECT 334.950 511.950 337.050 514.050 ;
        RECT 334.950 505.950 337.050 508.050 ;
        RECT 335.400 490.050 336.450 505.950 ;
        RECT 356.400 490.050 357.450 523.950 ;
        RECT 359.400 505.050 360.450 523.950 ;
        RECT 358.950 502.950 361.050 505.050 ;
        RECT 334.950 487.950 337.050 490.050 ;
        RECT 338.250 488.250 339.750 489.150 ;
        RECT 349.950 487.950 352.050 490.050 ;
        RECT 352.950 488.250 355.050 489.150 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 334.950 485.850 336.750 486.750 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 341.250 485.850 343.050 486.750 ;
        RECT 338.400 463.050 339.450 484.950 ;
        RECT 350.400 483.450 351.450 487.950 ;
        RECT 359.400 487.050 360.450 502.950 ;
        RECT 352.950 484.950 355.050 487.050 ;
        RECT 356.250 485.250 357.750 486.150 ;
        RECT 358.950 484.950 361.050 487.050 ;
        RECT 362.250 485.250 364.050 486.150 ;
        RECT 350.400 482.400 354.450 483.450 ;
        RECT 337.950 460.950 340.050 463.050 ;
        RECT 349.950 460.950 352.050 463.050 ;
        RECT 319.950 454.950 322.050 457.050 ;
        RECT 323.250 455.250 325.050 456.150 ;
        RECT 328.950 454.950 331.050 457.050 ;
        RECT 332.250 455.250 334.050 456.150 ;
        RECT 334.950 454.950 337.050 457.050 ;
        RECT 340.950 456.450 343.050 457.050 ;
        RECT 338.400 455.400 343.050 456.450 ;
        RECT 316.950 451.950 319.050 454.050 ;
        RECT 319.950 452.850 321.750 453.750 ;
        RECT 322.950 451.950 325.050 454.050 ;
        RECT 328.950 452.850 330.750 453.750 ;
        RECT 331.950 451.950 334.050 454.050 ;
        RECT 323.400 445.050 324.450 451.950 ;
        RECT 322.950 442.950 325.050 445.050 ;
        RECT 310.950 418.950 313.050 421.050 ;
        RECT 307.950 415.950 310.050 418.050 ;
        RECT 319.950 415.950 322.050 418.050 ;
        RECT 325.950 415.950 328.050 418.050 ;
        RECT 308.400 379.050 309.450 415.950 ;
        RECT 320.400 415.050 321.450 415.950 ;
        RECT 310.950 413.250 312.750 414.150 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 317.250 413.250 318.750 414.150 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 323.250 413.250 325.050 414.150 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 314.250 410.850 315.750 411.750 ;
        RECT 316.950 409.950 319.050 412.050 ;
        RECT 320.250 410.850 321.750 411.750 ;
        RECT 322.950 411.450 325.050 412.050 ;
        RECT 326.400 411.450 327.450 415.950 ;
        RECT 322.950 410.400 327.450 411.450 ;
        RECT 335.400 411.450 336.450 454.950 ;
        RECT 338.400 451.050 339.450 455.400 ;
        RECT 340.950 454.950 343.050 455.400 ;
        RECT 344.250 455.250 345.750 456.150 ;
        RECT 346.950 454.950 349.050 457.050 ;
        RECT 350.400 454.050 351.450 460.950 ;
        RECT 340.950 452.850 342.750 453.750 ;
        RECT 343.950 451.950 346.050 454.050 ;
        RECT 347.250 452.850 348.750 453.750 ;
        RECT 349.950 451.950 352.050 454.050 ;
        RECT 337.950 448.950 340.050 451.050 ;
        RECT 344.400 445.050 345.450 451.950 ;
        RECT 349.950 449.850 352.050 450.750 ;
        RECT 353.400 445.050 354.450 482.400 ;
        RECT 355.950 481.950 358.050 484.050 ;
        RECT 359.250 482.850 360.750 483.750 ;
        RECT 361.950 481.950 364.050 484.050 ;
        RECT 356.400 480.450 357.450 481.950 ;
        RECT 362.400 481.050 363.450 481.950 ;
        RECT 356.400 479.400 360.450 480.450 ;
        RECT 355.950 469.950 358.050 472.050 ;
        RECT 343.950 442.950 346.050 445.050 ;
        RECT 352.950 442.950 355.050 445.050 ;
        RECT 352.950 439.950 355.050 442.050 ;
        RECT 343.950 419.250 346.050 420.150 ;
        RECT 337.950 415.950 340.050 418.050 ;
        RECT 341.250 416.250 342.750 417.150 ;
        RECT 343.950 415.950 346.050 418.050 ;
        RECT 347.250 416.250 349.050 417.150 ;
        RECT 344.400 415.050 345.450 415.950 ;
        RECT 337.950 413.850 339.750 414.750 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 346.950 414.450 349.050 415.050 ;
        RECT 346.950 413.400 351.450 414.450 ;
        RECT 346.950 412.950 349.050 413.400 ;
        RECT 335.400 410.400 339.450 411.450 ;
        RECT 322.950 409.950 325.050 410.400 ;
        RECT 317.400 384.450 318.450 409.950 ;
        RECT 334.950 406.950 337.050 409.050 ;
        RECT 319.950 385.950 322.050 388.050 ;
        RECT 314.400 383.400 318.450 384.450 ;
        RECT 307.950 376.950 310.050 379.050 ;
        RECT 310.950 364.950 313.050 367.050 ;
        RECT 304.950 358.950 307.050 361.050 ;
        RECT 311.400 343.050 312.450 364.950 ;
        RECT 314.400 345.450 315.450 383.400 ;
        RECT 320.400 382.050 321.450 385.950 ;
        RECT 316.950 380.250 318.750 381.150 ;
        RECT 319.950 379.950 322.050 382.050 ;
        RECT 322.950 379.950 325.050 382.050 ;
        RECT 325.950 381.450 328.050 382.050 ;
        RECT 325.950 380.400 330.450 381.450 ;
        RECT 325.950 379.950 328.050 380.400 ;
        RECT 323.400 379.050 324.450 379.950 ;
        RECT 316.950 376.950 319.050 379.050 ;
        RECT 320.250 377.850 321.750 378.750 ;
        RECT 322.950 376.950 325.050 379.050 ;
        RECT 326.250 377.850 328.050 378.750 ;
        RECT 322.950 374.850 325.050 375.750 ;
        RECT 329.400 373.050 330.450 380.400 ;
        RECT 335.400 379.050 336.450 406.950 ;
        RECT 338.400 385.050 339.450 410.400 ;
        RECT 341.400 406.050 342.450 412.950 ;
        RECT 350.400 412.050 351.450 413.400 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 340.950 403.950 343.050 406.050 ;
        RECT 337.950 382.950 340.050 385.050 ;
        RECT 337.950 379.950 340.050 382.050 ;
        RECT 340.950 380.250 342.750 381.150 ;
        RECT 343.950 379.950 346.050 382.050 ;
        RECT 347.250 380.250 349.050 381.150 ;
        RECT 334.950 376.950 337.050 379.050 ;
        RECT 338.400 375.450 339.450 379.950 ;
        RECT 340.950 376.950 343.050 379.050 ;
        RECT 344.250 377.850 345.750 378.750 ;
        RECT 346.950 376.950 349.050 379.050 ;
        RECT 338.400 374.400 342.450 375.450 ;
        RECT 322.950 370.950 325.050 373.050 ;
        RECT 328.950 370.950 331.050 373.050 ;
        RECT 314.400 344.400 318.450 345.450 ;
        RECT 286.950 341.250 289.050 342.150 ;
        RECT 289.950 340.950 292.050 343.050 ;
        RECT 301.950 341.250 303.750 342.150 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 308.250 341.250 309.750 342.150 ;
        RECT 310.950 340.950 313.050 343.050 ;
        RECT 314.250 341.250 316.050 342.150 ;
        RECT 301.950 337.950 304.050 340.050 ;
        RECT 305.250 338.850 306.750 339.750 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 311.250 338.850 312.750 339.750 ;
        RECT 313.950 337.950 316.050 340.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 299.400 328.050 300.450 334.950 ;
        RECT 298.950 325.950 301.050 328.050 ;
        RECT 286.950 319.950 289.050 322.050 ;
        RECT 283.950 250.950 286.050 253.050 ;
        RECT 287.400 247.050 288.450 319.950 ;
        RECT 295.950 313.950 298.050 316.050 ;
        RECT 296.400 313.050 297.450 313.950 ;
        RECT 292.950 311.250 294.750 312.150 ;
        RECT 295.950 310.950 298.050 313.050 ;
        RECT 292.950 307.950 295.050 310.050 ;
        RECT 296.250 308.850 298.050 309.750 ;
        RECT 299.400 309.450 300.450 325.950 ;
        RECT 302.400 325.050 303.450 337.950 ;
        RECT 301.950 322.950 304.050 325.050 ;
        RECT 308.400 322.050 309.450 337.950 ;
        RECT 307.950 319.950 310.050 322.050 ;
        RECT 304.950 312.450 307.050 313.050 ;
        RECT 301.950 311.250 303.750 312.150 ;
        RECT 304.950 311.400 309.450 312.450 ;
        RECT 304.950 310.950 307.050 311.400 ;
        RECT 301.950 309.450 304.050 310.050 ;
        RECT 299.400 308.400 304.050 309.450 ;
        RECT 305.250 308.850 307.050 309.750 ;
        RECT 301.950 307.950 304.050 308.400 ;
        RECT 293.400 274.050 294.450 307.950 ;
        RECT 308.400 292.050 309.450 311.400 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 317.400 280.050 318.450 344.400 ;
        RECT 319.950 328.950 322.050 331.050 ;
        RECT 320.400 313.050 321.450 328.950 ;
        RECT 323.400 316.050 324.450 370.950 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 335.400 343.050 336.450 367.950 ;
        RECT 325.950 341.250 327.750 342.150 ;
        RECT 328.950 340.950 331.050 343.050 ;
        RECT 332.250 341.250 333.750 342.150 ;
        RECT 334.950 340.950 337.050 343.050 ;
        RECT 338.250 341.250 340.050 342.150 ;
        RECT 341.400 340.050 342.450 374.400 ;
        RECT 347.400 349.050 348.450 376.950 ;
        RECT 350.400 349.050 351.450 409.950 ;
        RECT 353.400 355.050 354.450 439.950 ;
        RECT 356.400 382.050 357.450 469.950 ;
        RECT 359.400 469.050 360.450 479.400 ;
        RECT 361.950 478.950 364.050 481.050 ;
        RECT 365.400 472.050 366.450 526.950 ;
        RECT 377.400 526.050 378.450 532.950 ;
        RECT 379.950 529.950 382.050 532.050 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 380.400 523.050 381.450 529.950 ;
        RECT 379.950 520.950 382.050 523.050 ;
        RECT 379.950 490.950 382.050 493.050 ;
        RECT 380.400 490.050 381.450 490.950 ;
        RECT 373.950 487.950 376.050 490.050 ;
        RECT 377.250 488.250 378.750 489.150 ;
        RECT 379.950 487.950 382.050 490.050 ;
        RECT 373.950 485.850 375.750 486.750 ;
        RECT 376.950 484.950 379.050 487.050 ;
        RECT 380.250 485.850 382.050 486.750 ;
        RECT 383.400 484.050 384.450 550.950 ;
        RECT 386.400 535.050 387.450 592.950 ;
        RECT 389.400 555.450 390.450 592.950 ;
        RECT 401.400 571.050 402.450 661.950 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 403.950 628.950 406.050 631.050 ;
        RECT 404.400 619.050 405.450 628.950 ;
        RECT 407.400 627.450 408.450 646.950 ;
        RECT 419.400 636.450 420.450 748.950 ;
        RECT 421.950 745.950 424.050 748.050 ;
        RECT 427.950 745.950 430.050 748.050 ;
        RECT 422.400 739.050 423.450 745.950 ;
        RECT 424.950 743.250 427.050 744.150 ;
        RECT 427.950 743.850 430.050 744.750 ;
        RECT 433.950 744.450 436.050 745.050 ;
        RECT 430.950 743.250 432.750 744.150 ;
        RECT 433.950 743.400 438.450 744.450 ;
        RECT 433.950 742.950 436.050 743.400 ;
        RECT 424.950 739.950 427.050 742.050 ;
        RECT 430.950 739.950 433.050 742.050 ;
        RECT 434.250 740.850 436.050 741.750 ;
        RECT 421.950 736.950 424.050 739.050 ;
        RECT 424.950 736.950 427.050 739.050 ;
        RECT 422.400 694.050 423.450 736.950 ;
        RECT 425.400 700.050 426.450 736.950 ;
        RECT 437.400 736.050 438.450 743.400 ;
        RECT 440.400 738.450 441.450 769.950 ;
        RECT 443.400 769.050 444.450 776.400 ;
        RECT 442.950 766.950 445.050 769.050 ;
        RECT 446.400 751.050 447.450 805.950 ;
        RECT 452.400 784.050 453.450 838.950 ;
        RECT 461.250 837.600 462.450 849.600 ;
        RECT 475.950 847.950 478.050 850.050 ;
        RECT 463.950 841.950 466.050 844.050 ;
        RECT 476.400 843.450 477.450 847.950 ;
        RECT 482.400 847.050 483.450 850.950 ;
        RECT 478.950 845.250 480.750 846.150 ;
        RECT 481.950 844.950 484.050 847.050 ;
        RECT 487.950 846.450 490.050 847.050 ;
        RECT 487.950 845.400 492.450 846.450 ;
        RECT 487.950 844.950 490.050 845.400 ;
        RECT 478.950 843.450 481.050 844.050 ;
        RECT 476.400 842.400 481.050 843.450 ;
        RECT 482.250 842.850 484.050 843.750 ;
        RECT 478.950 841.950 481.050 842.400 ;
        RECT 484.950 842.250 487.050 843.150 ;
        RECT 487.950 842.850 490.050 843.750 ;
        RECT 491.400 841.050 492.450 845.400 ;
        RECT 499.950 845.250 502.050 846.150 ;
        RECT 496.950 842.250 498.750 843.150 ;
        RECT 499.950 841.950 502.050 844.050 ;
        RECT 463.950 839.850 466.050 840.750 ;
        RECT 484.950 838.950 487.050 841.050 ;
        RECT 487.950 838.950 490.050 841.050 ;
        RECT 490.950 838.950 493.050 841.050 ;
        RECT 496.950 838.950 499.050 841.050 ;
        RECT 485.400 838.050 486.450 838.950 ;
        RECT 460.950 835.500 463.050 837.600 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 472.950 814.950 475.050 817.050 ;
        RECT 478.950 814.950 481.050 817.050 ;
        RECT 484.950 814.950 487.050 817.050 ;
        RECT 457.950 812.250 459.750 813.150 ;
        RECT 460.950 811.950 463.050 814.050 ;
        RECT 464.250 812.250 466.050 813.150 ;
        RECT 457.950 808.950 460.050 811.050 ;
        RECT 461.250 809.850 462.750 810.750 ;
        RECT 463.950 808.950 466.050 811.050 ;
        RECT 458.400 807.450 459.450 808.950 ;
        RECT 458.400 806.400 462.450 807.450 ;
        RECT 461.400 796.050 462.450 806.400 ;
        RECT 460.950 793.950 463.050 796.050 ;
        RECT 451.950 781.950 454.050 784.050 ;
        RECT 451.950 775.950 454.050 778.050 ;
        RECT 457.950 776.250 460.050 777.150 ;
        RECT 452.400 775.050 453.450 775.950 ;
        RECT 448.950 773.250 450.750 774.150 ;
        RECT 451.950 772.950 454.050 775.050 ;
        RECT 455.250 773.250 456.750 774.150 ;
        RECT 457.950 772.950 460.050 775.050 ;
        RECT 448.950 769.950 451.050 772.050 ;
        RECT 452.250 770.850 453.750 771.750 ;
        RECT 454.950 769.950 457.050 772.050 ;
        RECT 445.950 748.950 448.050 751.050 ;
        RECT 451.950 748.950 454.050 751.050 ;
        RECT 445.950 747.450 448.050 748.050 ;
        RECT 443.400 746.400 448.050 747.450 ;
        RECT 443.400 742.050 444.450 746.400 ;
        RECT 445.950 745.950 448.050 746.400 ;
        RECT 445.950 743.850 448.050 744.750 ;
        RECT 448.950 743.250 451.050 744.150 ;
        RECT 442.950 739.950 445.050 742.050 ;
        RECT 448.950 739.950 451.050 742.050 ;
        RECT 440.400 737.400 444.450 738.450 ;
        RECT 436.950 733.950 439.050 736.050 ;
        RECT 430.950 704.250 433.050 705.150 ;
        RECT 436.950 703.950 439.050 706.050 ;
        RECT 437.400 703.050 438.450 703.950 ;
        RECT 430.950 700.950 433.050 703.050 ;
        RECT 434.250 701.250 435.750 702.150 ;
        RECT 436.950 700.950 439.050 703.050 ;
        RECT 440.250 701.250 442.050 702.150 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 431.400 697.050 432.450 700.950 ;
        RECT 433.950 697.950 436.050 700.050 ;
        RECT 437.250 698.850 438.750 699.750 ;
        RECT 439.950 697.950 442.050 700.050 ;
        RECT 434.400 697.050 435.450 697.950 ;
        RECT 443.400 697.050 444.450 737.400 ;
        RECT 449.400 730.050 450.450 739.950 ;
        RECT 448.950 727.950 451.050 730.050 ;
        RECT 445.950 703.950 448.050 706.050 ;
        RECT 446.400 697.050 447.450 703.950 ;
        RECT 452.400 700.050 453.450 748.950 ;
        RECT 454.950 706.950 457.050 709.050 ;
        RECT 455.400 703.050 456.450 706.950 ;
        RECT 454.950 700.950 457.050 703.050 ;
        RECT 451.950 697.950 454.050 700.050 ;
        RECT 454.950 698.850 457.050 699.750 ;
        RECT 457.950 698.250 460.050 699.150 ;
        RECT 424.950 694.950 427.050 697.050 ;
        RECT 430.950 694.950 433.050 697.050 ;
        RECT 433.950 694.950 436.050 697.050 ;
        RECT 439.950 694.950 442.050 697.050 ;
        RECT 442.950 694.950 445.050 697.050 ;
        RECT 445.950 694.950 448.050 697.050 ;
        RECT 457.950 694.950 460.050 697.050 ;
        RECT 421.950 691.950 424.050 694.050 ;
        RECT 425.400 670.050 426.450 694.950 ;
        RECT 436.950 676.950 439.050 679.050 ;
        RECT 421.950 668.250 423.750 669.150 ;
        RECT 424.950 667.950 427.050 670.050 ;
        RECT 428.250 668.250 430.050 669.150 ;
        RECT 421.950 664.950 424.050 667.050 ;
        RECT 425.250 665.850 426.750 666.750 ;
        RECT 422.400 664.050 423.450 664.950 ;
        RECT 421.950 661.950 424.050 664.050 ;
        RECT 419.400 635.400 423.450 636.450 ;
        RECT 409.950 629.250 411.750 630.150 ;
        RECT 412.950 628.950 415.050 631.050 ;
        RECT 418.950 628.950 421.050 631.050 ;
        RECT 409.950 627.450 412.050 628.050 ;
        RECT 407.400 626.400 412.050 627.450 ;
        RECT 413.250 626.850 415.050 627.750 ;
        RECT 409.950 625.950 412.050 626.400 ;
        RECT 415.950 626.250 418.050 627.150 ;
        RECT 418.950 626.850 421.050 627.750 ;
        RECT 415.950 622.950 418.050 625.050 ;
        RECT 403.950 616.950 406.050 619.050 ;
        RECT 416.400 601.050 417.450 622.950 ;
        RECT 418.950 619.950 421.050 622.050 ;
        RECT 419.400 613.050 420.450 619.950 ;
        RECT 418.950 610.950 421.050 613.050 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 403.950 596.250 405.750 597.150 ;
        RECT 406.950 595.950 409.050 598.050 ;
        RECT 410.250 596.250 412.050 597.150 ;
        RECT 403.950 592.950 406.050 595.050 ;
        RECT 407.250 593.850 408.750 594.750 ;
        RECT 404.400 583.050 405.450 592.950 ;
        RECT 403.950 580.950 406.050 583.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 391.950 565.950 394.050 568.050 ;
        RECT 392.400 562.050 393.450 565.950 ;
        RECT 397.950 563.250 400.050 564.150 ;
        RECT 403.950 562.950 406.050 565.050 ;
        RECT 415.950 562.950 418.050 565.050 ;
        RECT 391.950 559.950 394.050 562.050 ;
        RECT 395.250 560.250 396.750 561.150 ;
        RECT 397.950 559.950 400.050 562.050 ;
        RECT 401.250 560.250 403.050 561.150 ;
        RECT 391.950 557.850 393.750 558.750 ;
        RECT 394.950 556.950 397.050 559.050 ;
        RECT 400.950 556.950 403.050 559.050 ;
        RECT 389.400 554.400 393.450 555.450 ;
        RECT 385.950 532.950 388.050 535.050 ;
        RECT 385.950 529.950 388.050 532.050 ;
        RECT 386.400 529.050 387.450 529.950 ;
        RECT 392.400 529.050 393.450 554.400 ;
        RECT 395.400 553.050 396.450 556.950 ;
        RECT 401.400 556.050 402.450 556.950 ;
        RECT 400.950 553.950 403.050 556.050 ;
        RECT 404.400 553.050 405.450 562.950 ;
        RECT 416.400 562.050 417.450 562.950 ;
        RECT 409.950 561.450 412.050 562.050 ;
        RECT 407.400 560.400 412.050 561.450 ;
        RECT 407.400 556.050 408.450 560.400 ;
        RECT 409.950 559.950 412.050 560.400 ;
        RECT 413.250 560.250 414.750 561.150 ;
        RECT 415.950 559.950 418.050 562.050 ;
        RECT 409.950 557.850 411.750 558.750 ;
        RECT 412.950 556.950 415.050 559.050 ;
        RECT 416.250 557.850 418.050 558.750 ;
        RECT 419.400 556.050 420.450 610.950 ;
        RECT 406.950 553.950 409.050 556.050 ;
        RECT 418.950 553.950 421.050 556.050 ;
        RECT 394.950 550.950 397.050 553.050 ;
        RECT 403.950 550.950 406.050 553.050 ;
        RECT 407.400 547.050 408.450 553.950 ;
        RECT 406.950 544.950 409.050 547.050 ;
        RECT 397.950 529.950 400.050 532.050 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 389.250 527.250 390.750 528.150 ;
        RECT 391.950 526.950 394.050 529.050 ;
        RECT 394.950 526.950 397.050 529.050 ;
        RECT 395.400 526.050 396.450 526.950 ;
        RECT 385.950 524.850 387.750 525.750 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 392.250 524.850 393.750 525.750 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 389.400 490.050 390.450 523.950 ;
        RECT 394.950 521.850 397.050 522.750 ;
        RECT 391.950 502.950 394.050 505.050 ;
        RECT 392.400 490.050 393.450 502.950 ;
        RECT 398.400 493.050 399.450 529.950 ;
        RECT 403.950 493.950 406.050 496.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 398.400 490.050 399.450 490.950 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 391.950 487.950 394.050 490.050 ;
        RECT 397.950 489.450 400.050 490.050 ;
        RECT 395.250 488.250 396.750 489.150 ;
        RECT 397.950 488.400 402.450 489.450 ;
        RECT 397.950 487.950 400.050 488.400 ;
        RECT 382.950 481.950 385.050 484.050 ;
        RECT 370.950 475.950 373.050 478.050 ;
        RECT 364.950 469.950 367.050 472.050 ;
        RECT 358.950 466.950 361.050 469.050 ;
        RECT 364.950 466.950 367.050 469.050 ;
        RECT 361.950 461.400 364.050 463.500 ;
        RECT 358.950 458.250 361.050 459.150 ;
        RECT 358.950 454.950 361.050 457.050 ;
        RECT 359.400 454.050 360.450 454.950 ;
        RECT 358.950 451.950 361.050 454.050 ;
        RECT 362.550 449.400 363.750 461.400 ;
        RECT 361.950 447.300 364.050 449.400 ;
        RECT 362.550 443.700 363.750 447.300 ;
        RECT 361.950 441.600 364.050 443.700 ;
        RECT 365.400 424.050 366.450 466.950 ;
        RECT 371.400 457.050 372.450 475.950 ;
        RECT 382.950 461.400 385.050 463.500 ;
        RECT 370.950 456.450 373.050 457.050 ;
        RECT 368.400 455.400 373.050 456.450 ;
        RECT 368.400 442.050 369.450 455.400 ;
        RECT 370.950 454.950 373.050 455.400 ;
        RECT 376.950 454.950 379.050 457.050 ;
        RECT 370.950 452.850 373.050 453.750 ;
        RECT 373.950 451.950 376.050 454.050 ;
        RECT 376.950 452.850 379.050 453.750 ;
        RECT 367.950 439.950 370.050 442.050 ;
        RECT 364.950 421.950 367.050 424.050 ;
        RECT 358.950 418.950 361.050 421.050 ;
        RECT 359.400 418.050 360.450 418.950 ;
        RECT 365.400 418.050 366.450 421.950 ;
        RECT 374.400 421.050 375.450 451.950 ;
        RECT 383.400 444.600 384.600 461.400 ;
        RECT 389.400 454.050 390.450 487.950 ;
        RECT 391.950 485.850 393.750 486.750 ;
        RECT 394.950 484.950 397.050 487.050 ;
        RECT 398.250 485.850 400.050 486.750 ;
        RECT 391.950 481.950 394.050 484.050 ;
        RECT 388.950 451.950 391.050 454.050 ;
        RECT 382.950 442.500 385.050 444.600 ;
        RECT 373.950 418.950 376.050 421.050 ;
        RECT 379.950 419.250 382.050 420.150 ;
        RECT 385.950 418.950 388.050 421.050 ;
        RECT 358.950 415.950 361.050 418.050 ;
        RECT 362.250 416.250 363.750 417.150 ;
        RECT 364.950 415.950 367.050 418.050 ;
        RECT 358.950 413.850 360.750 414.750 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 365.250 413.850 367.050 414.750 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 362.250 383.250 364.050 384.150 ;
        RECT 367.950 382.950 370.050 385.050 ;
        RECT 371.250 383.250 373.050 384.150 ;
        RECT 355.950 379.950 358.050 382.050 ;
        RECT 358.950 380.850 360.750 381.750 ;
        RECT 361.950 379.950 364.050 382.050 ;
        RECT 367.950 380.850 369.750 381.750 ;
        RECT 370.950 379.950 373.050 382.050 ;
        RECT 362.400 367.050 363.450 379.950 ;
        RECT 371.400 379.050 372.450 379.950 ;
        RECT 370.950 376.950 373.050 379.050 ;
        RECT 361.950 364.950 364.050 367.050 ;
        RECT 358.950 358.950 361.050 361.050 ;
        RECT 352.950 352.950 355.050 355.050 ;
        RECT 346.950 346.950 349.050 349.050 ;
        RECT 349.950 346.950 352.050 349.050 ;
        RECT 350.400 346.050 351.450 346.950 ;
        RECT 349.950 343.950 352.050 346.050 ;
        RECT 353.250 344.250 354.750 345.150 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 349.950 341.850 351.750 342.750 ;
        RECT 352.950 340.950 355.050 343.050 ;
        RECT 356.250 341.850 358.050 342.750 ;
        RECT 325.950 337.950 328.050 340.050 ;
        RECT 329.250 338.850 330.750 339.750 ;
        RECT 331.950 337.950 334.050 340.050 ;
        RECT 335.250 338.850 336.750 339.750 ;
        RECT 337.950 337.950 340.050 340.050 ;
        RECT 340.950 337.950 343.050 340.050 ;
        RECT 346.950 337.950 349.050 340.050 ;
        RECT 326.400 337.050 327.450 337.950 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 322.950 313.950 325.050 316.050 ;
        RECT 319.950 310.950 322.050 313.050 ;
        RECT 319.950 308.850 322.050 309.750 ;
        RECT 316.950 277.950 319.050 280.050 ;
        RECT 317.400 277.050 318.450 277.950 ;
        RECT 304.950 274.950 307.050 277.050 ;
        RECT 310.950 274.950 313.050 277.050 ;
        RECT 316.950 274.950 319.050 277.050 ;
        RECT 292.950 271.950 295.050 274.050 ;
        RECT 298.950 273.450 301.050 274.050 ;
        RECT 296.250 272.250 297.750 273.150 ;
        RECT 298.950 272.400 303.450 273.450 ;
        RECT 298.950 271.950 301.050 272.400 ;
        RECT 292.950 269.850 294.750 270.750 ;
        RECT 295.950 268.950 298.050 271.050 ;
        RECT 299.250 269.850 301.050 270.750 ;
        RECT 302.400 259.050 303.450 272.400 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 286.950 244.950 289.050 247.050 ;
        RECT 295.950 244.950 298.050 247.050 ;
        RECT 277.950 241.950 280.050 244.050 ;
        RECT 280.950 241.950 283.050 244.050 ;
        RECT 286.950 241.950 289.050 244.050 ;
        RECT 277.950 238.950 280.050 241.050 ;
        RECT 278.400 232.050 279.450 238.950 ;
        RECT 277.950 229.950 280.050 232.050 ;
        RECT 281.400 195.450 282.450 241.950 ;
        RECT 283.950 239.250 286.050 240.150 ;
        RECT 286.950 239.850 289.050 240.750 ;
        RECT 289.950 239.250 291.750 240.150 ;
        RECT 292.950 238.950 295.050 241.050 ;
        RECT 296.400 238.050 297.450 244.950 ;
        RECT 283.950 235.950 286.050 238.050 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 293.250 236.850 295.050 237.750 ;
        RECT 295.950 235.950 298.050 238.050 ;
        RECT 284.400 235.050 285.450 235.950 ;
        RECT 283.950 232.950 286.050 235.050 ;
        RECT 292.950 205.950 295.050 208.050 ;
        RECT 301.950 205.950 304.050 208.050 ;
        RECT 283.950 197.250 286.050 198.150 ;
        RECT 289.950 197.250 292.050 198.150 ;
        RECT 283.950 195.450 286.050 196.050 ;
        RECT 281.400 194.400 286.050 195.450 ;
        RECT 281.400 190.050 282.450 194.400 ;
        RECT 283.950 193.950 286.050 194.400 ;
        RECT 280.950 187.950 283.050 190.050 ;
        RECT 293.400 181.050 294.450 205.950 ;
        RECT 302.400 187.050 303.450 205.950 ;
        RECT 305.400 202.050 306.450 274.950 ;
        RECT 311.400 238.050 312.450 274.950 ;
        RECT 316.950 271.950 319.050 274.050 ;
        RECT 317.400 271.050 318.450 271.950 ;
        RECT 323.400 271.050 324.450 313.950 ;
        RECT 325.950 310.950 328.050 313.050 ;
        RECT 328.950 310.950 331.050 313.050 ;
        RECT 325.950 308.850 328.050 309.750 ;
        RECT 313.950 269.250 315.750 270.150 ;
        RECT 316.950 268.950 319.050 271.050 ;
        RECT 322.950 268.950 325.050 271.050 ;
        RECT 329.400 270.450 330.450 310.950 ;
        RECT 332.400 274.050 333.450 337.950 ;
        RECT 338.400 319.050 339.450 337.950 ;
        RECT 334.950 316.950 337.050 319.050 ;
        RECT 337.950 316.950 340.050 319.050 ;
        RECT 335.400 309.450 336.450 316.950 ;
        RECT 340.950 313.950 343.050 316.050 ;
        RECT 347.400 313.050 348.450 337.950 ;
        RECT 337.950 311.250 340.050 312.150 ;
        RECT 340.950 311.850 343.050 312.750 ;
        RECT 343.950 311.250 345.750 312.150 ;
        RECT 346.950 310.950 349.050 313.050 ;
        RECT 337.950 309.450 340.050 310.050 ;
        RECT 335.400 308.400 340.050 309.450 ;
        RECT 337.950 307.950 340.050 308.400 ;
        RECT 343.950 307.950 346.050 310.050 ;
        RECT 347.250 308.850 349.050 309.750 ;
        RECT 359.400 304.050 360.450 358.950 ;
        RECT 374.400 346.050 375.450 418.950 ;
        RECT 386.400 418.050 387.450 418.950 ;
        RECT 376.950 416.250 378.750 417.150 ;
        RECT 379.950 415.950 382.050 418.050 ;
        RECT 383.250 416.250 384.750 417.150 ;
        RECT 385.950 415.950 388.050 418.050 ;
        RECT 376.950 412.950 379.050 415.050 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 386.250 413.850 388.050 414.750 ;
        RECT 377.400 412.050 378.450 412.950 ;
        RECT 376.950 409.950 379.050 412.050 ;
        RECT 392.400 409.050 393.450 481.950 ;
        RECT 395.400 451.050 396.450 484.950 ;
        RECT 401.400 484.050 402.450 488.400 ;
        RECT 404.400 487.050 405.450 493.950 ;
        RECT 403.950 484.950 406.050 487.050 ;
        RECT 400.950 481.950 403.050 484.050 ;
        RECT 401.400 481.050 402.450 481.950 ;
        RECT 407.400 481.050 408.450 544.950 ;
        RECT 418.950 538.950 421.050 541.050 ;
        RECT 409.950 532.950 412.050 535.050 ;
        RECT 410.400 529.050 411.450 532.950 ;
        RECT 409.950 526.950 412.050 529.050 ;
        RECT 413.250 527.250 414.750 528.150 ;
        RECT 415.950 526.950 418.050 529.050 ;
        RECT 419.400 526.050 420.450 538.950 ;
        RECT 409.950 524.850 411.750 525.750 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 416.250 524.850 417.750 525.750 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 413.400 522.450 414.450 523.950 ;
        RECT 410.400 521.400 414.450 522.450 ;
        RECT 418.950 521.850 421.050 522.750 ;
        RECT 410.400 493.050 411.450 521.400 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 410.400 490.050 411.450 490.950 ;
        RECT 422.400 490.050 423.450 635.400 ;
        RECT 430.950 631.950 433.050 634.050 ;
        RECT 431.400 631.050 432.450 631.950 ;
        RECT 430.950 628.950 433.050 631.050 ;
        RECT 427.950 626.250 430.050 627.150 ;
        RECT 430.950 626.850 433.050 627.750 ;
        RECT 427.950 622.950 430.050 625.050 ;
        RECT 428.400 619.050 429.450 622.950 ;
        RECT 427.950 616.950 430.050 619.050 ;
        RECT 427.950 604.950 430.050 607.050 ;
        RECT 428.400 601.050 429.450 604.950 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 434.400 601.050 435.450 601.950 ;
        RECT 427.950 598.950 430.050 601.050 ;
        RECT 431.250 599.250 432.750 600.150 ;
        RECT 433.950 598.950 436.050 601.050 ;
        RECT 424.950 595.950 427.050 598.050 ;
        RECT 428.250 596.850 429.750 597.750 ;
        RECT 430.950 595.950 433.050 598.050 ;
        RECT 434.250 596.850 436.050 597.750 ;
        RECT 424.950 593.850 427.050 594.750 ;
        RECT 431.400 583.050 432.450 595.950 ;
        RECT 430.950 580.950 433.050 583.050 ;
        RECT 424.950 559.950 427.050 562.050 ;
        RECT 431.250 560.250 432.750 561.150 ;
        RECT 433.950 559.950 436.050 562.050 ;
        RECT 425.400 526.050 426.450 559.950 ;
        RECT 427.950 557.850 429.750 558.750 ;
        RECT 430.950 556.950 433.050 559.050 ;
        RECT 434.250 557.850 436.050 558.750 ;
        RECT 431.400 541.050 432.450 556.950 ;
        RECT 437.400 541.050 438.450 676.950 ;
        RECT 440.400 664.050 441.450 694.950 ;
        RECT 445.950 691.950 448.050 694.050 ;
        RECT 446.400 673.050 447.450 691.950 ;
        RECT 458.400 691.050 459.450 694.950 ;
        RECT 457.950 688.950 460.050 691.050 ;
        RECT 461.400 678.450 462.450 793.950 ;
        RECT 466.950 790.950 469.050 793.050 ;
        RECT 463.950 772.950 466.050 775.050 ;
        RECT 464.400 745.050 465.450 772.950 ;
        RECT 467.400 772.050 468.450 790.950 ;
        RECT 473.400 781.050 474.450 814.950 ;
        RECT 479.400 814.050 480.450 814.950 ;
        RECT 475.950 812.250 477.750 813.150 ;
        RECT 478.950 811.950 481.050 814.050 ;
        RECT 482.250 812.250 484.050 813.150 ;
        RECT 485.400 811.050 486.450 814.950 ;
        RECT 475.950 808.950 478.050 811.050 ;
        RECT 479.250 809.850 480.750 810.750 ;
        RECT 481.950 808.950 484.050 811.050 ;
        RECT 484.950 808.950 487.050 811.050 ;
        RECT 476.400 808.050 477.450 808.950 ;
        RECT 475.950 805.950 478.050 808.050 ;
        RECT 482.400 805.050 483.450 808.950 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 472.950 778.950 475.050 781.050 ;
        RECT 472.950 774.450 475.050 775.050 ;
        RECT 470.400 773.400 475.050 774.450 ;
        RECT 466.950 769.950 469.050 772.050 ;
        RECT 470.400 769.050 471.450 773.400 ;
        RECT 472.950 772.950 475.050 773.400 ;
        RECT 478.950 772.950 481.050 775.050 ;
        RECT 472.950 770.850 475.050 771.750 ;
        RECT 475.950 770.250 478.050 771.150 ;
        RECT 469.950 766.950 472.050 769.050 ;
        RECT 475.950 768.450 478.050 769.050 ;
        RECT 479.400 768.450 480.450 772.950 ;
        RECT 475.950 767.400 480.450 768.450 ;
        RECT 475.950 766.950 478.050 767.400 ;
        RECT 470.400 748.050 471.450 766.950 ;
        RECT 484.950 763.950 487.050 766.050 ;
        RECT 485.400 748.050 486.450 763.950 ;
        RECT 488.400 748.050 489.450 838.950 ;
        RECT 500.400 838.050 501.450 841.950 ;
        RECT 503.400 841.050 504.450 883.950 ;
        RECT 512.400 862.050 513.450 883.950 ;
        RECT 521.400 865.050 522.450 890.400 ;
        RECT 523.950 889.950 526.050 890.400 ;
        RECT 550.950 889.950 553.050 892.050 ;
        RECT 568.950 891.450 571.050 892.050 ;
        RECT 568.950 890.400 573.450 891.450 ;
        RECT 568.950 889.950 571.050 890.400 ;
        RECT 523.950 887.850 526.050 888.750 ;
        RECT 544.950 888.450 547.050 889.050 ;
        RECT 526.950 887.250 529.050 888.150 ;
        RECT 542.400 887.400 547.050 888.450 ;
        RECT 526.950 883.950 529.050 886.050 ;
        RECT 520.950 862.950 523.050 865.050 ;
        RECT 511.950 859.950 514.050 862.050 ;
        RECT 538.950 859.950 541.050 862.050 ;
        RECT 532.950 850.950 535.050 853.050 ;
        RECT 533.400 850.050 534.450 850.950 ;
        RECT 526.950 847.950 529.050 850.050 ;
        RECT 532.950 847.950 535.050 850.050 ;
        RECT 527.400 847.050 528.450 847.950 ;
        RECT 533.400 847.050 534.450 847.950 ;
        RECT 505.950 844.950 508.050 847.050 ;
        RECT 523.950 845.250 525.750 846.150 ;
        RECT 526.950 844.950 529.050 847.050 ;
        RECT 530.250 845.250 531.750 846.150 ;
        RECT 532.950 844.950 535.050 847.050 ;
        RECT 536.250 845.250 538.050 846.150 ;
        RECT 539.400 844.050 540.450 859.950 ;
        RECT 542.400 859.050 543.450 887.400 ;
        RECT 544.950 886.950 547.050 887.400 ;
        RECT 548.250 887.250 550.050 888.150 ;
        RECT 550.950 887.850 553.050 888.750 ;
        RECT 553.950 887.250 556.050 888.150 ;
        RECT 565.950 887.250 568.050 888.150 ;
        RECT 568.950 887.850 571.050 888.750 ;
        RECT 544.950 884.850 546.750 885.750 ;
        RECT 547.950 883.950 550.050 886.050 ;
        RECT 553.950 883.950 556.050 886.050 ;
        RECT 565.950 883.950 568.050 886.050 ;
        RECT 554.400 883.050 555.450 883.950 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 572.400 880.050 573.450 890.400 ;
        RECT 574.950 889.950 577.050 892.050 ;
        RECT 580.950 889.950 583.050 892.050 ;
        RECT 586.950 889.950 589.050 892.050 ;
        RECT 598.950 889.950 601.050 892.050 ;
        RECT 607.950 889.950 610.050 892.050 ;
        RECT 613.950 889.950 616.050 892.050 ;
        RECT 637.950 889.950 640.050 892.050 ;
        RECT 575.400 888.450 576.450 889.950 ;
        RECT 577.950 888.450 580.050 889.050 ;
        RECT 575.400 887.400 580.050 888.450 ;
        RECT 581.250 887.850 582.750 888.750 ;
        RECT 583.950 888.450 586.050 889.050 ;
        RECT 587.400 888.450 588.450 889.950 ;
        RECT 575.400 886.050 576.450 887.400 ;
        RECT 577.950 886.950 580.050 887.400 ;
        RECT 583.950 887.400 588.450 888.450 ;
        RECT 598.950 887.850 601.050 888.750 ;
        RECT 583.950 886.950 586.050 887.400 ;
        RECT 574.950 883.950 577.050 886.050 ;
        RECT 577.950 884.850 580.050 885.750 ;
        RECT 583.950 884.850 586.050 885.750 ;
        RECT 587.400 883.050 588.450 887.400 ;
        RECT 601.950 887.250 604.050 888.150 ;
        RECT 601.950 883.950 604.050 886.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 571.950 877.950 574.050 880.050 ;
        RECT 565.950 862.950 568.050 865.050 ;
        RECT 541.950 856.950 544.050 859.050 ;
        RECT 566.400 850.050 567.450 862.950 ;
        RECT 574.950 853.950 577.050 856.050 ;
        RECT 568.950 850.950 571.050 853.050 ;
        RECT 569.400 850.050 570.450 850.950 ;
        RECT 575.400 850.050 576.450 853.950 ;
        RECT 553.950 848.250 556.050 849.150 ;
        RECT 562.950 847.950 565.050 850.050 ;
        RECT 565.950 847.950 568.050 850.050 ;
        RECT 568.950 847.950 571.050 850.050 ;
        RECT 572.250 848.250 573.750 849.150 ;
        RECT 574.950 847.950 577.050 850.050 ;
        RECT 541.950 844.950 544.050 847.050 ;
        RECT 544.950 845.250 546.750 846.150 ;
        RECT 547.950 844.950 550.050 847.050 ;
        RECT 551.250 845.250 552.750 846.150 ;
        RECT 553.950 844.950 556.050 847.050 ;
        RECT 505.950 842.850 508.050 843.750 ;
        RECT 523.950 841.950 526.050 844.050 ;
        RECT 527.250 842.850 528.750 843.750 ;
        RECT 529.950 841.950 532.050 844.050 ;
        RECT 533.250 842.850 534.750 843.750 ;
        RECT 535.950 841.950 538.050 844.050 ;
        RECT 538.950 841.950 541.050 844.050 ;
        RECT 530.400 841.050 531.450 841.950 ;
        RECT 502.950 838.950 505.050 841.050 ;
        RECT 529.950 838.950 532.050 841.050 ;
        RECT 542.400 838.050 543.450 844.950 ;
        RECT 544.950 841.950 547.050 844.050 ;
        RECT 548.250 842.850 549.750 843.750 ;
        RECT 550.950 841.950 553.050 844.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 493.950 823.950 496.050 826.050 ;
        RECT 494.400 814.050 495.450 823.950 ;
        RECT 490.950 812.250 492.750 813.150 ;
        RECT 493.950 811.950 496.050 814.050 ;
        RECT 497.250 812.250 499.050 813.150 ;
        RECT 490.950 808.950 493.050 811.050 ;
        RECT 494.250 809.850 495.750 810.750 ;
        RECT 496.950 808.950 499.050 811.050 ;
        RECT 500.400 775.050 501.450 835.950 ;
        RECT 520.950 823.950 523.050 826.050 ;
        RECT 521.400 817.050 522.450 823.950 ;
        RECT 542.400 820.050 543.450 835.950 ;
        RECT 541.950 817.950 544.050 820.050 ;
        RECT 514.950 814.950 517.050 817.050 ;
        RECT 518.250 815.250 519.750 816.150 ;
        RECT 520.950 814.950 523.050 817.050 ;
        RECT 532.950 814.950 535.050 817.050 ;
        RECT 538.950 814.950 541.050 817.050 ;
        RECT 511.950 811.950 514.050 814.050 ;
        RECT 515.250 812.850 516.750 813.750 ;
        RECT 517.950 811.950 520.050 814.050 ;
        RECT 521.250 812.850 523.050 813.750 ;
        RECT 511.950 809.850 514.050 810.750 ;
        RECT 518.400 778.050 519.450 811.950 ;
        RECT 533.400 808.050 534.450 814.950 ;
        RECT 539.400 814.050 540.450 814.950 ;
        RECT 535.950 812.250 537.750 813.150 ;
        RECT 538.950 811.950 541.050 814.050 ;
        RECT 542.250 812.250 544.050 813.150 ;
        RECT 553.950 812.250 555.750 813.150 ;
        RECT 556.950 811.950 559.050 814.050 ;
        RECT 560.250 812.250 562.050 813.150 ;
        RECT 535.950 808.950 538.050 811.050 ;
        RECT 539.250 809.850 540.750 810.750 ;
        RECT 541.950 808.950 544.050 811.050 ;
        RECT 553.950 808.950 556.050 811.050 ;
        RECT 557.250 809.850 558.750 810.750 ;
        RECT 559.950 808.950 562.050 811.050 ;
        RECT 532.950 805.950 535.050 808.050 ;
        RECT 536.400 796.050 537.450 808.950 ;
        RECT 542.400 801.450 543.450 808.950 ;
        RECT 539.400 800.400 543.450 801.450 ;
        RECT 535.950 793.950 538.050 796.050 ;
        RECT 529.950 787.950 532.050 790.050 ;
        RECT 517.950 775.950 520.050 778.050 ;
        RECT 530.400 775.050 531.450 787.950 ;
        RECT 490.950 772.950 493.050 775.050 ;
        RECT 496.950 773.250 499.050 774.150 ;
        RECT 499.950 772.950 502.050 775.050 ;
        RECT 514.950 772.950 517.050 775.050 ;
        RECT 529.950 772.950 532.050 775.050 ;
        RECT 539.400 772.050 540.450 800.400 ;
        RECT 554.400 790.050 555.450 808.950 ;
        RECT 560.400 805.050 561.450 808.950 ;
        RECT 563.400 805.050 564.450 847.950 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 544.950 787.950 547.050 790.050 ;
        RECT 553.950 787.950 556.050 790.050 ;
        RECT 541.950 783.300 544.050 785.400 ;
        RECT 542.550 779.700 543.750 783.300 ;
        RECT 541.950 777.600 544.050 779.700 ;
        RECT 490.950 770.850 493.050 771.750 ;
        RECT 496.950 769.950 499.050 772.050 ;
        RECT 500.250 770.250 502.050 771.150 ;
        RECT 514.950 770.850 517.050 771.750 ;
        RECT 517.950 770.250 520.050 771.150 ;
        RECT 529.950 770.850 532.050 771.750 ;
        RECT 538.950 771.450 541.050 772.050 ;
        RECT 532.950 770.250 535.050 771.150 ;
        RECT 536.400 770.400 541.050 771.450 ;
        RECT 499.950 766.950 502.050 769.050 ;
        RECT 517.950 768.450 520.050 769.050 ;
        RECT 532.950 768.450 535.050 769.050 ;
        RECT 536.400 768.450 537.450 770.400 ;
        RECT 538.950 769.950 541.050 770.400 ;
        RECT 517.950 767.400 522.450 768.450 ;
        RECT 517.950 766.950 520.050 767.400 ;
        RECT 469.950 745.950 472.050 748.050 ;
        RECT 484.950 745.950 487.050 748.050 ;
        RECT 487.950 745.950 490.050 748.050 ;
        RECT 463.950 742.950 466.050 745.050 ;
        RECT 467.250 743.250 469.050 744.150 ;
        RECT 469.950 743.850 472.050 744.750 ;
        RECT 472.950 743.250 475.050 744.150 ;
        RECT 481.950 743.250 484.050 744.150 ;
        RECT 484.950 743.850 487.050 744.750 ;
        RECT 490.950 744.450 493.050 745.050 ;
        RECT 487.950 743.250 489.750 744.150 ;
        RECT 490.950 743.400 495.450 744.450 ;
        RECT 490.950 742.950 493.050 743.400 ;
        RECT 463.950 740.850 465.750 741.750 ;
        RECT 466.950 739.950 469.050 742.050 ;
        RECT 472.950 739.950 475.050 742.050 ;
        RECT 481.950 739.950 484.050 742.050 ;
        RECT 487.950 739.950 490.050 742.050 ;
        RECT 491.250 740.850 493.050 741.750 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 464.400 703.050 465.450 724.950 ;
        RECT 463.950 700.950 466.050 703.050 ;
        RECT 467.400 700.050 468.450 739.950 ;
        RECT 473.400 739.050 474.450 739.950 ;
        RECT 472.950 736.950 475.050 739.050 ;
        RECT 469.950 704.250 472.050 705.150 ;
        RECT 469.950 700.950 472.050 703.050 ;
        RECT 473.250 701.250 474.750 702.150 ;
        RECT 475.950 700.950 478.050 703.050 ;
        RECT 479.250 701.250 481.050 702.150 ;
        RECT 466.950 697.950 469.050 700.050 ;
        RECT 470.400 691.050 471.450 700.950 ;
        RECT 472.950 697.950 475.050 700.050 ;
        RECT 476.250 698.850 477.750 699.750 ;
        RECT 478.950 697.950 481.050 700.050 ;
        RECT 469.950 688.950 472.050 691.050 ;
        RECT 479.400 685.050 480.450 697.950 ;
        RECT 478.950 682.950 481.050 685.050 ;
        RECT 482.400 679.050 483.450 739.950 ;
        RECT 488.400 739.050 489.450 739.950 ;
        RECT 487.950 736.950 490.050 739.050 ;
        RECT 490.950 736.950 493.050 739.050 ;
        RECT 491.400 735.450 492.450 736.950 ;
        RECT 488.400 734.400 492.450 735.450 ;
        RECT 488.400 700.050 489.450 734.400 ;
        RECT 494.400 730.050 495.450 743.400 ;
        RECT 496.950 742.950 499.050 745.050 ;
        RECT 497.400 736.050 498.450 742.950 ;
        RECT 500.400 738.450 501.450 766.950 ;
        RECT 508.950 745.950 511.050 748.050 ;
        RECT 509.400 745.050 510.450 745.950 ;
        RECT 502.950 742.950 505.050 745.050 ;
        RECT 506.250 743.250 507.750 744.150 ;
        RECT 508.950 742.950 511.050 745.050 ;
        RECT 502.950 740.850 504.750 741.750 ;
        RECT 505.950 739.950 508.050 742.050 ;
        RECT 509.250 740.850 510.750 741.750 ;
        RECT 511.950 739.950 514.050 742.050 ;
        RECT 500.400 737.400 504.450 738.450 ;
        RECT 496.950 733.950 499.050 736.050 ;
        RECT 493.950 727.950 496.050 730.050 ;
        RECT 494.400 705.450 495.450 727.950 ;
        RECT 503.400 724.050 504.450 737.400 ;
        RECT 506.400 733.050 507.450 739.950 ;
        RECT 511.950 737.850 514.050 738.750 ;
        RECT 505.950 730.950 508.050 733.050 ;
        RECT 502.950 721.950 505.050 724.050 ;
        RECT 490.950 704.250 493.050 705.150 ;
        RECT 494.400 704.400 498.450 705.450 ;
        RECT 497.400 703.050 498.450 704.400 ;
        RECT 490.950 700.950 493.050 703.050 ;
        RECT 494.250 701.250 495.750 702.150 ;
        RECT 496.950 700.950 499.050 703.050 ;
        RECT 500.250 701.250 502.050 702.150 ;
        RECT 487.950 697.950 490.050 700.050 ;
        RECT 491.400 697.050 492.450 700.950 ;
        RECT 493.950 697.950 496.050 700.050 ;
        RECT 497.250 698.850 498.750 699.750 ;
        RECT 499.950 699.450 502.050 700.050 ;
        RECT 503.400 699.450 504.450 721.950 ;
        RECT 508.950 706.950 511.050 709.050 ;
        RECT 499.950 698.400 504.450 699.450 ;
        RECT 509.400 699.450 510.450 706.950 ;
        RECT 511.950 701.250 514.050 702.150 ;
        RECT 517.950 701.250 520.050 702.150 ;
        RECT 511.950 699.450 514.050 700.050 ;
        RECT 509.400 698.400 514.050 699.450 ;
        RECT 499.950 697.950 502.050 698.400 ;
        RECT 490.950 694.950 493.050 697.050 ;
        RECT 496.950 694.950 499.050 697.050 ;
        RECT 458.400 677.400 462.450 678.450 ;
        RECT 445.950 670.950 448.050 673.050 ;
        RECT 449.250 671.250 450.750 672.150 ;
        RECT 451.950 670.950 454.050 673.050 ;
        RECT 442.950 667.950 445.050 670.050 ;
        RECT 446.250 668.850 447.750 669.750 ;
        RECT 448.950 667.950 451.050 670.050 ;
        RECT 452.250 668.850 454.050 669.750 ;
        RECT 442.950 665.850 445.050 666.750 ;
        RECT 449.400 666.450 450.450 667.950 ;
        RECT 449.400 665.400 453.450 666.450 ;
        RECT 439.950 661.950 442.050 664.050 ;
        RECT 442.950 633.450 445.050 634.050 ;
        RECT 440.400 632.400 445.050 633.450 ;
        RECT 440.400 625.050 441.450 632.400 ;
        RECT 442.950 631.950 445.050 632.400 ;
        RECT 446.250 632.250 447.750 633.150 ;
        RECT 448.950 631.950 451.050 634.050 ;
        RECT 442.950 629.850 444.750 630.750 ;
        RECT 445.950 628.950 448.050 631.050 ;
        RECT 449.250 629.850 451.050 630.750 ;
        RECT 439.950 622.950 442.050 625.050 ;
        RECT 452.400 622.050 453.450 665.400 ;
        RECT 451.950 619.950 454.050 622.050 ;
        RECT 458.400 613.050 459.450 677.400 ;
        RECT 481.950 676.950 484.050 679.050 ;
        RECT 466.950 673.950 469.050 676.050 ;
        RECT 487.950 673.950 490.050 676.050 ;
        RECT 460.950 672.450 463.050 673.050 ;
        RECT 463.950 672.450 466.050 673.050 ;
        RECT 460.950 671.400 466.050 672.450 ;
        RECT 467.250 671.850 468.750 672.750 ;
        RECT 460.950 670.950 463.050 671.400 ;
        RECT 463.950 670.950 466.050 671.400 ;
        RECT 469.950 670.950 472.050 673.050 ;
        RECT 457.950 610.950 460.050 613.050 ;
        RECT 442.950 605.400 445.050 607.500 ;
        RECT 443.400 588.600 444.600 605.400 ;
        RECT 448.950 604.950 451.050 607.050 ;
        RECT 449.400 601.050 450.450 604.950 ;
        RECT 445.950 598.950 448.050 601.050 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 454.950 598.950 457.050 601.050 ;
        RECT 442.950 586.500 445.050 588.600 ;
        RECT 430.950 538.950 433.050 541.050 ;
        RECT 436.950 538.950 439.050 541.050 ;
        RECT 430.950 533.400 433.050 535.500 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 409.950 487.950 412.050 490.050 ;
        RECT 413.250 488.250 414.750 489.150 ;
        RECT 421.950 487.950 424.050 490.050 ;
        RECT 409.950 485.850 411.750 486.750 ;
        RECT 412.950 484.950 415.050 487.050 ;
        RECT 416.250 485.850 418.050 486.750 ;
        RECT 428.400 484.050 429.450 523.950 ;
        RECT 431.400 516.600 432.600 533.400 ;
        RECT 446.400 532.050 447.450 598.950 ;
        RECT 448.950 596.850 451.050 597.750 ;
        RECT 454.950 596.850 457.050 597.750 ;
        RECT 451.950 557.250 454.050 558.150 ;
        RECT 457.950 557.250 460.050 558.150 ;
        RECT 451.950 553.950 454.050 556.050 ;
        RECT 457.950 553.950 460.050 556.050 ;
        RECT 458.400 550.050 459.450 553.950 ;
        RECT 457.950 547.950 460.050 550.050 ;
        RECT 457.950 538.950 460.050 541.050 ;
        RECT 451.950 533.400 454.050 535.500 ;
        RECT 445.950 529.950 448.050 532.050 ;
        RECT 436.950 526.950 439.050 529.050 ;
        RECT 442.950 528.450 445.050 529.050 ;
        RECT 446.400 528.450 447.450 529.950 ;
        RECT 442.950 527.400 447.450 528.450 ;
        RECT 442.950 526.950 445.050 527.400 ;
        RECT 436.950 524.850 439.050 525.750 ;
        RECT 442.950 524.850 445.050 525.750 ;
        RECT 442.950 520.950 445.050 523.050 ;
        RECT 430.950 514.500 433.050 516.600 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 430.950 488.250 433.050 489.150 ;
        RECT 437.400 487.050 438.450 490.950 ;
        RECT 430.950 484.950 433.050 487.050 ;
        RECT 434.250 485.250 435.750 486.150 ;
        RECT 436.950 484.950 439.050 487.050 ;
        RECT 440.250 485.250 442.050 486.150 ;
        RECT 412.950 481.950 415.050 484.050 ;
        RECT 427.950 481.950 430.050 484.050 ;
        RECT 433.950 481.950 436.050 484.050 ;
        RECT 437.250 482.850 438.750 483.750 ;
        RECT 439.950 481.950 442.050 484.050 ;
        RECT 400.950 478.950 403.050 481.050 ;
        RECT 406.950 478.950 409.050 481.050 ;
        RECT 400.950 451.950 403.050 454.050 ;
        RECT 406.950 451.950 409.050 454.050 ;
        RECT 410.250 452.250 412.050 453.150 ;
        RECT 413.400 451.050 414.450 481.950 ;
        RECT 433.950 478.950 436.050 481.050 ;
        RECT 418.950 469.950 421.050 472.050 ;
        RECT 419.400 460.050 420.450 469.950 ;
        RECT 418.950 457.950 421.050 460.050 ;
        RECT 430.950 457.950 433.050 460.050 ;
        RECT 394.950 448.950 397.050 451.050 ;
        RECT 400.950 449.850 402.750 450.750 ;
        RECT 403.950 448.950 406.050 451.050 ;
        RECT 407.250 449.850 408.750 450.750 ;
        RECT 409.950 448.950 412.050 451.050 ;
        RECT 412.950 448.950 415.050 451.050 ;
        RECT 419.400 450.450 420.450 457.950 ;
        RECT 431.400 457.050 432.450 457.950 ;
        RECT 430.950 454.950 433.050 457.050 ;
        RECT 421.950 452.250 423.750 453.150 ;
        RECT 424.950 451.950 427.050 454.050 ;
        RECT 428.250 452.250 430.050 453.150 ;
        RECT 421.950 450.450 424.050 451.050 ;
        RECT 419.400 449.400 424.050 450.450 ;
        RECT 425.250 449.850 426.750 450.750 ;
        RECT 427.950 450.450 430.050 451.050 ;
        RECT 431.400 450.450 432.450 454.950 ;
        RECT 421.950 448.950 424.050 449.400 ;
        RECT 427.950 449.400 432.450 450.450 ;
        RECT 427.950 448.950 430.050 449.400 ;
        RECT 403.950 446.850 406.050 447.750 ;
        RECT 410.400 421.050 411.450 448.950 ;
        RECT 434.400 447.450 435.450 478.950 ;
        RECT 440.400 460.050 441.450 481.950 ;
        RECT 439.950 457.950 442.050 460.050 ;
        RECT 443.400 456.450 444.450 520.950 ;
        RECT 446.400 478.050 447.450 527.400 ;
        RECT 452.250 521.400 453.450 533.400 ;
        RECT 454.950 530.250 457.050 531.150 ;
        RECT 454.950 526.950 457.050 529.050 ;
        RECT 455.400 523.050 456.450 526.950 ;
        RECT 451.950 519.300 454.050 521.400 ;
        RECT 454.950 520.950 457.050 523.050 ;
        RECT 452.250 515.700 453.450 519.300 ;
        RECT 451.950 513.600 454.050 515.700 ;
        RECT 451.950 486.450 454.050 487.050 ;
        RECT 449.400 485.400 454.050 486.450 ;
        RECT 449.400 484.050 450.450 485.400 ;
        RECT 451.950 484.950 454.050 485.400 ;
        RECT 448.950 481.950 451.050 484.050 ;
        RECT 451.950 482.850 454.050 483.750 ;
        RECT 454.950 482.250 457.050 483.150 ;
        RECT 454.950 478.950 457.050 481.050 ;
        RECT 445.950 475.950 448.050 478.050 ;
        RECT 451.950 457.950 454.050 460.050 ;
        RECT 440.400 455.400 444.450 456.450 ;
        RECT 440.400 450.450 441.450 455.400 ;
        RECT 442.950 452.250 444.750 453.150 ;
        RECT 445.950 451.950 448.050 454.050 ;
        RECT 449.250 452.250 451.050 453.150 ;
        RECT 442.950 450.450 445.050 451.050 ;
        RECT 440.400 449.400 445.050 450.450 ;
        RECT 446.250 449.850 447.750 450.750 ;
        RECT 442.950 448.950 445.050 449.400 ;
        RECT 448.950 448.950 451.050 451.050 ;
        RECT 431.400 446.400 435.450 447.450 ;
        RECT 412.950 442.950 415.050 445.050 ;
        RECT 409.950 418.950 412.050 421.050 ;
        RECT 397.950 415.950 400.050 418.050 ;
        RECT 403.950 417.450 406.050 418.050 ;
        RECT 401.250 416.250 402.750 417.150 ;
        RECT 403.950 416.400 408.450 417.450 ;
        RECT 403.950 415.950 406.050 416.400 ;
        RECT 397.950 413.850 399.750 414.750 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 404.250 413.850 406.050 414.750 ;
        RECT 376.950 406.950 379.050 409.050 ;
        RECT 391.950 406.950 394.050 409.050 ;
        RECT 367.950 343.950 370.050 346.050 ;
        RECT 373.950 343.950 376.050 346.050 ;
        RECT 361.950 340.950 364.050 343.050 ;
        RECT 364.950 341.250 367.050 342.150 ;
        RECT 362.400 316.050 363.450 340.950 ;
        RECT 368.400 339.450 369.450 343.950 ;
        RECT 370.950 341.250 373.050 342.150 ;
        RECT 377.400 340.050 378.450 406.950 ;
        RECT 401.400 406.050 402.450 412.950 ;
        RECT 407.400 406.050 408.450 416.400 ;
        RECT 409.950 415.950 412.050 418.050 ;
        RECT 410.400 412.050 411.450 415.950 ;
        RECT 409.950 409.950 412.050 412.050 ;
        RECT 413.400 411.450 414.450 442.950 ;
        RECT 415.950 415.950 418.050 418.050 ;
        RECT 421.950 417.450 424.050 418.050 ;
        RECT 419.250 416.250 420.750 417.150 ;
        RECT 421.950 416.400 426.450 417.450 ;
        RECT 421.950 415.950 424.050 416.400 ;
        RECT 415.950 413.850 417.750 414.750 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 422.250 413.850 424.050 414.750 ;
        RECT 413.400 410.400 417.450 411.450 ;
        RECT 400.950 403.950 403.050 406.050 ;
        RECT 406.950 403.950 409.050 406.050 ;
        RECT 406.950 385.950 409.050 388.050 ;
        RECT 407.400 385.050 408.450 385.950 ;
        RECT 382.950 384.450 385.050 385.050 ;
        RECT 391.950 384.450 394.050 385.050 ;
        RECT 379.950 383.250 381.750 384.150 ;
        RECT 382.950 383.400 387.450 384.450 ;
        RECT 382.950 382.950 385.050 383.400 ;
        RECT 379.950 379.950 382.050 382.050 ;
        RECT 383.250 380.850 385.050 381.750 ;
        RECT 386.400 367.050 387.450 383.400 ;
        RECT 388.950 383.250 390.750 384.150 ;
        RECT 391.950 383.400 396.450 384.450 ;
        RECT 391.950 382.950 394.050 383.400 ;
        RECT 388.950 379.950 391.050 382.050 ;
        RECT 392.250 380.850 394.050 381.750 ;
        RECT 385.950 364.950 388.050 367.050 ;
        RECT 385.950 346.950 388.050 349.050 ;
        RECT 379.950 340.950 382.050 343.050 ;
        RECT 382.950 341.250 385.050 342.150 ;
        RECT 370.950 339.450 373.050 340.050 ;
        RECT 368.400 338.400 373.050 339.450 ;
        RECT 370.950 337.950 373.050 338.400 ;
        RECT 376.950 337.950 379.050 340.050 ;
        RECT 380.400 334.050 381.450 340.950 ;
        RECT 382.950 337.950 385.050 340.050 ;
        RECT 386.400 339.450 387.450 346.950 ;
        RECT 389.400 345.450 390.450 379.950 ;
        RECT 395.400 373.050 396.450 383.400 ;
        RECT 406.950 382.950 409.050 385.050 ;
        RECT 410.400 384.450 411.450 409.950 ;
        RECT 412.950 384.450 415.050 385.050 ;
        RECT 410.400 383.400 415.050 384.450 ;
        RECT 410.400 382.050 411.450 383.400 ;
        RECT 412.950 382.950 415.050 383.400 ;
        RECT 406.950 380.850 409.050 381.750 ;
        RECT 409.950 379.950 412.050 382.050 ;
        RECT 412.950 380.850 415.050 381.750 ;
        RECT 394.950 370.950 397.050 373.050 ;
        RECT 412.950 364.950 415.050 367.050 ;
        RECT 394.950 352.950 397.050 355.050 ;
        RECT 389.400 344.400 393.450 345.450 ;
        RECT 388.950 341.250 391.050 342.150 ;
        RECT 388.950 339.450 391.050 340.050 ;
        RECT 386.400 338.400 391.050 339.450 ;
        RECT 388.950 337.950 391.050 338.400 ;
        RECT 379.950 331.950 382.050 334.050 ;
        RECT 383.400 325.050 384.450 337.950 ;
        RECT 373.950 322.950 376.050 325.050 ;
        RECT 382.950 322.950 385.050 325.050 ;
        RECT 361.950 313.950 364.050 316.050 ;
        RECT 361.950 311.850 364.050 312.750 ;
        RECT 364.950 311.250 367.050 312.150 ;
        RECT 364.950 307.950 367.050 310.050 ;
        RECT 365.400 307.050 366.450 307.950 ;
        RECT 364.950 304.950 367.050 307.050 ;
        RECT 340.950 301.950 343.050 304.050 ;
        RECT 358.950 301.950 361.050 304.050 ;
        RECT 331.950 271.950 334.050 274.050 ;
        RECT 341.400 271.050 342.450 301.950 ;
        RECT 370.950 274.950 373.050 277.050 ;
        RECT 331.950 270.450 334.050 271.050 ;
        RECT 329.400 269.400 334.050 270.450 ;
        RECT 331.950 268.950 334.050 269.400 ;
        RECT 335.250 269.250 337.050 270.150 ;
        RECT 340.950 268.950 343.050 271.050 ;
        RECT 344.250 269.250 346.050 270.150 ;
        RECT 361.950 269.250 364.050 270.150 ;
        RECT 367.950 269.250 370.050 270.150 ;
        RECT 313.950 265.950 316.050 268.050 ;
        RECT 317.250 266.850 319.050 267.750 ;
        RECT 319.950 266.250 322.050 267.150 ;
        RECT 322.950 266.850 325.050 267.750 ;
        RECT 331.950 266.850 333.750 267.750 ;
        RECT 334.950 265.950 337.050 268.050 ;
        RECT 340.950 266.850 342.750 267.750 ;
        RECT 343.950 265.950 346.050 268.050 ;
        RECT 361.950 265.950 364.050 268.050 ;
        RECT 367.950 267.450 370.050 268.050 ;
        RECT 371.400 267.450 372.450 274.950 ;
        RECT 374.400 268.050 375.450 322.950 ;
        RECT 382.950 310.950 385.050 313.050 ;
        RECT 388.950 310.950 391.050 313.050 ;
        RECT 383.400 310.050 384.450 310.950 ;
        RECT 379.950 308.250 381.750 309.150 ;
        RECT 382.950 307.950 385.050 310.050 ;
        RECT 386.250 308.250 388.050 309.150 ;
        RECT 389.400 307.050 390.450 310.950 ;
        RECT 379.950 304.950 382.050 307.050 ;
        RECT 383.250 305.850 384.750 306.750 ;
        RECT 385.950 304.950 388.050 307.050 ;
        RECT 388.950 304.950 391.050 307.050 ;
        RECT 380.400 283.050 381.450 304.950 ;
        RECT 386.400 292.050 387.450 304.950 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 379.950 280.950 382.050 283.050 ;
        RECT 392.400 274.050 393.450 344.400 ;
        RECT 395.400 313.050 396.450 352.950 ;
        RECT 400.950 340.950 403.050 343.050 ;
        RECT 406.950 340.950 409.050 343.050 ;
        RECT 410.250 341.250 412.050 342.150 ;
        RECT 400.950 338.850 403.050 339.750 ;
        RECT 403.950 338.250 406.050 339.150 ;
        RECT 406.950 338.850 408.750 339.750 ;
        RECT 409.950 339.450 412.050 340.050 ;
        RECT 413.400 339.450 414.450 364.950 ;
        RECT 409.950 338.400 414.450 339.450 ;
        RECT 409.950 337.950 412.050 338.400 ;
        RECT 416.400 337.050 417.450 410.400 ;
        RECT 425.400 403.050 426.450 416.400 ;
        RECT 424.950 400.950 427.050 403.050 ;
        RECT 418.950 385.950 421.050 388.050 ;
        RECT 421.950 385.950 424.050 388.050 ;
        RECT 427.950 385.950 430.050 388.050 ;
        RECT 403.950 334.950 406.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 404.400 322.050 405.450 334.950 ;
        RECT 415.950 331.950 418.050 334.050 ;
        RECT 403.950 319.950 406.050 322.050 ;
        RECT 394.950 310.950 397.050 313.050 ;
        RECT 394.950 308.250 396.750 309.150 ;
        RECT 397.950 307.950 400.050 310.050 ;
        RECT 401.250 308.250 403.050 309.150 ;
        RECT 394.950 304.950 397.050 307.050 ;
        RECT 398.250 305.850 399.750 306.750 ;
        RECT 400.950 304.950 403.050 307.050 ;
        RECT 394.950 301.950 397.050 304.050 ;
        RECT 391.950 271.950 394.050 274.050 ;
        RECT 395.400 271.050 396.450 301.950 ;
        RECT 401.400 301.050 402.450 304.950 ;
        RECT 404.400 304.050 405.450 319.950 ;
        RECT 416.400 310.050 417.450 331.950 ;
        RECT 419.400 331.050 420.450 385.950 ;
        RECT 422.400 370.050 423.450 385.950 ;
        RECT 428.400 385.050 429.450 385.950 ;
        RECT 424.950 383.250 426.750 384.150 ;
        RECT 427.950 382.950 430.050 385.050 ;
        RECT 424.950 379.950 427.050 382.050 ;
        RECT 428.250 380.850 430.050 381.750 ;
        RECT 421.950 367.950 424.050 370.050 ;
        RECT 431.400 367.050 432.450 446.400 ;
        RECT 443.400 439.050 444.450 448.950 ;
        RECT 442.950 436.950 445.050 439.050 ;
        RECT 442.950 421.950 445.050 424.050 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 440.250 413.250 442.050 414.150 ;
        RECT 436.950 410.850 438.750 411.750 ;
        RECT 439.950 411.450 442.050 412.050 ;
        RECT 443.400 411.450 444.450 421.950 ;
        RECT 445.950 415.950 448.050 418.050 ;
        RECT 446.400 415.050 447.450 415.950 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 449.250 413.250 451.050 414.150 ;
        RECT 452.400 412.050 453.450 457.950 ;
        RECT 458.400 445.050 459.450 538.950 ;
        RECT 461.400 484.050 462.450 670.950 ;
        RECT 488.400 670.050 489.450 673.950 ;
        RECT 493.950 670.950 496.050 673.050 ;
        RECT 463.950 668.850 466.050 669.750 ;
        RECT 469.950 668.850 472.050 669.750 ;
        RECT 484.950 668.250 486.750 669.150 ;
        RECT 487.950 667.950 490.050 670.050 ;
        RECT 491.250 668.250 493.050 669.150 ;
        RECT 484.950 664.950 487.050 667.050 ;
        RECT 488.250 665.850 489.750 666.750 ;
        RECT 490.950 666.450 493.050 667.050 ;
        RECT 494.400 666.450 495.450 670.950 ;
        RECT 497.400 667.050 498.450 694.950 ;
        RECT 503.400 670.050 504.450 698.400 ;
        RECT 511.950 697.950 514.050 698.400 ;
        RECT 515.250 698.250 516.750 699.150 ;
        RECT 517.950 697.950 520.050 700.050 ;
        RECT 514.950 694.950 517.050 697.050 ;
        RECT 518.400 685.050 519.450 697.950 ;
        RECT 521.400 697.050 522.450 767.400 ;
        RECT 532.950 767.400 537.450 768.450 ;
        RECT 538.950 767.850 541.050 768.750 ;
        RECT 532.950 766.950 535.050 767.400 ;
        RECT 542.550 765.600 543.750 777.600 ;
        RECT 541.950 763.500 544.050 765.600 ;
        RECT 532.950 754.950 535.050 757.050 ;
        RECT 533.400 745.050 534.450 754.950 ;
        RECT 545.400 745.050 546.450 787.950 ;
        RECT 547.950 781.950 550.050 784.050 ;
        RECT 548.400 771.450 549.450 781.950 ;
        RECT 550.950 773.250 553.050 774.150 ;
        RECT 556.950 773.250 559.050 774.150 ;
        RECT 550.950 771.450 553.050 772.050 ;
        RECT 548.400 770.400 553.050 771.450 ;
        RECT 550.950 769.950 553.050 770.400 ;
        RECT 556.950 769.950 559.050 772.050 ;
        RECT 547.950 749.400 550.050 751.500 ;
        RECT 532.950 742.950 535.050 745.050 ;
        RECT 536.250 743.250 537.750 744.150 ;
        RECT 538.950 742.950 541.050 745.050 ;
        RECT 544.950 742.950 547.050 745.050 ;
        RECT 529.950 741.450 532.050 742.050 ;
        RECT 527.400 740.400 532.050 741.450 ;
        RECT 533.250 740.850 534.750 741.750 ;
        RECT 527.400 727.050 528.450 740.400 ;
        RECT 529.950 739.950 532.050 740.400 ;
        RECT 535.950 739.950 538.050 742.050 ;
        RECT 539.250 740.850 541.050 741.750 ;
        RECT 529.950 737.850 532.050 738.750 ;
        RECT 532.950 730.950 535.050 733.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 533.400 706.050 534.450 730.950 ;
        RECT 536.400 721.050 537.450 739.950 ;
        RECT 544.950 733.950 547.050 736.050 ;
        RECT 535.950 718.950 538.050 721.050 ;
        RECT 532.950 703.950 535.050 706.050 ;
        RECT 536.250 704.250 537.750 705.150 ;
        RECT 545.400 703.050 546.450 733.950 ;
        RECT 548.400 732.600 549.600 749.400 ;
        RECT 551.400 745.050 552.450 769.950 ;
        RECT 557.400 757.050 558.450 769.950 ;
        RECT 560.400 759.450 561.450 802.950 ;
        RECT 562.950 782.400 565.050 784.500 ;
        RECT 563.400 765.600 564.600 782.400 ;
        RECT 566.400 775.050 567.450 847.950 ;
        RECT 568.950 845.850 570.750 846.750 ;
        RECT 571.950 844.950 574.050 847.050 ;
        RECT 575.250 845.850 577.050 846.750 ;
        RECT 568.950 814.950 571.050 817.050 ;
        RECT 569.400 810.450 570.450 814.950 ;
        RECT 571.950 812.250 573.750 813.150 ;
        RECT 574.950 811.950 577.050 814.050 ;
        RECT 587.400 813.450 588.450 880.950 ;
        RECT 608.400 880.050 609.450 889.950 ;
        RECT 614.400 889.050 615.450 889.950 ;
        RECT 638.400 889.050 639.450 889.950 ;
        RECT 613.950 886.950 616.050 889.050 ;
        RECT 617.250 887.250 618.750 888.150 ;
        RECT 619.950 886.950 622.050 889.050 ;
        RECT 637.950 886.950 640.050 889.050 ;
        RECT 641.250 887.250 642.750 888.150 ;
        RECT 643.950 886.950 646.050 889.050 ;
        RECT 661.950 888.450 664.050 889.050 ;
        RECT 661.950 887.400 666.450 888.450 ;
        RECT 661.950 886.950 664.050 887.400 ;
        RECT 613.950 884.850 615.750 885.750 ;
        RECT 616.950 883.950 619.050 886.050 ;
        RECT 620.250 884.850 621.750 885.750 ;
        RECT 622.950 883.950 625.050 886.050 ;
        RECT 637.950 884.850 639.750 885.750 ;
        RECT 640.950 883.950 643.050 886.050 ;
        RECT 644.250 884.850 645.750 885.750 ;
        RECT 646.950 883.950 649.050 886.050 ;
        RECT 661.950 884.850 664.050 885.750 ;
        RECT 665.400 883.050 666.450 887.400 ;
        RECT 667.950 884.850 670.050 885.750 ;
        RECT 622.950 881.850 625.050 882.750 ;
        RECT 646.950 881.850 649.050 882.750 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 607.950 877.950 610.050 880.050 ;
        RECT 589.950 853.950 592.050 856.050 ;
        RECT 590.400 844.050 591.450 853.950 ;
        RECT 592.950 847.950 595.050 850.050 ;
        RECT 598.950 849.450 601.050 850.050 ;
        RECT 596.250 848.250 597.750 849.150 ;
        RECT 598.950 848.400 603.450 849.450 ;
        RECT 598.950 847.950 601.050 848.400 ;
        RECT 592.950 845.850 594.750 846.750 ;
        RECT 595.950 844.950 598.050 847.050 ;
        RECT 599.250 845.850 601.050 846.750 ;
        RECT 589.950 841.950 592.050 844.050 ;
        RECT 592.950 841.950 595.050 844.050 ;
        RECT 593.400 820.050 594.450 841.950 ;
        RECT 596.400 841.050 597.450 844.950 ;
        RECT 595.950 838.950 598.050 841.050 ;
        RECT 592.950 817.950 595.050 820.050 ;
        RECT 598.950 817.950 601.050 820.050 ;
        RECT 599.400 817.050 600.450 817.950 ;
        RECT 589.950 815.250 592.050 816.150 ;
        RECT 592.950 815.850 595.050 816.750 ;
        RECT 595.950 815.250 597.750 816.150 ;
        RECT 598.950 814.950 601.050 817.050 ;
        RECT 589.950 813.450 592.050 814.050 ;
        RECT 578.250 812.250 580.050 813.150 ;
        RECT 587.400 812.400 592.050 813.450 ;
        RECT 589.950 811.950 592.050 812.400 ;
        RECT 595.950 811.950 598.050 814.050 ;
        RECT 599.250 812.850 601.050 813.750 ;
        RECT 571.950 810.450 574.050 811.050 ;
        RECT 569.400 809.400 574.050 810.450 ;
        RECT 575.250 809.850 576.750 810.750 ;
        RECT 571.950 808.950 574.050 809.400 ;
        RECT 577.950 808.950 580.050 811.050 ;
        RECT 590.400 793.050 591.450 811.950 ;
        RECT 596.400 808.050 597.450 811.950 ;
        RECT 595.950 805.950 598.050 808.050 ;
        RECT 589.950 790.950 592.050 793.050 ;
        RECT 577.950 777.450 580.050 778.050 ;
        RECT 575.400 776.400 580.050 777.450 ;
        RECT 565.950 772.950 568.050 775.050 ;
        RECT 575.400 766.050 576.450 776.400 ;
        RECT 577.950 775.950 580.050 776.400 ;
        RECT 581.250 776.250 582.750 777.150 ;
        RECT 583.950 775.950 586.050 778.050 ;
        RECT 598.950 775.950 601.050 778.050 ;
        RECT 599.400 775.050 600.450 775.950 ;
        RECT 602.400 775.050 603.450 848.400 ;
        RECT 608.400 841.050 609.450 877.950 ;
        RECT 643.950 856.950 646.050 859.050 ;
        RECT 610.950 844.950 613.050 847.050 ;
        RECT 616.950 844.950 619.050 847.050 ;
        RECT 628.950 845.250 631.050 846.150 ;
        RECT 634.950 844.950 637.050 847.050 ;
        RECT 610.950 842.850 613.050 843.750 ;
        RECT 613.950 842.250 616.050 843.150 ;
        RECT 607.950 838.950 610.050 841.050 ;
        RECT 613.950 840.450 616.050 841.050 ;
        RECT 617.400 840.450 618.450 844.950 ;
        RECT 625.950 842.250 627.750 843.150 ;
        RECT 628.950 841.950 631.050 844.050 ;
        RECT 634.950 842.850 637.050 843.750 ;
        RECT 644.400 843.450 645.450 856.950 ;
        RECT 652.950 849.450 655.050 850.050 ;
        RECT 650.400 848.400 655.050 849.450 ;
        RECT 646.950 845.250 649.050 846.150 ;
        RECT 646.950 843.450 649.050 844.050 ;
        RECT 644.400 842.400 649.050 843.450 ;
        RECT 646.950 841.950 649.050 842.400 ;
        RECT 613.950 839.400 618.450 840.450 ;
        RECT 613.950 838.950 616.050 839.400 ;
        RECT 625.950 838.950 628.050 841.050 ;
        RECT 629.400 826.050 630.450 841.950 ;
        RECT 650.400 826.050 651.450 848.400 ;
        RECT 652.950 847.950 655.050 848.400 ;
        RECT 665.400 847.050 666.450 880.950 ;
        RECT 680.400 876.600 681.600 893.400 ;
        RECT 685.950 886.950 688.050 889.050 ;
        RECT 691.950 886.950 694.050 889.050 ;
        RECT 685.950 884.850 688.050 885.750 ;
        RECT 691.950 884.850 694.050 885.750 ;
        RECT 701.250 881.400 702.450 893.400 ;
        RECT 745.950 892.950 748.050 895.050 ;
        RECT 772.950 893.400 775.050 895.500 ;
        RECT 793.950 893.400 796.050 895.500 ;
        RECT 703.950 890.250 706.050 891.150 ;
        RECT 703.950 886.950 706.050 889.050 ;
        RECT 704.400 883.050 705.450 886.950 ;
        RECT 715.950 884.250 717.750 885.150 ;
        RECT 718.950 883.950 721.050 886.050 ;
        RECT 722.250 884.250 724.050 885.150 ;
        RECT 736.950 884.250 738.750 885.150 ;
        RECT 739.950 883.950 742.050 886.050 ;
        RECT 743.250 884.250 745.050 885.150 ;
        RECT 700.950 879.300 703.050 881.400 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 715.950 880.950 718.050 883.050 ;
        RECT 719.250 881.850 720.750 882.750 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 736.950 880.950 739.050 883.050 ;
        RECT 740.250 881.850 741.750 882.750 ;
        RECT 742.950 880.950 745.050 883.050 ;
        RECT 679.950 874.500 682.050 876.600 ;
        RECT 701.250 875.700 702.450 879.300 ;
        RECT 700.950 873.600 703.050 875.700 ;
        RECT 722.400 865.050 723.450 880.950 ;
        RECT 715.950 862.950 718.050 865.050 ;
        RECT 721.950 862.950 724.050 865.050 ;
        RECT 673.950 856.950 676.050 859.050 ;
        RECT 674.400 847.050 675.450 856.950 ;
        RECT 716.400 850.050 717.450 862.950 ;
        RECT 730.950 854.400 733.050 856.500 ;
        RECT 724.950 850.950 727.050 853.050 ;
        RECT 679.950 848.250 682.050 849.150 ;
        RECT 700.950 848.250 703.050 849.150 ;
        RECT 703.950 847.950 706.050 850.050 ;
        RECT 715.950 847.950 718.050 850.050 ;
        RECT 719.250 848.250 720.750 849.150 ;
        RECT 721.950 847.950 724.050 850.050 ;
        RECT 652.950 845.850 655.050 846.750 ;
        RECT 655.950 845.250 658.050 846.150 ;
        RECT 664.950 844.950 667.050 847.050 ;
        RECT 670.950 845.250 672.750 846.150 ;
        RECT 673.950 844.950 676.050 847.050 ;
        RECT 677.250 845.250 678.750 846.150 ;
        RECT 679.950 844.950 682.050 847.050 ;
        RECT 691.950 845.250 693.750 846.150 ;
        RECT 694.950 844.950 697.050 847.050 ;
        RECT 698.250 845.250 699.750 846.150 ;
        RECT 700.950 844.950 703.050 847.050 ;
        RECT 655.950 841.950 658.050 844.050 ;
        RECT 670.950 841.950 673.050 844.050 ;
        RECT 674.250 842.850 675.750 843.750 ;
        RECT 676.950 841.950 679.050 844.050 ;
        RECT 671.400 826.050 672.450 841.950 ;
        RECT 677.400 841.050 678.450 841.950 ;
        RECT 676.950 838.950 679.050 841.050 ;
        RECT 676.950 829.950 679.050 832.050 ;
        RECT 628.950 823.950 631.050 826.050 ;
        RECT 649.950 823.950 652.050 826.050 ;
        RECT 670.950 823.950 673.050 826.050 ;
        RECT 625.950 819.450 628.050 820.050 ;
        RECT 620.400 818.400 628.050 819.450 ;
        RECT 620.400 817.050 621.450 818.400 ;
        RECT 625.950 817.950 628.050 818.400 ;
        RECT 631.950 817.950 634.050 820.050 ;
        RECT 634.950 817.950 637.050 820.050 ;
        RECT 670.950 817.950 673.050 820.050 ;
        RECT 616.950 814.950 619.050 817.050 ;
        RECT 619.950 814.950 622.050 817.050 ;
        RECT 625.950 816.450 628.050 817.050 ;
        RECT 628.950 816.450 631.050 817.050 ;
        RECT 623.250 815.250 624.750 816.150 ;
        RECT 625.950 815.400 631.050 816.450 ;
        RECT 625.950 814.950 628.050 815.400 ;
        RECT 628.950 814.950 631.050 815.400 ;
        RECT 617.400 814.050 618.450 814.950 ;
        RECT 616.950 811.950 619.050 814.050 ;
        RECT 620.250 812.850 621.750 813.750 ;
        RECT 622.950 811.950 625.050 814.050 ;
        RECT 626.250 812.850 628.050 813.750 ;
        RECT 629.400 811.050 630.450 814.950 ;
        RECT 616.950 809.850 619.050 810.750 ;
        RECT 628.950 808.950 631.050 811.050 ;
        RECT 632.400 808.050 633.450 817.950 ;
        RECT 635.400 817.050 636.450 817.950 ;
        RECT 634.950 814.950 637.050 817.050 ;
        RECT 643.950 816.450 646.050 817.050 ;
        RECT 643.950 815.400 648.450 816.450 ;
        RECT 643.950 814.950 646.050 815.400 ;
        RECT 634.950 812.850 637.050 813.750 ;
        RECT 640.950 812.250 643.050 813.150 ;
        RECT 643.950 812.850 646.050 813.750 ;
        RECT 640.950 808.950 643.050 811.050 ;
        RECT 631.950 805.950 634.050 808.050 ;
        RECT 643.950 784.950 646.050 787.050 ;
        RECT 616.950 775.950 619.050 778.050 ;
        RECT 625.950 775.950 628.050 778.050 ;
        RECT 628.950 775.950 631.050 778.050 ;
        RECT 634.950 777.450 637.050 778.050 ;
        RECT 632.250 776.250 633.750 777.150 ;
        RECT 634.950 776.400 639.450 777.450 ;
        RECT 634.950 775.950 637.050 776.400 ;
        RECT 617.400 775.050 618.450 775.950 ;
        RECT 577.950 773.850 579.750 774.750 ;
        RECT 580.950 772.950 583.050 775.050 ;
        RECT 584.250 773.850 586.050 774.750 ;
        RECT 598.950 772.950 601.050 775.050 ;
        RECT 601.950 772.950 604.050 775.050 ;
        RECT 616.950 772.950 619.050 775.050 ;
        RECT 598.950 770.850 601.050 771.750 ;
        RECT 601.950 770.250 604.050 771.150 ;
        RECT 613.950 770.250 616.050 771.150 ;
        RECT 616.950 770.850 619.050 771.750 ;
        RECT 601.950 766.950 604.050 769.050 ;
        RECT 613.950 766.950 616.050 769.050 ;
        RECT 562.950 763.500 565.050 765.600 ;
        RECT 574.950 763.950 577.050 766.050 ;
        RECT 577.950 763.950 580.050 766.050 ;
        RECT 560.400 758.400 564.450 759.450 ;
        RECT 556.950 754.950 559.050 757.050 ;
        RECT 553.950 745.950 556.050 748.050 ;
        RECT 554.400 745.050 555.450 745.950 ;
        RECT 550.950 742.950 553.050 745.050 ;
        RECT 553.950 742.950 556.050 745.050 ;
        RECT 559.950 742.950 562.050 745.050 ;
        RECT 553.950 740.850 556.050 741.750 ;
        RECT 559.950 740.850 562.050 741.750 ;
        RECT 547.950 730.500 550.050 732.600 ;
        RECT 532.950 701.850 534.750 702.750 ;
        RECT 535.950 700.950 538.050 703.050 ;
        RECT 539.250 701.850 541.050 702.750 ;
        RECT 544.950 700.950 547.050 703.050 ;
        RECT 550.950 700.950 553.050 703.050 ;
        RECT 547.950 698.250 550.050 699.150 ;
        RECT 550.950 698.850 553.050 699.750 ;
        RECT 520.950 694.950 523.050 697.050 ;
        RECT 547.950 694.950 550.050 697.050 ;
        RECT 548.400 694.050 549.450 694.950 ;
        RECT 547.950 691.950 550.050 694.050 ;
        RECT 517.950 682.950 520.050 685.050 ;
        RECT 563.400 682.050 564.450 758.400 ;
        RECT 568.950 749.400 571.050 751.500 ;
        RECT 569.250 737.400 570.450 749.400 ;
        RECT 571.950 746.250 574.050 747.150 ;
        RECT 571.950 742.950 574.050 745.050 ;
        RECT 578.400 744.450 579.450 763.950 ;
        RECT 583.950 749.400 586.050 751.500 ;
        RECT 580.950 746.250 583.050 747.150 ;
        RECT 580.950 744.450 583.050 745.050 ;
        RECT 578.400 743.400 583.050 744.450 ;
        RECT 580.950 742.950 583.050 743.400 ;
        RECT 572.400 739.050 573.450 742.950 ;
        RECT 568.950 735.300 571.050 737.400 ;
        RECT 571.950 736.950 574.050 739.050 ;
        RECT 584.550 737.400 585.750 749.400 ;
        RECT 592.950 742.950 595.050 745.050 ;
        RECT 598.950 742.950 601.050 745.050 ;
        RECT 592.950 740.850 595.050 741.750 ;
        RECT 598.950 740.850 601.050 741.750 ;
        RECT 583.950 735.300 586.050 737.400 ;
        RECT 569.250 731.700 570.450 735.300 ;
        RECT 584.550 731.700 585.750 735.300 ;
        RECT 568.950 729.600 571.050 731.700 ;
        RECT 583.950 729.600 586.050 731.700 ;
        RECT 602.400 726.450 603.450 766.950 ;
        RECT 614.400 766.050 615.450 766.950 ;
        RECT 613.950 763.950 616.050 766.050 ;
        RECT 604.950 749.400 607.050 751.500 ;
        RECT 605.400 732.600 606.600 749.400 ;
        RECT 626.400 748.050 627.450 775.950 ;
        RECT 628.950 773.850 630.750 774.750 ;
        RECT 631.950 772.950 634.050 775.050 ;
        RECT 635.250 773.850 637.050 774.750 ;
        RECT 638.400 769.050 639.450 776.400 ;
        RECT 644.400 771.450 645.450 784.950 ;
        RECT 647.400 778.050 648.450 815.400 ;
        RECT 658.950 814.950 661.050 817.050 ;
        RECT 662.250 815.250 663.750 816.150 ;
        RECT 664.950 814.950 667.050 817.050 ;
        RECT 658.950 812.850 660.750 813.750 ;
        RECT 661.950 811.950 664.050 814.050 ;
        RECT 665.250 812.850 666.750 813.750 ;
        RECT 667.950 813.450 670.050 814.050 ;
        RECT 671.400 813.450 672.450 817.950 ;
        RECT 677.400 814.050 678.450 829.950 ;
        RECT 680.400 820.050 681.450 844.950 ;
        RECT 691.950 841.950 694.050 844.050 ;
        RECT 695.250 842.850 696.750 843.750 ;
        RECT 697.950 841.950 700.050 844.050 ;
        RECT 692.400 841.050 693.450 841.950 ;
        RECT 691.950 838.950 694.050 841.050 ;
        RECT 682.950 823.950 685.050 826.050 ;
        RECT 679.950 817.950 682.050 820.050 ;
        RECT 683.400 817.050 684.450 823.950 ;
        RECT 688.950 817.950 691.050 820.050 ;
        RECT 689.400 817.050 690.450 817.950 ;
        RECT 704.400 817.050 705.450 847.950 ;
        RECT 715.950 845.850 717.750 846.750 ;
        RECT 718.950 844.950 721.050 847.050 ;
        RECT 722.250 845.850 724.050 846.750 ;
        RECT 715.950 820.950 718.050 823.050 ;
        RECT 682.950 816.450 685.050 817.050 ;
        RECT 680.400 815.400 685.050 816.450 ;
        RECT 667.950 812.400 672.450 813.450 ;
        RECT 667.950 811.950 670.050 812.400 ;
        RECT 664.950 808.950 667.050 811.050 ;
        RECT 667.950 809.850 670.050 810.750 ;
        RECT 649.950 778.950 652.050 781.050 ;
        RECT 658.950 778.950 661.050 781.050 ;
        RECT 646.950 775.950 649.050 778.050 ;
        RECT 650.400 775.050 651.450 778.950 ;
        RECT 655.950 776.250 658.050 777.150 ;
        RECT 646.950 773.250 648.750 774.150 ;
        RECT 649.950 772.950 652.050 775.050 ;
        RECT 653.250 773.250 654.750 774.150 ;
        RECT 655.950 772.950 658.050 775.050 ;
        RECT 646.950 771.450 649.050 772.050 ;
        RECT 644.400 770.400 649.050 771.450 ;
        RECT 650.250 770.850 651.750 771.750 ;
        RECT 646.950 769.950 649.050 770.400 ;
        RECT 652.950 769.950 655.050 772.050 ;
        RECT 637.950 766.950 640.050 769.050 ;
        RECT 625.950 745.950 628.050 748.050 ;
        RECT 631.950 745.950 634.050 748.050 ;
        RECT 649.950 745.950 652.050 748.050 ;
        RECT 632.400 745.050 633.450 745.950 ;
        RECT 625.950 742.950 628.050 745.050 ;
        RECT 629.250 743.250 630.750 744.150 ;
        RECT 631.950 742.950 634.050 745.050 ;
        RECT 622.950 741.450 625.050 742.050 ;
        RECT 620.400 740.400 625.050 741.450 ;
        RECT 626.250 740.850 627.750 741.750 ;
        RECT 620.400 736.050 621.450 740.400 ;
        RECT 622.950 739.950 625.050 740.400 ;
        RECT 628.950 739.950 631.050 742.050 ;
        RECT 632.250 740.850 634.050 741.750 ;
        RECT 640.950 740.250 642.750 741.150 ;
        RECT 643.950 739.950 646.050 742.050 ;
        RECT 647.250 740.250 649.050 741.150 ;
        RECT 622.950 737.850 625.050 738.750 ;
        RECT 619.950 733.950 622.050 736.050 ;
        RECT 629.400 733.050 630.450 739.950 ;
        RECT 640.950 736.950 643.050 739.050 ;
        RECT 644.250 737.850 645.750 738.750 ;
        RECT 646.950 738.450 649.050 739.050 ;
        RECT 650.400 738.450 651.450 745.950 ;
        RECT 646.950 737.400 651.450 738.450 ;
        RECT 646.950 736.950 649.050 737.400 ;
        RECT 604.950 730.500 607.050 732.600 ;
        RECT 628.950 730.950 631.050 733.050 ;
        RECT 602.400 725.400 606.450 726.450 ;
        RECT 589.950 703.950 592.050 706.050 ;
        RECT 595.950 704.250 598.050 705.150 ;
        RECT 590.400 703.050 591.450 703.950 ;
        RECT 565.950 701.250 568.050 702.150 ;
        RECT 571.950 701.250 574.050 702.150 ;
        RECT 586.950 701.250 588.750 702.150 ;
        RECT 589.950 700.950 592.050 703.050 ;
        RECT 593.250 701.250 594.750 702.150 ;
        RECT 595.950 700.950 598.050 703.050 ;
        RECT 565.950 697.950 568.050 700.050 ;
        RECT 571.950 699.450 574.050 700.050 ;
        RECT 569.250 698.250 570.750 699.150 ;
        RECT 571.950 698.400 576.450 699.450 ;
        RECT 571.950 697.950 574.050 698.400 ;
        RECT 568.950 694.950 571.050 697.050 ;
        RECT 568.950 682.950 571.050 685.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 514.950 676.950 517.050 679.050 ;
        RECT 499.950 668.250 501.750 669.150 ;
        RECT 502.950 667.950 505.050 670.050 ;
        RECT 506.250 668.250 508.050 669.150 ;
        RECT 490.950 665.400 495.450 666.450 ;
        RECT 490.950 664.950 493.050 665.400 ;
        RECT 496.950 664.950 499.050 667.050 ;
        RECT 499.950 664.950 502.050 667.050 ;
        RECT 503.250 665.850 504.750 666.750 ;
        RECT 505.950 664.950 508.050 667.050 ;
        RECT 485.400 664.050 486.450 664.950 ;
        RECT 484.950 661.950 487.050 664.050 ;
        RECT 481.950 643.950 484.050 646.050 ;
        RECT 463.950 631.950 466.050 634.050 ;
        RECT 472.950 631.950 475.050 634.050 ;
        RECT 475.950 631.950 478.050 634.050 ;
        RECT 464.400 631.050 465.450 631.950 ;
        RECT 463.950 628.950 466.050 631.050 ;
        RECT 463.950 626.850 466.050 627.750 ;
        RECT 466.950 626.250 469.050 627.150 ;
        RECT 473.400 625.050 474.450 631.950 ;
        RECT 476.400 628.050 477.450 631.950 ;
        RECT 482.400 631.050 483.450 643.950 ;
        RECT 485.400 631.050 486.450 661.950 ;
        RECT 491.400 646.050 492.450 664.950 ;
        RECT 490.950 643.950 493.050 646.050 ;
        RECT 493.950 637.950 496.050 640.050 ;
        RECT 481.950 628.950 484.050 631.050 ;
        RECT 484.950 628.950 487.050 631.050 ;
        RECT 494.400 628.050 495.450 637.950 ;
        RECT 475.950 625.950 478.050 628.050 ;
        RECT 478.950 626.250 481.050 627.150 ;
        RECT 481.950 626.850 484.050 627.750 ;
        RECT 493.950 625.950 496.050 628.050 ;
        RECT 466.950 624.450 469.050 625.050 ;
        RECT 466.950 623.400 471.450 624.450 ;
        RECT 466.950 622.950 469.050 623.400 ;
        RECT 463.950 605.400 466.050 607.500 ;
        RECT 464.250 593.400 465.450 605.400 ;
        RECT 466.950 602.250 469.050 603.150 ;
        RECT 466.950 598.950 469.050 601.050 ;
        RECT 467.400 595.050 468.450 598.950 ;
        RECT 470.400 595.050 471.450 623.400 ;
        RECT 472.950 622.950 475.050 625.050 ;
        RECT 476.400 624.450 477.450 625.950 ;
        RECT 478.950 624.450 481.050 625.050 ;
        RECT 476.400 623.400 481.050 624.450 ;
        RECT 478.950 622.950 481.050 623.400 ;
        RECT 473.400 604.050 474.450 622.950 ;
        RECT 497.400 622.050 498.450 664.950 ;
        RECT 500.400 640.050 501.450 664.950 ;
        RECT 499.950 637.950 502.050 640.050 ;
        RECT 499.950 632.250 502.050 633.150 ;
        RECT 511.950 631.950 514.050 634.050 ;
        RECT 499.950 628.950 502.050 631.050 ;
        RECT 503.250 629.250 504.750 630.150 ;
        RECT 505.950 628.950 508.050 631.050 ;
        RECT 509.250 629.250 511.050 630.150 ;
        RECT 500.400 625.050 501.450 628.950 ;
        RECT 512.400 628.050 513.450 631.950 ;
        RECT 502.950 625.950 505.050 628.050 ;
        RECT 506.250 626.850 507.750 627.750 ;
        RECT 508.950 625.950 511.050 628.050 ;
        RECT 511.950 625.950 514.050 628.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 484.950 619.950 487.050 622.050 ;
        RECT 496.950 619.950 499.050 622.050 ;
        RECT 502.950 619.950 505.050 622.050 ;
        RECT 485.400 604.050 486.450 619.950 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 481.950 600.450 484.050 601.050 ;
        RECT 479.400 599.400 484.050 600.450 ;
        RECT 485.250 599.850 486.750 600.750 ;
        RECT 463.950 591.300 466.050 593.400 ;
        RECT 466.950 592.950 469.050 595.050 ;
        RECT 469.950 592.950 472.050 595.050 ;
        RECT 464.250 587.700 465.450 591.300 ;
        RECT 479.400 589.050 480.450 599.400 ;
        RECT 481.950 598.950 484.050 599.400 ;
        RECT 487.950 598.950 490.050 601.050 ;
        RECT 496.950 598.950 499.050 601.050 ;
        RECT 497.400 598.050 498.450 598.950 ;
        RECT 503.400 598.050 504.450 619.950 ;
        RECT 509.400 607.050 510.450 625.950 ;
        RECT 508.950 604.950 511.050 607.050 ;
        RECT 508.950 601.950 511.050 604.050 ;
        RECT 481.950 596.850 484.050 597.750 ;
        RECT 487.950 596.850 490.050 597.750 ;
        RECT 496.950 595.950 499.050 598.050 ;
        RECT 499.950 596.250 501.750 597.150 ;
        RECT 502.950 595.950 505.050 598.050 ;
        RECT 506.250 596.250 508.050 597.150 ;
        RECT 463.950 585.600 466.050 587.700 ;
        RECT 478.950 586.950 481.050 589.050 ;
        RECT 479.400 562.050 480.450 586.950 ;
        RECT 481.950 580.950 484.050 583.050 ;
        RECT 478.950 559.950 481.050 562.050 ;
        RECT 466.950 557.250 469.050 558.150 ;
        RECT 472.950 557.250 475.050 558.150 ;
        RECT 466.950 553.950 469.050 556.050 ;
        RECT 472.950 553.950 475.050 556.050 ;
        RECT 463.950 538.950 466.050 541.050 ;
        RECT 460.950 481.950 463.050 484.050 ;
        RECT 464.400 481.050 465.450 538.950 ;
        RECT 473.400 538.050 474.450 553.950 ;
        RECT 472.950 535.950 475.050 538.050 ;
        RECT 466.950 533.400 469.050 535.500 ;
        RECT 467.400 516.600 468.600 533.400 ;
        RECT 473.400 531.450 474.450 535.950 ;
        RECT 470.400 530.400 474.450 531.450 ;
        RECT 466.950 514.500 469.050 516.600 ;
        RECT 470.400 487.050 471.450 530.400 ;
        RECT 478.950 529.950 481.050 532.050 ;
        RECT 479.400 529.050 480.450 529.950 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 478.950 526.950 481.050 529.050 ;
        RECT 472.950 524.850 475.050 525.750 ;
        RECT 478.950 524.850 481.050 525.750 ;
        RECT 482.400 517.050 483.450 580.950 ;
        RECT 487.950 559.950 490.050 562.050 ;
        RECT 484.950 557.250 487.050 558.150 ;
        RECT 484.950 553.950 487.050 556.050 ;
        RECT 488.400 555.450 489.450 559.950 ;
        RECT 490.950 557.250 493.050 558.150 ;
        RECT 490.950 555.450 493.050 556.050 ;
        RECT 488.400 554.400 493.050 555.450 ;
        RECT 490.950 553.950 493.050 554.400 ;
        RECT 485.400 544.050 486.450 553.950 ;
        RECT 484.950 541.950 487.050 544.050 ;
        RECT 493.950 538.950 496.050 541.050 ;
        RECT 487.950 533.400 490.050 535.500 ;
        RECT 488.250 521.400 489.450 533.400 ;
        RECT 490.950 530.250 493.050 531.150 ;
        RECT 490.950 528.450 493.050 529.050 ;
        RECT 494.400 528.450 495.450 538.950 ;
        RECT 490.950 527.400 495.450 528.450 ;
        RECT 490.950 526.950 493.050 527.400 ;
        RECT 487.950 519.300 490.050 521.400 ;
        RECT 481.950 514.950 484.050 517.050 ;
        RECT 488.250 515.700 489.450 519.300 ;
        RECT 466.950 485.250 468.750 486.150 ;
        RECT 469.950 484.950 472.050 487.050 ;
        RECT 475.950 484.950 478.050 487.050 ;
        RECT 466.950 481.950 469.050 484.050 ;
        RECT 470.250 482.850 472.050 483.750 ;
        RECT 472.950 482.250 475.050 483.150 ;
        RECT 475.950 482.850 478.050 483.750 ;
        RECT 463.950 478.950 466.050 481.050 ;
        RECT 472.950 478.950 475.050 481.050 ;
        RECT 464.400 478.050 465.450 478.950 ;
        RECT 463.950 475.950 466.050 478.050 ;
        RECT 482.400 466.050 483.450 514.950 ;
        RECT 487.950 513.600 490.050 515.700 ;
        RECT 497.400 511.050 498.450 595.950 ;
        RECT 499.950 592.950 502.050 595.050 ;
        RECT 503.250 593.850 504.750 594.750 ;
        RECT 505.950 594.450 508.050 595.050 ;
        RECT 509.400 594.450 510.450 601.950 ;
        RECT 505.950 593.400 510.450 594.450 ;
        RECT 505.950 592.950 508.050 593.400 ;
        RECT 515.400 580.050 516.450 676.950 ;
        RECT 569.400 676.050 570.450 682.950 ;
        RECT 575.400 676.050 576.450 698.400 ;
        RECT 586.950 697.950 589.050 700.050 ;
        RECT 590.250 698.850 591.750 699.750 ;
        RECT 592.950 697.950 595.050 700.050 ;
        RECT 587.400 697.050 588.450 697.950 ;
        RECT 586.950 694.950 589.050 697.050 ;
        RECT 583.950 688.950 586.050 691.050 ;
        RECT 520.950 675.450 523.050 676.050 ;
        RECT 518.400 674.400 523.050 675.450 ;
        RECT 518.400 664.050 519.450 674.400 ;
        RECT 520.950 673.950 523.050 674.400 ;
        RECT 544.950 673.950 547.050 676.050 ;
        RECT 568.950 673.950 571.050 676.050 ;
        RECT 574.950 673.950 577.050 676.050 ;
        RECT 520.950 671.850 522.750 672.750 ;
        RECT 523.950 670.950 526.050 673.050 ;
        RECT 529.950 671.250 532.050 672.150 ;
        RECT 541.950 671.250 544.050 672.150 ;
        RECT 544.950 671.850 547.050 672.750 ;
        RECT 550.950 672.450 553.050 673.050 ;
        RECT 565.950 672.450 568.050 673.050 ;
        RECT 547.950 671.250 549.750 672.150 ;
        RECT 550.950 671.400 555.450 672.450 ;
        RECT 550.950 670.950 553.050 671.400 ;
        RECT 523.950 668.850 526.050 669.750 ;
        RECT 529.950 667.950 532.050 670.050 ;
        RECT 541.950 667.950 544.050 670.050 ;
        RECT 547.950 667.950 550.050 670.050 ;
        RECT 551.250 668.850 553.050 669.750 ;
        RECT 548.400 667.050 549.450 667.950 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 517.950 661.950 520.050 664.050 ;
        RECT 554.400 658.050 555.450 671.400 ;
        RECT 563.400 671.400 568.050 672.450 ;
        RECT 569.250 671.850 570.750 672.750 ;
        RECT 563.400 664.050 564.450 671.400 ;
        RECT 565.950 670.950 568.050 671.400 ;
        RECT 571.950 670.950 574.050 673.050 ;
        RECT 565.950 668.850 568.050 669.750 ;
        RECT 571.950 668.850 574.050 669.750 ;
        RECT 562.950 661.950 565.050 664.050 ;
        RECT 553.950 655.950 556.050 658.050 ;
        RECT 523.950 631.950 526.050 634.050 ;
        RECT 538.950 632.250 541.050 633.150 ;
        RECT 565.950 631.950 568.050 634.050 ;
        RECT 524.400 631.050 525.450 631.950 ;
        RECT 520.950 628.950 523.050 631.050 ;
        RECT 523.950 628.950 526.050 631.050 ;
        RECT 538.950 628.950 541.050 631.050 ;
        RECT 542.250 629.250 543.750 630.150 ;
        RECT 544.950 628.950 547.050 631.050 ;
        RECT 548.250 629.250 550.050 630.150 ;
        RECT 556.950 629.250 559.050 630.150 ;
        RECT 562.950 629.250 565.050 630.150 ;
        RECT 521.400 610.050 522.450 628.950 ;
        RECT 523.950 626.850 526.050 627.750 ;
        RECT 526.950 626.250 529.050 627.150 ;
        RECT 539.400 625.050 540.450 628.950 ;
        RECT 541.950 625.950 544.050 628.050 ;
        RECT 545.250 626.850 546.750 627.750 ;
        RECT 547.950 625.950 550.050 628.050 ;
        RECT 556.950 625.950 559.050 628.050 ;
        RECT 562.950 627.450 565.050 628.050 ;
        RECT 566.400 627.450 567.450 631.950 ;
        RECT 560.250 626.250 561.750 627.150 ;
        RECT 562.950 626.400 567.450 627.450 ;
        RECT 562.950 625.950 565.050 626.400 ;
        RECT 526.950 622.950 529.050 625.050 ;
        RECT 538.950 622.950 541.050 625.050 ;
        RECT 520.950 607.950 523.050 610.050 ;
        RECT 526.950 607.950 529.050 610.050 ;
        RECT 520.950 604.950 523.050 607.050 ;
        RECT 521.400 601.050 522.450 604.950 ;
        RECT 523.950 601.950 526.050 604.050 ;
        RECT 527.400 601.050 528.450 607.950 ;
        RECT 520.950 598.950 523.050 601.050 ;
        RECT 524.250 599.850 525.750 600.750 ;
        RECT 526.950 598.950 529.050 601.050 ;
        RECT 535.950 598.950 538.050 601.050 ;
        RECT 520.950 596.850 523.050 597.750 ;
        RECT 526.950 596.850 529.050 597.750 ;
        RECT 514.950 577.950 517.050 580.050 ;
        RECT 505.950 562.950 508.050 565.050 ;
        RECT 506.400 559.050 507.450 562.950 ;
        RECT 520.950 559.950 523.050 562.050 ;
        RECT 532.950 560.250 535.050 561.150 ;
        RECT 502.950 557.250 505.050 558.150 ;
        RECT 505.950 556.950 508.050 559.050 ;
        RECT 508.950 557.250 511.050 558.150 ;
        RECT 502.950 553.950 505.050 556.050 ;
        RECT 487.950 508.950 490.050 511.050 ;
        RECT 496.950 508.950 499.050 511.050 ;
        RECT 488.400 484.050 489.450 508.950 ;
        RECT 503.400 489.450 504.450 553.950 ;
        RECT 506.400 529.050 507.450 556.950 ;
        RECT 508.950 553.950 511.050 556.050 ;
        RECT 521.400 555.450 522.450 559.950 ;
        RECT 523.950 557.250 525.750 558.150 ;
        RECT 526.950 556.950 529.050 559.050 ;
        RECT 530.250 557.250 531.750 558.150 ;
        RECT 532.950 556.950 535.050 559.050 ;
        RECT 523.950 555.450 526.050 556.050 ;
        RECT 521.400 554.400 526.050 555.450 ;
        RECT 527.250 554.850 528.750 555.750 ;
        RECT 523.950 553.950 526.050 554.400 ;
        RECT 529.950 553.950 532.050 556.050 ;
        RECT 509.400 553.050 510.450 553.950 ;
        RECT 508.950 550.950 511.050 553.050 ;
        RECT 533.400 550.050 534.450 556.950 ;
        RECT 532.950 547.950 535.050 550.050 ;
        RECT 533.400 547.050 534.450 547.950 ;
        RECT 532.950 544.950 535.050 547.050 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 526.950 529.950 529.050 532.050 ;
        RECT 505.950 526.950 508.050 529.050 ;
        RECT 509.250 527.250 511.050 528.150 ;
        RECT 511.950 527.850 514.050 528.750 ;
        RECT 523.950 528.450 526.050 529.050 ;
        RECT 514.950 527.250 517.050 528.150 ;
        RECT 521.400 527.400 526.050 528.450 ;
        RECT 521.400 526.050 522.450 527.400 ;
        RECT 523.950 526.950 526.050 527.400 ;
        RECT 505.950 524.850 507.750 525.750 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 523.950 524.850 526.050 525.750 ;
        RECT 509.400 523.050 510.450 523.950 ;
        RECT 508.950 520.950 511.050 523.050 ;
        RECT 515.400 490.050 516.450 523.950 ;
        RECT 527.400 522.450 528.450 529.950 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 529.950 524.250 532.050 525.150 ;
        RECT 532.950 524.850 535.050 525.750 ;
        RECT 529.950 522.450 532.050 523.050 ;
        RECT 527.400 521.400 532.050 522.450 ;
        RECT 523.950 517.950 526.050 520.050 ;
        RECT 517.950 493.950 520.050 496.050 ;
        RECT 490.950 488.250 493.050 489.150 ;
        RECT 503.400 488.400 507.450 489.450 ;
        RECT 490.950 484.950 493.050 487.050 ;
        RECT 494.250 485.250 495.750 486.150 ;
        RECT 496.950 484.950 499.050 487.050 ;
        RECT 500.250 485.250 502.050 486.150 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 487.950 481.950 490.050 484.050 ;
        RECT 491.400 469.050 492.450 484.950 ;
        RECT 493.950 481.950 496.050 484.050 ;
        RECT 497.250 482.850 498.750 483.750 ;
        RECT 499.950 481.950 502.050 484.050 ;
        RECT 500.400 481.050 501.450 481.950 ;
        RECT 493.950 478.950 496.050 481.050 ;
        RECT 499.950 478.950 502.050 481.050 ;
        RECT 490.950 466.950 493.050 469.050 ;
        RECT 481.950 463.950 484.050 466.050 ;
        RECT 484.950 460.950 487.050 463.050 ;
        RECT 466.950 457.950 469.050 460.050 ;
        RECT 467.400 457.050 468.450 457.950 ;
        RECT 485.400 457.050 486.450 460.950 ;
        RECT 466.950 454.950 469.050 457.050 ;
        RECT 470.250 455.250 471.750 456.150 ;
        RECT 472.950 454.950 475.050 457.050 ;
        RECT 475.950 454.950 478.050 457.050 ;
        RECT 478.950 454.950 481.050 457.050 ;
        RECT 484.950 454.950 487.050 457.050 ;
        RECT 463.950 451.950 466.050 454.050 ;
        RECT 467.250 452.850 468.750 453.750 ;
        RECT 469.950 451.950 472.050 454.050 ;
        RECT 473.250 452.850 475.050 453.750 ;
        RECT 463.950 449.850 466.050 450.750 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 457.950 442.950 460.050 445.050 ;
        RECT 454.950 436.950 457.050 439.050 ;
        RECT 439.950 410.400 444.450 411.450 ;
        RECT 445.950 410.850 447.750 411.750 ;
        RECT 439.950 409.950 442.050 410.400 ;
        RECT 448.950 409.950 451.050 412.050 ;
        RECT 451.950 409.950 454.050 412.050 ;
        RECT 445.950 406.950 448.050 409.050 ;
        RECT 436.950 384.450 439.050 385.050 ;
        RECT 433.950 383.250 435.750 384.150 ;
        RECT 436.950 383.400 441.450 384.450 ;
        RECT 436.950 382.950 439.050 383.400 ;
        RECT 440.400 382.050 441.450 383.400 ;
        RECT 433.950 379.950 436.050 382.050 ;
        RECT 437.250 380.850 439.050 381.750 ;
        RECT 439.950 379.950 442.050 382.050 ;
        RECT 430.950 364.950 433.050 367.050 ;
        RECT 424.950 349.950 427.050 352.050 ;
        RECT 425.400 339.450 426.450 349.950 ;
        RECT 434.400 346.050 435.450 379.950 ;
        RECT 442.950 364.950 445.050 367.050 ;
        RECT 433.950 343.950 436.050 346.050 ;
        RECT 430.950 342.450 433.050 343.050 ;
        RECT 439.950 342.450 442.050 343.050 ;
        RECT 443.400 342.450 444.450 364.950 ;
        RECT 427.950 341.250 429.750 342.150 ;
        RECT 430.950 341.400 435.450 342.450 ;
        RECT 430.950 340.950 433.050 341.400 ;
        RECT 427.950 339.450 430.050 340.050 ;
        RECT 425.400 338.400 430.050 339.450 ;
        RECT 431.250 338.850 433.050 339.750 ;
        RECT 427.950 337.950 430.050 338.400 ;
        RECT 434.400 336.450 435.450 341.400 ;
        RECT 436.950 341.250 438.750 342.150 ;
        RECT 439.950 341.400 444.450 342.450 ;
        RECT 439.950 340.950 442.050 341.400 ;
        RECT 436.950 337.950 439.050 340.050 ;
        RECT 440.250 338.850 442.050 339.750 ;
        RECT 434.400 335.400 438.450 336.450 ;
        RECT 418.950 328.950 421.050 331.050 ;
        RECT 430.950 316.950 433.050 319.050 ;
        RECT 431.400 316.050 432.450 316.950 ;
        RECT 430.950 313.950 433.050 316.050 ;
        RECT 427.950 310.950 430.050 313.050 ;
        RECT 430.950 311.850 433.050 312.750 ;
        RECT 433.950 311.250 436.050 312.150 ;
        RECT 412.950 308.250 414.750 309.150 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 419.250 308.250 421.050 309.150 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 412.950 304.950 415.050 307.050 ;
        RECT 416.250 305.850 417.750 306.750 ;
        RECT 418.950 306.450 421.050 307.050 ;
        RECT 422.400 306.450 423.450 307.950 ;
        RECT 418.950 305.400 423.450 306.450 ;
        RECT 418.950 304.950 421.050 305.400 ;
        RECT 403.950 301.950 406.050 304.050 ;
        RECT 400.950 298.950 403.050 301.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 397.950 271.950 400.050 274.050 ;
        RECT 385.950 270.450 388.050 271.050 ;
        RECT 382.950 269.250 384.750 270.150 ;
        RECT 385.950 269.400 390.450 270.450 ;
        RECT 385.950 268.950 388.050 269.400 ;
        RECT 367.950 266.400 372.450 267.450 ;
        RECT 367.950 265.950 370.050 266.400 ;
        RECT 373.950 265.950 376.050 268.050 ;
        RECT 382.950 265.950 385.050 268.050 ;
        RECT 386.250 266.850 388.050 267.750 ;
        RECT 314.400 244.050 315.450 265.950 ;
        RECT 319.950 262.950 322.050 265.050 ;
        RECT 320.400 256.050 321.450 262.950 ;
        RECT 335.400 259.050 336.450 265.950 ;
        RECT 344.400 259.050 345.450 265.950 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 335.400 256.050 336.450 256.950 ;
        RECT 319.950 253.950 322.050 256.050 ;
        RECT 334.950 253.950 337.050 256.050 ;
        RECT 343.950 253.950 346.050 256.050 ;
        RECT 337.950 244.950 340.050 247.050 ;
        RECT 313.950 241.950 316.050 244.050 ;
        RECT 307.950 236.250 309.750 237.150 ;
        RECT 310.950 235.950 313.050 238.050 ;
        RECT 314.400 237.450 315.450 241.950 ;
        RECT 338.400 241.050 339.450 244.950 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 328.950 238.950 331.050 241.050 ;
        RECT 331.950 238.950 334.050 241.050 ;
        RECT 335.250 239.250 336.750 240.150 ;
        RECT 337.950 238.950 340.050 241.050 ;
        RECT 316.950 237.450 319.050 238.050 ;
        RECT 314.400 236.400 319.050 237.450 ;
        RECT 316.950 235.950 319.050 236.400 ;
        RECT 320.400 235.050 321.450 238.950 ;
        RECT 329.400 238.050 330.450 238.950 ;
        RECT 328.950 235.950 331.050 238.050 ;
        RECT 332.250 236.850 333.750 237.750 ;
        RECT 334.950 235.950 337.050 238.050 ;
        RECT 338.250 236.850 340.050 237.750 ;
        RECT 307.950 232.950 310.050 235.050 ;
        RECT 311.250 233.850 312.750 234.750 ;
        RECT 313.950 232.950 316.050 235.050 ;
        RECT 317.250 233.850 319.050 234.750 ;
        RECT 319.950 232.950 322.050 235.050 ;
        RECT 328.950 233.850 331.050 234.750 ;
        RECT 308.400 208.050 309.450 232.950 ;
        RECT 313.950 230.850 316.050 231.750 ;
        RECT 307.950 205.950 310.050 208.050 ;
        RECT 340.950 206.400 343.050 208.500 ;
        RECT 304.950 199.950 307.050 202.050 ;
        RECT 308.250 200.250 309.750 201.150 ;
        RECT 322.950 200.250 325.050 201.150 ;
        RECT 328.950 199.950 331.050 202.050 ;
        RECT 329.400 199.050 330.450 199.950 ;
        RECT 304.950 197.850 306.750 198.750 ;
        RECT 307.950 196.950 310.050 199.050 ;
        RECT 311.250 197.850 313.050 198.750 ;
        RECT 322.950 196.950 325.050 199.050 ;
        RECT 326.250 197.250 327.750 198.150 ;
        RECT 328.950 196.950 331.050 199.050 ;
        RECT 332.250 197.250 334.050 198.150 ;
        RECT 325.950 193.950 328.050 196.050 ;
        RECT 329.250 194.850 330.750 195.750 ;
        RECT 331.950 193.950 334.050 196.050 ;
        RECT 301.950 184.950 304.050 187.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 293.400 169.050 294.450 178.950 ;
        RECT 295.950 172.950 298.050 175.050 ;
        RECT 238.950 166.950 241.050 169.050 ;
        RECT 250.950 166.950 253.050 169.050 ;
        RECT 274.950 166.950 277.050 169.050 ;
        RECT 278.250 167.250 279.750 168.150 ;
        RECT 280.950 166.950 283.050 169.050 ;
        RECT 292.950 166.950 295.050 169.050 ;
        RECT 229.950 164.250 231.750 165.150 ;
        RECT 232.950 163.950 235.050 166.050 ;
        RECT 236.250 164.250 238.050 165.150 ;
        RECT 229.950 160.950 232.050 163.050 ;
        RECT 233.250 161.850 234.750 162.750 ;
        RECT 235.950 162.450 238.050 163.050 ;
        RECT 239.400 162.450 240.450 166.950 ;
        RECT 250.950 164.850 253.050 165.750 ;
        RECT 256.950 164.850 259.050 165.750 ;
        RECT 271.950 163.950 274.050 166.050 ;
        RECT 275.250 164.850 276.750 165.750 ;
        RECT 277.950 163.950 280.050 166.050 ;
        RECT 281.250 164.850 283.050 165.750 ;
        RECT 292.950 164.850 295.050 165.750 ;
        RECT 296.400 165.450 297.450 172.950 ;
        RECT 302.400 169.050 303.450 184.950 ;
        RECT 332.400 180.450 333.450 193.950 ;
        RECT 341.400 189.600 342.600 206.400 ;
        RECT 340.950 187.500 343.050 189.600 ;
        RECT 332.400 179.400 336.450 180.450 ;
        RECT 322.950 172.950 325.050 175.050 ;
        RECT 323.400 172.050 324.450 172.950 ;
        RECT 322.950 169.950 325.050 172.050 ;
        RECT 331.950 169.950 334.050 172.050 ;
        RECT 298.950 167.250 300.750 168.150 ;
        RECT 301.950 166.950 304.050 169.050 ;
        RECT 307.950 167.250 310.050 168.150 ;
        RECT 322.950 167.850 325.050 168.750 ;
        RECT 325.950 167.250 328.050 168.150 ;
        RECT 298.950 165.450 301.050 166.050 ;
        RECT 296.400 164.400 301.050 165.450 ;
        RECT 302.250 164.850 304.050 165.750 ;
        RECT 298.950 163.950 301.050 164.400 ;
        RECT 307.950 163.950 310.050 166.050 ;
        RECT 325.950 163.950 328.050 166.050 ;
        RECT 235.950 161.400 240.450 162.450 ;
        RECT 271.950 161.850 274.050 162.750 ;
        RECT 235.950 160.950 238.050 161.400 ;
        RECT 278.400 160.050 279.450 163.950 ;
        RECT 277.950 157.950 280.050 160.050 ;
        RECT 308.400 136.050 309.450 163.950 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 326.400 133.050 327.450 163.950 ;
        RECT 223.950 130.950 226.050 133.050 ;
        RECT 271.950 131.250 274.050 132.150 ;
        RECT 307.950 131.250 310.050 132.150 ;
        RECT 325.950 130.950 328.050 133.050 ;
        RECT 224.400 126.450 225.450 130.950 ;
        RECT 265.950 129.450 268.050 130.050 ;
        RECT 226.950 128.250 229.050 129.150 ;
        RECT 263.400 128.400 268.050 129.450 ;
        RECT 226.950 126.450 229.050 127.050 ;
        RECT 224.400 125.400 229.050 126.450 ;
        RECT 226.950 124.950 229.050 125.400 ;
        RECT 230.250 125.250 231.750 126.150 ;
        RECT 232.950 124.950 235.050 127.050 ;
        RECT 236.250 125.250 238.050 126.150 ;
        RECT 247.950 124.950 250.050 127.050 ;
        RECT 229.950 121.950 232.050 124.050 ;
        RECT 233.250 122.850 234.750 123.750 ;
        RECT 235.950 121.950 238.050 124.050 ;
        RECT 244.950 122.250 247.050 123.150 ;
        RECT 247.950 122.850 250.050 123.750 ;
        RECT 220.950 97.950 223.050 100.050 ;
        RECT 226.950 96.450 229.050 97.050 ;
        RECT 230.400 96.450 231.450 121.950 ;
        RECT 263.400 121.050 264.450 128.400 ;
        RECT 265.950 127.950 268.050 128.400 ;
        RECT 269.250 128.250 270.750 129.150 ;
        RECT 271.950 127.950 274.050 130.050 ;
        RECT 275.250 128.250 277.050 129.150 ;
        RECT 283.950 127.950 286.050 130.050 ;
        RECT 304.950 128.250 306.750 129.150 ;
        RECT 307.950 127.950 310.050 130.050 ;
        RECT 313.950 129.450 316.050 130.050 ;
        RECT 311.250 128.250 312.750 129.150 ;
        RECT 313.950 128.400 318.450 129.450 ;
        RECT 313.950 127.950 316.050 128.400 ;
        RECT 265.950 125.850 267.750 126.750 ;
        RECT 268.950 124.950 271.050 127.050 ;
        RECT 244.950 118.950 247.050 121.050 ;
        RECT 262.950 118.950 265.050 121.050 ;
        RECT 269.400 118.050 270.450 124.950 ;
        RECT 268.950 115.950 271.050 118.050 ;
        RECT 269.400 115.050 270.450 115.950 ;
        RECT 268.950 112.950 271.050 115.050 ;
        RECT 265.950 109.950 268.050 112.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 226.950 95.400 231.450 96.450 ;
        RECT 235.950 96.450 238.050 97.050 ;
        RECT 235.950 95.400 240.450 96.450 ;
        RECT 226.950 94.950 229.050 95.400 ;
        RECT 235.950 94.950 238.050 95.400 ;
        RECT 217.950 91.950 220.050 94.050 ;
        RECT 226.950 92.850 229.050 93.750 ;
        RECT 232.950 92.250 235.050 93.150 ;
        RECT 235.950 92.850 238.050 93.750 ;
        RECT 169.950 88.950 172.050 91.050 ;
        RECT 184.950 88.950 187.050 91.050 ;
        RECT 188.250 89.850 189.750 90.750 ;
        RECT 190.950 88.950 193.050 91.050 ;
        RECT 194.250 89.850 196.050 90.750 ;
        RECT 208.950 88.950 211.050 91.050 ;
        RECT 212.250 89.850 213.750 90.750 ;
        RECT 214.950 88.950 217.050 91.050 ;
        RECT 218.250 89.850 220.050 90.750 ;
        RECT 232.950 88.950 235.050 91.050 ;
        RECT 155.400 77.400 159.450 78.450 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 149.250 56.250 150.750 57.150 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 145.950 53.850 147.750 54.750 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 152.250 53.850 154.050 54.750 ;
        RECT 145.950 31.950 148.050 34.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 139.950 21.450 142.050 22.050 ;
        RECT 143.400 21.450 144.450 22.950 ;
        RECT 146.400 22.050 147.450 31.950 ;
        RECT 149.400 24.450 150.450 52.950 ;
        RECT 155.400 37.050 156.450 77.400 ;
        RECT 157.950 73.950 160.050 76.050 ;
        RECT 158.400 52.050 159.450 73.950 ;
        RECT 163.950 57.450 166.050 58.050 ;
        RECT 166.950 57.450 169.050 58.050 ;
        RECT 163.950 56.400 169.050 57.450 ;
        RECT 163.950 55.950 166.050 56.400 ;
        RECT 166.950 55.950 169.050 56.400 ;
        RECT 160.950 53.250 163.050 54.150 ;
        RECT 157.950 49.950 160.050 52.050 ;
        RECT 160.950 49.950 163.050 52.050 ;
        RECT 161.400 49.050 162.450 49.950 ;
        RECT 160.950 46.950 163.050 49.050 ;
        RECT 164.400 46.050 165.450 55.950 ;
        RECT 166.950 53.850 169.050 54.750 ;
        RECT 169.950 53.250 172.050 54.150 ;
        RECT 169.950 49.950 172.050 52.050 ;
        RECT 163.950 43.950 166.050 46.050 ;
        RECT 154.950 34.950 157.050 37.050 ;
        RECT 160.950 31.950 163.050 34.050 ;
        RECT 149.400 23.400 153.450 24.450 ;
        RECT 139.950 20.400 144.450 21.450 ;
        RECT 139.950 19.950 142.050 20.400 ;
        RECT 145.950 19.950 148.050 22.050 ;
        RECT 149.250 20.250 151.050 21.150 ;
        RECT 49.950 17.850 52.050 18.750 ;
        RECT 97.950 16.950 100.050 19.050 ;
        RECT 103.950 17.850 106.050 18.750 ;
        RECT 106.950 16.950 109.050 19.050 ;
        RECT 118.950 17.850 120.750 18.750 ;
        RECT 121.950 16.950 124.050 19.050 ;
        RECT 125.250 17.850 126.750 18.750 ;
        RECT 127.950 16.950 130.050 19.050 ;
        RECT 136.950 16.950 139.050 19.050 ;
        RECT 139.950 17.850 141.750 18.750 ;
        RECT 142.950 16.950 145.050 19.050 ;
        RECT 146.250 17.850 147.750 18.750 ;
        RECT 148.950 16.950 151.050 19.050 ;
        RECT 121.950 14.850 124.050 15.750 ;
        RECT 142.950 14.850 145.050 15.750 ;
        RECT 152.400 13.050 153.450 23.400 ;
        RECT 161.400 21.450 162.450 31.950 ;
        RECT 185.400 31.050 186.450 88.950 ;
        RECT 190.950 86.850 193.050 87.750 ;
        RECT 187.950 52.950 190.050 55.050 ;
        RECT 202.950 54.450 205.050 55.050 ;
        RECT 202.950 53.400 207.450 54.450 ;
        RECT 202.950 52.950 205.050 53.400 ;
        RECT 187.950 50.850 190.050 51.750 ;
        RECT 190.950 50.250 193.050 51.150 ;
        RECT 199.950 50.250 202.050 51.150 ;
        RECT 202.950 50.850 205.050 51.750 ;
        RECT 190.950 46.950 193.050 49.050 ;
        RECT 199.950 46.950 202.050 49.050 ;
        RECT 191.400 46.050 192.450 46.950 ;
        RECT 190.950 43.950 193.050 46.050 ;
        RECT 206.400 34.050 207.450 53.400 ;
        RECT 209.400 49.050 210.450 88.950 ;
        RECT 214.950 86.850 217.050 87.750 ;
        RECT 229.950 58.950 232.050 61.050 ;
        RECT 214.950 52.950 217.050 55.050 ;
        RECT 217.950 53.250 219.750 54.150 ;
        RECT 220.950 52.950 223.050 55.050 ;
        RECT 226.950 52.950 229.050 55.050 ;
        RECT 208.950 46.950 211.050 49.050 ;
        RECT 215.400 46.050 216.450 52.950 ;
        RECT 230.400 52.050 231.450 58.950 ;
        RECT 239.400 58.050 240.450 95.400 ;
        RECT 245.400 90.450 246.450 100.950 ;
        RECT 248.400 97.050 249.450 100.950 ;
        RECT 266.400 100.050 267.450 109.950 ;
        RECT 272.400 109.050 273.450 127.950 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 275.400 124.050 276.450 124.950 ;
        RECT 274.950 121.950 277.050 124.050 ;
        RECT 271.950 106.950 274.050 109.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 269.400 100.050 270.450 100.950 ;
        RECT 265.950 97.950 268.050 100.050 ;
        RECT 268.950 97.950 271.050 100.050 ;
        RECT 271.950 97.950 274.050 100.050 ;
        RECT 266.400 97.050 267.450 97.950 ;
        RECT 272.400 97.050 273.450 97.950 ;
        RECT 247.950 94.950 250.050 97.050 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 265.950 94.950 268.050 97.050 ;
        RECT 269.250 95.850 270.750 96.750 ;
        RECT 271.950 94.950 274.050 97.050 ;
        RECT 247.950 92.250 249.750 93.150 ;
        RECT 250.950 91.950 253.050 94.050 ;
        RECT 254.250 92.250 256.050 93.150 ;
        RECT 247.950 90.450 250.050 91.050 ;
        RECT 245.400 89.400 250.050 90.450 ;
        RECT 251.250 89.850 252.750 90.750 ;
        RECT 253.950 90.450 256.050 91.050 ;
        RECT 257.400 90.450 258.450 94.950 ;
        RECT 265.950 92.850 268.050 93.750 ;
        RECT 271.950 92.850 274.050 93.750 ;
        RECT 247.950 88.950 250.050 89.400 ;
        RECT 253.950 89.400 258.450 90.450 ;
        RECT 253.950 88.950 256.050 89.400 ;
        RECT 253.950 85.950 256.050 88.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 244.950 56.250 247.050 57.150 ;
        RECT 217.950 49.950 220.050 52.050 ;
        RECT 221.250 50.850 223.050 51.750 ;
        RECT 223.950 50.250 226.050 51.150 ;
        RECT 226.950 50.850 229.050 51.750 ;
        RECT 229.950 49.950 232.050 52.050 ;
        RECT 223.950 46.950 226.050 49.050 ;
        RECT 214.950 43.950 217.050 46.050 ;
        RECT 205.950 31.950 208.050 34.050 ;
        RECT 184.950 28.950 187.050 31.050 ;
        RECT 166.950 25.950 169.050 28.050 ;
        RECT 175.950 25.950 178.050 28.050 ;
        RECT 193.950 25.950 196.050 28.050 ;
        RECT 163.950 23.250 166.050 24.150 ;
        RECT 166.950 23.850 169.050 24.750 ;
        RECT 169.950 23.250 171.750 24.150 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 163.950 21.450 166.050 22.050 ;
        RECT 161.400 20.400 166.050 21.450 ;
        RECT 163.950 19.950 166.050 20.400 ;
        RECT 166.950 19.950 169.050 22.050 ;
        RECT 169.950 19.950 172.050 22.050 ;
        RECT 173.250 20.850 175.050 21.750 ;
        RECT 167.400 18.450 168.450 19.950 ;
        RECT 176.400 18.450 177.450 25.950 ;
        RECT 187.950 24.450 190.050 25.050 ;
        RECT 167.400 17.400 177.450 18.450 ;
        RECT 185.400 23.400 190.050 24.450 ;
        RECT 185.400 16.050 186.450 23.400 ;
        RECT 187.950 22.950 190.050 23.400 ;
        RECT 191.250 23.250 193.050 24.150 ;
        RECT 193.950 23.850 196.050 24.750 ;
        RECT 196.950 23.250 199.050 24.150 ;
        RECT 206.400 22.050 207.450 31.950 ;
        RECT 233.400 31.050 234.450 55.950 ;
        RECT 235.950 53.250 237.750 54.150 ;
        RECT 238.950 52.950 241.050 55.050 ;
        RECT 242.250 53.250 243.750 54.150 ;
        RECT 244.950 52.950 247.050 55.050 ;
        RECT 235.950 49.950 238.050 52.050 ;
        RECT 239.250 50.850 240.750 51.750 ;
        RECT 241.950 49.950 244.050 52.050 ;
        RECT 236.400 49.050 237.450 49.950 ;
        RECT 235.950 46.950 238.050 49.050 ;
        RECT 245.400 43.050 246.450 52.950 ;
        RECT 254.400 49.050 255.450 85.950 ;
        RECT 262.950 58.950 265.050 61.050 ;
        RECT 263.400 55.050 264.450 58.950 ;
        RECT 284.400 58.050 285.450 127.950 ;
        RECT 289.950 125.250 292.050 126.150 ;
        RECT 295.950 125.250 298.050 126.150 ;
        RECT 304.950 124.950 307.050 127.050 ;
        RECT 286.950 121.950 289.050 124.050 ;
        RECT 289.950 121.950 292.050 124.050 ;
        RECT 295.950 121.950 298.050 124.050 ;
        RECT 287.400 94.050 288.450 121.950 ;
        RECT 290.400 121.050 291.450 121.950 ;
        RECT 289.950 118.950 292.050 121.050 ;
        RECT 296.400 106.050 297.450 121.950 ;
        RECT 295.950 103.950 298.050 106.050 ;
        RECT 305.400 103.050 306.450 124.950 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 304.950 99.450 307.050 100.050 ;
        RECT 308.400 99.450 309.450 127.950 ;
        RECT 310.950 124.950 313.050 127.050 ;
        RECT 314.250 125.850 316.050 126.750 ;
        RECT 317.400 118.050 318.450 128.400 ;
        RECT 328.950 127.950 331.050 130.050 ;
        RECT 329.400 127.050 330.450 127.950 ;
        RECT 322.950 124.950 325.050 127.050 ;
        RECT 328.950 124.950 331.050 127.050 ;
        RECT 316.950 115.950 319.050 118.050 ;
        RECT 304.950 98.400 309.450 99.450 ;
        RECT 304.950 97.950 307.050 98.400 ;
        RECT 323.400 97.050 324.450 124.950 ;
        RECT 332.400 124.050 333.450 169.950 ;
        RECT 335.400 157.050 336.450 179.400 ;
        RECT 344.400 169.050 345.450 253.950 ;
        RECT 362.400 247.050 363.450 265.950 ;
        RECT 383.400 262.050 384.450 265.950 ;
        RECT 382.950 259.950 385.050 262.050 ;
        RECT 389.400 247.050 390.450 269.400 ;
        RECT 391.950 269.250 393.750 270.150 ;
        RECT 394.950 268.950 397.050 271.050 ;
        RECT 398.400 268.050 399.450 271.950 ;
        RECT 391.950 265.950 394.050 268.050 ;
        RECT 395.250 266.850 397.050 267.750 ;
        RECT 397.950 265.950 400.050 268.050 ;
        RECT 401.400 264.450 402.450 289.950 ;
        RECT 409.950 280.950 412.050 283.050 ;
        RECT 410.400 274.050 411.450 280.950 ;
        RECT 403.950 271.950 406.050 274.050 ;
        RECT 407.250 272.250 408.750 273.150 ;
        RECT 409.950 271.950 412.050 274.050 ;
        RECT 413.400 271.050 414.450 304.950 ;
        RECT 415.950 271.950 418.050 274.050 ;
        RECT 403.950 269.850 405.750 270.750 ;
        RECT 406.950 268.950 409.050 271.050 ;
        RECT 410.250 269.850 412.050 270.750 ;
        RECT 412.950 268.950 415.050 271.050 ;
        RECT 398.400 263.400 402.450 264.450 ;
        RECT 394.950 250.950 397.050 253.050 ;
        RECT 361.950 244.950 364.050 247.050 ;
        RECT 367.950 244.950 370.050 247.050 ;
        RECT 376.950 244.950 379.050 247.050 ;
        RECT 388.950 244.950 391.050 247.050 ;
        RECT 352.950 243.450 355.050 244.050 ;
        RECT 352.950 242.400 357.450 243.450 ;
        RECT 352.950 241.950 355.050 242.400 ;
        RECT 356.400 241.050 357.450 242.400 ;
        RECT 346.950 238.950 349.050 241.050 ;
        RECT 349.950 239.250 352.050 240.150 ;
        RECT 352.950 239.850 355.050 240.750 ;
        RECT 355.950 238.950 358.050 241.050 ;
        RECT 347.400 229.050 348.450 238.950 ;
        RECT 349.950 235.950 352.050 238.050 ;
        RECT 346.950 226.950 349.050 229.050 ;
        RECT 362.400 214.050 363.450 244.950 ;
        RECT 368.400 244.050 369.450 244.950 ;
        RECT 367.950 241.950 370.050 244.050 ;
        RECT 364.950 238.950 367.050 241.050 ;
        RECT 368.250 239.850 369.750 240.750 ;
        RECT 370.950 240.450 373.050 241.050 ;
        RECT 370.950 239.400 375.450 240.450 ;
        RECT 370.950 238.950 373.050 239.400 ;
        RECT 364.950 236.850 367.050 237.750 ;
        RECT 370.950 236.850 373.050 237.750 ;
        RECT 374.400 235.050 375.450 239.400 ;
        RECT 373.950 232.950 376.050 235.050 ;
        RECT 374.400 232.050 375.450 232.950 ;
        RECT 373.950 229.950 376.050 232.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 346.950 197.250 349.050 198.150 ;
        RECT 352.950 197.250 355.050 198.150 ;
        RECT 346.950 193.950 349.050 196.050 ;
        RECT 352.950 193.950 355.050 196.050 ;
        RECT 353.400 193.050 354.450 193.950 ;
        RECT 352.950 190.950 355.050 193.050 ;
        RECT 337.950 166.950 340.050 169.050 ;
        RECT 341.250 167.250 342.750 168.150 ;
        RECT 343.950 166.950 346.050 169.050 ;
        RECT 337.950 164.850 339.750 165.750 ;
        RECT 340.950 163.950 343.050 166.050 ;
        RECT 344.250 164.850 345.750 165.750 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 341.400 157.050 342.450 163.950 ;
        RECT 346.950 161.850 349.050 162.750 ;
        RECT 334.950 154.950 337.050 157.050 ;
        RECT 340.950 154.950 343.050 157.050 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 334.950 127.950 337.050 130.050 ;
        RECT 325.950 122.250 328.050 123.150 ;
        RECT 328.950 122.850 331.050 123.750 ;
        RECT 331.950 121.950 334.050 124.050 ;
        RECT 325.950 118.950 328.050 121.050 ;
        RECT 326.400 112.050 327.450 118.950 ;
        RECT 325.950 109.950 328.050 112.050 ;
        RECT 335.400 103.050 336.450 127.950 ;
        RECT 347.400 127.050 348.450 133.950 ;
        RECT 352.950 128.250 355.050 129.150 ;
        RECT 343.950 125.250 345.750 126.150 ;
        RECT 346.950 124.950 349.050 127.050 ;
        RECT 350.250 125.250 351.750 126.150 ;
        RECT 352.950 124.950 355.050 127.050 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 347.250 122.850 348.750 123.750 ;
        RECT 349.950 121.950 352.050 124.050 ;
        RECT 344.400 118.050 345.450 121.950 ;
        RECT 343.950 115.950 346.050 118.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 289.950 94.950 292.050 97.050 ;
        RECT 293.250 95.250 294.750 96.150 ;
        RECT 295.950 94.950 298.050 97.050 ;
        RECT 304.950 95.850 307.050 96.750 ;
        RECT 307.950 95.250 310.050 96.150 ;
        RECT 322.950 94.950 325.050 97.050 ;
        RECT 286.950 91.950 289.050 94.050 ;
        RECT 290.250 92.850 291.750 93.750 ;
        RECT 292.950 91.950 295.050 94.050 ;
        RECT 296.250 92.850 298.050 93.750 ;
        RECT 304.950 91.950 307.050 94.050 ;
        RECT 307.950 91.950 310.050 94.050 ;
        RECT 293.400 91.050 294.450 91.950 ;
        RECT 286.950 89.850 289.050 90.750 ;
        RECT 292.950 88.950 295.050 91.050 ;
        RECT 295.950 88.950 298.050 91.050 ;
        RECT 292.950 79.950 295.050 82.050 ;
        RECT 268.950 56.250 271.050 57.150 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 293.400 55.050 294.450 79.950 ;
        RECT 296.400 55.050 297.450 88.950 ;
        RECT 305.400 64.050 306.450 91.950 ;
        RECT 308.400 67.050 309.450 91.950 ;
        RECT 323.400 90.450 324.450 94.950 ;
        RECT 325.950 92.250 327.750 93.150 ;
        RECT 328.950 91.950 331.050 94.050 ;
        RECT 332.250 92.250 334.050 93.150 ;
        RECT 325.950 90.450 328.050 91.050 ;
        RECT 323.400 89.400 328.050 90.450 ;
        RECT 329.250 89.850 330.750 90.750 ;
        RECT 331.950 90.450 334.050 91.050 ;
        RECT 335.400 90.450 336.450 100.950 ;
        RECT 344.400 97.050 345.450 115.950 ;
        RECT 353.400 112.050 354.450 124.950 ;
        RECT 356.400 118.050 357.450 211.950 ;
        RECT 361.950 207.300 364.050 209.400 ;
        RECT 362.250 203.700 363.450 207.300 ;
        RECT 361.950 201.600 364.050 203.700 ;
        RECT 362.250 189.600 363.450 201.600 ;
        RECT 364.950 193.950 367.050 196.050 ;
        RECT 364.950 191.850 367.050 192.750 ;
        RECT 361.950 187.500 364.050 189.600 ;
        RECT 377.400 184.050 378.450 244.950 ;
        RECT 382.950 238.950 385.050 241.050 ;
        RECT 383.400 238.050 384.450 238.950 ;
        RECT 382.950 235.950 385.050 238.050 ;
        RECT 388.950 235.950 391.050 238.050 ;
        RECT 392.250 236.250 394.050 237.150 ;
        RECT 382.950 233.850 384.750 234.750 ;
        RECT 385.950 232.950 388.050 235.050 ;
        RECT 389.250 233.850 390.750 234.750 ;
        RECT 391.950 232.950 394.050 235.050 ;
        RECT 385.950 230.850 388.050 231.750 ;
        RECT 382.950 201.450 385.050 202.050 ;
        RECT 380.400 200.400 385.050 201.450 ;
        RECT 388.950 201.450 391.050 202.050 ;
        RECT 380.400 196.050 381.450 200.400 ;
        RECT 382.950 199.950 385.050 200.400 ;
        RECT 386.250 200.250 387.750 201.150 ;
        RECT 388.950 200.400 393.450 201.450 ;
        RECT 388.950 199.950 391.050 200.400 ;
        RECT 382.950 197.850 384.750 198.750 ;
        RECT 385.950 196.950 388.050 199.050 ;
        RECT 389.250 197.850 391.050 198.750 ;
        RECT 379.950 193.950 382.050 196.050 ;
        RECT 376.950 181.950 379.050 184.050 ;
        RECT 380.400 172.050 381.450 193.950 ;
        RECT 392.400 178.050 393.450 200.400 ;
        RECT 391.950 175.950 394.050 178.050 ;
        RECT 379.950 171.450 382.050 172.050 ;
        RECT 377.400 170.400 382.050 171.450 ;
        RECT 358.950 166.950 361.050 169.050 ;
        RECT 359.400 162.450 360.450 166.950 ;
        RECT 361.950 164.250 363.750 165.150 ;
        RECT 364.950 163.950 367.050 166.050 ;
        RECT 368.250 164.250 370.050 165.150 ;
        RECT 361.950 162.450 364.050 163.050 ;
        RECT 359.400 161.400 364.050 162.450 ;
        RECT 365.250 161.850 366.750 162.750 ;
        RECT 361.950 160.950 364.050 161.400 ;
        RECT 367.950 160.950 370.050 163.050 ;
        RECT 367.950 131.250 370.050 132.150 ;
        RECT 364.950 128.250 366.750 129.150 ;
        RECT 367.950 127.950 370.050 130.050 ;
        RECT 371.250 128.250 372.750 129.150 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 377.400 127.050 378.450 170.400 ;
        RECT 379.950 169.950 382.050 170.400 ;
        RECT 392.400 169.050 393.450 175.950 ;
        RECT 395.400 172.050 396.450 250.950 ;
        RECT 398.400 196.050 399.450 263.400 ;
        RECT 416.400 259.050 417.450 271.950 ;
        RECT 428.400 271.050 429.450 310.950 ;
        RECT 433.950 307.950 436.050 310.050 ;
        RECT 434.400 307.050 435.450 307.950 ;
        RECT 433.950 304.950 436.050 307.050 ;
        RECT 418.950 268.950 421.050 271.050 ;
        RECT 424.950 269.250 427.050 270.150 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 430.950 269.250 433.050 270.150 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 400.950 235.950 403.050 238.050 ;
        RECT 406.950 236.250 408.750 237.150 ;
        RECT 409.950 235.950 412.050 238.050 ;
        RECT 413.250 236.250 415.050 237.150 ;
        RECT 401.400 232.050 402.450 235.950 ;
        RECT 406.950 232.950 409.050 235.050 ;
        RECT 410.250 233.850 411.750 234.750 ;
        RECT 412.950 232.950 415.050 235.050 ;
        RECT 400.950 229.950 403.050 232.050 ;
        RECT 413.400 229.050 414.450 232.950 ;
        RECT 412.950 226.950 415.050 229.050 ;
        RECT 416.400 225.450 417.450 256.950 ;
        RECT 413.400 224.400 417.450 225.450 ;
        RECT 400.950 200.250 403.050 201.150 ;
        RECT 400.950 196.950 403.050 199.050 ;
        RECT 404.250 197.250 405.750 198.150 ;
        RECT 406.950 196.950 409.050 199.050 ;
        RECT 410.250 197.250 412.050 198.150 ;
        RECT 413.400 196.050 414.450 224.400 ;
        RECT 415.950 196.950 418.050 199.050 ;
        RECT 397.950 193.950 400.050 196.050 ;
        RECT 403.950 193.950 406.050 196.050 ;
        RECT 407.250 194.850 408.750 195.750 ;
        RECT 409.950 193.950 412.050 196.050 ;
        RECT 412.950 193.950 415.050 196.050 ;
        RECT 410.400 178.050 411.450 193.950 ;
        RECT 409.950 175.950 412.050 178.050 ;
        RECT 410.400 175.050 411.450 175.950 ;
        RECT 409.950 172.950 412.050 175.050 ;
        RECT 412.950 173.400 415.050 175.500 ;
        RECT 394.950 169.950 397.050 172.050 ;
        RECT 400.950 169.950 403.050 172.050 ;
        RECT 409.950 170.250 412.050 171.150 ;
        RECT 395.400 169.050 396.450 169.950 ;
        RECT 401.400 169.050 402.450 169.950 ;
        RECT 379.950 167.850 382.050 168.750 ;
        RECT 382.950 167.250 385.050 168.150 ;
        RECT 391.950 166.950 394.050 169.050 ;
        RECT 394.950 166.950 397.050 169.050 ;
        RECT 400.950 166.950 403.050 169.050 ;
        RECT 409.950 166.950 412.050 169.050 ;
        RECT 382.950 163.950 385.050 166.050 ;
        RECT 394.950 164.850 397.050 165.750 ;
        RECT 400.950 164.850 403.050 165.750 ;
        RECT 383.400 157.050 384.450 163.950 ;
        RECT 410.400 163.050 411.450 166.950 ;
        RECT 409.950 160.950 412.050 163.050 ;
        RECT 413.550 161.400 414.750 173.400 ;
        RECT 416.400 166.050 417.450 196.950 ;
        RECT 419.400 193.050 420.450 268.950 ;
        RECT 430.950 265.950 433.050 268.050 ;
        RECT 433.950 244.950 436.050 247.050 ;
        RECT 434.400 238.050 435.450 244.950 ;
        RECT 430.950 236.250 432.750 237.150 ;
        RECT 433.950 235.950 436.050 238.050 ;
        RECT 437.400 235.050 438.450 335.400 ;
        RECT 443.400 322.050 444.450 341.400 ;
        RECT 446.400 340.050 447.450 406.950 ;
        RECT 449.400 406.050 450.450 409.950 ;
        RECT 448.950 403.950 451.050 406.050 ;
        RECT 449.400 397.050 450.450 403.950 ;
        RECT 448.950 394.950 451.050 397.050 ;
        RECT 455.400 387.450 456.450 436.950 ;
        RECT 461.400 424.050 462.450 445.950 ;
        RECT 460.950 421.950 463.050 424.050 ;
        RECT 461.400 415.050 462.450 421.950 ;
        RECT 460.950 414.450 463.050 415.050 ;
        RECT 452.400 386.400 456.450 387.450 ;
        RECT 458.400 413.400 463.050 414.450 ;
        RECT 452.400 385.050 453.450 386.400 ;
        RECT 451.950 382.950 454.050 385.050 ;
        RECT 455.250 383.250 457.050 384.150 ;
        RECT 451.950 380.850 453.750 381.750 ;
        RECT 454.950 379.950 457.050 382.050 ;
        RECT 455.400 370.050 456.450 379.950 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 458.400 361.050 459.450 413.400 ;
        RECT 460.950 412.950 463.050 413.400 ;
        RECT 464.250 413.250 466.050 414.150 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 473.250 413.250 475.050 414.150 ;
        RECT 460.950 410.850 462.750 411.750 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 466.950 409.950 469.050 412.050 ;
        RECT 469.950 410.850 471.750 411.750 ;
        RECT 472.950 409.950 475.050 412.050 ;
        RECT 460.950 385.950 463.050 388.050 ;
        RECT 461.400 385.050 462.450 385.950 ;
        RECT 460.950 382.950 463.050 385.050 ;
        RECT 464.250 383.250 466.050 384.150 ;
        RECT 460.950 380.850 462.750 381.750 ;
        RECT 463.950 381.450 466.050 382.050 ;
        RECT 467.400 381.450 468.450 409.950 ;
        RECT 473.400 403.050 474.450 409.950 ;
        RECT 472.950 400.950 475.050 403.050 ;
        RECT 476.400 387.450 477.450 454.950 ;
        RECT 479.400 453.450 480.450 454.950 ;
        RECT 481.950 453.450 484.050 454.050 ;
        RECT 479.400 452.400 484.050 453.450 ;
        RECT 479.400 451.050 480.450 452.400 ;
        RECT 481.950 451.950 484.050 452.400 ;
        RECT 485.400 451.050 486.450 454.950 ;
        RECT 487.950 451.950 490.050 454.050 ;
        RECT 491.250 452.250 493.050 453.150 ;
        RECT 478.950 448.950 481.050 451.050 ;
        RECT 481.950 449.850 483.750 450.750 ;
        RECT 484.950 448.950 487.050 451.050 ;
        RECT 488.250 449.850 489.750 450.750 ;
        RECT 490.950 450.450 493.050 451.050 ;
        RECT 494.400 450.450 495.450 478.950 ;
        RECT 503.400 472.050 504.450 484.950 ;
        RECT 502.950 469.950 505.050 472.050 ;
        RECT 503.400 463.050 504.450 469.950 ;
        RECT 502.950 460.950 505.050 463.050 ;
        RECT 499.950 454.950 502.050 457.050 ;
        RECT 506.400 456.450 507.450 488.400 ;
        RECT 508.950 487.950 511.050 490.050 ;
        RECT 511.950 488.250 514.050 489.150 ;
        RECT 514.950 487.950 517.050 490.050 ;
        RECT 509.400 486.450 510.450 487.950 ;
        RECT 518.400 487.050 519.450 493.950 ;
        RECT 511.950 486.450 514.050 487.050 ;
        RECT 509.400 485.400 514.050 486.450 ;
        RECT 511.950 484.950 514.050 485.400 ;
        RECT 515.250 485.250 516.750 486.150 ;
        RECT 517.950 484.950 520.050 487.050 ;
        RECT 521.250 485.250 523.050 486.150 ;
        RECT 508.950 472.950 511.050 475.050 ;
        RECT 503.400 455.400 507.450 456.450 ;
        RECT 490.950 449.400 495.450 450.450 ;
        RECT 490.950 448.950 493.050 449.400 ;
        RECT 479.400 412.050 480.450 448.950 ;
        RECT 484.950 446.850 487.050 447.750 ;
        RECT 484.950 418.950 487.050 421.050 ;
        RECT 481.950 415.950 484.050 418.050 ;
        RECT 478.950 409.950 481.050 412.050 ;
        RECT 463.950 380.400 468.450 381.450 ;
        RECT 473.400 386.400 477.450 387.450 ;
        RECT 463.950 379.950 466.050 380.400 ;
        RECT 464.400 379.050 465.450 379.950 ;
        RECT 463.950 376.950 466.050 379.050 ;
        RECT 457.950 358.950 460.050 361.050 ;
        RECT 469.950 358.950 472.050 361.050 ;
        RECT 448.950 355.950 451.050 358.050 ;
        RECT 445.950 337.950 448.050 340.050 ;
        RECT 449.400 339.450 450.450 355.950 ;
        RECT 454.950 343.950 457.050 346.050 ;
        RECT 455.400 343.050 456.450 343.950 ;
        RECT 451.950 341.250 453.750 342.150 ;
        RECT 454.950 340.950 457.050 343.050 ;
        RECT 457.950 340.950 460.050 343.050 ;
        RECT 463.950 342.450 466.050 343.050 ;
        RECT 460.950 341.250 462.750 342.150 ;
        RECT 463.950 341.400 468.450 342.450 ;
        RECT 463.950 340.950 466.050 341.400 ;
        RECT 451.950 339.450 454.050 340.050 ;
        RECT 449.400 338.400 454.050 339.450 ;
        RECT 455.250 338.850 457.050 339.750 ;
        RECT 451.950 337.950 454.050 338.400 ;
        RECT 445.950 328.950 448.050 331.050 ;
        RECT 442.950 319.950 445.050 322.050 ;
        RECT 439.950 316.950 442.050 319.050 ;
        RECT 440.400 277.050 441.450 316.950 ;
        RECT 446.400 313.050 447.450 328.950 ;
        RECT 445.950 310.950 448.050 313.050 ;
        RECT 451.950 310.950 454.050 313.050 ;
        RECT 445.950 308.850 448.050 309.750 ;
        RECT 451.950 308.850 454.050 309.750 ;
        RECT 439.950 274.950 442.050 277.050 ;
        RECT 448.950 268.950 451.050 271.050 ;
        RECT 448.950 266.850 451.050 267.750 ;
        RECT 451.950 244.950 454.050 247.050 ;
        RECT 439.950 241.950 442.050 244.050 ;
        RECT 440.400 238.050 441.450 241.950 ;
        RECT 439.950 235.950 442.050 238.050 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 448.950 235.950 451.050 238.050 ;
        RECT 430.950 232.950 433.050 235.050 ;
        RECT 434.250 233.850 435.750 234.750 ;
        RECT 436.950 232.950 439.050 235.050 ;
        RECT 440.250 233.850 442.050 234.750 ;
        RECT 431.400 232.050 432.450 232.950 ;
        RECT 430.950 229.950 433.050 232.050 ;
        RECT 436.950 230.850 439.050 231.750 ;
        RECT 446.400 208.050 447.450 235.950 ;
        RECT 449.400 229.050 450.450 235.950 ;
        RECT 452.400 234.450 453.450 244.950 ;
        RECT 458.400 241.050 459.450 340.950 ;
        RECT 467.400 340.050 468.450 341.400 ;
        RECT 460.950 337.950 463.050 340.050 ;
        RECT 464.250 338.850 466.050 339.750 ;
        RECT 466.950 337.950 469.050 340.050 ;
        RECT 470.400 313.050 471.450 358.950 ;
        RECT 473.400 349.050 474.450 386.400 ;
        RECT 478.950 384.450 481.050 385.050 ;
        RECT 482.400 384.450 483.450 415.950 ;
        RECT 485.400 388.050 486.450 418.950 ;
        RECT 487.950 413.250 490.050 414.150 ;
        RECT 493.950 413.250 496.050 414.150 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 487.950 388.950 490.050 391.050 ;
        RECT 490.950 388.950 493.050 391.050 ;
        RECT 484.950 385.950 487.050 388.050 ;
        RECT 488.400 385.050 489.450 388.950 ;
        RECT 475.950 383.250 477.750 384.150 ;
        RECT 478.950 383.400 483.450 384.450 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 484.950 383.250 486.750 384.150 ;
        RECT 487.950 382.950 490.050 385.050 ;
        RECT 475.950 379.950 478.050 382.050 ;
        RECT 479.250 380.850 481.050 381.750 ;
        RECT 484.950 379.950 487.050 382.050 ;
        RECT 488.250 380.850 490.050 381.750 ;
        RECT 476.400 367.050 477.450 379.950 ;
        RECT 475.950 364.950 478.050 367.050 ;
        RECT 472.950 346.950 475.050 349.050 ;
        RECT 472.950 341.250 475.050 342.150 ;
        RECT 478.950 341.250 481.050 342.150 ;
        RECT 478.950 337.950 481.050 340.050 ;
        RECT 485.400 331.050 486.450 379.950 ;
        RECT 491.400 348.450 492.450 388.950 ;
        RECT 500.400 388.050 501.450 454.950 ;
        RECT 503.400 391.050 504.450 455.400 ;
        RECT 509.400 454.050 510.450 472.950 ;
        RECT 512.400 457.050 513.450 484.950 ;
        RECT 524.400 484.050 525.450 517.950 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 518.250 482.850 519.750 483.750 ;
        RECT 520.950 481.950 523.050 484.050 ;
        RECT 523.950 481.950 526.050 484.050 ;
        RECT 521.400 481.050 522.450 481.950 ;
        RECT 514.950 478.950 517.050 481.050 ;
        RECT 520.950 478.950 523.050 481.050 ;
        RECT 527.400 480.450 528.450 521.400 ;
        RECT 529.950 520.950 532.050 521.400 ;
        RECT 536.400 520.050 537.450 598.950 ;
        RECT 539.400 574.050 540.450 622.950 ;
        RECT 541.950 610.950 544.050 613.050 ;
        RECT 542.400 601.050 543.450 610.950 ;
        RECT 544.950 604.950 547.050 607.050 ;
        RECT 545.400 604.050 546.450 604.950 ;
        RECT 548.400 604.050 549.450 625.950 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 541.950 598.950 544.050 601.050 ;
        RECT 545.250 599.850 546.750 600.750 ;
        RECT 547.950 598.950 550.050 601.050 ;
        RECT 541.950 596.850 544.050 597.750 ;
        RECT 547.950 596.850 550.050 597.750 ;
        RECT 538.950 571.950 541.050 574.050 ;
        RECT 557.400 562.050 558.450 625.950 ;
        RECT 575.400 625.050 576.450 673.950 ;
        RECT 577.950 670.950 580.050 673.050 ;
        RECT 578.400 666.450 579.450 670.950 ;
        RECT 584.400 670.050 585.450 688.950 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 580.950 668.250 582.750 669.150 ;
        RECT 583.950 667.950 586.050 670.050 ;
        RECT 587.250 668.250 589.050 669.150 ;
        RECT 580.950 666.450 583.050 667.050 ;
        RECT 578.400 665.400 583.050 666.450 ;
        RECT 584.250 665.850 585.750 666.750 ;
        RECT 559.950 622.950 562.050 625.050 ;
        RECT 574.950 622.950 577.050 625.050 ;
        RECT 562.950 610.950 565.050 613.050 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 559.950 596.850 562.050 597.750 ;
        RECT 563.400 594.450 564.450 610.950 ;
        RECT 568.950 607.950 571.050 610.050 ;
        RECT 569.400 601.050 570.450 607.950 ;
        RECT 568.950 598.950 571.050 601.050 ;
        RECT 565.950 596.250 568.050 597.150 ;
        RECT 568.950 596.850 571.050 597.750 ;
        RECT 565.950 594.450 568.050 595.050 ;
        RECT 563.400 593.400 568.050 594.450 ;
        RECT 565.950 592.950 568.050 593.400 ;
        RECT 574.950 571.950 577.050 574.050 ;
        RECT 568.950 563.250 571.050 564.150 ;
        RECT 575.400 562.050 576.450 571.950 ;
        RECT 556.950 559.950 559.050 562.050 ;
        RECT 565.950 560.250 567.750 561.150 ;
        RECT 568.950 559.950 571.050 562.050 ;
        RECT 572.250 560.250 573.750 561.150 ;
        RECT 574.950 559.950 577.050 562.050 ;
        RECT 547.950 557.250 549.750 558.150 ;
        RECT 550.950 556.950 553.050 559.050 ;
        RECT 556.950 556.950 559.050 559.050 ;
        RECT 565.950 556.950 568.050 559.050 ;
        RECT 566.400 556.050 567.450 556.950 ;
        RECT 544.950 553.950 547.050 556.050 ;
        RECT 547.950 553.950 550.050 556.050 ;
        RECT 551.250 554.850 553.050 555.750 ;
        RECT 553.950 554.250 556.050 555.150 ;
        RECT 556.950 554.850 559.050 555.750 ;
        RECT 565.950 553.950 568.050 556.050 ;
        RECT 545.400 547.050 546.450 553.950 ;
        RECT 553.950 550.950 556.050 553.050 ;
        RECT 554.400 547.050 555.450 550.950 ;
        RECT 544.950 544.950 547.050 547.050 ;
        RECT 553.950 544.950 556.050 547.050 ;
        RECT 553.950 541.950 556.050 544.050 ;
        RECT 550.950 535.950 553.050 538.050 ;
        RECT 544.950 532.950 547.050 535.050 ;
        RECT 535.950 517.950 538.050 520.050 ;
        RECT 532.950 487.950 535.050 490.050 ;
        RECT 538.950 488.250 541.050 489.150 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 533.400 487.050 534.450 487.950 ;
        RECT 529.950 485.250 531.750 486.150 ;
        RECT 532.950 484.950 535.050 487.050 ;
        RECT 536.250 485.250 537.750 486.150 ;
        RECT 538.950 484.950 541.050 487.050 ;
        RECT 529.950 481.950 532.050 484.050 ;
        RECT 533.250 482.850 534.750 483.750 ;
        RECT 535.950 481.950 538.050 484.050 ;
        RECT 524.400 479.400 528.450 480.450 ;
        RECT 515.400 457.050 516.450 478.950 ;
        RECT 524.400 475.050 525.450 479.400 ;
        RECT 526.950 475.950 529.050 478.050 ;
        RECT 523.950 472.950 526.050 475.050 ;
        RECT 511.950 454.950 514.050 457.050 ;
        RECT 514.950 454.950 517.050 457.050 ;
        RECT 505.950 452.250 507.750 453.150 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 512.250 452.250 514.050 453.150 ;
        RECT 505.950 448.950 508.050 451.050 ;
        RECT 509.250 449.850 510.750 450.750 ;
        RECT 511.950 448.950 514.050 451.050 ;
        RECT 506.400 448.050 507.450 448.950 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 505.950 442.950 508.050 445.050 ;
        RECT 506.400 415.050 507.450 442.950 ;
        RECT 512.400 430.050 513.450 448.950 ;
        RECT 515.400 448.050 516.450 454.950 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 511.950 427.950 514.050 430.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 505.950 410.850 508.050 411.750 ;
        RECT 508.950 410.250 511.050 411.150 ;
        RECT 508.950 406.950 511.050 409.050 ;
        RECT 509.400 406.050 510.450 406.950 ;
        RECT 508.950 403.950 511.050 406.050 ;
        RECT 508.950 391.950 511.050 394.050 ;
        RECT 502.950 388.950 505.050 391.050 ;
        RECT 499.950 385.950 502.050 388.050 ;
        RECT 500.400 349.050 501.450 385.950 ;
        RECT 509.400 385.050 510.450 391.950 ;
        RECT 508.950 382.950 511.050 385.050 ;
        RECT 502.950 380.850 505.050 381.750 ;
        RECT 508.950 380.850 511.050 381.750 ;
        RECT 512.400 378.450 513.450 412.950 ;
        RECT 515.400 409.050 516.450 445.950 ;
        RECT 517.950 424.950 520.050 427.050 ;
        RECT 518.400 414.450 519.450 424.950 ;
        RECT 527.400 421.050 528.450 475.950 ;
        RECT 530.400 460.050 531.450 481.950 ;
        RECT 529.950 457.950 532.050 460.050 ;
        RECT 532.950 459.450 535.050 460.050 ;
        RECT 532.950 458.400 537.450 459.450 ;
        RECT 532.950 457.950 535.050 458.400 ;
        RECT 529.950 455.250 532.050 456.150 ;
        RECT 532.950 455.850 535.050 456.750 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 536.400 451.050 537.450 458.400 ;
        RECT 539.400 451.050 540.450 484.950 ;
        RECT 542.400 454.050 543.450 487.950 ;
        RECT 545.400 484.050 546.450 532.950 ;
        RECT 547.950 526.950 550.050 529.050 ;
        RECT 548.400 523.050 549.450 526.950 ;
        RECT 551.400 526.050 552.450 535.950 ;
        RECT 554.400 529.050 555.450 541.950 ;
        RECT 566.400 541.050 567.450 553.950 ;
        RECT 569.400 547.050 570.450 559.950 ;
        RECT 571.950 556.950 574.050 559.050 ;
        RECT 575.250 557.850 577.050 558.750 ;
        RECT 568.950 544.950 571.050 547.050 ;
        RECT 565.950 538.950 568.050 541.050 ;
        RECT 574.950 538.950 577.050 541.050 ;
        RECT 568.950 535.950 571.050 538.050 ;
        RECT 559.950 529.950 562.050 532.050 ;
        RECT 560.400 529.050 561.450 529.950 ;
        RECT 553.950 526.950 556.050 529.050 ;
        RECT 557.250 527.250 558.750 528.150 ;
        RECT 559.950 526.950 562.050 529.050 ;
        RECT 550.950 523.950 553.050 526.050 ;
        RECT 554.250 524.850 555.750 525.750 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 560.250 524.850 562.050 525.750 ;
        RECT 547.950 520.950 550.050 523.050 ;
        RECT 550.950 521.850 553.050 522.750 ;
        RECT 548.400 484.050 549.450 520.950 ;
        RECT 553.950 493.950 556.050 496.050 ;
        RECT 554.400 486.450 555.450 493.950 ;
        RECT 556.950 488.250 559.050 489.150 ;
        RECT 556.950 486.450 559.050 487.050 ;
        RECT 554.400 485.400 559.050 486.450 ;
        RECT 556.950 484.950 559.050 485.400 ;
        RECT 560.250 485.250 561.750 486.150 ;
        RECT 562.950 484.950 565.050 487.050 ;
        RECT 566.250 485.250 568.050 486.150 ;
        RECT 544.950 481.950 547.050 484.050 ;
        RECT 547.950 481.950 550.050 484.050 ;
        RECT 556.950 481.950 559.050 484.050 ;
        RECT 559.950 481.950 562.050 484.050 ;
        RECT 563.250 482.850 564.750 483.750 ;
        RECT 565.950 481.950 568.050 484.050 ;
        RECT 547.950 466.950 550.050 469.050 ;
        RECT 548.400 457.050 549.450 466.950 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 547.950 454.950 550.050 457.050 ;
        RECT 551.250 455.250 552.750 456.150 ;
        RECT 553.950 454.950 556.050 457.050 ;
        RECT 545.400 454.050 546.450 454.950 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 544.950 451.950 547.050 454.050 ;
        RECT 548.250 452.850 549.750 453.750 ;
        RECT 550.950 451.950 553.050 454.050 ;
        RECT 554.250 452.850 556.050 453.750 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 538.950 448.950 541.050 451.050 ;
        RECT 544.950 449.850 547.050 450.750 ;
        RECT 553.950 448.950 556.050 451.050 ;
        RECT 526.950 418.950 529.050 421.050 ;
        RECT 544.950 418.950 547.050 421.050 ;
        RECT 547.950 418.950 550.050 421.050 ;
        RECT 545.400 418.050 546.450 418.950 ;
        RECT 520.950 416.250 523.050 417.150 ;
        RECT 526.950 415.950 529.050 418.050 ;
        RECT 538.950 417.450 541.050 418.050 ;
        RECT 536.400 416.400 541.050 417.450 ;
        RECT 527.400 415.050 528.450 415.950 ;
        RECT 520.950 414.450 523.050 415.050 ;
        RECT 518.400 413.400 523.050 414.450 ;
        RECT 520.950 412.950 523.050 413.400 ;
        RECT 524.250 413.250 525.750 414.150 ;
        RECT 526.950 412.950 529.050 415.050 ;
        RECT 530.250 413.250 532.050 414.150 ;
        RECT 520.950 409.950 523.050 412.050 ;
        RECT 523.950 409.950 526.050 412.050 ;
        RECT 527.250 410.850 528.750 411.750 ;
        RECT 529.950 409.950 532.050 412.050 ;
        RECT 514.950 406.950 517.050 409.050 ;
        RECT 509.400 377.400 513.450 378.450 ;
        RECT 488.400 347.400 492.450 348.450 ;
        RECT 488.400 336.450 489.450 347.400 ;
        RECT 493.950 347.250 496.050 348.150 ;
        RECT 499.950 346.950 502.050 349.050 ;
        RECT 490.950 344.250 492.750 345.150 ;
        RECT 493.950 343.950 496.050 346.050 ;
        RECT 499.950 345.450 502.050 346.050 ;
        RECT 497.250 344.250 498.750 345.150 ;
        RECT 499.950 344.400 504.450 345.450 ;
        RECT 499.950 343.950 502.050 344.400 ;
        RECT 490.950 340.950 493.050 343.050 ;
        RECT 496.950 340.950 499.050 343.050 ;
        RECT 500.250 341.850 502.050 342.750 ;
        RECT 488.400 335.400 492.450 336.450 ;
        RECT 484.950 328.950 487.050 331.050 ;
        RECT 491.400 319.050 492.450 335.400 ;
        RECT 497.400 331.050 498.450 340.950 ;
        RECT 496.950 328.950 499.050 331.050 ;
        RECT 503.400 322.050 504.450 344.400 ;
        RECT 509.400 342.450 510.450 377.400 ;
        RECT 511.950 346.950 514.050 349.050 ;
        RECT 506.400 341.400 510.450 342.450 ;
        RECT 502.950 319.950 505.050 322.050 ;
        RECT 490.950 316.950 493.050 319.050 ;
        RECT 499.950 313.950 502.050 316.050 ;
        RECT 469.950 310.950 472.050 313.050 ;
        RECT 469.950 308.250 471.750 309.150 ;
        RECT 472.950 307.950 475.050 310.050 ;
        RECT 476.250 308.250 478.050 309.150 ;
        RECT 478.950 307.950 481.050 310.050 ;
        RECT 490.950 308.250 492.750 309.150 ;
        RECT 493.950 307.950 496.050 310.050 ;
        RECT 497.250 308.250 499.050 309.150 ;
        RECT 469.950 304.950 472.050 307.050 ;
        RECT 473.250 305.850 474.750 306.750 ;
        RECT 475.950 304.950 478.050 307.050 ;
        RECT 476.400 304.050 477.450 304.950 ;
        RECT 475.950 301.950 478.050 304.050 ;
        RECT 479.400 301.050 480.450 307.950 ;
        RECT 490.950 304.950 493.050 307.050 ;
        RECT 494.250 305.850 495.750 306.750 ;
        RECT 496.950 304.950 499.050 307.050 ;
        RECT 478.950 298.950 481.050 301.050 ;
        RECT 497.400 289.050 498.450 304.950 ;
        RECT 496.950 286.950 499.050 289.050 ;
        RECT 500.400 276.450 501.450 313.950 ;
        RECT 506.400 307.050 507.450 341.400 ;
        RECT 508.950 316.950 511.050 319.050 ;
        RECT 509.400 313.050 510.450 316.950 ;
        RECT 512.400 316.050 513.450 346.950 ;
        RECT 515.400 340.050 516.450 406.950 ;
        RECT 521.400 343.050 522.450 409.950 ;
        RECT 524.400 406.050 525.450 409.950 ;
        RECT 523.950 403.950 526.050 406.050 ;
        RECT 530.400 400.050 531.450 409.950 ;
        RECT 529.950 397.950 532.050 400.050 ;
        RECT 532.950 397.950 535.050 400.050 ;
        RECT 526.950 385.950 529.050 388.050 ;
        RECT 527.400 382.050 528.450 385.950 ;
        RECT 523.950 380.250 525.750 381.150 ;
        RECT 526.950 379.950 529.050 382.050 ;
        RECT 530.250 380.250 532.050 381.150 ;
        RECT 523.950 376.950 526.050 379.050 ;
        RECT 527.250 377.850 528.750 378.750 ;
        RECT 529.950 378.450 532.050 379.050 ;
        RECT 533.400 378.450 534.450 397.950 ;
        RECT 536.400 394.050 537.450 416.400 ;
        RECT 538.950 415.950 541.050 416.400 ;
        RECT 542.250 416.250 543.750 417.150 ;
        RECT 544.950 415.950 547.050 418.050 ;
        RECT 538.950 413.850 540.750 414.750 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 545.250 413.850 547.050 414.750 ;
        RECT 535.950 391.950 538.050 394.050 ;
        RECT 548.400 385.050 549.450 418.950 ;
        RECT 547.950 382.950 550.050 385.050 ;
        RECT 551.250 383.250 553.050 384.150 ;
        RECT 547.950 380.850 549.750 381.750 ;
        RECT 550.950 379.950 553.050 382.050 ;
        RECT 529.950 377.400 534.450 378.450 ;
        RECT 529.950 376.950 532.050 377.400 ;
        RECT 524.400 352.050 525.450 376.950 ;
        RECT 551.400 373.050 552.450 379.950 ;
        RECT 550.950 370.950 553.050 373.050 ;
        RECT 523.950 349.950 526.050 352.050 ;
        RECT 554.400 343.050 555.450 448.950 ;
        RECT 557.400 412.050 558.450 481.950 ;
        RECT 566.400 460.050 567.450 481.950 ;
        RECT 569.400 465.450 570.450 535.950 ;
        RECT 575.400 532.050 576.450 538.950 ;
        RECT 574.950 529.950 577.050 532.050 ;
        RECT 571.950 527.250 574.050 528.150 ;
        RECT 574.950 527.850 577.050 528.750 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 572.400 523.050 573.450 523.950 ;
        RECT 571.950 520.950 574.050 523.050 ;
        RECT 571.950 517.950 574.050 520.050 ;
        RECT 572.400 484.050 573.450 517.950 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 575.400 483.450 576.450 523.950 ;
        RECT 578.400 490.050 579.450 665.400 ;
        RECT 580.950 664.950 583.050 665.400 ;
        RECT 586.950 664.950 589.050 667.050 ;
        RECT 587.400 664.050 588.450 664.950 ;
        RECT 586.950 661.950 589.050 664.050 ;
        RECT 580.950 628.950 583.050 631.050 ;
        RECT 580.950 626.850 583.050 627.750 ;
        RECT 583.950 626.250 586.050 627.150 ;
        RECT 583.950 622.950 586.050 625.050 ;
        RECT 584.400 607.050 585.450 622.950 ;
        RECT 583.950 604.950 586.050 607.050 ;
        RECT 593.400 601.050 594.450 679.950 ;
        RECT 598.950 673.950 601.050 676.050 ;
        RECT 598.950 671.850 601.050 672.750 ;
        RECT 601.950 671.250 604.050 672.150 ;
        RECT 601.950 667.950 604.050 670.050 ;
        RECT 605.400 661.050 606.450 725.400 ;
        RECT 622.950 715.950 625.050 718.050 ;
        RECT 607.950 710.400 610.050 712.500 ;
        RECT 608.400 693.600 609.600 710.400 ;
        RECT 616.950 703.950 619.050 706.050 ;
        RECT 613.950 701.250 616.050 702.150 ;
        RECT 613.950 697.950 616.050 700.050 ;
        RECT 607.950 691.500 610.050 693.600 ;
        RECT 610.950 691.950 613.050 694.050 ;
        RECT 611.400 672.450 612.450 691.950 ;
        RECT 617.400 687.450 618.450 703.950 ;
        RECT 619.950 701.250 622.050 702.150 ;
        RECT 619.950 697.950 622.050 700.050 ;
        RECT 620.400 691.050 621.450 697.950 ;
        RECT 619.950 688.950 622.050 691.050 ;
        RECT 617.400 686.400 621.450 687.450 ;
        RECT 620.400 673.050 621.450 686.400 ;
        RECT 613.950 672.450 616.050 673.050 ;
        RECT 611.400 671.400 616.050 672.450 ;
        RECT 604.950 658.950 607.050 661.050 ;
        RECT 595.950 632.250 598.050 633.150 ;
        RECT 595.950 628.950 598.050 631.050 ;
        RECT 599.250 629.250 600.750 630.150 ;
        RECT 601.950 628.950 604.050 631.050 ;
        RECT 605.250 629.250 607.050 630.150 ;
        RECT 598.950 625.950 601.050 628.050 ;
        RECT 602.250 626.850 603.750 627.750 ;
        RECT 604.950 625.950 607.050 628.050 ;
        RECT 605.400 613.050 606.450 625.950 ;
        RECT 604.950 610.950 607.050 613.050 ;
        RECT 611.400 612.450 612.450 671.400 ;
        RECT 613.950 670.950 616.050 671.400 ;
        RECT 617.250 671.250 618.750 672.150 ;
        RECT 619.950 670.950 622.050 673.050 ;
        RECT 623.400 670.050 624.450 715.950 ;
        RECT 628.950 711.300 631.050 713.400 ;
        RECT 629.250 707.700 630.450 711.300 ;
        RECT 628.950 705.600 631.050 707.700 ;
        RECT 650.400 706.050 651.450 737.400 ;
        RECT 656.400 736.050 657.450 772.950 ;
        RECT 659.400 772.050 660.450 778.950 ;
        RECT 665.400 772.050 666.450 808.950 ;
        RECT 671.400 784.050 672.450 812.400 ;
        RECT 676.950 811.950 679.050 814.050 ;
        RECT 680.400 787.050 681.450 815.400 ;
        RECT 682.950 814.950 685.050 815.400 ;
        RECT 686.250 815.250 687.750 816.150 ;
        RECT 688.950 814.950 691.050 817.050 ;
        RECT 703.950 816.450 706.050 817.050 ;
        RECT 701.400 815.400 706.050 816.450 ;
        RECT 682.950 812.850 684.750 813.750 ;
        RECT 685.950 811.950 688.050 814.050 ;
        RECT 689.250 812.850 690.750 813.750 ;
        RECT 691.950 811.950 694.050 814.050 ;
        RECT 697.950 811.950 700.050 814.050 ;
        RECT 691.950 809.850 694.050 810.750 ;
        RECT 688.950 796.950 691.050 799.050 ;
        RECT 679.950 784.950 682.050 787.050 ;
        RECT 670.950 781.950 673.050 784.050 ;
        RECT 679.950 781.950 682.050 784.050 ;
        RECT 673.950 775.950 676.050 778.050 ;
        RECT 674.400 775.050 675.450 775.950 ;
        RECT 680.400 775.050 681.450 781.950 ;
        RECT 670.950 773.250 672.750 774.150 ;
        RECT 673.950 772.950 676.050 775.050 ;
        RECT 677.250 773.250 678.750 774.150 ;
        RECT 679.950 772.950 682.050 775.050 ;
        RECT 683.250 773.250 685.050 774.150 ;
        RECT 685.950 772.950 688.050 775.050 ;
        RECT 658.950 769.950 661.050 772.050 ;
        RECT 664.950 769.950 667.050 772.050 ;
        RECT 670.950 769.950 673.050 772.050 ;
        RECT 674.250 770.850 675.750 771.750 ;
        RECT 676.950 769.950 679.050 772.050 ;
        RECT 680.250 770.850 681.750 771.750 ;
        RECT 682.950 771.450 685.050 772.050 ;
        RECT 686.400 771.450 687.450 772.950 ;
        RECT 682.950 770.400 687.450 771.450 ;
        RECT 682.950 769.950 685.050 770.400 ;
        RECT 677.400 769.050 678.450 769.950 ;
        RECT 676.950 766.950 679.050 769.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 664.950 751.950 667.050 754.050 ;
        RECT 665.400 742.050 666.450 751.950 ;
        RECT 661.950 740.250 663.750 741.150 ;
        RECT 664.950 739.950 667.050 742.050 ;
        RECT 668.250 740.250 670.050 741.150 ;
        RECT 661.950 736.950 664.050 739.050 ;
        RECT 665.250 737.850 666.750 738.750 ;
        RECT 667.950 736.950 670.050 739.050 ;
        RECT 655.950 733.950 658.050 736.050 ;
        RECT 661.950 733.950 664.050 736.050 ;
        RECT 629.250 693.600 630.450 705.600 ;
        RECT 631.950 703.950 634.050 706.050 ;
        RECT 643.950 703.950 646.050 706.050 ;
        RECT 647.250 704.250 648.750 705.150 ;
        RECT 649.950 703.950 652.050 706.050 ;
        RECT 632.400 700.050 633.450 703.950 ;
        RECT 643.950 701.850 645.750 702.750 ;
        RECT 646.950 700.950 649.050 703.050 ;
        RECT 650.250 701.850 652.050 702.750 ;
        RECT 631.950 697.950 634.050 700.050 ;
        RECT 652.950 697.950 655.050 700.050 ;
        RECT 655.950 697.950 658.050 700.050 ;
        RECT 631.950 695.850 634.050 696.750 ;
        RECT 628.950 691.500 631.050 693.600 ;
        RECT 625.950 673.950 628.050 676.050 ;
        RECT 637.950 673.950 640.050 676.050 ;
        RECT 613.950 668.850 615.750 669.750 ;
        RECT 616.950 667.950 619.050 670.050 ;
        RECT 620.250 668.850 621.750 669.750 ;
        RECT 622.950 667.950 625.050 670.050 ;
        RECT 622.950 665.850 625.050 666.750 ;
        RECT 622.950 658.950 625.050 661.050 ;
        RECT 616.950 628.950 619.050 631.050 ;
        RECT 616.950 626.850 619.050 627.750 ;
        RECT 619.950 626.250 622.050 627.150 ;
        RECT 619.950 622.950 622.050 625.050 ;
        RECT 613.950 616.950 616.050 619.050 ;
        RECT 608.400 611.400 612.450 612.450 ;
        RECT 608.400 604.050 609.450 611.400 ;
        RECT 614.400 609.450 615.450 616.950 ;
        RECT 611.400 608.400 615.450 609.450 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 611.400 601.050 612.450 608.400 ;
        RECT 586.950 598.950 589.050 601.050 ;
        RECT 590.250 599.250 591.750 600.150 ;
        RECT 592.950 598.950 595.050 601.050 ;
        RECT 601.950 600.450 604.050 601.050 ;
        RECT 604.950 600.450 607.050 601.050 ;
        RECT 601.950 599.400 607.050 600.450 ;
        RECT 601.950 598.950 604.050 599.400 ;
        RECT 604.950 598.950 607.050 599.400 ;
        RECT 608.250 599.250 609.750 600.150 ;
        RECT 610.950 598.950 613.050 601.050 ;
        RECT 583.950 595.950 586.050 598.050 ;
        RECT 587.250 596.850 588.750 597.750 ;
        RECT 589.950 595.950 592.050 598.050 ;
        RECT 593.250 596.850 595.050 597.750 ;
        RECT 583.950 593.850 586.050 594.750 ;
        RECT 590.400 592.050 591.450 595.950 ;
        RECT 583.950 589.950 586.050 592.050 ;
        RECT 589.950 589.950 592.050 592.050 ;
        RECT 584.400 520.050 585.450 589.950 ;
        RECT 589.950 557.250 592.050 558.150 ;
        RECT 595.950 556.950 598.050 559.050 ;
        RECT 586.950 554.250 588.750 555.150 ;
        RECT 589.950 553.950 592.050 556.050 ;
        RECT 595.950 554.850 598.050 555.750 ;
        RECT 586.950 550.950 589.050 553.050 ;
        RECT 587.400 544.050 588.450 550.950 ;
        RECT 590.400 550.050 591.450 553.950 ;
        RECT 602.400 553.050 603.450 598.950 ;
        RECT 604.950 596.850 606.750 597.750 ;
        RECT 607.950 595.950 610.050 598.050 ;
        RECT 611.250 596.850 612.750 597.750 ;
        RECT 613.950 595.950 616.050 598.050 ;
        RECT 608.400 595.050 609.450 595.950 ;
        RECT 607.950 592.950 610.050 595.050 ;
        RECT 613.950 593.850 616.050 594.750 ;
        RECT 616.950 560.250 619.050 561.150 ;
        RECT 604.950 556.950 607.050 559.050 ;
        RECT 607.950 557.250 609.750 558.150 ;
        RECT 610.950 556.950 613.050 559.050 ;
        RECT 614.250 557.250 615.750 558.150 ;
        RECT 616.950 556.950 619.050 559.050 ;
        RECT 601.950 550.950 604.050 553.050 ;
        RECT 589.950 547.950 592.050 550.050 ;
        RECT 598.950 547.950 601.050 550.050 ;
        RECT 586.950 541.950 589.050 544.050 ;
        RECT 586.950 535.950 589.050 538.050 ;
        RECT 587.400 526.050 588.450 535.950 ;
        RECT 586.950 523.950 589.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 596.250 524.250 598.050 525.150 ;
        RECT 586.950 521.850 588.750 522.750 ;
        RECT 589.950 520.950 592.050 523.050 ;
        RECT 593.250 521.850 594.750 522.750 ;
        RECT 595.950 522.450 598.050 523.050 ;
        RECT 599.400 522.450 600.450 547.950 ;
        RECT 605.400 535.050 606.450 556.950 ;
        RECT 607.950 553.950 610.050 556.050 ;
        RECT 611.250 554.850 612.750 555.750 ;
        RECT 613.950 553.950 616.050 556.050 ;
        RECT 608.400 553.050 609.450 553.950 ;
        RECT 607.950 550.950 610.050 553.050 ;
        RECT 613.950 541.950 616.050 544.050 ;
        RECT 604.950 532.950 607.050 535.050 ;
        RECT 614.400 532.050 615.450 541.950 ;
        RECT 617.400 541.050 618.450 556.950 ;
        RECT 616.950 538.950 619.050 541.050 ;
        RECT 616.950 532.950 619.050 535.050 ;
        RECT 619.950 532.950 622.050 535.050 ;
        RECT 613.950 529.950 616.050 532.050 ;
        RECT 617.400 529.050 618.450 532.950 ;
        RECT 610.950 526.950 613.050 529.050 ;
        RECT 614.250 527.850 615.750 528.750 ;
        RECT 616.950 526.950 619.050 529.050 ;
        RECT 620.400 526.050 621.450 532.950 ;
        RECT 610.950 524.850 613.050 525.750 ;
        RECT 613.950 523.950 616.050 526.050 ;
        RECT 616.950 524.850 619.050 525.750 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 595.950 521.400 600.450 522.450 ;
        RECT 595.950 520.950 598.050 521.400 ;
        RECT 583.950 517.950 586.050 520.050 ;
        RECT 589.950 518.850 592.050 519.750 ;
        RECT 586.950 499.950 589.050 502.050 ;
        RECT 577.950 487.950 580.050 490.050 ;
        RECT 577.950 485.250 580.050 486.150 ;
        RECT 583.950 485.250 586.050 486.150 ;
        RECT 577.950 483.450 580.050 484.050 ;
        RECT 575.400 482.400 580.050 483.450 ;
        RECT 577.950 481.950 580.050 482.400 ;
        RECT 581.250 482.250 582.750 483.150 ;
        RECT 583.950 481.950 586.050 484.050 ;
        RECT 584.400 481.050 585.450 481.950 ;
        RECT 577.950 478.950 580.050 481.050 ;
        RECT 580.950 478.950 583.050 481.050 ;
        RECT 583.950 478.950 586.050 481.050 ;
        RECT 569.400 464.400 573.450 465.450 ;
        RECT 568.950 460.950 571.050 463.050 ;
        RECT 565.950 457.950 568.050 460.050 ;
        RECT 566.400 454.050 567.450 457.950 ;
        RECT 569.400 454.050 570.450 460.950 ;
        RECT 572.400 454.050 573.450 464.400 ;
        RECT 565.950 451.950 568.050 454.050 ;
        RECT 568.950 451.950 571.050 454.050 ;
        RECT 571.950 451.950 574.050 454.050 ;
        RECT 575.250 452.250 577.050 453.150 ;
        RECT 569.400 451.050 570.450 451.950 ;
        RECT 565.950 449.850 567.750 450.750 ;
        RECT 568.950 448.950 571.050 451.050 ;
        RECT 572.250 449.850 573.750 450.750 ;
        RECT 574.950 448.950 577.050 451.050 ;
        RECT 575.400 448.050 576.450 448.950 ;
        RECT 568.950 446.850 571.050 447.750 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 574.950 442.950 577.050 445.050 ;
        RECT 559.950 416.250 562.050 417.150 ;
        RECT 565.950 415.950 568.050 418.050 ;
        RECT 566.400 415.050 567.450 415.950 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 563.250 413.250 564.750 414.150 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 569.250 413.250 571.050 414.150 ;
        RECT 575.400 412.050 576.450 442.950 ;
        RECT 578.400 430.050 579.450 478.950 ;
        RECT 581.400 475.050 582.450 478.950 ;
        RECT 580.950 472.950 583.050 475.050 ;
        RECT 577.950 427.950 580.050 430.050 ;
        RECT 556.950 409.950 559.050 412.050 ;
        RECT 562.950 409.950 565.050 412.050 ;
        RECT 566.250 410.850 567.750 411.750 ;
        RECT 568.950 409.950 571.050 412.050 ;
        RECT 574.950 409.950 577.050 412.050 ;
        RECT 563.400 397.050 564.450 409.950 ;
        RECT 562.950 394.950 565.050 397.050 ;
        RECT 569.400 394.050 570.450 409.950 ;
        RECT 562.950 391.950 565.050 394.050 ;
        RECT 568.950 391.950 571.050 394.050 ;
        RECT 556.950 388.950 559.050 391.050 ;
        RECT 557.400 385.050 558.450 388.950 ;
        RECT 556.950 382.950 559.050 385.050 ;
        RECT 560.250 383.250 562.050 384.150 ;
        RECT 556.950 380.850 558.750 381.750 ;
        RECT 559.950 381.450 562.050 382.050 ;
        RECT 563.400 381.450 564.450 391.950 ;
        RECT 574.950 388.950 577.050 391.050 ;
        RECT 575.400 385.050 576.450 388.950 ;
        RECT 578.400 388.050 579.450 427.950 ;
        RECT 587.400 418.050 588.450 499.950 ;
        RECT 614.400 487.050 615.450 523.950 ;
        RECT 623.400 523.050 624.450 658.950 ;
        RECT 626.400 589.050 627.450 673.950 ;
        RECT 637.950 671.850 640.050 672.750 ;
        RECT 640.950 671.250 643.050 672.150 ;
        RECT 649.950 670.950 652.050 673.050 ;
        RECT 640.950 667.950 643.050 670.050 ;
        RECT 643.950 667.950 646.050 670.050 ;
        RECT 637.950 664.950 640.050 667.050 ;
        RECT 638.400 634.050 639.450 664.950 ;
        RECT 641.400 664.050 642.450 667.950 ;
        RECT 640.950 661.950 643.050 664.050 ;
        RECT 628.950 631.950 631.050 634.050 ;
        RECT 637.950 631.950 640.050 634.050 ;
        RECT 625.950 586.950 628.050 589.050 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 622.950 520.950 625.050 523.050 ;
        RECT 626.400 502.050 627.450 553.950 ;
        RECT 625.950 499.950 628.050 502.050 ;
        RECT 625.950 495.300 628.050 497.400 ;
        RECT 626.550 491.700 627.750 495.300 ;
        RECT 622.950 487.950 625.050 490.050 ;
        RECT 625.950 489.600 628.050 491.700 ;
        RECT 595.950 485.250 598.050 486.150 ;
        RECT 601.950 485.250 604.050 486.150 ;
        RECT 604.950 484.950 607.050 487.050 ;
        RECT 613.950 484.950 616.050 487.050 ;
        RECT 595.950 481.950 598.050 484.050 ;
        RECT 599.250 482.250 600.750 483.150 ;
        RECT 601.950 481.950 604.050 484.050 ;
        RECT 596.400 469.050 597.450 481.950 ;
        RECT 598.950 478.950 601.050 481.050 ;
        RECT 599.400 478.050 600.450 478.950 ;
        RECT 598.950 475.950 601.050 478.050 ;
        RECT 595.950 466.950 598.050 469.050 ;
        RECT 596.400 466.050 597.450 466.950 ;
        RECT 595.950 463.950 598.050 466.050 ;
        RECT 592.950 457.950 595.050 460.050 ;
        RECT 593.400 454.050 594.450 457.950 ;
        RECT 605.400 457.050 606.450 484.950 ;
        RECT 623.400 484.050 624.450 487.950 ;
        RECT 610.950 482.250 613.050 483.150 ;
        RECT 613.950 482.850 616.050 483.750 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 610.950 478.950 613.050 481.050 ;
        RECT 622.950 479.850 625.050 480.750 ;
        RECT 626.550 477.600 627.750 489.600 ;
        RECT 625.950 475.500 628.050 477.600 ;
        RECT 613.950 463.950 616.050 466.050 ;
        RECT 614.400 457.050 615.450 463.950 ;
        RECT 619.950 460.950 622.050 463.050 ;
        RECT 620.400 457.050 621.450 460.950 ;
        RECT 601.950 454.950 604.050 457.050 ;
        RECT 604.950 454.950 607.050 457.050 ;
        RECT 613.950 454.950 616.050 457.050 ;
        RECT 617.250 455.250 618.750 456.150 ;
        RECT 619.950 454.950 622.050 457.050 ;
        RECT 589.950 452.250 591.750 453.150 ;
        RECT 592.950 451.950 595.050 454.050 ;
        RECT 596.250 452.250 598.050 453.150 ;
        RECT 598.950 451.950 601.050 454.050 ;
        RECT 589.950 448.950 592.050 451.050 ;
        RECT 593.250 449.850 594.750 450.750 ;
        RECT 595.950 450.450 598.050 451.050 ;
        RECT 599.400 450.450 600.450 451.950 ;
        RECT 595.950 449.400 600.450 450.450 ;
        RECT 595.950 448.950 598.050 449.400 ;
        RECT 590.400 445.050 591.450 448.950 ;
        RECT 589.950 442.950 592.050 445.050 ;
        RECT 595.950 439.950 598.050 442.050 ;
        RECT 589.950 421.950 592.050 424.050 ;
        RECT 580.950 415.950 583.050 418.050 ;
        RECT 583.950 416.250 586.050 417.150 ;
        RECT 586.950 415.950 589.050 418.050 ;
        RECT 577.950 385.950 580.050 388.050 ;
        RECT 574.950 382.950 577.050 385.050 ;
        RECT 578.250 383.250 580.050 384.150 ;
        RECT 581.400 382.050 582.450 415.950 ;
        RECT 590.400 415.050 591.450 421.950 ;
        RECT 583.950 412.950 586.050 415.050 ;
        RECT 587.250 413.250 588.750 414.150 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 593.250 413.250 595.050 414.150 ;
        RECT 584.400 409.050 585.450 412.950 ;
        RECT 586.950 409.950 589.050 412.050 ;
        RECT 590.250 410.850 591.750 411.750 ;
        RECT 592.950 409.950 595.050 412.050 ;
        RECT 583.950 406.950 586.050 409.050 ;
        RECT 593.400 394.050 594.450 409.950 ;
        RECT 589.950 391.950 592.050 394.050 ;
        RECT 592.950 391.950 595.050 394.050 ;
        RECT 583.950 385.950 586.050 388.050 ;
        RECT 584.400 385.050 585.450 385.950 ;
        RECT 583.950 382.950 586.050 385.050 ;
        RECT 587.250 383.250 589.050 384.150 ;
        RECT 559.950 380.400 564.450 381.450 ;
        RECT 574.950 380.850 576.750 381.750 ;
        RECT 559.950 379.950 562.050 380.400 ;
        RECT 577.950 379.950 580.050 382.050 ;
        RECT 580.950 379.950 583.050 382.050 ;
        RECT 583.950 380.850 585.750 381.750 ;
        RECT 586.950 381.450 589.050 382.050 ;
        RECT 590.400 381.450 591.450 391.950 ;
        RECT 596.400 385.050 597.450 439.950 ;
        RECT 599.400 427.050 600.450 449.400 ;
        RECT 602.400 442.050 603.450 454.950 ;
        RECT 604.950 451.950 607.050 454.050 ;
        RECT 610.950 451.950 613.050 454.050 ;
        RECT 614.250 452.850 615.750 453.750 ;
        RECT 616.950 451.950 619.050 454.050 ;
        RECT 620.250 452.850 622.050 453.750 ;
        RECT 601.950 439.950 604.050 442.050 ;
        RECT 598.950 424.950 601.050 427.050 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 595.950 382.950 598.050 385.050 ;
        RECT 586.950 380.400 591.450 381.450 ;
        RECT 586.950 379.950 589.050 380.400 ;
        RECT 590.400 379.050 591.450 380.400 ;
        RECT 589.950 376.950 592.050 379.050 ;
        RECT 556.950 349.950 559.050 352.050 ;
        RECT 592.950 349.950 595.050 352.050 ;
        RECT 557.400 346.050 558.450 349.950 ;
        RECT 580.950 346.950 583.050 349.050 ;
        RECT 556.950 343.950 559.050 346.050 ;
        RECT 562.950 345.450 565.050 346.050 ;
        RECT 560.250 344.250 561.750 345.150 ;
        RECT 562.950 344.400 567.450 345.450 ;
        RECT 562.950 343.950 565.050 344.400 ;
        RECT 517.950 341.250 519.750 342.150 ;
        RECT 520.950 340.950 523.050 343.050 ;
        RECT 526.950 341.250 528.750 342.150 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 538.950 341.250 541.050 342.150 ;
        RECT 544.950 341.250 547.050 342.150 ;
        RECT 553.950 340.950 556.050 343.050 ;
        RECT 556.950 341.850 558.750 342.750 ;
        RECT 559.950 340.950 562.050 343.050 ;
        RECT 563.250 341.850 565.050 342.750 ;
        RECT 514.950 337.950 517.050 340.050 ;
        RECT 517.950 337.950 520.050 340.050 ;
        RECT 521.250 338.850 523.050 339.750 ;
        RECT 526.950 337.950 529.050 340.050 ;
        RECT 530.250 338.850 532.050 339.750 ;
        RECT 544.950 337.950 547.050 340.050 ;
        RECT 518.400 328.050 519.450 337.950 ;
        RECT 517.950 325.950 520.050 328.050 ;
        RECT 514.950 322.950 517.050 325.050 ;
        RECT 511.950 313.950 514.050 316.050 ;
        RECT 515.400 313.050 516.450 322.950 ;
        RECT 527.400 321.450 528.450 337.950 ;
        RECT 524.400 320.400 528.450 321.450 ;
        RECT 508.950 310.950 511.050 313.050 ;
        RECT 514.950 312.450 517.050 313.050 ;
        RECT 512.400 311.400 517.050 312.450 ;
        RECT 508.950 308.850 511.050 309.750 ;
        RECT 505.950 304.950 508.050 307.050 ;
        RECT 505.950 277.950 508.050 280.050 ;
        RECT 497.400 275.400 501.450 276.450 ;
        RECT 487.950 271.950 490.050 274.050 ;
        RECT 484.950 268.950 487.050 271.050 ;
        RECT 469.950 266.850 472.050 267.750 ;
        RECT 481.950 266.250 484.050 267.150 ;
        RECT 484.950 266.850 487.050 267.750 ;
        RECT 481.950 262.950 484.050 265.050 ;
        RECT 482.400 244.050 483.450 262.950 ;
        RECT 475.950 241.950 478.050 244.050 ;
        RECT 481.950 241.950 484.050 244.050 ;
        RECT 457.950 238.950 460.050 241.050 ;
        RECT 463.950 238.950 466.050 241.050 ;
        RECT 469.950 238.950 472.050 241.050 ;
        RECT 464.400 238.050 465.450 238.950 ;
        RECT 454.950 236.250 456.750 237.150 ;
        RECT 457.950 235.950 460.050 238.050 ;
        RECT 461.250 236.250 463.050 237.150 ;
        RECT 463.950 235.950 466.050 238.050 ;
        RECT 454.950 234.450 457.050 235.050 ;
        RECT 452.400 233.400 457.050 234.450 ;
        RECT 458.250 233.850 459.750 234.750 ;
        RECT 454.950 232.950 457.050 233.400 ;
        RECT 460.950 232.950 463.050 235.050 ;
        RECT 464.400 232.050 465.450 235.950 ;
        RECT 457.950 229.950 460.050 232.050 ;
        RECT 463.950 229.950 466.050 232.050 ;
        RECT 448.950 226.950 451.050 229.050 ;
        RECT 445.950 205.950 448.050 208.050 ;
        RECT 424.950 199.950 427.050 202.050 ;
        RECT 430.950 200.250 433.050 201.150 ;
        RECT 446.250 200.250 447.750 201.150 ;
        RECT 448.950 199.950 451.050 202.050 ;
        RECT 425.400 199.050 426.450 199.950 ;
        RECT 421.950 197.250 423.750 198.150 ;
        RECT 424.950 196.950 427.050 199.050 ;
        RECT 428.250 197.250 429.750 198.150 ;
        RECT 430.950 196.950 433.050 199.050 ;
        RECT 442.950 197.850 444.750 198.750 ;
        RECT 445.950 196.950 448.050 199.050 ;
        RECT 449.250 197.850 451.050 198.750 ;
        RECT 421.950 193.950 424.050 196.050 ;
        RECT 425.250 194.850 426.750 195.750 ;
        RECT 427.950 193.950 430.050 196.050 ;
        RECT 422.400 193.050 423.450 193.950 ;
        RECT 418.950 190.950 421.050 193.050 ;
        RECT 421.950 190.950 424.050 193.050 ;
        RECT 419.400 168.450 420.450 190.950 ;
        RECT 428.400 169.050 429.450 193.950 ;
        RECT 439.950 190.950 442.050 193.050 ;
        RECT 430.950 181.950 433.050 184.050 ;
        RECT 421.950 168.450 424.050 169.050 ;
        RECT 419.400 167.400 424.050 168.450 ;
        RECT 421.950 166.950 424.050 167.400 ;
        RECT 427.950 166.950 430.050 169.050 ;
        RECT 415.950 163.950 418.050 166.050 ;
        RECT 421.950 164.850 424.050 165.750 ;
        RECT 427.950 164.850 430.050 165.750 ;
        RECT 412.950 159.300 415.050 161.400 ;
        RECT 424.950 160.950 427.050 163.050 ;
        RECT 382.950 154.950 385.050 157.050 ;
        RECT 413.550 155.700 414.750 159.300 ;
        RECT 364.950 124.950 367.050 127.050 ;
        RECT 370.950 124.950 373.050 127.050 ;
        RECT 374.250 125.850 376.050 126.750 ;
        RECT 376.950 124.950 379.050 127.050 ;
        RECT 365.400 121.050 366.450 124.950 ;
        RECT 364.950 118.950 367.050 121.050 ;
        RECT 371.400 118.050 372.450 124.950 ;
        RECT 373.950 118.950 376.050 121.050 ;
        RECT 355.950 115.950 358.050 118.050 ;
        RECT 361.950 115.950 364.050 118.050 ;
        RECT 370.950 115.950 373.050 118.050 ;
        RECT 356.400 112.050 357.450 115.950 ;
        RECT 352.950 109.950 355.050 112.050 ;
        RECT 355.950 109.950 358.050 112.050 ;
        RECT 353.400 109.050 354.450 109.950 ;
        RECT 352.950 106.950 355.050 109.050 ;
        RECT 349.950 103.950 352.050 106.050 ;
        RECT 350.400 97.050 351.450 103.950 ;
        RECT 352.950 100.950 355.050 103.050 ;
        RECT 343.950 96.450 346.050 97.050 ;
        RECT 325.950 88.950 328.050 89.400 ;
        RECT 331.950 89.400 336.450 90.450 ;
        RECT 341.400 95.400 346.050 96.450 ;
        RECT 331.950 88.950 334.050 89.400 ;
        RECT 341.400 76.050 342.450 95.400 ;
        RECT 343.950 94.950 346.050 95.400 ;
        RECT 347.250 95.250 348.750 96.150 ;
        RECT 349.950 94.950 352.050 97.050 ;
        RECT 353.400 94.050 354.450 100.950 ;
        RECT 362.400 100.050 363.450 115.950 ;
        RECT 364.950 106.950 367.050 109.050 ;
        RECT 361.950 97.950 364.050 100.050 ;
        RECT 362.400 94.050 363.450 97.950 ;
        RECT 365.400 97.050 366.450 106.950 ;
        RECT 364.950 94.950 367.050 97.050 ;
        RECT 368.250 95.250 369.750 96.150 ;
        RECT 370.950 94.950 373.050 97.050 ;
        RECT 374.400 94.050 375.450 118.950 ;
        RECT 383.400 97.050 384.450 154.950 ;
        RECT 412.950 153.600 415.050 155.700 ;
        RECT 388.950 131.250 391.050 132.150 ;
        RECT 403.950 130.950 406.050 133.050 ;
        RECT 415.950 131.250 418.050 132.150 ;
        RECT 385.950 128.250 387.750 129.150 ;
        RECT 388.950 127.950 391.050 130.050 ;
        RECT 392.250 128.250 393.750 129.150 ;
        RECT 394.950 127.950 397.050 130.050 ;
        RECT 400.950 127.950 403.050 130.050 ;
        RECT 385.950 124.950 388.050 127.050 ;
        RECT 391.950 124.950 394.050 127.050 ;
        RECT 395.250 125.850 397.050 126.750 ;
        RECT 392.400 124.050 393.450 124.950 ;
        RECT 391.950 121.950 394.050 124.050 ;
        RECT 391.950 106.950 394.050 109.050 ;
        RECT 379.950 94.950 382.050 97.050 ;
        RECT 382.950 94.950 385.050 97.050 ;
        RECT 343.950 92.850 345.750 93.750 ;
        RECT 346.950 91.950 349.050 94.050 ;
        RECT 350.250 92.850 351.750 93.750 ;
        RECT 352.950 91.950 355.050 94.050 ;
        RECT 361.950 91.950 364.050 94.050 ;
        RECT 364.950 92.850 366.750 93.750 ;
        RECT 367.950 91.950 370.050 94.050 ;
        RECT 371.250 92.850 372.750 93.750 ;
        RECT 373.950 91.950 376.050 94.050 ;
        RECT 352.950 89.850 355.050 90.750 ;
        RECT 373.950 89.850 376.050 90.750 ;
        RECT 340.950 73.950 343.050 76.050 ;
        RECT 361.950 70.950 364.050 73.050 ;
        RECT 307.950 64.950 310.050 67.050 ;
        RECT 352.950 64.950 355.050 67.050 ;
        RECT 304.950 61.950 307.050 64.050 ;
        RECT 325.950 61.950 328.050 64.050 ;
        RECT 256.950 52.950 259.050 55.050 ;
        RECT 259.950 53.250 261.750 54.150 ;
        RECT 262.950 52.950 265.050 55.050 ;
        RECT 266.250 53.250 267.750 54.150 ;
        RECT 268.950 52.950 271.050 55.050 ;
        RECT 286.950 53.250 289.050 54.150 ;
        RECT 292.950 52.950 295.050 55.050 ;
        RECT 295.950 52.950 298.050 55.050 ;
        RECT 305.400 54.450 306.450 61.950 ;
        RECT 310.950 59.250 313.050 60.150 ;
        RECT 307.950 56.250 309.750 57.150 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 316.950 57.450 319.050 58.050 ;
        RECT 314.250 56.250 315.750 57.150 ;
        RECT 316.950 56.400 321.450 57.450 ;
        RECT 316.950 55.950 319.050 56.400 ;
        RECT 307.950 54.450 310.050 55.050 ;
        RECT 305.400 53.400 310.050 54.450 ;
        RECT 307.950 52.950 310.050 53.400 ;
        RECT 313.950 52.950 316.050 55.050 ;
        RECT 317.250 53.850 319.050 54.750 ;
        RECT 253.950 46.950 256.050 49.050 ;
        RECT 244.950 40.950 247.050 43.050 ;
        RECT 217.950 28.950 220.050 31.050 ;
        RECT 232.950 28.950 235.050 31.050 ;
        RECT 208.950 25.950 211.050 28.050 ;
        RECT 209.400 25.050 210.450 25.950 ;
        RECT 218.400 25.050 219.450 28.950 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 187.950 20.850 189.750 21.750 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 196.950 19.950 199.050 22.050 ;
        RECT 205.950 19.950 208.050 22.050 ;
        RECT 208.950 20.850 211.050 21.750 ;
        RECT 211.950 20.250 214.050 21.150 ;
        RECT 217.950 20.850 220.050 21.750 ;
        RECT 229.950 19.950 232.050 22.050 ;
        RECT 233.400 21.450 234.450 28.950 ;
        RECT 257.400 25.050 258.450 52.950 ;
        RECT 259.950 49.950 262.050 52.050 ;
        RECT 263.250 50.850 264.750 51.750 ;
        RECT 265.950 49.950 268.050 52.050 ;
        RECT 260.400 49.050 261.450 49.950 ;
        RECT 259.950 46.950 262.050 49.050 ;
        RECT 260.400 37.050 261.450 46.950 ;
        RECT 259.950 34.950 262.050 37.050 ;
        RECT 250.950 24.450 253.050 25.050 ;
        RECT 248.400 23.400 253.050 24.450 ;
        RECT 235.950 21.450 238.050 22.050 ;
        RECT 233.400 20.400 238.050 21.450 ;
        RECT 235.950 19.950 238.050 20.400 ;
        RECT 239.250 20.250 241.050 21.150 ;
        RECT 248.400 19.050 249.450 23.400 ;
        RECT 250.950 22.950 253.050 23.400 ;
        RECT 254.250 23.250 255.750 24.150 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 250.950 20.850 252.750 21.750 ;
        RECT 253.950 19.950 256.050 22.050 ;
        RECT 257.250 20.850 258.750 21.750 ;
        RECT 259.950 21.450 262.050 22.050 ;
        RECT 259.950 20.400 264.450 21.450 ;
        RECT 259.950 19.950 262.050 20.400 ;
        RECT 263.400 19.050 264.450 20.400 ;
        RECT 211.950 16.950 214.050 19.050 ;
        RECT 229.950 17.850 231.750 18.750 ;
        RECT 232.950 16.950 235.050 19.050 ;
        RECT 236.250 17.850 237.750 18.750 ;
        RECT 238.950 16.950 241.050 19.050 ;
        RECT 247.950 16.950 250.050 19.050 ;
        RECT 259.950 17.850 262.050 18.750 ;
        RECT 262.950 16.950 265.050 19.050 ;
        RECT 263.400 16.050 264.450 16.950 ;
        RECT 266.400 16.050 267.450 49.950 ;
        RECT 269.400 43.050 270.450 52.950 ;
        RECT 320.400 52.050 321.450 56.400 ;
        RECT 326.400 54.450 327.450 61.950 ;
        RECT 331.950 59.250 334.050 60.150 ;
        RECT 353.400 58.050 354.450 64.950 ;
        RECT 328.950 56.250 330.750 57.150 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 337.950 57.450 340.050 58.050 ;
        RECT 335.250 56.250 336.750 57.150 ;
        RECT 337.950 56.400 342.450 57.450 ;
        RECT 337.950 55.950 340.050 56.400 ;
        RECT 328.950 54.450 331.050 55.050 ;
        RECT 326.400 53.400 331.050 54.450 ;
        RECT 328.950 52.950 331.050 53.400 ;
        RECT 334.950 52.950 337.050 55.050 ;
        RECT 338.250 53.850 340.050 54.750 ;
        RECT 280.950 49.950 283.050 52.050 ;
        RECT 283.950 50.250 285.750 51.150 ;
        RECT 286.950 49.950 289.050 52.050 ;
        RECT 292.950 50.850 295.050 51.750 ;
        RECT 319.950 49.950 322.050 52.050 ;
        RECT 271.950 46.950 274.050 49.050 ;
        RECT 281.400 48.450 282.450 49.950 ;
        RECT 283.950 48.450 286.050 49.050 ;
        RECT 281.400 47.400 286.050 48.450 ;
        RECT 283.950 46.950 286.050 47.400 ;
        RECT 268.950 40.950 271.050 43.050 ;
        RECT 272.400 22.050 273.450 46.950 ;
        RECT 287.400 40.050 288.450 49.950 ;
        RECT 289.950 46.950 292.050 49.050 ;
        RECT 277.950 37.950 280.050 40.050 ;
        RECT 286.950 37.950 289.050 40.050 ;
        RECT 278.400 25.050 279.450 37.950 ;
        RECT 290.400 37.050 291.450 46.950 ;
        RECT 341.400 46.050 342.450 56.400 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 356.250 56.250 357.750 57.150 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 352.950 53.850 354.750 54.750 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 359.250 53.850 361.050 54.750 ;
        RECT 316.950 43.950 319.050 46.050 ;
        RECT 340.950 43.950 343.050 46.050 ;
        RECT 286.950 34.950 289.050 37.050 ;
        RECT 289.950 34.950 292.050 37.050 ;
        RECT 287.400 30.450 288.450 34.950 ;
        RECT 289.950 30.450 292.050 31.050 ;
        RECT 287.400 29.400 292.050 30.450 ;
        RECT 289.950 28.950 292.050 29.400 ;
        RECT 298.950 28.950 301.050 31.050 ;
        RECT 299.400 28.050 300.450 28.950 ;
        RECT 283.950 25.950 286.050 28.050 ;
        RECT 289.950 25.950 292.050 28.050 ;
        RECT 298.950 25.950 301.050 28.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 281.250 23.250 283.050 24.150 ;
        RECT 283.950 23.850 286.050 24.750 ;
        RECT 286.950 23.250 289.050 24.150 ;
        RECT 271.950 19.950 274.050 22.050 ;
        RECT 277.950 20.850 279.750 21.750 ;
        RECT 280.950 19.950 283.050 22.050 ;
        RECT 286.950 19.950 289.050 22.050 ;
        RECT 184.950 13.950 187.050 16.050 ;
        RECT 232.950 14.850 235.050 15.750 ;
        RECT 262.950 13.950 265.050 16.050 ;
        RECT 265.950 13.950 268.050 16.050 ;
        RECT 281.400 13.050 282.450 19.950 ;
        RECT 286.950 18.450 289.050 19.050 ;
        RECT 290.400 18.450 291.450 25.950 ;
        RECT 317.400 25.050 318.450 43.950 ;
        RECT 325.950 37.950 328.050 40.050 ;
        RECT 326.400 25.050 327.450 37.950 ;
        RECT 298.950 23.850 301.050 24.750 ;
        RECT 301.950 23.250 304.050 24.150 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 322.950 23.250 324.750 24.150 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 331.950 23.250 334.050 24.150 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 350.250 23.250 351.750 24.150 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 362.400 22.050 363.450 70.950 ;
        RECT 373.950 58.950 376.050 61.050 ;
        RECT 374.400 58.050 375.450 58.950 ;
        RECT 380.400 58.050 381.450 94.950 ;
        RECT 388.950 91.950 391.050 94.050 ;
        RECT 392.400 91.050 393.450 106.950 ;
        RECT 394.950 91.950 397.050 94.050 ;
        RECT 398.250 92.250 400.050 93.150 ;
        RECT 388.950 89.850 390.750 90.750 ;
        RECT 391.950 88.950 394.050 91.050 ;
        RECT 395.250 89.850 396.750 90.750 ;
        RECT 397.950 88.950 400.050 91.050 ;
        RECT 391.950 86.850 394.050 87.750 ;
        RECT 397.950 61.950 400.050 64.050 ;
        RECT 398.400 58.050 399.450 61.950 ;
        RECT 401.400 61.050 402.450 127.950 ;
        RECT 404.400 124.050 405.450 130.950 ;
        RECT 409.950 129.450 412.050 130.050 ;
        RECT 407.400 128.400 412.050 129.450 ;
        RECT 403.950 121.950 406.050 124.050 ;
        RECT 407.400 118.050 408.450 128.400 ;
        RECT 409.950 127.950 412.050 128.400 ;
        RECT 413.250 128.250 414.750 129.150 ;
        RECT 415.950 127.950 418.050 130.050 ;
        RECT 419.250 128.250 421.050 129.150 ;
        RECT 409.950 125.850 411.750 126.750 ;
        RECT 412.950 124.950 415.050 127.050 ;
        RECT 416.400 124.050 417.450 127.950 ;
        RECT 418.950 124.950 421.050 127.050 ;
        RECT 415.950 121.950 418.050 124.050 ;
        RECT 406.950 115.950 409.050 118.050 ;
        RECT 407.400 94.050 408.450 115.950 ;
        RECT 415.950 103.950 418.050 106.050 ;
        RECT 409.950 94.950 412.050 97.050 ;
        RECT 410.400 94.050 411.450 94.950 ;
        RECT 416.400 94.050 417.450 103.950 ;
        RECT 425.400 100.050 426.450 160.950 ;
        RECT 431.400 130.050 432.450 181.950 ;
        RECT 433.950 173.400 436.050 175.500 ;
        RECT 434.400 156.600 435.600 173.400 ;
        RECT 440.400 160.050 441.450 190.950 ;
        RECT 454.950 184.950 457.050 187.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 448.950 169.950 451.050 172.050 ;
        RECT 449.400 166.050 450.450 169.950 ;
        RECT 448.950 163.950 451.050 166.050 ;
        RECT 452.400 163.050 453.450 178.950 ;
        RECT 455.400 166.050 456.450 184.950 ;
        RECT 458.400 172.050 459.450 229.950 ;
        RECT 470.400 229.050 471.450 238.950 ;
        RECT 472.950 235.950 475.050 238.050 ;
        RECT 476.400 235.050 477.450 241.950 ;
        RECT 478.950 238.950 481.050 241.050 ;
        RECT 484.950 238.950 487.050 241.050 ;
        RECT 479.400 238.050 480.450 238.950 ;
        RECT 478.950 235.950 481.050 238.050 ;
        RECT 482.250 236.250 484.050 237.150 ;
        RECT 472.950 233.850 474.750 234.750 ;
        RECT 475.950 232.950 478.050 235.050 ;
        RECT 479.250 233.850 480.750 234.750 ;
        RECT 481.950 234.450 484.050 235.050 ;
        RECT 485.400 234.450 486.450 238.950 ;
        RECT 488.400 235.050 489.450 271.950 ;
        RECT 493.950 236.850 496.050 237.750 ;
        RECT 481.950 233.400 486.450 234.450 ;
        RECT 481.950 232.950 484.050 233.400 ;
        RECT 487.950 232.950 490.050 235.050 ;
        RECT 475.950 230.850 478.050 231.750 ;
        RECT 469.950 226.950 472.050 229.050 ;
        RECT 493.950 208.950 496.050 211.050 ;
        RECT 494.400 202.050 495.450 208.950 ;
        RECT 463.950 199.950 466.050 202.050 ;
        RECT 469.950 200.250 472.050 201.150 ;
        RECT 472.950 199.950 475.050 202.050 ;
        RECT 475.950 199.950 478.050 202.050 ;
        RECT 487.950 199.950 490.050 202.050 ;
        RECT 491.250 200.250 492.750 201.150 ;
        RECT 493.950 199.950 496.050 202.050 ;
        RECT 464.400 199.050 465.450 199.950 ;
        RECT 460.950 197.250 462.750 198.150 ;
        RECT 463.950 196.950 466.050 199.050 ;
        RECT 467.250 197.250 468.750 198.150 ;
        RECT 469.950 196.950 472.050 199.050 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 464.250 194.850 465.750 195.750 ;
        RECT 466.950 193.950 469.050 196.050 ;
        RECT 461.400 175.050 462.450 193.950 ;
        RECT 473.400 181.050 474.450 199.950 ;
        RECT 472.950 178.950 475.050 181.050 ;
        RECT 460.950 172.950 463.050 175.050 ;
        RECT 476.400 172.050 477.450 199.950 ;
        RECT 487.950 197.850 489.750 198.750 ;
        RECT 490.950 196.950 493.050 199.050 ;
        RECT 494.250 197.850 496.050 198.750 ;
        RECT 493.950 190.950 496.050 193.050 ;
        RECT 487.950 184.950 490.050 187.050 ;
        RECT 484.950 173.400 487.050 175.500 ;
        RECT 457.950 169.950 460.050 172.050 ;
        RECT 466.950 169.950 469.050 172.050 ;
        RECT 475.950 171.450 478.050 172.050 ;
        RECT 475.950 170.400 480.450 171.450 ;
        RECT 475.950 169.950 478.050 170.400 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 458.250 164.250 460.050 165.150 ;
        RECT 448.950 161.850 450.750 162.750 ;
        RECT 451.950 160.950 454.050 163.050 ;
        RECT 455.250 161.850 456.750 162.750 ;
        RECT 457.950 160.950 460.050 163.050 ;
        RECT 439.950 157.950 442.050 160.050 ;
        RECT 451.950 158.850 454.050 159.750 ;
        RECT 433.950 154.500 436.050 156.600 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 436.950 128.250 439.050 129.150 ;
        RECT 431.400 127.050 432.450 127.950 ;
        RECT 427.950 125.250 429.750 126.150 ;
        RECT 430.950 124.950 433.050 127.050 ;
        RECT 434.250 125.250 435.750 126.150 ;
        RECT 436.950 124.950 439.050 127.050 ;
        RECT 427.950 121.950 430.050 124.050 ;
        RECT 431.250 122.850 432.750 123.750 ;
        RECT 433.950 121.950 436.050 124.050 ;
        RECT 428.400 112.050 429.450 121.950 ;
        RECT 434.400 118.050 435.450 121.950 ;
        RECT 433.950 115.950 436.050 118.050 ;
        RECT 427.950 109.950 430.050 112.050 ;
        RECT 421.950 97.950 424.050 100.050 ;
        RECT 424.950 97.950 427.050 100.050 ;
        RECT 430.950 97.950 433.050 100.050 ;
        RECT 406.950 91.950 409.050 94.050 ;
        RECT 409.950 91.950 412.050 94.050 ;
        RECT 415.950 91.950 418.050 94.050 ;
        RECT 419.250 92.250 421.050 93.150 ;
        RECT 409.950 89.850 411.750 90.750 ;
        RECT 412.950 88.950 415.050 91.050 ;
        RECT 416.250 89.850 417.750 90.750 ;
        RECT 418.950 88.950 421.050 91.050 ;
        RECT 412.950 86.850 415.050 87.750 ;
        RECT 419.400 67.050 420.450 88.950 ;
        RECT 418.950 64.950 421.050 67.050 ;
        RECT 400.950 58.950 403.050 61.050 ;
        RECT 403.950 59.250 406.050 60.150 ;
        RECT 422.400 58.050 423.450 97.950 ;
        RECT 430.950 95.850 433.050 96.750 ;
        RECT 433.950 95.250 436.050 96.150 ;
        RECT 440.400 94.050 441.450 157.950 ;
        RECT 458.400 130.050 459.450 160.950 ;
        RECT 457.950 127.950 460.050 130.050 ;
        RECT 454.950 124.950 457.050 127.050 ;
        RECT 467.400 126.450 468.450 169.950 ;
        RECT 472.950 167.250 475.050 168.150 ;
        RECT 475.950 167.850 478.050 168.750 ;
        RECT 479.400 168.450 480.450 170.400 ;
        RECT 481.950 170.250 484.050 171.150 ;
        RECT 481.950 168.450 484.050 169.050 ;
        RECT 479.400 167.400 484.050 168.450 ;
        RECT 481.950 166.950 484.050 167.400 ;
        RECT 472.950 163.950 475.050 166.050 ;
        RECT 469.950 128.250 472.050 129.150 ;
        RECT 469.950 126.450 472.050 127.050 ;
        RECT 467.400 125.400 472.050 126.450 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 473.250 125.250 474.750 126.150 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 479.250 125.250 481.050 126.150 ;
        RECT 448.950 121.950 451.050 124.050 ;
        RECT 454.950 122.850 457.050 123.750 ;
        RECT 457.950 122.250 460.050 123.150 ;
        RECT 460.950 121.950 463.050 124.050 ;
        RECT 449.400 97.050 450.450 121.950 ;
        RECT 457.950 120.450 460.050 121.050 ;
        RECT 461.400 120.450 462.450 121.950 ;
        RECT 470.400 121.050 471.450 124.950 ;
        RECT 472.950 121.950 475.050 124.050 ;
        RECT 476.250 122.850 477.750 123.750 ;
        RECT 478.950 121.950 481.050 124.050 ;
        RECT 457.950 119.400 462.450 120.450 ;
        RECT 457.950 118.950 460.050 119.400 ;
        RECT 469.950 118.950 472.050 121.050 ;
        RECT 451.950 106.950 454.050 109.050 ;
        RECT 452.400 100.050 453.450 106.950 ;
        RECT 473.400 103.050 474.450 121.950 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 451.950 97.950 454.050 100.050 ;
        RECT 455.400 97.050 456.450 100.950 ;
        RECT 448.950 94.950 451.050 97.050 ;
        RECT 452.250 95.850 453.750 96.750 ;
        RECT 454.950 94.950 457.050 97.050 ;
        RECT 433.950 91.950 436.050 94.050 ;
        RECT 439.950 91.950 442.050 94.050 ;
        RECT 448.950 92.850 451.050 93.750 ;
        RECT 454.950 92.850 457.050 93.750 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 377.250 56.250 378.750 57.150 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 401.250 56.250 402.750 57.150 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 407.250 56.250 409.050 57.150 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 373.950 53.850 375.750 54.750 ;
        RECT 376.950 52.950 379.050 55.050 ;
        RECT 380.250 53.850 382.050 54.750 ;
        RECT 397.950 53.850 399.750 54.750 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 377.400 49.050 378.450 52.950 ;
        RECT 404.400 52.050 405.450 55.950 ;
        RECT 406.950 54.450 409.050 55.050 ;
        RECT 410.400 54.450 411.450 55.950 ;
        RECT 406.950 53.400 411.450 54.450 ;
        RECT 406.950 52.950 409.050 53.400 ;
        RECT 403.950 49.950 406.050 52.050 ;
        RECT 413.400 49.050 414.450 55.950 ;
        RECT 422.400 55.050 423.450 55.950 ;
        RECT 434.400 55.050 435.450 91.950 ;
        RECT 464.400 91.050 465.450 100.950 ;
        RECT 472.950 97.950 475.050 100.050 ;
        RECT 466.950 94.950 469.050 97.050 ;
        RECT 463.950 88.950 466.050 91.050 ;
        RECT 467.400 90.450 468.450 94.950 ;
        RECT 473.400 94.050 474.450 97.950 ;
        RECT 482.400 94.050 483.450 166.950 ;
        RECT 485.550 161.400 486.750 173.400 ;
        RECT 484.950 159.300 487.050 161.400 ;
        RECT 485.550 155.700 486.750 159.300 ;
        RECT 484.950 153.600 487.050 155.700 ;
        RECT 488.400 127.050 489.450 184.950 ;
        RECT 494.400 169.050 495.450 190.950 ;
        RECT 493.950 166.950 496.050 169.050 ;
        RECT 493.950 164.850 496.050 165.750 ;
        RECT 497.400 163.050 498.450 275.400 ;
        RECT 499.950 272.250 502.050 273.150 ;
        RECT 506.400 271.050 507.450 277.950 ;
        RECT 499.950 268.950 502.050 271.050 ;
        RECT 503.250 269.250 504.750 270.150 ;
        RECT 505.950 268.950 508.050 271.050 ;
        RECT 509.250 269.250 511.050 270.150 ;
        RECT 512.400 268.050 513.450 311.400 ;
        RECT 514.950 310.950 517.050 311.400 ;
        RECT 517.950 310.950 520.050 313.050 ;
        RECT 514.950 308.850 517.050 309.750 ;
        RECT 518.400 307.050 519.450 310.950 ;
        RECT 524.400 310.050 525.450 320.400 ;
        RECT 541.950 316.950 544.050 319.050 ;
        RECT 542.400 313.050 543.450 316.950 ;
        RECT 566.400 316.050 567.450 344.400 ;
        RECT 581.400 343.050 582.450 346.950 ;
        RECT 586.950 344.250 589.050 345.150 ;
        RECT 593.400 343.050 594.450 349.950 ;
        RECT 574.950 340.950 577.050 343.050 ;
        RECT 577.950 341.250 579.750 342.150 ;
        RECT 580.950 340.950 583.050 343.050 ;
        RECT 584.250 341.250 585.750 342.150 ;
        RECT 586.950 340.950 589.050 343.050 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 565.950 313.950 568.050 316.050 ;
        RECT 526.950 310.950 529.050 313.050 ;
        RECT 529.950 311.250 531.750 312.150 ;
        RECT 532.950 310.950 535.050 313.050 ;
        RECT 538.950 311.250 540.750 312.150 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 559.950 312.450 562.050 313.050 ;
        RECT 556.950 311.250 558.750 312.150 ;
        RECT 559.950 311.400 564.450 312.450 ;
        RECT 559.950 310.950 562.050 311.400 ;
        RECT 523.950 307.950 526.050 310.050 ;
        RECT 517.950 304.950 520.050 307.050 ;
        RECT 527.400 289.050 528.450 310.950 ;
        RECT 529.950 307.950 532.050 310.050 ;
        RECT 533.250 308.850 535.050 309.750 ;
        RECT 538.950 307.950 541.050 310.050 ;
        RECT 542.250 308.850 544.050 309.750 ;
        RECT 556.950 307.950 559.050 310.050 ;
        RECT 560.250 308.850 562.050 309.750 ;
        RECT 530.400 307.050 531.450 307.950 ;
        RECT 557.400 307.050 558.450 307.950 ;
        RECT 529.950 304.950 532.050 307.050 ;
        RECT 556.950 304.950 559.050 307.050 ;
        RECT 563.400 304.050 564.450 311.400 ;
        RECT 565.950 311.250 567.750 312.150 ;
        RECT 568.950 310.950 571.050 313.050 ;
        RECT 565.950 307.950 568.050 310.050 ;
        RECT 569.250 308.850 571.050 309.750 ;
        RECT 571.950 307.950 574.050 310.050 ;
        RECT 538.950 301.950 541.050 304.050 ;
        RECT 562.950 301.950 565.050 304.050 ;
        RECT 526.950 286.950 529.050 289.050 ;
        RECT 535.950 286.950 538.050 289.050 ;
        RECT 526.950 274.950 529.050 277.050 ;
        RECT 527.400 274.050 528.450 274.950 ;
        RECT 520.950 272.250 523.050 273.150 ;
        RECT 526.950 271.950 529.050 274.050 ;
        RECT 527.400 271.050 528.450 271.950 ;
        RECT 520.950 268.950 523.050 271.050 ;
        RECT 524.250 269.250 525.750 270.150 ;
        RECT 526.950 268.950 529.050 271.050 ;
        RECT 530.250 269.250 532.050 270.150 ;
        RECT 502.950 265.950 505.050 268.050 ;
        RECT 506.250 266.850 507.750 267.750 ;
        RECT 508.950 267.450 511.050 268.050 ;
        RECT 511.950 267.450 514.050 268.050 ;
        RECT 508.950 266.400 514.050 267.450 ;
        RECT 508.950 265.950 511.050 266.400 ;
        RECT 511.950 265.950 514.050 266.400 ;
        RECT 503.400 250.050 504.450 265.950 ;
        RECT 502.950 247.950 505.050 250.050 ;
        RECT 521.400 247.050 522.450 268.950 ;
        RECT 523.950 265.950 526.050 268.050 ;
        RECT 527.250 266.850 528.750 267.750 ;
        RECT 529.950 265.950 532.050 268.050 ;
        RECT 524.400 265.050 525.450 265.950 ;
        RECT 523.950 262.950 526.050 265.050 ;
        RECT 536.400 264.450 537.450 286.950 ;
        RECT 539.400 268.050 540.450 301.950 ;
        RECT 562.950 298.950 565.050 301.050 ;
        RECT 563.400 274.050 564.450 298.950 ;
        RECT 562.950 273.450 565.050 274.050 ;
        RECT 541.950 272.250 544.050 273.150 ;
        RECT 560.400 272.400 565.050 273.450 ;
        RECT 541.950 268.950 544.050 271.050 ;
        RECT 545.250 269.250 546.750 270.150 ;
        RECT 547.950 268.950 550.050 271.050 ;
        RECT 551.250 269.250 553.050 270.150 ;
        RECT 538.950 265.950 541.050 268.050 ;
        RECT 536.400 263.400 540.450 264.450 ;
        RECT 520.950 244.950 523.050 247.050 ;
        RECT 499.950 241.950 502.050 244.050 ;
        RECT 532.950 241.950 535.050 244.050 ;
        RECT 500.400 241.050 501.450 241.950 ;
        RECT 499.950 238.950 502.050 241.050 ;
        RECT 499.950 236.850 502.050 237.750 ;
        RECT 508.950 235.950 511.050 238.050 ;
        RECT 514.950 236.250 516.750 237.150 ;
        RECT 517.950 235.950 520.050 238.050 ;
        RECT 521.250 236.250 523.050 237.150 ;
        RECT 505.950 202.950 508.050 205.050 ;
        RECT 506.400 199.050 507.450 202.950 ;
        RECT 509.400 202.050 510.450 235.950 ;
        RECT 514.950 232.950 517.050 235.050 ;
        RECT 518.250 233.850 519.750 234.750 ;
        RECT 515.400 205.050 516.450 232.950 ;
        RECT 533.400 211.050 534.450 241.950 ;
        RECT 539.400 241.050 540.450 263.400 ;
        RECT 542.400 262.050 543.450 268.950 ;
        RECT 560.400 268.050 561.450 272.400 ;
        RECT 562.950 271.950 565.050 272.400 ;
        RECT 566.250 272.250 567.750 273.150 ;
        RECT 568.950 271.950 571.050 274.050 ;
        RECT 562.950 269.850 564.750 270.750 ;
        RECT 565.950 268.950 568.050 271.050 ;
        RECT 569.250 269.850 571.050 270.750 ;
        RECT 566.400 268.050 567.450 268.950 ;
        RECT 572.400 268.050 573.450 307.950 ;
        RECT 544.950 265.950 547.050 268.050 ;
        RECT 548.250 266.850 549.750 267.750 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 559.950 265.950 562.050 268.050 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 571.950 265.950 574.050 268.050 ;
        RECT 541.950 259.950 544.050 262.050 ;
        RECT 547.950 259.950 550.050 262.050 ;
        RECT 544.950 241.950 547.050 244.050 ;
        RECT 545.400 241.050 546.450 241.950 ;
        RECT 538.950 238.950 541.050 241.050 ;
        RECT 542.250 239.250 543.750 240.150 ;
        RECT 544.950 238.950 547.050 241.050 ;
        RECT 535.950 235.950 538.050 238.050 ;
        RECT 539.250 236.850 540.750 237.750 ;
        RECT 541.950 235.950 544.050 238.050 ;
        RECT 545.250 236.850 547.050 237.750 ;
        RECT 535.950 233.850 538.050 234.750 ;
        RECT 538.950 232.950 541.050 235.050 ;
        RECT 532.950 208.950 535.050 211.050 ;
        RECT 514.950 202.950 517.050 205.050 ;
        RECT 533.400 202.050 534.450 208.950 ;
        RECT 508.950 199.950 511.050 202.050 ;
        RECT 511.950 200.250 514.050 201.150 ;
        RECT 526.950 199.950 529.050 202.050 ;
        RECT 530.250 200.250 531.750 201.150 ;
        RECT 532.950 199.950 535.050 202.050 ;
        RECT 535.950 199.950 538.050 202.050 ;
        RECT 502.950 197.250 504.750 198.150 ;
        RECT 505.950 196.950 508.050 199.050 ;
        RECT 509.250 197.250 510.750 198.150 ;
        RECT 511.950 196.950 514.050 199.050 ;
        RECT 526.950 197.850 528.750 198.750 ;
        RECT 529.950 196.950 532.050 199.050 ;
        RECT 533.250 197.850 535.050 198.750 ;
        RECT 502.950 193.950 505.050 196.050 ;
        RECT 506.250 194.850 507.750 195.750 ;
        RECT 508.950 193.950 511.050 196.050 ;
        RECT 536.400 195.450 537.450 199.950 ;
        RECT 539.400 199.050 540.450 232.950 ;
        RECT 542.400 217.050 543.450 235.950 ;
        RECT 548.400 229.050 549.450 259.950 ;
        RECT 551.400 244.050 552.450 265.950 ;
        RECT 559.950 247.950 562.050 250.050 ;
        RECT 550.950 241.950 553.050 244.050 ;
        RECT 560.400 238.050 561.450 247.950 ;
        RECT 565.950 244.950 568.050 247.050 ;
        RECT 562.950 241.950 565.050 244.050 ;
        RECT 563.400 241.050 564.450 241.950 ;
        RECT 562.950 238.950 565.050 241.050 ;
        RECT 556.950 236.250 558.750 237.150 ;
        RECT 559.950 235.950 562.050 238.050 ;
        RECT 563.400 235.050 564.450 238.950 ;
        RECT 566.400 238.050 567.450 244.950 ;
        RECT 565.950 235.950 568.050 238.050 ;
        RECT 556.950 232.950 559.050 235.050 ;
        RECT 560.250 233.850 561.750 234.750 ;
        RECT 562.950 232.950 565.050 235.050 ;
        RECT 566.250 233.850 568.050 234.750 ;
        RECT 557.400 232.050 558.450 232.950 ;
        RECT 556.950 229.950 559.050 232.050 ;
        RECT 562.950 230.850 565.050 231.750 ;
        RECT 547.950 226.950 550.050 229.050 ;
        RECT 541.950 214.950 544.050 217.050 ;
        RECT 541.950 207.300 544.050 209.400 ;
        RECT 542.550 203.700 543.750 207.300 ;
        RECT 562.950 206.400 565.050 208.500 ;
        RECT 541.950 201.600 544.050 203.700 ;
        RECT 538.950 196.950 541.050 199.050 ;
        RECT 538.950 195.450 541.050 196.050 ;
        RECT 536.400 194.400 541.050 195.450 ;
        RECT 503.400 181.050 504.450 193.950 ;
        RECT 517.950 184.950 520.050 187.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 499.950 172.950 502.050 175.050 ;
        RECT 500.400 169.050 501.450 172.950 ;
        RECT 499.950 166.950 502.050 169.050 ;
        RECT 499.950 164.850 502.050 165.750 ;
        RECT 493.950 160.950 496.050 163.050 ;
        RECT 496.950 160.950 499.050 163.050 ;
        RECT 494.400 127.050 495.450 160.950 ;
        RECT 503.400 127.050 504.450 178.950 ;
        RECT 505.950 173.400 508.050 175.500 ;
        RECT 506.400 156.600 507.600 173.400 ;
        RECT 518.400 166.050 519.450 184.950 ;
        RECT 536.400 181.050 537.450 194.400 ;
        RECT 538.950 193.950 541.050 194.400 ;
        RECT 538.950 191.850 541.050 192.750 ;
        RECT 542.550 189.600 543.750 201.600 ;
        RECT 544.950 196.950 547.050 199.050 ;
        RECT 550.950 197.250 553.050 198.150 ;
        RECT 556.950 197.250 559.050 198.150 ;
        RECT 541.950 187.500 544.050 189.600 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 535.950 178.950 538.050 181.050 ;
        RECT 517.950 163.950 520.050 166.050 ;
        RECT 521.400 165.450 522.450 178.950 ;
        RECT 527.400 172.050 528.450 178.950 ;
        RECT 526.950 169.950 529.050 172.050 ;
        RECT 535.950 169.950 538.050 172.050 ;
        RECT 541.950 169.950 544.050 172.050 ;
        RECT 536.400 169.050 537.450 169.950 ;
        RECT 542.400 169.050 543.450 169.950 ;
        RECT 523.950 167.250 526.050 168.150 ;
        RECT 526.950 167.850 529.050 168.750 ;
        RECT 532.950 166.950 535.050 169.050 ;
        RECT 535.950 166.950 538.050 169.050 ;
        RECT 539.250 167.250 540.750 168.150 ;
        RECT 541.950 166.950 544.050 169.050 ;
        RECT 523.950 165.450 526.050 166.050 ;
        RECT 521.400 164.400 526.050 165.450 ;
        RECT 523.950 163.950 526.050 164.400 ;
        RECT 523.950 160.950 526.050 163.050 ;
        RECT 505.950 154.500 508.050 156.600 ;
        RECT 511.950 131.250 514.050 132.150 ;
        RECT 508.950 128.250 510.750 129.150 ;
        RECT 511.950 127.950 514.050 130.050 ;
        RECT 517.950 129.450 520.050 130.050 ;
        RECT 515.250 128.250 516.750 129.150 ;
        RECT 517.950 128.400 522.450 129.450 ;
        RECT 517.950 127.950 520.050 128.400 ;
        RECT 487.950 124.950 490.050 127.050 ;
        RECT 493.950 124.950 496.050 127.050 ;
        RECT 497.250 125.250 499.050 126.150 ;
        RECT 502.950 124.950 505.050 127.050 ;
        RECT 508.950 124.950 511.050 127.050 ;
        RECT 487.950 122.850 490.050 123.750 ;
        RECT 490.950 122.250 493.050 123.150 ;
        RECT 493.950 122.850 495.750 123.750 ;
        RECT 496.950 121.950 499.050 124.050 ;
        RECT 512.400 121.050 513.450 127.950 ;
        RECT 514.950 124.950 517.050 127.050 ;
        RECT 518.250 125.850 520.050 126.750 ;
        RECT 490.950 118.950 493.050 121.050 ;
        RECT 511.950 118.950 514.050 121.050 ;
        RECT 515.400 118.050 516.450 124.950 ;
        RECT 514.950 115.950 517.050 118.050 ;
        RECT 502.950 112.950 505.050 115.050 ;
        RECT 503.400 109.050 504.450 112.950 ;
        RECT 502.950 106.950 505.050 109.050 ;
        RECT 496.950 103.950 499.050 106.050 ;
        RECT 497.400 97.050 498.450 103.950 ;
        RECT 503.400 97.050 504.450 106.950 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 496.950 94.950 499.050 97.050 ;
        RECT 500.250 95.250 501.750 96.150 ;
        RECT 502.950 94.950 505.050 97.050 ;
        RECT 514.950 95.250 517.050 96.150 ;
        RECT 517.950 95.850 520.050 96.750 ;
        RECT 469.950 92.250 471.750 93.150 ;
        RECT 472.950 91.950 475.050 94.050 ;
        RECT 476.250 92.250 478.050 93.150 ;
        RECT 481.950 91.950 484.050 94.050 ;
        RECT 493.950 91.950 496.050 94.050 ;
        RECT 497.250 92.850 498.750 93.750 ;
        RECT 499.950 91.950 502.050 94.050 ;
        RECT 503.250 92.850 505.050 93.750 ;
        RECT 514.950 91.950 517.050 94.050 ;
        RECT 469.950 90.450 472.050 91.050 ;
        RECT 467.400 89.400 472.050 90.450 ;
        RECT 473.250 89.850 474.750 90.750 ;
        RECT 469.950 88.950 472.050 89.400 ;
        RECT 475.950 88.950 478.050 91.050 ;
        RECT 493.950 89.850 496.050 90.750 ;
        RECT 521.400 88.050 522.450 128.400 ;
        RECT 524.400 93.450 525.450 160.950 ;
        RECT 529.950 97.950 532.050 100.050 ;
        RECT 530.400 97.050 531.450 97.950 ;
        RECT 526.950 95.250 528.750 96.150 ;
        RECT 529.950 94.950 532.050 97.050 ;
        RECT 526.950 93.450 529.050 94.050 ;
        RECT 524.400 92.400 529.050 93.450 ;
        RECT 530.250 92.850 532.050 93.750 ;
        RECT 520.950 85.950 523.050 88.050 ;
        RECT 493.950 82.950 496.050 85.050 ;
        RECT 478.950 64.950 481.050 67.050 ;
        RECT 479.400 64.050 480.450 64.950 ;
        RECT 475.950 61.950 478.050 64.050 ;
        RECT 478.950 61.950 481.050 64.050 ;
        RECT 463.950 59.250 466.050 60.150 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 460.950 56.250 462.750 57.150 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 467.250 56.250 468.750 57.150 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 437.400 55.050 438.450 55.950 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 421.950 52.950 424.050 55.050 ;
        RECT 425.250 53.250 427.050 54.150 ;
        RECT 433.950 52.950 436.050 55.050 ;
        RECT 436.950 52.950 439.050 55.050 ;
        RECT 442.950 52.950 445.050 55.050 ;
        RECT 446.250 53.250 448.050 54.150 ;
        RECT 460.950 52.950 463.050 55.050 ;
        RECT 415.950 50.850 418.050 51.750 ;
        RECT 418.950 50.250 421.050 51.150 ;
        RECT 421.950 50.850 423.750 51.750 ;
        RECT 424.950 49.950 427.050 52.050 ;
        RECT 436.950 50.850 439.050 51.750 ;
        RECT 439.950 50.250 442.050 51.150 ;
        RECT 442.950 50.850 444.750 51.750 ;
        RECT 445.950 49.950 448.050 52.050 ;
        RECT 376.950 46.950 379.050 49.050 ;
        RECT 412.950 46.950 415.050 49.050 ;
        RECT 418.950 46.950 421.050 49.050 ;
        RECT 425.400 40.050 426.450 49.950 ;
        RECT 439.950 46.950 442.050 49.050 ;
        RECT 440.400 46.050 441.450 46.950 ;
        RECT 446.400 46.050 447.450 49.950 ;
        RECT 464.400 49.050 465.450 55.950 ;
        RECT 476.400 55.050 477.450 61.950 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 470.250 53.850 472.050 54.750 ;
        RECT 475.950 52.950 478.050 55.050 ;
        RECT 479.400 51.450 480.450 61.950 ;
        RECT 487.950 58.950 490.050 61.050 ;
        RECT 488.400 58.050 489.450 58.950 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 481.950 53.250 484.050 54.150 ;
        RECT 487.950 53.850 490.050 54.750 ;
        RECT 490.950 53.250 493.050 54.150 ;
        RECT 481.950 51.450 484.050 52.050 ;
        RECT 479.400 50.400 484.050 51.450 ;
        RECT 481.950 49.950 484.050 50.400 ;
        RECT 490.950 49.950 493.050 52.050 ;
        RECT 463.950 46.950 466.050 49.050 ;
        RECT 439.950 43.950 442.050 46.050 ;
        RECT 445.950 43.950 448.050 46.050 ;
        RECT 439.950 40.950 442.050 43.050 ;
        RECT 457.950 40.950 460.050 43.050 ;
        RECT 424.950 37.950 427.050 40.050 ;
        RECT 412.950 31.950 415.050 34.050 ;
        RECT 415.950 31.950 418.050 34.050 ;
        RECT 379.950 28.950 382.050 31.050 ;
        RECT 394.950 28.950 397.050 31.050 ;
        RECT 376.950 25.950 379.050 28.050 ;
        RECT 301.950 19.950 304.050 22.050 ;
        RECT 316.950 20.850 319.050 21.750 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 326.250 20.850 328.050 21.750 ;
        RECT 331.950 19.950 334.050 22.050 ;
        RECT 346.950 20.850 348.750 21.750 ;
        RECT 349.950 19.950 352.050 22.050 ;
        RECT 353.250 20.850 354.750 21.750 ;
        RECT 355.950 19.950 358.050 22.050 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 370.950 20.250 372.750 21.150 ;
        RECT 373.950 19.950 376.050 22.050 ;
        RECT 286.950 17.400 291.450 18.450 ;
        RECT 286.950 16.950 289.050 17.400 ;
        RECT 350.400 16.050 351.450 19.950 ;
        RECT 377.400 19.050 378.450 25.950 ;
        RECT 380.400 22.050 381.450 28.950 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 379.950 19.950 382.050 22.050 ;
        RECT 355.950 17.850 358.050 18.750 ;
        RECT 370.950 16.950 373.050 19.050 ;
        RECT 374.250 17.850 375.750 18.750 ;
        RECT 376.950 16.950 379.050 19.050 ;
        RECT 380.250 17.850 382.050 18.750 ;
        RECT 349.950 13.950 352.050 16.050 ;
        RECT 376.950 14.850 379.050 15.750 ;
        RECT 389.400 13.050 390.450 22.950 ;
        RECT 391.950 20.850 394.050 21.750 ;
        RECT 395.400 18.450 396.450 28.950 ;
        RECT 413.400 25.050 414.450 31.950 ;
        RECT 416.400 28.050 417.450 31.950 ;
        RECT 430.950 28.950 433.050 31.050 ;
        RECT 436.950 28.950 439.050 31.050 ;
        RECT 415.950 25.950 418.050 28.050 ;
        RECT 431.400 25.050 432.450 28.950 ;
        RECT 437.400 25.050 438.450 28.950 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 416.250 23.850 417.750 24.750 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 434.250 23.250 435.750 24.150 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 440.400 22.050 441.450 40.950 ;
        RECT 458.400 31.050 459.450 40.950 ;
        RECT 472.950 31.950 475.050 34.050 ;
        RECT 454.950 28.950 457.050 31.050 ;
        RECT 457.950 28.950 460.050 31.050 ;
        RECT 451.950 27.450 454.050 28.050 ;
        RECT 449.400 26.400 454.050 27.450 ;
        RECT 449.400 25.050 450.450 26.400 ;
        RECT 451.950 25.950 454.050 26.400 ;
        RECT 455.400 25.050 456.450 28.950 ;
        RECT 473.400 25.050 474.450 31.950 ;
        RECT 475.950 25.950 478.050 28.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 451.950 23.850 453.750 24.750 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 460.950 23.250 463.050 24.150 ;
        RECT 472.950 22.950 475.050 25.050 ;
        RECT 397.950 20.250 400.050 21.150 ;
        RECT 400.950 20.850 403.050 21.750 ;
        RECT 412.950 20.850 415.050 21.750 ;
        RECT 418.950 20.850 421.050 21.750 ;
        RECT 430.950 20.850 432.750 21.750 ;
        RECT 433.950 19.950 436.050 22.050 ;
        RECT 437.250 20.850 438.750 21.750 ;
        RECT 439.950 19.950 442.050 22.050 ;
        RECT 454.950 20.850 457.050 21.750 ;
        RECT 460.950 19.950 463.050 22.050 ;
        RECT 472.950 20.850 475.050 21.750 ;
        RECT 434.400 19.050 435.450 19.950 ;
        RECT 397.950 18.450 400.050 19.050 ;
        RECT 395.400 17.400 400.050 18.450 ;
        RECT 397.950 16.950 400.050 17.400 ;
        RECT 433.950 16.950 436.050 19.050 ;
        RECT 439.950 17.850 442.050 18.750 ;
        RECT 476.400 18.450 477.450 25.950 ;
        RECT 481.950 24.450 484.050 25.050 ;
        RECT 481.950 23.400 486.450 24.450 ;
        RECT 481.950 22.950 484.050 23.400 ;
        RECT 478.950 20.250 481.050 21.150 ;
        RECT 481.950 20.850 484.050 21.750 ;
        RECT 478.950 18.450 481.050 19.050 ;
        RECT 476.400 17.400 481.050 18.450 ;
        RECT 478.950 16.950 481.050 17.400 ;
        RECT 485.400 16.050 486.450 23.400 ;
        RECT 494.400 22.050 495.450 82.950 ;
        RECT 524.400 69.450 525.450 92.400 ;
        RECT 526.950 91.950 529.050 92.400 ;
        RECT 533.400 85.050 534.450 166.950 ;
        RECT 545.400 166.050 546.450 196.950 ;
        RECT 550.950 193.950 553.050 196.050 ;
        RECT 556.950 193.950 559.050 196.050 ;
        RECT 551.400 193.050 552.450 193.950 ;
        RECT 550.950 190.950 553.050 193.050 ;
        RECT 563.400 189.600 564.600 206.400 ;
        RECT 575.400 199.050 576.450 340.950 ;
        RECT 596.400 340.050 597.450 382.950 ;
        RECT 602.400 382.050 603.450 412.950 ;
        RECT 605.400 397.050 606.450 451.950 ;
        RECT 610.950 449.850 613.050 450.750 ;
        RECT 617.400 424.050 618.450 451.950 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 620.400 424.050 621.450 445.950 ;
        RECT 629.400 427.050 630.450 631.950 ;
        RECT 638.400 631.050 639.450 631.950 ;
        RECT 631.950 628.950 634.050 631.050 ;
        RECT 637.950 628.950 640.050 631.050 ;
        RECT 641.250 629.250 643.050 630.150 ;
        RECT 631.950 626.850 634.050 627.750 ;
        RECT 634.950 626.250 637.050 627.150 ;
        RECT 637.950 626.850 639.750 627.750 ;
        RECT 640.950 625.950 643.050 628.050 ;
        RECT 634.950 622.950 637.050 625.050 ;
        RECT 637.950 622.950 640.050 625.050 ;
        RECT 635.400 622.050 636.450 622.950 ;
        RECT 634.950 619.950 637.050 622.050 ;
        RECT 638.400 604.050 639.450 622.950 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 632.400 601.050 633.450 601.950 ;
        RECT 631.950 598.950 634.050 601.050 ;
        RECT 635.250 599.250 637.050 600.150 ;
        RECT 637.950 599.850 640.050 600.750 ;
        RECT 640.950 599.250 643.050 600.150 ;
        RECT 631.950 596.850 633.750 597.750 ;
        RECT 634.950 595.950 637.050 598.050 ;
        RECT 640.950 595.950 643.050 598.050 ;
        RECT 635.400 586.050 636.450 595.950 ;
        RECT 640.950 592.950 643.050 595.050 ;
        RECT 634.950 583.950 637.050 586.050 ;
        RECT 634.950 563.250 637.050 564.150 ;
        RECT 641.400 562.050 642.450 592.950 ;
        RECT 631.950 560.250 633.750 561.150 ;
        RECT 634.950 559.950 637.050 562.050 ;
        RECT 638.250 560.250 639.750 561.150 ;
        RECT 640.950 559.950 643.050 562.050 ;
        RECT 631.950 556.950 634.050 559.050 ;
        RECT 632.400 556.050 633.450 556.950 ;
        RECT 631.950 553.950 634.050 556.050 ;
        RECT 635.400 550.050 636.450 559.950 ;
        RECT 637.950 556.950 640.050 559.050 ;
        RECT 641.250 557.850 643.050 558.750 ;
        RECT 644.400 555.450 645.450 667.950 ;
        RECT 650.400 625.050 651.450 670.950 ;
        RECT 653.400 670.050 654.450 697.950 ;
        RECT 656.400 673.050 657.450 697.950 ;
        RECT 662.400 673.050 663.450 733.950 ;
        RECT 664.950 703.950 667.050 706.050 ;
        RECT 668.250 704.250 669.750 705.150 ;
        RECT 670.950 703.950 673.050 706.050 ;
        RECT 664.950 701.850 666.750 702.750 ;
        RECT 667.950 700.950 670.050 703.050 ;
        RECT 671.250 701.850 673.050 702.750 ;
        RECT 668.400 676.050 669.450 700.950 ;
        RECT 670.950 691.950 673.050 694.050 ;
        RECT 667.950 673.950 670.050 676.050 ;
        RECT 655.950 670.950 658.050 673.050 ;
        RECT 659.250 671.250 660.750 672.150 ;
        RECT 661.950 670.950 664.050 673.050 ;
        RECT 667.950 672.450 670.050 673.050 ;
        RECT 671.400 672.450 672.450 691.950 ;
        RECT 665.250 671.250 666.750 672.150 ;
        RECT 667.950 671.400 672.450 672.450 ;
        RECT 667.950 670.950 670.050 671.400 ;
        RECT 652.950 667.950 655.050 670.050 ;
        RECT 655.950 668.850 657.750 669.750 ;
        RECT 658.950 667.950 661.050 670.050 ;
        RECT 662.250 668.850 663.750 669.750 ;
        RECT 664.950 667.950 667.050 670.050 ;
        RECT 668.250 668.850 670.050 669.750 ;
        RECT 665.400 657.450 666.450 667.950 ;
        RECT 665.400 656.400 669.450 657.450 ;
        RECT 662.250 632.250 663.750 633.150 ;
        RECT 664.950 631.950 667.050 634.050 ;
        RECT 658.950 629.850 660.750 630.750 ;
        RECT 661.950 628.950 664.050 631.050 ;
        RECT 665.250 629.850 667.050 630.750 ;
        RECT 649.950 622.950 652.050 625.050 ;
        RECT 661.950 619.950 664.050 622.050 ;
        RECT 646.950 604.950 649.050 607.050 ;
        RECT 647.400 598.050 648.450 604.950 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 646.950 597.450 649.050 598.050 ;
        RECT 649.950 597.450 652.050 598.050 ;
        RECT 646.950 596.400 652.050 597.450 ;
        RECT 646.950 595.950 649.050 596.400 ;
        RECT 649.950 595.950 652.050 596.400 ;
        RECT 641.400 554.400 645.450 555.450 ;
        RECT 634.950 547.950 637.050 550.050 ;
        RECT 631.950 526.950 634.050 529.050 ;
        RECT 635.250 527.250 636.750 528.150 ;
        RECT 637.950 526.950 640.050 529.050 ;
        RECT 641.400 526.050 642.450 554.400 ;
        RECT 647.400 544.050 648.450 595.950 ;
        RECT 653.400 595.050 654.450 601.950 ;
        RECT 655.950 595.950 658.050 598.050 ;
        RECT 659.250 596.250 661.050 597.150 ;
        RECT 649.950 593.850 651.750 594.750 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 656.250 593.850 657.750 594.750 ;
        RECT 658.950 594.450 661.050 595.050 ;
        RECT 662.400 594.450 663.450 619.950 ;
        RECT 664.950 610.950 667.050 613.050 ;
        RECT 665.400 604.050 666.450 610.950 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 658.950 593.400 663.450 594.450 ;
        RECT 658.950 592.950 661.050 593.400 ;
        RECT 652.950 590.850 655.050 591.750 ;
        RECT 665.400 586.050 666.450 601.950 ;
        RECT 664.950 583.950 667.050 586.050 ;
        RECT 652.950 559.950 655.050 562.050 ;
        RECT 653.400 559.050 654.450 559.950 ;
        RECT 652.950 556.950 655.050 559.050 ;
        RECT 658.950 556.950 661.050 559.050 ;
        RECT 662.250 557.250 664.050 558.150 ;
        RECT 652.950 554.850 655.050 555.750 ;
        RECT 655.950 554.250 658.050 555.150 ;
        RECT 658.950 554.850 660.750 555.750 ;
        RECT 661.950 555.450 664.050 556.050 ;
        RECT 665.400 555.450 666.450 583.950 ;
        RECT 661.950 554.400 666.450 555.450 ;
        RECT 668.400 555.450 669.450 656.400 ;
        RECT 671.400 634.050 672.450 671.400 ;
        RECT 670.950 631.950 673.050 634.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 674.400 603.450 675.450 757.950 ;
        RECT 685.950 748.950 688.050 751.050 ;
        RECT 686.400 745.050 687.450 748.950 ;
        RECT 676.950 744.450 679.050 745.050 ;
        RECT 676.950 743.400 681.450 744.450 ;
        RECT 676.950 742.950 679.050 743.400 ;
        RECT 676.950 740.850 679.050 741.750 ;
        RECT 680.400 730.050 681.450 743.400 ;
        RECT 685.950 742.950 688.050 745.050 ;
        RECT 682.950 740.250 685.050 741.150 ;
        RECT 685.950 740.850 688.050 741.750 ;
        RECT 682.950 736.950 685.050 739.050 ;
        RECT 679.950 727.950 682.050 730.050 ;
        RECT 683.400 724.050 684.450 736.950 ;
        RECT 689.400 733.050 690.450 796.950 ;
        RECT 694.950 773.250 697.050 774.150 ;
        RECT 694.950 769.950 697.050 772.050 ;
        RECT 694.950 742.950 697.050 745.050 ;
        RECT 688.950 730.950 691.050 733.050 ;
        RECT 695.400 724.050 696.450 742.950 ;
        RECT 682.950 721.950 685.050 724.050 ;
        RECT 694.950 721.950 697.050 724.050 ;
        RECT 679.950 703.950 682.050 706.050 ;
        RECT 685.950 703.950 688.050 706.050 ;
        RECT 680.400 670.050 681.450 703.950 ;
        RECT 686.400 703.050 687.450 703.950 ;
        RECT 682.950 701.250 684.750 702.150 ;
        RECT 685.950 700.950 688.050 703.050 ;
        RECT 689.250 701.250 690.750 702.150 ;
        RECT 691.950 700.950 694.050 703.050 ;
        RECT 695.250 701.250 697.050 702.150 ;
        RECT 698.400 700.050 699.450 811.950 ;
        RECT 701.400 811.050 702.450 815.400 ;
        RECT 703.950 814.950 706.050 815.400 ;
        RECT 707.250 815.250 708.750 816.150 ;
        RECT 709.950 814.950 712.050 817.050 ;
        RECT 703.950 812.850 705.750 813.750 ;
        RECT 706.950 811.950 709.050 814.050 ;
        RECT 710.250 812.850 711.750 813.750 ;
        RECT 712.950 811.950 715.050 814.050 ;
        RECT 700.950 808.950 703.050 811.050 ;
        RECT 707.400 808.050 708.450 811.950 ;
        RECT 712.950 809.850 715.050 810.750 ;
        RECT 716.400 808.050 717.450 820.950 ;
        RECT 706.950 805.950 709.050 808.050 ;
        RECT 715.950 805.950 718.050 808.050 ;
        RECT 725.400 805.050 726.450 850.950 ;
        RECT 731.400 837.600 732.600 854.400 ;
        RECT 736.950 845.250 739.050 846.150 ;
        RECT 742.950 845.250 745.050 846.150 ;
        RECT 736.950 841.950 739.050 844.050 ;
        RECT 742.950 841.950 745.050 844.050 ;
        RECT 730.950 835.500 733.050 837.600 ;
        RECT 743.400 829.050 744.450 841.950 ;
        RECT 742.950 826.950 745.050 829.050 ;
        RECT 742.950 821.400 745.050 823.500 ;
        RECT 727.950 812.250 729.750 813.150 ;
        RECT 730.950 811.950 733.050 814.050 ;
        RECT 734.250 812.250 736.050 813.150 ;
        RECT 727.950 808.950 730.050 811.050 ;
        RECT 731.250 809.850 732.750 810.750 ;
        RECT 733.950 808.950 736.050 811.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 700.950 773.250 703.050 774.150 ;
        RECT 700.950 769.950 703.050 772.050 ;
        RECT 713.400 771.450 714.450 802.950 ;
        RECT 715.950 773.250 718.050 774.150 ;
        RECT 721.950 773.250 724.050 774.150 ;
        RECT 715.950 771.450 718.050 772.050 ;
        RECT 713.400 770.400 718.050 771.450 ;
        RECT 715.950 769.950 718.050 770.400 ;
        RECT 721.950 769.950 724.050 772.050 ;
        RECT 701.400 760.050 702.450 769.950 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 722.400 745.050 723.450 769.950 ;
        RECT 728.400 748.050 729.450 808.950 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 743.400 804.600 744.600 821.400 ;
        RECT 730.950 782.400 733.050 784.500 ;
        RECT 731.400 765.600 732.600 782.400 ;
        RECT 730.950 763.500 733.050 765.600 ;
        RECT 727.950 745.950 730.050 748.050 ;
        RECT 728.400 745.050 729.450 745.950 ;
        RECT 700.950 742.950 703.050 745.050 ;
        RECT 704.250 743.250 705.750 744.150 ;
        RECT 706.950 742.950 709.050 745.050 ;
        RECT 721.950 744.450 724.050 745.050 ;
        RECT 721.950 743.400 726.450 744.450 ;
        RECT 721.950 742.950 724.050 743.400 ;
        RECT 700.950 740.850 702.750 741.750 ;
        RECT 703.950 739.950 706.050 742.050 ;
        RECT 707.250 740.850 708.750 741.750 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 721.950 740.850 724.050 741.750 ;
        RECT 704.400 730.050 705.450 739.950 ;
        RECT 709.950 737.850 712.050 738.750 ;
        RECT 725.400 730.050 726.450 743.400 ;
        RECT 727.950 742.950 730.050 745.050 ;
        RECT 727.950 740.850 730.050 741.750 ;
        RECT 734.400 739.050 735.450 802.950 ;
        RECT 742.950 802.500 745.050 804.600 ;
        RECT 746.400 781.050 747.450 892.950 ;
        RECT 769.950 890.250 772.050 891.150 ;
        RECT 763.950 888.450 766.050 889.050 ;
        RECT 763.950 887.400 768.450 888.450 ;
        RECT 763.950 886.950 766.050 887.400 ;
        RECT 757.950 884.850 760.050 885.750 ;
        RECT 763.950 884.850 766.050 885.750 ;
        RECT 751.950 855.300 754.050 857.400 ;
        RECT 752.250 851.700 753.450 855.300 ;
        RECT 751.950 849.600 754.050 851.700 ;
        RECT 752.250 837.600 753.450 849.600 ;
        RECT 754.950 847.950 757.050 850.050 ;
        RECT 755.400 844.050 756.450 847.950 ;
        RECT 754.950 841.950 757.050 844.050 ;
        RECT 757.950 841.950 760.050 844.050 ;
        RECT 754.950 839.850 757.050 840.750 ;
        RECT 751.950 835.500 754.050 837.600 ;
        RECT 758.400 835.050 759.450 841.950 ;
        RECT 757.950 832.950 760.050 835.050 ;
        RECT 754.950 826.950 757.050 829.050 ;
        RECT 755.400 817.050 756.450 826.950 ;
        RECT 748.950 814.950 751.050 817.050 ;
        RECT 754.950 814.950 757.050 817.050 ;
        RECT 748.950 812.850 751.050 813.750 ;
        RECT 754.950 812.850 757.050 813.750 ;
        RECT 751.950 783.300 754.050 785.400 ;
        RECT 745.950 778.950 748.050 781.050 ;
        RECT 752.250 779.700 753.450 783.300 ;
        RECT 751.950 777.600 754.050 779.700 ;
        RECT 736.950 773.250 739.050 774.150 ;
        RECT 742.950 773.250 745.050 774.150 ;
        RECT 736.950 769.950 739.050 772.050 ;
        RECT 742.950 769.950 745.050 772.050 ;
        RECT 737.400 769.050 738.450 769.950 ;
        RECT 736.950 766.950 739.050 769.050 ;
        RECT 743.400 763.050 744.450 769.950 ;
        RECT 752.250 765.600 753.450 777.600 ;
        RECT 754.950 769.950 757.050 772.050 ;
        RECT 754.950 767.850 757.050 768.750 ;
        RECT 758.400 766.050 759.450 832.950 ;
        RECT 763.950 821.400 766.050 823.500 ;
        RECT 767.400 822.450 768.450 887.400 ;
        RECT 769.950 886.950 772.050 889.050 ;
        RECT 770.400 883.050 771.450 886.950 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 773.550 881.400 774.750 893.400 ;
        RECT 781.950 888.450 784.050 889.050 ;
        RECT 781.950 887.400 786.450 888.450 ;
        RECT 781.950 886.950 784.050 887.400 ;
        RECT 781.950 884.850 784.050 885.750 ;
        RECT 772.950 879.300 775.050 881.400 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 773.550 875.700 774.750 879.300 ;
        RECT 772.950 873.600 775.050 875.700 ;
        RECT 779.400 850.050 780.450 880.950 ;
        RECT 772.950 847.950 775.050 850.050 ;
        RECT 778.950 849.450 781.050 850.050 ;
        RECT 776.250 848.250 777.750 849.150 ;
        RECT 778.950 848.400 783.450 849.450 ;
        RECT 778.950 847.950 781.050 848.400 ;
        RECT 772.950 845.850 774.750 846.750 ;
        RECT 775.950 844.950 778.050 847.050 ;
        RECT 779.250 845.850 781.050 846.750 ;
        RECT 782.400 844.050 783.450 848.400 ;
        RECT 781.950 841.950 784.050 844.050 ;
        RECT 785.400 829.050 786.450 887.400 ;
        RECT 787.950 886.950 790.050 889.050 ;
        RECT 787.950 884.850 790.050 885.750 ;
        RECT 794.400 876.600 795.600 893.400 ;
        RECT 862.950 892.950 865.050 895.050 ;
        RECT 835.950 889.950 838.050 892.050 ;
        RECT 856.950 889.950 859.050 892.050 ;
        RECT 817.950 888.450 820.050 889.050 ;
        RECT 817.950 887.400 822.450 888.450 ;
        RECT 817.950 886.950 820.050 887.400 ;
        RECT 805.950 883.950 808.050 886.050 ;
        RECT 811.950 884.850 814.050 885.750 ;
        RECT 817.950 884.850 820.050 885.750 ;
        RECT 793.950 874.500 796.050 876.600 ;
        RECT 787.950 847.950 790.050 850.050 ;
        RECT 790.950 848.250 793.050 849.150 ;
        RECT 796.950 847.950 799.050 850.050 ;
        RECT 784.950 826.950 787.050 829.050 ;
        RECT 767.400 821.400 771.450 822.450 ;
        RECT 764.250 809.400 765.450 821.400 ;
        RECT 766.950 818.250 769.050 819.150 ;
        RECT 766.950 814.950 769.050 817.050 ;
        RECT 767.400 811.050 768.450 814.950 ;
        RECT 763.950 807.300 766.050 809.400 ;
        RECT 766.950 808.950 769.050 811.050 ;
        RECT 764.250 803.700 765.450 807.300 ;
        RECT 763.950 801.600 766.050 803.700 ;
        RECT 770.400 778.050 771.450 821.400 ;
        RECT 772.950 817.950 775.050 820.050 ;
        RECT 778.950 817.950 781.050 820.050 ;
        RECT 784.950 817.950 787.050 820.050 ;
        RECT 773.400 811.050 774.450 817.950 ;
        RECT 778.950 815.850 781.050 816.750 ;
        RECT 781.950 815.250 784.050 816.150 ;
        RECT 781.950 811.950 784.050 814.050 ;
        RECT 772.950 808.950 775.050 811.050 ;
        RECT 775.950 808.950 778.050 811.050 ;
        RECT 769.950 775.950 772.050 778.050 ;
        RECT 772.950 772.950 775.050 775.050 ;
        RECT 769.950 770.250 772.050 771.150 ;
        RECT 772.950 770.850 775.050 771.750 ;
        RECT 769.950 766.950 772.050 769.050 ;
        RECT 751.950 763.500 754.050 765.600 ;
        RECT 757.950 763.950 760.050 766.050 ;
        RECT 742.950 760.950 745.050 763.050 ;
        RECT 739.950 748.950 742.050 751.050 ;
        RECT 740.400 739.050 741.450 748.950 ;
        RECT 748.950 745.950 751.050 748.050 ;
        RECT 749.400 745.050 750.450 745.950 ;
        RECT 742.950 742.950 745.050 745.050 ;
        RECT 746.250 743.250 747.750 744.150 ;
        RECT 748.950 742.950 751.050 745.050 ;
        RECT 752.250 743.250 753.750 744.150 ;
        RECT 754.950 742.950 757.050 745.050 ;
        RECT 742.950 740.850 744.750 741.750 ;
        RECT 745.950 739.950 748.050 742.050 ;
        RECT 749.250 740.850 750.750 741.750 ;
        RECT 751.950 739.950 754.050 742.050 ;
        RECT 755.250 740.850 757.050 741.750 ;
        RECT 746.400 739.050 747.450 739.950 ;
        RECT 730.950 736.950 733.050 739.050 ;
        RECT 733.950 736.950 736.050 739.050 ;
        RECT 739.950 736.950 742.050 739.050 ;
        RECT 745.950 736.950 748.050 739.050 ;
        RECT 703.950 727.950 706.050 730.050 ;
        RECT 724.950 727.950 727.050 730.050 ;
        RECT 703.950 711.300 706.050 713.400 ;
        RECT 704.550 707.700 705.750 711.300 ;
        RECT 724.950 710.400 727.050 712.500 ;
        RECT 703.950 705.600 706.050 707.700 ;
        RECT 700.950 700.950 703.050 703.050 ;
        RECT 701.400 700.050 702.450 700.950 ;
        RECT 682.950 697.950 685.050 700.050 ;
        RECT 686.250 698.850 687.750 699.750 ;
        RECT 688.950 697.950 691.050 700.050 ;
        RECT 692.250 698.850 693.750 699.750 ;
        RECT 694.950 697.950 697.050 700.050 ;
        RECT 697.950 697.950 700.050 700.050 ;
        RECT 700.950 697.950 703.050 700.050 ;
        RECT 683.400 697.050 684.450 697.950 ;
        RECT 682.950 694.950 685.050 697.050 ;
        RECT 695.400 694.050 696.450 697.950 ;
        RECT 700.950 695.850 703.050 696.750 ;
        RECT 694.950 691.950 697.050 694.050 ;
        RECT 704.550 693.600 705.750 705.600 ;
        RECT 712.950 701.250 715.050 702.150 ;
        RECT 718.950 701.250 721.050 702.150 ;
        RECT 706.950 697.950 709.050 700.050 ;
        RECT 712.950 697.950 715.050 700.050 ;
        RECT 718.950 697.950 721.050 700.050 ;
        RECT 703.950 691.500 706.050 693.600 ;
        RECT 700.950 677.400 703.050 679.500 ;
        RECT 682.950 673.950 685.050 676.050 ;
        RECT 685.950 673.950 688.050 676.050 ;
        RECT 697.950 674.250 700.050 675.150 ;
        RECT 683.400 670.050 684.450 673.950 ;
        RECT 686.400 673.050 687.450 673.950 ;
        RECT 685.950 670.950 688.050 673.050 ;
        RECT 689.250 671.250 690.750 672.150 ;
        RECT 691.950 670.950 694.050 673.050 ;
        RECT 697.950 670.950 700.050 673.050 ;
        RECT 698.400 670.050 699.450 670.950 ;
        RECT 679.950 667.950 682.050 670.050 ;
        RECT 682.950 667.950 685.050 670.050 ;
        RECT 686.250 668.850 687.750 669.750 ;
        RECT 688.950 667.950 691.050 670.050 ;
        RECT 692.250 668.850 694.050 669.750 ;
        RECT 697.950 667.950 700.050 670.050 ;
        RECT 682.950 665.850 685.050 666.750 ;
        RECT 689.400 658.050 690.450 667.950 ;
        RECT 701.550 665.400 702.750 677.400 ;
        RECT 707.400 667.050 708.450 697.950 ;
        RECT 713.400 691.050 714.450 697.950 ;
        RECT 712.950 688.950 715.050 691.050 ;
        RECT 709.950 672.450 712.050 673.050 ;
        RECT 713.400 672.450 714.450 688.950 ;
        RECT 719.400 685.050 720.450 697.950 ;
        RECT 725.400 693.600 726.600 710.400 ;
        RECT 724.950 691.500 727.050 693.600 ;
        RECT 718.950 682.950 721.050 685.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 721.950 677.400 724.050 679.500 ;
        RECT 715.950 673.950 718.050 676.050 ;
        RECT 716.400 673.050 717.450 673.950 ;
        RECT 709.950 671.400 714.450 672.450 ;
        RECT 709.950 670.950 712.050 671.400 ;
        RECT 715.950 670.950 718.050 673.050 ;
        RECT 709.950 668.850 712.050 669.750 ;
        RECT 715.950 668.850 718.050 669.750 ;
        RECT 700.950 663.300 703.050 665.400 ;
        RECT 706.950 664.950 709.050 667.050 ;
        RECT 701.550 659.700 702.750 663.300 ;
        RECT 709.950 661.950 712.050 664.050 ;
        RECT 688.950 655.950 691.050 658.050 ;
        RECT 700.950 657.600 703.050 659.700 ;
        RECT 676.950 632.250 679.050 633.150 ;
        RECT 688.950 631.950 691.050 634.050 ;
        RECT 700.950 631.950 703.050 634.050 ;
        RECT 676.950 628.950 679.050 631.050 ;
        RECT 680.250 629.250 681.750 630.150 ;
        RECT 682.950 628.950 685.050 631.050 ;
        RECT 686.250 629.250 688.050 630.150 ;
        RECT 679.950 625.950 682.050 628.050 ;
        RECT 683.250 626.850 684.750 627.750 ;
        RECT 685.950 627.450 688.050 628.050 ;
        RECT 689.400 627.450 690.450 631.950 ;
        RECT 694.950 629.250 697.050 630.150 ;
        RECT 700.950 629.850 703.050 630.750 ;
        RECT 703.950 629.250 706.050 630.150 ;
        RECT 710.400 628.050 711.450 661.950 ;
        RECT 715.950 658.950 718.050 661.050 ;
        RECT 722.400 660.600 723.600 677.400 ;
        RECT 712.950 631.950 715.050 634.050 ;
        RECT 685.950 626.400 690.450 627.450 ;
        RECT 685.950 625.950 688.050 626.400 ;
        RECT 674.400 602.400 678.450 603.450 ;
        RECT 670.950 599.850 673.050 600.750 ;
        RECT 673.950 599.250 676.050 600.150 ;
        RECT 673.950 595.950 676.050 598.050 ;
        RECT 673.950 567.300 676.050 569.400 ;
        RECT 674.550 563.700 675.750 567.300 ;
        RECT 673.950 561.600 676.050 563.700 ;
        RECT 670.950 555.450 673.050 556.050 ;
        RECT 668.400 554.400 673.050 555.450 ;
        RECT 661.950 553.950 664.050 554.400 ;
        RECT 655.950 550.950 658.050 553.050 ;
        RECT 656.400 550.050 657.450 550.950 ;
        RECT 655.950 547.950 658.050 550.050 ;
        RECT 646.950 541.950 649.050 544.050 ;
        RECT 658.950 541.950 661.050 544.050 ;
        RECT 659.400 529.050 660.450 541.950 ;
        RECT 664.950 538.950 667.050 541.050 ;
        RECT 652.950 526.950 655.050 529.050 ;
        RECT 656.250 527.250 657.750 528.150 ;
        RECT 658.950 526.950 661.050 529.050 ;
        RECT 631.950 524.850 633.750 525.750 ;
        RECT 634.950 523.950 637.050 526.050 ;
        RECT 638.250 524.850 639.750 525.750 ;
        RECT 640.950 525.450 643.050 526.050 ;
        RECT 640.950 524.400 645.450 525.450 ;
        RECT 652.950 524.850 654.750 525.750 ;
        RECT 640.950 523.950 643.050 524.400 ;
        RECT 637.950 520.950 640.050 523.050 ;
        RECT 640.950 521.850 643.050 522.750 ;
        RECT 631.950 484.950 634.050 487.050 ;
        RECT 634.950 485.250 637.050 486.150 ;
        RECT 625.950 424.950 628.050 427.050 ;
        RECT 628.950 424.950 631.050 427.050 ;
        RECT 616.950 421.950 619.050 424.050 ;
        RECT 619.950 421.950 622.050 424.050 ;
        RECT 613.950 418.950 616.050 421.050 ;
        RECT 607.950 416.250 610.050 417.150 ;
        RECT 614.400 415.050 615.450 418.950 ;
        RECT 626.400 418.050 627.450 424.950 ;
        RECT 632.400 421.050 633.450 484.950 ;
        RECT 634.950 481.950 637.050 484.050 ;
        RECT 635.400 481.050 636.450 481.950 ;
        RECT 634.950 478.950 637.050 481.050 ;
        RECT 638.400 454.050 639.450 520.950 ;
        RECT 644.400 517.050 645.450 524.400 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 659.250 524.850 660.750 525.750 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 643.950 514.950 646.050 517.050 ;
        RECT 646.950 494.400 649.050 496.500 ;
        RECT 640.950 485.250 643.050 486.150 ;
        RECT 640.950 481.950 643.050 484.050 ;
        RECT 647.400 477.600 648.600 494.400 ;
        RECT 646.950 475.500 649.050 477.600 ;
        RECT 656.400 475.050 657.450 523.950 ;
        RECT 661.950 521.850 664.050 522.750 ;
        RECT 661.950 514.950 664.050 517.050 ;
        RECT 658.950 484.950 661.050 487.050 ;
        RECT 659.400 478.050 660.450 484.950 ;
        RECT 658.950 475.950 661.050 478.050 ;
        RECT 655.950 472.950 658.050 475.050 ;
        RECT 662.400 460.050 663.450 514.950 ;
        RECT 665.400 481.050 666.450 538.950 ;
        RECT 668.400 523.050 669.450 554.400 ;
        RECT 670.950 553.950 673.050 554.400 ;
        RECT 670.950 551.850 673.050 552.750 ;
        RECT 674.550 549.600 675.750 561.600 ;
        RECT 673.950 547.500 676.050 549.600 ;
        RECT 670.950 544.950 673.050 547.050 ;
        RECT 667.950 520.950 670.050 523.050 ;
        RECT 671.400 499.050 672.450 544.950 ;
        RECT 677.400 535.050 678.450 602.400 ;
        RECT 680.400 601.050 681.450 625.950 ;
        RECT 689.400 613.050 690.450 626.400 ;
        RECT 694.950 625.950 697.050 628.050 ;
        RECT 703.950 625.950 706.050 628.050 ;
        RECT 709.950 625.950 712.050 628.050 ;
        RECT 688.950 610.950 691.050 613.050 ;
        RECT 685.950 605.400 688.050 607.500 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 679.950 586.950 682.050 589.050 ;
        RECT 686.400 588.600 687.600 605.400 ;
        RECT 689.400 589.050 690.450 610.950 ;
        RECT 695.400 610.050 696.450 625.950 ;
        RECT 704.400 622.050 705.450 625.950 ;
        RECT 703.950 619.950 706.050 622.050 ;
        RECT 694.950 607.950 697.050 610.050 ;
        RECT 691.950 598.950 694.050 601.050 ;
        RECT 691.950 596.850 694.050 597.750 ;
        RECT 695.400 592.050 696.450 607.950 ;
        RECT 697.950 604.950 700.050 607.050 ;
        RECT 706.950 605.400 709.050 607.500 ;
        RECT 698.400 601.050 699.450 604.950 ;
        RECT 697.950 598.950 700.050 601.050 ;
        RECT 697.950 596.850 700.050 597.750 ;
        RECT 707.250 593.400 708.450 605.400 ;
        RECT 709.950 602.250 712.050 603.150 ;
        RECT 709.950 598.950 712.050 601.050 ;
        RECT 713.400 598.050 714.450 631.950 ;
        RECT 712.950 595.950 715.050 598.050 ;
        RECT 694.950 589.950 697.050 592.050 ;
        RECT 706.950 591.300 709.050 593.400 ;
        RECT 680.400 552.450 681.450 586.950 ;
        RECT 685.950 586.500 688.050 588.600 ;
        RECT 688.950 586.950 691.050 589.050 ;
        RECT 707.250 587.700 708.450 591.300 ;
        RECT 706.950 585.600 709.050 587.700 ;
        RECT 709.950 586.950 712.050 589.050 ;
        RECT 706.950 577.950 709.050 580.050 ;
        RECT 685.950 574.950 688.050 577.050 ;
        RECT 682.950 557.250 685.050 558.150 ;
        RECT 682.950 553.950 685.050 556.050 ;
        RECT 680.400 551.400 684.450 552.450 ;
        RECT 676.950 532.950 679.050 535.050 ;
        RECT 673.950 524.250 675.750 525.150 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 680.250 524.250 682.050 525.150 ;
        RECT 673.950 520.950 676.050 523.050 ;
        RECT 677.250 521.850 678.750 522.750 ;
        RECT 679.950 520.950 682.050 523.050 ;
        RECT 679.950 517.950 682.050 520.050 ;
        RECT 670.950 496.950 673.050 499.050 ;
        RECT 667.950 485.250 669.750 486.150 ;
        RECT 670.950 484.950 673.050 487.050 ;
        RECT 676.950 484.950 679.050 487.050 ;
        RECT 667.950 481.950 670.050 484.050 ;
        RECT 671.250 482.850 673.050 483.750 ;
        RECT 673.950 482.250 676.050 483.150 ;
        RECT 676.950 482.850 679.050 483.750 ;
        RECT 664.950 478.950 667.050 481.050 ;
        RECT 673.950 478.950 676.050 481.050 ;
        RECT 664.950 475.950 667.050 478.050 ;
        RECT 661.950 457.950 664.050 460.050 ;
        RECT 646.950 454.950 649.050 457.050 ;
        RECT 655.950 454.950 658.050 457.050 ;
        RECT 659.250 455.250 660.750 456.150 ;
        RECT 661.950 454.950 664.050 457.050 ;
        RECT 634.950 452.250 636.750 453.150 ;
        RECT 637.950 451.950 640.050 454.050 ;
        RECT 641.250 452.250 643.050 453.150 ;
        RECT 634.950 448.950 637.050 451.050 ;
        RECT 638.250 449.850 639.750 450.750 ;
        RECT 640.950 448.950 643.050 451.050 ;
        RECT 635.400 444.450 636.450 448.950 ;
        RECT 647.400 448.050 648.450 454.950 ;
        RECT 652.950 451.950 655.050 454.050 ;
        RECT 656.250 452.850 657.750 453.750 ;
        RECT 658.950 451.950 661.050 454.050 ;
        RECT 662.250 452.850 664.050 453.750 ;
        RECT 652.950 449.850 655.050 450.750 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 635.400 443.400 639.450 444.450 ;
        RECT 634.950 421.950 637.050 424.050 ;
        RECT 631.950 418.950 634.050 421.050 ;
        RECT 625.950 415.950 628.050 418.050 ;
        RECT 629.250 416.250 630.750 417.150 ;
        RECT 631.950 415.950 634.050 418.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 611.250 413.250 612.750 414.150 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 617.250 413.250 619.050 414.150 ;
        RECT 625.950 413.850 627.750 414.750 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 632.250 413.850 634.050 414.750 ;
        RECT 610.950 409.950 613.050 412.050 ;
        RECT 614.250 410.850 615.750 411.750 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 611.400 403.050 612.450 409.950 ;
        RECT 613.950 403.950 616.050 406.050 ;
        RECT 610.950 400.950 613.050 403.050 ;
        RECT 604.950 394.950 607.050 397.050 ;
        RECT 610.950 394.950 613.050 397.050 ;
        RECT 598.950 380.250 600.750 381.150 ;
        RECT 601.950 379.950 604.050 382.050 ;
        RECT 605.250 380.250 607.050 381.150 ;
        RECT 598.950 376.950 601.050 379.050 ;
        RECT 602.250 377.850 603.750 378.750 ;
        RECT 604.950 376.950 607.050 379.050 ;
        RECT 601.950 341.250 604.050 342.150 ;
        RECT 607.950 341.250 610.050 342.150 ;
        RECT 577.950 337.950 580.050 340.050 ;
        RECT 581.250 338.850 582.750 339.750 ;
        RECT 583.950 337.950 586.050 340.050 ;
        RECT 595.950 337.950 598.050 340.050 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 605.250 338.250 606.750 339.150 ;
        RECT 607.950 337.950 610.050 340.050 ;
        RECT 584.400 328.050 585.450 337.950 ;
        RECT 583.950 325.950 586.050 328.050 ;
        RECT 602.400 316.050 603.450 337.950 ;
        RECT 608.400 337.050 609.450 337.950 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 601.950 313.950 604.050 316.050 ;
        RECT 586.950 310.950 589.050 313.050 ;
        RECT 592.950 312.450 595.050 313.050 ;
        RECT 595.950 312.450 598.050 313.050 ;
        RECT 605.400 312.450 606.450 334.950 ;
        RECT 611.400 325.050 612.450 394.950 ;
        RECT 610.950 322.950 613.050 325.050 ;
        RECT 614.400 316.050 615.450 403.950 ;
        RECT 617.400 394.050 618.450 409.950 ;
        RECT 619.950 397.950 622.050 400.050 ;
        RECT 616.950 391.950 619.050 394.050 ;
        RECT 620.400 388.050 621.450 397.950 ;
        RECT 622.950 391.950 625.050 394.050 ;
        RECT 619.950 385.950 622.050 388.050 ;
        RECT 623.400 385.050 624.450 391.950 ;
        RECT 625.950 388.950 628.050 391.050 ;
        RECT 626.400 385.050 627.450 388.950 ;
        RECT 616.950 382.950 619.050 385.050 ;
        RECT 620.250 383.850 621.750 384.750 ;
        RECT 622.950 382.950 625.050 385.050 ;
        RECT 625.950 382.950 628.050 385.050 ;
        RECT 616.950 380.850 619.050 381.750 ;
        RECT 622.950 380.850 625.050 381.750 ;
        RECT 626.400 379.050 627.450 382.950 ;
        RECT 625.950 376.950 628.050 379.050 ;
        RECT 635.400 349.050 636.450 421.950 ;
        RECT 638.400 415.050 639.450 443.400 ;
        RECT 647.400 415.050 648.450 445.950 ;
        RECT 659.400 442.050 660.450 451.950 ;
        RECT 658.950 439.950 661.050 442.050 ;
        RECT 665.400 418.050 666.450 475.950 ;
        RECT 674.400 469.050 675.450 478.950 ;
        RECT 673.950 466.950 676.050 469.050 ;
        RECT 673.950 460.950 676.050 463.050 ;
        RECT 670.950 457.950 673.050 460.050 ;
        RECT 664.950 415.950 667.050 418.050 ;
        RECT 667.950 416.250 670.050 417.150 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 658.950 413.250 660.750 414.150 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 665.250 413.250 666.750 414.150 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 643.950 410.250 646.050 411.150 ;
        RECT 646.950 410.850 649.050 411.750 ;
        RECT 643.950 406.950 646.050 409.050 ;
        RECT 644.400 400.050 645.450 406.950 ;
        RECT 643.950 397.950 646.050 400.050 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 637.950 383.250 640.050 384.150 ;
        RECT 640.950 383.850 643.050 384.750 ;
        RECT 637.950 379.950 640.050 382.050 ;
        RECT 638.400 379.050 639.450 379.950 ;
        RECT 637.950 376.950 640.050 379.050 ;
        RECT 634.950 346.950 637.050 349.050 ;
        RECT 653.400 346.050 654.450 412.950 ;
        RECT 658.950 409.950 661.050 412.050 ;
        RECT 662.250 410.850 663.750 411.750 ;
        RECT 664.950 409.950 667.050 412.050 ;
        RECT 659.400 403.050 660.450 409.950 ;
        RECT 658.950 400.950 661.050 403.050 ;
        RECT 668.400 397.050 669.450 412.950 ;
        RECT 667.950 394.950 670.050 397.050 ;
        RECT 664.950 388.950 667.050 391.050 ;
        RECT 655.950 380.250 657.750 381.150 ;
        RECT 658.950 379.950 661.050 382.050 ;
        RECT 662.250 380.250 664.050 381.150 ;
        RECT 659.250 377.850 660.750 378.750 ;
        RECT 661.950 378.450 664.050 379.050 ;
        RECT 665.400 378.450 666.450 388.950 ;
        RECT 661.950 377.400 666.450 378.450 ;
        RECT 661.950 376.950 664.050 377.400 ;
        RECT 625.950 343.950 628.050 346.050 ;
        RECT 631.950 345.450 634.050 346.050 ;
        RECT 629.250 344.250 630.750 345.150 ;
        RECT 631.950 344.400 636.450 345.450 ;
        RECT 631.950 343.950 634.050 344.400 ;
        RECT 625.950 341.850 627.750 342.750 ;
        RECT 628.950 340.950 631.050 343.050 ;
        RECT 632.250 341.850 634.050 342.750 ;
        RECT 629.400 325.050 630.450 340.950 ;
        RECT 635.400 340.050 636.450 344.400 ;
        RECT 640.950 343.950 643.050 346.050 ;
        RECT 652.950 343.950 655.050 346.050 ;
        RECT 667.950 344.250 670.050 345.150 ;
        RECT 634.950 337.950 637.050 340.050 ;
        RECT 641.400 339.450 642.450 343.950 ;
        RECT 643.950 341.250 646.050 342.150 ;
        RECT 649.950 341.250 652.050 342.150 ;
        RECT 658.950 341.250 660.750 342.150 ;
        RECT 661.950 340.950 664.050 343.050 ;
        RECT 667.950 342.450 670.050 343.050 ;
        RECT 671.400 342.450 672.450 457.950 ;
        RECT 674.400 457.050 675.450 460.950 ;
        RECT 680.400 457.050 681.450 517.950 ;
        RECT 683.400 478.050 684.450 551.400 ;
        RECT 686.400 523.050 687.450 574.950 ;
        RECT 694.950 566.400 697.050 568.500 ;
        RECT 688.950 557.250 691.050 558.150 ;
        RECT 688.950 553.950 691.050 556.050 ;
        RECT 689.400 544.050 690.450 553.950 ;
        RECT 695.400 549.600 696.600 566.400 ;
        RECT 707.400 556.050 708.450 577.950 ;
        RECT 703.950 553.950 706.050 556.050 ;
        RECT 706.950 553.950 709.050 556.050 ;
        RECT 710.400 555.450 711.450 586.950 ;
        RECT 712.950 557.250 715.050 558.150 ;
        RECT 712.950 555.450 715.050 556.050 ;
        RECT 710.400 554.400 715.050 555.450 ;
        RECT 712.950 553.950 715.050 554.400 ;
        RECT 694.950 547.500 697.050 549.600 ;
        RECT 688.950 541.950 691.050 544.050 ;
        RECT 704.400 541.050 705.450 553.950 ;
        RECT 716.400 550.050 717.450 658.950 ;
        RECT 721.950 658.500 724.050 660.600 ;
        RECT 721.950 629.250 724.050 630.150 ;
        RECT 718.950 626.250 720.750 627.150 ;
        RECT 721.950 625.950 724.050 628.050 ;
        RECT 718.950 622.950 721.050 625.050 ;
        RECT 719.400 622.050 720.450 622.950 ;
        RECT 718.950 619.950 721.050 622.050 ;
        RECT 725.400 606.450 726.450 679.950 ;
        RECT 727.950 655.950 730.050 658.050 ;
        RECT 728.400 631.050 729.450 655.950 ;
        RECT 727.950 628.950 730.050 631.050 ;
        RECT 727.950 626.850 730.050 627.750 ;
        RECT 722.400 605.400 726.450 606.450 ;
        RECT 722.400 558.450 723.450 605.400 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 724.950 599.850 727.050 600.750 ;
        RECT 727.950 599.250 730.050 600.150 ;
        RECT 727.950 595.950 730.050 598.050 ;
        RECT 731.400 571.050 732.450 736.950 ;
        RECT 733.950 730.950 736.050 733.050 ;
        RECT 734.400 661.050 735.450 730.950 ;
        RECT 742.950 705.450 745.050 706.050 ;
        RECT 740.400 704.400 745.050 705.450 ;
        RECT 740.400 688.050 741.450 704.400 ;
        RECT 742.950 703.950 745.050 704.400 ;
        RECT 746.250 704.250 747.750 705.150 ;
        RECT 748.950 703.950 751.050 706.050 ;
        RECT 742.950 701.850 744.750 702.750 ;
        RECT 745.950 700.950 748.050 703.050 ;
        RECT 749.250 701.850 751.050 702.750 ;
        RECT 754.950 688.950 757.050 691.050 ;
        RECT 739.950 685.950 742.050 688.050 ;
        RECT 742.950 682.950 745.050 685.050 ;
        RECT 743.400 673.050 744.450 682.950 ;
        RECT 751.950 673.950 754.050 676.050 ;
        RECT 736.950 670.950 739.050 673.050 ;
        RECT 740.250 671.250 741.750 672.150 ;
        RECT 742.950 670.950 745.050 673.050 ;
        RECT 748.950 670.950 751.050 673.050 ;
        RECT 736.950 668.850 738.750 669.750 ;
        RECT 739.950 667.950 742.050 670.050 ;
        RECT 743.250 668.850 744.750 669.750 ;
        RECT 745.950 667.950 748.050 670.050 ;
        RECT 740.400 664.050 741.450 667.950 ;
        RECT 745.950 665.850 748.050 666.750 ;
        RECT 739.950 661.950 742.050 664.050 ;
        RECT 733.950 658.950 736.050 661.050 ;
        RECT 736.950 658.950 739.050 661.050 ;
        RECT 737.400 583.050 738.450 658.950 ;
        RECT 739.950 638.400 742.050 640.500 ;
        RECT 740.400 621.600 741.600 638.400 ;
        RECT 745.950 629.250 748.050 630.150 ;
        RECT 742.950 625.950 745.050 628.050 ;
        RECT 745.950 625.950 748.050 628.050 ;
        RECT 739.950 619.500 742.050 621.600 ;
        RECT 743.400 616.050 744.450 625.950 ;
        RECT 742.950 613.950 745.050 616.050 ;
        RECT 743.400 604.050 744.450 613.950 ;
        RECT 745.950 607.950 748.050 610.050 ;
        RECT 742.950 601.950 745.050 604.050 ;
        RECT 746.400 601.050 747.450 607.950 ;
        RECT 739.950 598.950 742.050 601.050 ;
        RECT 743.250 599.850 744.750 600.750 ;
        RECT 745.950 598.950 748.050 601.050 ;
        RECT 739.950 596.850 742.050 597.750 ;
        RECT 745.950 596.850 748.050 597.750 ;
        RECT 736.950 580.950 739.050 583.050 ;
        RECT 745.950 580.950 748.050 583.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 727.950 562.950 730.050 565.050 ;
        RECT 728.400 558.450 729.450 562.950 ;
        RECT 730.950 560.250 733.050 561.150 ;
        RECT 736.950 559.950 739.050 562.050 ;
        RECT 737.400 559.050 738.450 559.950 ;
        RECT 730.950 558.450 733.050 559.050 ;
        RECT 718.950 557.250 721.050 558.150 ;
        RECT 722.400 557.400 726.450 558.450 ;
        RECT 728.400 557.400 733.050 558.450 ;
        RECT 718.950 553.950 721.050 556.050 ;
        RECT 715.950 547.950 718.050 550.050 ;
        RECT 719.400 547.050 720.450 553.950 ;
        RECT 718.950 544.950 721.050 547.050 ;
        RECT 703.950 538.950 706.050 541.050 ;
        RECT 691.950 533.400 694.050 535.500 ;
        RECT 685.950 520.950 688.050 523.050 ;
        RECT 682.950 475.950 685.050 478.050 ;
        RECT 682.950 457.950 685.050 460.050 ;
        RECT 673.950 454.950 676.050 457.050 ;
        RECT 677.250 455.250 678.750 456.150 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 683.400 454.050 684.450 457.950 ;
        RECT 673.950 452.850 675.750 453.750 ;
        RECT 676.950 451.950 679.050 454.050 ;
        RECT 680.250 452.850 681.750 453.750 ;
        RECT 682.950 451.950 685.050 454.050 ;
        RECT 682.950 449.850 685.050 450.750 ;
        RECT 686.400 442.050 687.450 520.950 ;
        RECT 692.400 516.600 693.600 533.400 ;
        RECT 704.400 529.050 705.450 538.950 ;
        RECT 712.950 533.400 715.050 535.500 ;
        RECT 697.950 528.450 700.050 529.050 ;
        RECT 697.950 527.400 702.450 528.450 ;
        RECT 697.950 526.950 700.050 527.400 ;
        RECT 697.950 524.850 700.050 525.750 ;
        RECT 701.400 522.450 702.450 527.400 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 703.950 524.850 706.050 525.750 ;
        RECT 698.400 521.400 702.450 522.450 ;
        RECT 713.250 521.400 714.450 533.400 ;
        RECT 718.950 532.950 721.050 535.050 ;
        RECT 715.950 530.250 718.050 531.150 ;
        RECT 715.950 526.950 718.050 529.050 ;
        RECT 691.950 514.500 694.050 516.600 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 688.950 482.850 691.050 483.750 ;
        RECT 691.950 482.250 694.050 483.150 ;
        RECT 698.400 481.050 699.450 521.400 ;
        RECT 712.950 519.300 715.050 521.400 ;
        RECT 713.250 515.700 714.450 519.300 ;
        RECT 712.950 513.600 715.050 515.700 ;
        RECT 712.950 505.950 715.050 508.050 ;
        RECT 709.950 488.250 712.050 489.150 ;
        RECT 700.950 485.250 702.750 486.150 ;
        RECT 703.950 484.950 706.050 487.050 ;
        RECT 707.250 485.250 708.750 486.150 ;
        RECT 709.950 484.950 712.050 487.050 ;
        RECT 710.400 484.050 711.450 484.950 ;
        RECT 700.950 481.950 703.050 484.050 ;
        RECT 704.250 482.850 705.750 483.750 ;
        RECT 706.950 481.950 709.050 484.050 ;
        RECT 709.950 481.950 712.050 484.050 ;
        RECT 707.400 481.050 708.450 481.950 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 706.950 478.950 709.050 481.050 ;
        RECT 700.950 463.950 703.050 466.050 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 692.400 453.450 693.450 454.950 ;
        RECT 701.400 454.050 702.450 463.950 ;
        RECT 694.950 453.450 697.050 454.050 ;
        RECT 692.400 452.400 697.050 453.450 ;
        RECT 685.950 439.950 688.050 442.050 ;
        RECT 682.950 421.950 685.050 424.050 ;
        RECT 683.400 418.050 684.450 421.950 ;
        RECT 673.950 415.950 676.050 418.050 ;
        RECT 682.950 415.950 685.050 418.050 ;
        RECT 686.250 416.250 687.750 417.150 ;
        RECT 688.950 415.950 691.050 418.050 ;
        RECT 674.400 412.050 675.450 415.950 ;
        RECT 682.950 413.850 684.750 414.750 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 689.250 413.850 691.050 414.750 ;
        RECT 673.950 409.950 676.050 412.050 ;
        RECT 682.950 406.950 685.050 409.050 ;
        RECT 683.400 391.050 684.450 406.950 ;
        RECT 692.400 403.050 693.450 452.400 ;
        RECT 694.950 451.950 697.050 452.400 ;
        RECT 700.950 451.950 703.050 454.050 ;
        RECT 704.250 452.250 706.050 453.150 ;
        RECT 694.950 449.850 696.750 450.750 ;
        RECT 697.950 448.950 700.050 451.050 ;
        RECT 701.250 449.850 702.750 450.750 ;
        RECT 703.950 448.950 706.050 451.050 ;
        RECT 697.950 446.850 700.050 447.750 ;
        RECT 694.950 424.950 697.050 427.050 ;
        RECT 691.950 400.950 694.050 403.050 ;
        RECT 682.950 388.950 685.050 391.050 ;
        RECT 691.950 389.400 694.050 391.500 ;
        RECT 676.950 385.950 679.050 388.050 ;
        RECT 677.400 385.050 678.450 385.950 ;
        RECT 683.400 385.050 684.450 388.950 ;
        RECT 688.950 386.250 691.050 387.150 ;
        RECT 676.950 382.950 679.050 385.050 ;
        RECT 680.250 383.250 681.750 384.150 ;
        RECT 682.950 382.950 685.050 385.050 ;
        RECT 688.950 382.950 691.050 385.050 ;
        RECT 673.950 379.950 676.050 382.050 ;
        RECT 677.250 380.850 678.750 381.750 ;
        RECT 679.950 379.950 682.050 382.050 ;
        RECT 683.250 380.850 685.050 381.750 ;
        RECT 680.400 379.050 681.450 379.950 ;
        RECT 673.950 377.850 676.050 378.750 ;
        RECT 679.950 376.950 682.050 379.050 ;
        RECT 692.550 377.400 693.750 389.400 ;
        RECT 676.950 373.950 679.050 376.050 ;
        RECT 691.950 375.300 694.050 377.400 ;
        RECT 665.250 341.250 666.750 342.150 ;
        RECT 667.950 341.400 672.450 342.450 ;
        RECT 667.950 340.950 670.050 341.400 ;
        RECT 643.950 339.450 646.050 340.050 ;
        RECT 641.400 338.400 646.050 339.450 ;
        RECT 649.950 339.450 652.050 340.050 ;
        RECT 643.950 337.950 646.050 338.400 ;
        RECT 647.250 338.250 648.750 339.150 ;
        RECT 649.950 338.400 654.450 339.450 ;
        RECT 649.950 337.950 652.050 338.400 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 647.400 331.050 648.450 334.950 ;
        RECT 646.950 328.950 649.050 331.050 ;
        RECT 628.950 322.950 631.050 325.050 ;
        RECT 643.950 319.950 646.050 322.050 ;
        RECT 625.950 316.950 628.050 319.050 ;
        RECT 613.950 313.950 616.050 316.050 ;
        RECT 590.250 311.250 591.750 312.150 ;
        RECT 592.950 311.400 598.050 312.450 ;
        RECT 592.950 310.950 595.050 311.400 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 602.400 311.400 606.450 312.450 ;
        RECT 583.950 307.950 586.050 310.050 ;
        RECT 587.250 308.850 588.750 309.750 ;
        RECT 589.950 307.950 592.050 310.050 ;
        RECT 593.250 308.850 595.050 309.750 ;
        RECT 583.950 305.850 586.050 306.750 ;
        RECT 586.950 301.950 589.050 304.050 ;
        RECT 580.950 279.300 583.050 281.400 ;
        RECT 581.550 275.700 582.750 279.300 ;
        RECT 577.950 271.950 580.050 274.050 ;
        RECT 580.950 273.600 583.050 275.700 ;
        RECT 578.400 268.050 579.450 271.950 ;
        RECT 577.950 265.950 580.050 268.050 ;
        RECT 577.950 263.850 580.050 264.750 ;
        RECT 581.550 261.600 582.750 273.600 ;
        RECT 587.400 265.050 588.450 301.950 ;
        RECT 590.400 283.050 591.450 307.950 ;
        RECT 596.400 301.050 597.450 310.950 ;
        RECT 595.950 298.950 598.050 301.050 ;
        RECT 602.400 286.050 603.450 311.400 ;
        RECT 604.950 308.250 606.750 309.150 ;
        RECT 607.950 307.950 610.050 310.050 ;
        RECT 611.250 308.250 613.050 309.150 ;
        RECT 604.950 304.950 607.050 307.050 ;
        RECT 608.250 305.850 609.750 306.750 ;
        RECT 610.950 304.950 613.050 307.050 ;
        RECT 601.950 283.950 604.050 286.050 ;
        RECT 589.950 280.950 592.050 283.050 ;
        RECT 601.950 278.400 604.050 280.500 ;
        RECT 592.950 271.950 595.050 274.050 ;
        RECT 589.950 269.250 592.050 270.150 ;
        RECT 589.950 265.950 592.050 268.050 ;
        RECT 586.950 262.950 589.050 265.050 ;
        RECT 580.950 259.500 583.050 261.600 ;
        RECT 586.950 247.950 589.050 250.050 ;
        RECT 580.950 241.950 583.050 244.050 ;
        RECT 587.400 241.050 588.450 247.950 ;
        RECT 590.400 241.050 591.450 265.950 ;
        RECT 593.400 265.050 594.450 271.950 ;
        RECT 595.950 269.250 598.050 270.150 ;
        RECT 598.950 268.950 601.050 271.050 ;
        RECT 595.950 265.950 598.050 268.050 ;
        RECT 592.950 262.950 595.050 265.050 ;
        RECT 599.400 244.050 600.450 268.950 ;
        RECT 602.400 261.600 603.600 278.400 ;
        RECT 601.950 259.500 604.050 261.600 ;
        RECT 605.400 247.050 606.450 304.950 ;
        RECT 611.400 301.050 612.450 304.950 ;
        RECT 610.950 298.950 613.050 301.050 ;
        RECT 607.950 283.950 610.050 286.050 ;
        RECT 604.950 244.950 607.050 247.050 ;
        RECT 605.400 244.050 606.450 244.950 ;
        RECT 598.950 241.950 601.050 244.050 ;
        RECT 604.950 241.950 607.050 244.050 ;
        RECT 577.950 239.250 580.050 240.150 ;
        RECT 580.950 239.850 583.050 240.750 ;
        RECT 583.950 239.250 585.750 240.150 ;
        RECT 586.950 238.950 589.050 241.050 ;
        RECT 589.950 238.950 592.050 241.050 ;
        RECT 577.950 235.950 580.050 238.050 ;
        RECT 583.950 235.950 586.050 238.050 ;
        RECT 587.250 236.850 589.050 237.750 ;
        RECT 578.400 235.050 579.450 235.950 ;
        RECT 577.950 232.950 580.050 235.050 ;
        RECT 580.950 202.950 583.050 205.050 ;
        RECT 581.400 199.050 582.450 202.950 ;
        RECT 586.950 200.250 589.050 201.150 ;
        RECT 571.950 196.950 574.050 199.050 ;
        RECT 574.950 196.950 577.050 199.050 ;
        RECT 577.950 197.250 579.750 198.150 ;
        RECT 580.950 196.950 583.050 199.050 ;
        RECT 584.250 197.250 585.750 198.150 ;
        RECT 586.950 196.950 589.050 199.050 ;
        RECT 562.950 187.500 565.050 189.600 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 535.950 164.850 537.750 165.750 ;
        RECT 538.950 163.950 541.050 166.050 ;
        RECT 542.250 164.850 543.750 165.750 ;
        RECT 544.950 163.950 547.050 166.050 ;
        RECT 539.400 163.050 540.450 163.950 ;
        RECT 538.950 160.950 541.050 163.050 ;
        RECT 544.950 161.850 547.050 162.750 ;
        RECT 554.400 130.050 555.450 178.950 ;
        RECT 556.950 169.950 559.050 172.050 ;
        RECT 556.950 167.850 559.050 168.750 ;
        RECT 559.950 167.250 562.050 168.150 ;
        RECT 559.950 163.950 562.050 166.050 ;
        RECT 572.400 136.050 573.450 196.950 ;
        RECT 577.950 193.950 580.050 196.050 ;
        RECT 581.250 194.850 582.750 195.750 ;
        RECT 583.950 193.950 586.050 196.050 ;
        RECT 578.400 187.050 579.450 193.950 ;
        RECT 574.950 184.950 577.050 187.050 ;
        RECT 577.950 184.950 580.050 187.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 575.400 130.050 576.450 184.950 ;
        RECT 584.400 175.050 585.450 193.950 ;
        RECT 590.400 193.050 591.450 238.950 ;
        RECT 599.400 237.450 600.450 241.950 ;
        RECT 601.950 239.250 604.050 240.150 ;
        RECT 604.950 239.850 607.050 240.750 ;
        RECT 601.950 237.450 604.050 238.050 ;
        RECT 599.400 236.400 604.050 237.450 ;
        RECT 601.950 235.950 604.050 236.400 ;
        RECT 608.400 205.050 609.450 283.950 ;
        RECT 614.400 252.450 615.450 313.950 ;
        RECT 626.400 313.050 627.450 316.950 ;
        RECT 644.400 316.050 645.450 319.950 ;
        RECT 649.950 316.950 652.050 319.050 ;
        RECT 643.950 313.950 646.050 316.050 ;
        RECT 650.400 313.050 651.450 316.950 ;
        RECT 619.950 310.950 622.050 313.050 ;
        RECT 623.250 311.250 624.750 312.150 ;
        RECT 625.950 310.950 628.050 313.050 ;
        RECT 640.950 311.250 643.050 312.150 ;
        RECT 643.950 311.850 646.050 312.750 ;
        RECT 646.950 311.250 648.750 312.150 ;
        RECT 649.950 310.950 652.050 313.050 ;
        RECT 619.950 308.850 621.750 309.750 ;
        RECT 622.950 307.950 625.050 310.050 ;
        RECT 626.250 308.850 627.750 309.750 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 640.950 307.950 643.050 310.050 ;
        RECT 646.950 307.950 649.050 310.050 ;
        RECT 650.250 308.850 652.050 309.750 ;
        RECT 623.400 307.050 624.450 307.950 ;
        RECT 619.950 304.950 622.050 307.050 ;
        RECT 622.950 304.950 625.050 307.050 ;
        RECT 628.950 305.850 631.050 306.750 ;
        RECT 620.400 271.050 621.450 304.950 ;
        RECT 641.400 304.050 642.450 307.950 ;
        RECT 647.400 307.050 648.450 307.950 ;
        RECT 646.950 304.950 649.050 307.050 ;
        RECT 640.950 301.950 643.050 304.050 ;
        RECT 653.400 283.050 654.450 338.400 ;
        RECT 658.950 337.950 661.050 340.050 ;
        RECT 662.250 338.850 663.750 339.750 ;
        RECT 664.950 337.950 667.050 340.050 ;
        RECT 659.400 331.050 660.450 337.950 ;
        RECT 677.400 334.050 678.450 373.950 ;
        RECT 692.550 371.700 693.750 375.300 ;
        RECT 691.950 369.600 694.050 371.700 ;
        RECT 695.400 349.050 696.450 424.950 ;
        RECT 706.950 417.450 709.050 418.050 ;
        RECT 704.250 416.250 705.750 417.150 ;
        RECT 706.950 416.400 711.450 417.450 ;
        RECT 706.950 415.950 709.050 416.400 ;
        RECT 700.950 413.850 702.750 414.750 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 707.250 413.850 709.050 414.750 ;
        RECT 710.400 409.050 711.450 416.400 ;
        RECT 709.950 406.950 712.050 409.050 ;
        RECT 713.400 406.050 714.450 505.950 ;
        RECT 719.400 460.050 720.450 532.950 ;
        RECT 725.400 499.050 726.450 557.400 ;
        RECT 730.950 556.950 733.050 557.400 ;
        RECT 734.250 557.250 735.750 558.150 ;
        RECT 736.950 556.950 739.050 559.050 ;
        RECT 740.250 557.250 742.050 558.150 ;
        RECT 733.950 553.950 736.050 556.050 ;
        RECT 737.250 554.850 738.750 555.750 ;
        RECT 739.950 553.950 742.050 556.050 ;
        RECT 746.400 553.050 747.450 580.950 ;
        RECT 749.400 577.050 750.450 670.950 ;
        RECT 752.400 661.050 753.450 673.950 ;
        RECT 751.950 658.950 754.050 661.050 ;
        RECT 751.950 629.250 754.050 630.150 ;
        RECT 751.950 627.450 754.050 628.050 ;
        RECT 755.400 627.450 756.450 688.950 ;
        RECT 758.400 682.050 759.450 763.950 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 766.950 751.950 769.050 754.050 ;
        RECT 767.400 742.050 768.450 751.950 ;
        RECT 770.400 745.050 771.450 757.950 ;
        RECT 776.400 745.050 777.450 808.950 ;
        RECT 778.950 805.950 781.050 808.050 ;
        RECT 769.950 742.950 772.050 745.050 ;
        RECT 773.250 743.250 774.750 744.150 ;
        RECT 775.950 742.950 778.050 745.050 ;
        RECT 766.950 739.950 769.050 742.050 ;
        RECT 770.250 740.850 771.750 741.750 ;
        RECT 772.950 739.950 775.050 742.050 ;
        RECT 776.250 740.850 778.050 741.750 ;
        RECT 773.400 739.050 774.450 739.950 ;
        RECT 760.950 736.950 763.050 739.050 ;
        RECT 766.950 737.850 769.050 738.750 ;
        RECT 772.950 736.950 775.050 739.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 761.400 676.050 762.450 736.950 ;
        RECT 763.950 704.250 766.050 705.150 ;
        RECT 763.950 700.950 766.050 703.050 ;
        RECT 767.250 701.250 768.750 702.150 ;
        RECT 769.950 700.950 772.050 703.050 ;
        RECT 773.250 701.250 775.050 702.150 ;
        RECT 775.950 700.950 778.050 703.050 ;
        RECT 766.950 697.950 769.050 700.050 ;
        RECT 770.250 698.850 771.750 699.750 ;
        RECT 772.950 697.950 775.050 700.050 ;
        RECT 773.400 688.050 774.450 697.950 ;
        RECT 772.950 685.950 775.050 688.050 ;
        RECT 760.950 673.950 763.050 676.050 ;
        RECT 769.950 670.950 772.050 673.050 ;
        RECT 773.400 672.450 774.450 685.950 ;
        RECT 776.400 676.050 777.450 700.950 ;
        RECT 779.400 688.050 780.450 805.950 ;
        RECT 781.950 775.950 784.050 778.050 ;
        RECT 782.400 769.050 783.450 775.950 ;
        RECT 781.950 766.950 784.050 769.050 ;
        RECT 785.400 768.450 786.450 817.950 ;
        RECT 788.400 814.050 789.450 847.950 ;
        RECT 797.400 847.050 798.450 847.950 ;
        RECT 790.950 844.950 793.050 847.050 ;
        RECT 794.250 845.250 795.750 846.150 ;
        RECT 796.950 844.950 799.050 847.050 ;
        RECT 800.250 845.250 802.050 846.150 ;
        RECT 793.950 841.950 796.050 844.050 ;
        RECT 797.250 842.850 798.750 843.750 ;
        RECT 799.950 841.950 802.050 844.050 ;
        RECT 794.400 841.050 795.450 841.950 ;
        RECT 793.950 838.950 796.050 841.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 791.400 814.050 792.450 835.950 ;
        RECT 793.950 817.950 796.050 820.050 ;
        RECT 793.950 815.850 796.050 816.750 ;
        RECT 796.950 815.250 799.050 816.150 ;
        RECT 787.950 811.950 790.050 814.050 ;
        RECT 790.950 811.950 793.050 814.050 ;
        RECT 796.950 811.950 799.050 814.050 ;
        RECT 799.950 811.950 802.050 814.050 ;
        RECT 797.400 811.050 798.450 811.950 ;
        RECT 796.950 808.950 799.050 811.050 ;
        RECT 787.950 776.250 790.050 777.150 ;
        RECT 793.950 775.950 796.050 778.050 ;
        RECT 794.400 775.050 795.450 775.950 ;
        RECT 787.950 772.950 790.050 775.050 ;
        RECT 791.250 773.250 792.750 774.150 ;
        RECT 793.950 772.950 796.050 775.050 ;
        RECT 797.250 773.250 799.050 774.150 ;
        RECT 788.400 772.050 789.450 772.950 ;
        RECT 787.950 769.950 790.050 772.050 ;
        RECT 790.950 769.950 793.050 772.050 ;
        RECT 794.250 770.850 795.750 771.750 ;
        RECT 796.950 769.950 799.050 772.050 ;
        RECT 791.400 769.050 792.450 769.950 ;
        RECT 785.400 767.400 789.450 768.450 ;
        RECT 784.950 749.400 787.050 751.500 ;
        RECT 781.950 746.250 784.050 747.150 ;
        RECT 781.950 742.950 784.050 745.050 ;
        RECT 785.550 737.400 786.750 749.400 ;
        RECT 788.400 745.050 789.450 767.400 ;
        RECT 790.950 766.950 793.050 769.050 ;
        RECT 793.950 760.950 796.050 763.050 ;
        RECT 790.950 754.950 793.050 757.050 ;
        RECT 787.950 742.950 790.050 745.050 ;
        RECT 784.950 735.300 787.050 737.400 ;
        RECT 785.550 731.700 786.750 735.300 ;
        RECT 784.950 729.600 787.050 731.700 ;
        RECT 781.950 710.400 784.050 712.500 ;
        RECT 782.400 693.600 783.600 710.400 ;
        RECT 787.950 701.250 790.050 702.150 ;
        RECT 787.950 697.950 790.050 700.050 ;
        RECT 781.950 691.500 784.050 693.600 ;
        RECT 778.950 685.950 781.050 688.050 ;
        RECT 775.950 673.950 778.050 676.050 ;
        RECT 775.950 672.450 778.050 673.050 ;
        RECT 773.400 671.400 778.050 672.450 ;
        RECT 757.950 668.250 759.750 669.150 ;
        RECT 760.950 667.950 763.050 670.050 ;
        RECT 764.250 668.250 766.050 669.150 ;
        RECT 757.950 664.950 760.050 667.050 ;
        RECT 761.250 665.850 762.750 666.750 ;
        RECT 763.950 664.950 766.050 667.050 ;
        RECT 763.950 661.950 766.050 664.050 ;
        RECT 760.950 639.300 763.050 641.400 ;
        RECT 761.250 635.700 762.450 639.300 ;
        RECT 760.950 633.600 763.050 635.700 ;
        RECT 764.400 634.050 765.450 661.950 ;
        RECT 751.950 626.400 756.450 627.450 ;
        RECT 751.950 625.950 754.050 626.400 ;
        RECT 752.400 607.050 753.450 625.950 ;
        RECT 761.250 621.600 762.450 633.600 ;
        RECT 763.950 631.950 766.050 634.050 ;
        RECT 764.400 628.050 765.450 631.950 ;
        RECT 770.400 628.050 771.450 670.950 ;
        RECT 773.400 667.050 774.450 671.400 ;
        RECT 775.950 670.950 778.050 671.400 ;
        RECT 779.250 671.250 780.750 672.150 ;
        RECT 781.950 670.950 784.050 673.050 ;
        RECT 775.950 668.850 777.750 669.750 ;
        RECT 778.950 667.950 781.050 670.050 ;
        RECT 782.250 668.850 783.750 669.750 ;
        RECT 784.950 667.950 787.050 670.050 ;
        RECT 772.950 664.950 775.050 667.050 ;
        RECT 772.950 663.450 775.050 664.050 ;
        RECT 772.950 662.400 777.450 663.450 ;
        RECT 772.950 661.950 775.050 662.400 ;
        RECT 772.950 658.950 775.050 661.050 ;
        RECT 763.950 625.950 766.050 628.050 ;
        RECT 769.950 625.950 772.050 628.050 ;
        RECT 763.950 623.850 766.050 624.750 ;
        RECT 760.950 619.500 763.050 621.600 ;
        RECT 751.950 604.950 754.050 607.050 ;
        RECT 757.950 599.850 760.050 600.750 ;
        RECT 760.950 599.250 763.050 600.150 ;
        RECT 773.400 598.050 774.450 658.950 ;
        RECT 776.400 654.450 777.450 662.400 ;
        RECT 779.400 658.050 780.450 667.950 ;
        RECT 784.950 665.850 787.050 666.750 ;
        RECT 791.400 661.050 792.450 754.950 ;
        RECT 794.400 745.050 795.450 760.950 ;
        RECT 797.400 757.050 798.450 769.950 ;
        RECT 800.400 759.450 801.450 811.950 ;
        RECT 806.400 778.050 807.450 883.950 ;
        RECT 817.950 853.950 820.050 856.050 ;
        RECT 818.400 847.050 819.450 853.950 ;
        RECT 821.400 853.050 822.450 887.400 ;
        RECT 823.950 886.950 826.050 889.050 ;
        RECT 832.950 887.250 835.050 888.150 ;
        RECT 835.950 887.850 838.050 888.750 ;
        RECT 820.950 850.950 823.050 853.050 ;
        RECT 811.950 846.450 814.050 847.050 ;
        RECT 809.400 845.400 814.050 846.450 ;
        RECT 809.400 823.050 810.450 845.400 ;
        RECT 811.950 844.950 814.050 845.400 ;
        RECT 817.950 844.950 820.050 847.050 ;
        RECT 821.250 845.250 823.050 846.150 ;
        RECT 824.400 844.050 825.450 886.950 ;
        RECT 832.950 883.950 835.050 886.050 ;
        RECT 844.950 884.250 846.750 885.150 ;
        RECT 847.950 883.950 850.050 886.050 ;
        RECT 851.250 884.250 853.050 885.150 ;
        RECT 833.400 883.050 834.450 883.950 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 844.950 880.950 847.050 883.050 ;
        RECT 848.250 881.850 849.750 882.750 ;
        RECT 850.950 880.950 853.050 883.050 ;
        RECT 832.950 850.950 835.050 853.050 ;
        RECT 826.950 847.950 829.050 850.050 ;
        RECT 811.950 842.850 814.050 843.750 ;
        RECT 814.950 842.250 817.050 843.150 ;
        RECT 817.950 842.850 819.750 843.750 ;
        RECT 820.950 841.950 823.050 844.050 ;
        RECT 823.950 841.950 826.050 844.050 ;
        RECT 821.400 841.050 822.450 841.950 ;
        RECT 814.950 838.950 817.050 841.050 ;
        RECT 820.950 838.950 823.050 841.050 ;
        RECT 814.950 832.950 817.050 835.050 ;
        RECT 808.950 820.950 811.050 823.050 ;
        RECT 811.950 820.950 814.050 823.050 ;
        RECT 808.950 814.950 811.050 817.050 ;
        RECT 809.400 805.050 810.450 814.950 ;
        RECT 812.400 811.050 813.450 820.950 ;
        RECT 815.400 817.050 816.450 832.950 ;
        RECT 817.950 820.950 820.050 823.050 ;
        RECT 818.400 820.050 819.450 820.950 ;
        RECT 817.950 817.950 820.050 820.050 ;
        RECT 814.950 814.950 817.050 817.050 ;
        RECT 818.250 815.850 819.750 816.750 ;
        RECT 820.950 816.450 823.050 817.050 ;
        RECT 824.400 816.450 825.450 841.950 ;
        RECT 827.400 841.050 828.450 847.950 ;
        RECT 829.950 844.950 832.050 847.050 ;
        RECT 826.950 838.950 829.050 841.050 ;
        RECT 830.400 837.450 831.450 844.950 ;
        RECT 833.400 843.450 834.450 850.950 ;
        RECT 835.950 848.250 838.050 849.150 ;
        RECT 841.950 847.950 844.050 850.050 ;
        RECT 845.400 849.450 846.450 880.950 ;
        RECT 853.950 855.300 856.050 857.400 ;
        RECT 854.550 851.700 855.750 855.300 ;
        RECT 853.950 849.600 856.050 851.700 ;
        RECT 845.400 848.400 849.450 849.450 ;
        RECT 842.400 847.050 843.450 847.950 ;
        RECT 835.950 844.950 838.050 847.050 ;
        RECT 839.250 845.250 840.750 846.150 ;
        RECT 841.950 844.950 844.050 847.050 ;
        RECT 845.250 845.250 847.050 846.150 ;
        RECT 838.950 843.450 841.050 844.050 ;
        RECT 833.400 842.400 841.050 843.450 ;
        RECT 842.250 842.850 843.750 843.750 ;
        RECT 838.950 841.950 841.050 842.400 ;
        RECT 844.950 841.950 847.050 844.050 ;
        RECT 841.950 838.950 844.050 841.050 ;
        RECT 820.950 815.400 825.450 816.450 ;
        RECT 820.950 814.950 823.050 815.400 ;
        RECT 814.950 812.850 817.050 813.750 ;
        RECT 820.950 812.850 823.050 813.750 ;
        RECT 824.400 811.050 825.450 815.400 ;
        RECT 827.400 836.400 831.450 837.450 ;
        RECT 811.950 808.950 814.050 811.050 ;
        RECT 820.950 808.950 823.050 811.050 ;
        RECT 823.950 808.950 826.050 811.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 802.950 775.950 805.050 778.050 ;
        RECT 805.950 775.950 808.050 778.050 ;
        RECT 814.950 776.250 817.050 777.150 ;
        RECT 803.400 763.050 804.450 775.950 ;
        RECT 805.950 773.250 807.750 774.150 ;
        RECT 808.950 772.950 811.050 775.050 ;
        RECT 812.250 773.250 813.750 774.150 ;
        RECT 814.950 772.950 817.050 775.050 ;
        RECT 805.950 769.950 808.050 772.050 ;
        RECT 809.250 770.850 810.750 771.750 ;
        RECT 811.950 769.950 814.050 772.050 ;
        RECT 814.950 769.950 817.050 772.050 ;
        RECT 806.400 766.050 807.450 769.950 ;
        RECT 808.950 766.950 811.050 769.050 ;
        RECT 805.950 763.950 808.050 766.050 ;
        RECT 802.950 760.950 805.050 763.050 ;
        RECT 800.400 758.400 804.450 759.450 ;
        RECT 796.950 754.950 799.050 757.050 ;
        RECT 799.950 745.950 802.050 748.050 ;
        RECT 800.400 745.050 801.450 745.950 ;
        RECT 793.950 744.450 796.050 745.050 ;
        RECT 793.950 743.400 798.450 744.450 ;
        RECT 793.950 742.950 796.050 743.400 ;
        RECT 793.950 740.850 796.050 741.750 ;
        RECT 793.950 701.250 796.050 702.150 ;
        RECT 793.950 697.950 796.050 700.050 ;
        RECT 794.400 691.050 795.450 697.950 ;
        RECT 797.400 691.050 798.450 743.400 ;
        RECT 799.950 742.950 802.050 745.050 ;
        RECT 799.950 740.850 802.050 741.750 ;
        RECT 803.400 739.050 804.450 758.400 ;
        RECT 805.950 749.400 808.050 751.500 ;
        RECT 802.950 736.950 805.050 739.050 ;
        RECT 806.400 732.600 807.600 749.400 ;
        RECT 805.950 730.500 808.050 732.600 ;
        RECT 802.950 711.300 805.050 713.400 ;
        RECT 803.250 707.700 804.450 711.300 ;
        RECT 802.950 705.600 805.050 707.700 ;
        RECT 803.250 693.600 804.450 705.600 ;
        RECT 805.950 703.950 808.050 706.050 ;
        RECT 806.400 703.050 807.450 703.950 ;
        RECT 805.950 700.950 808.050 703.050 ;
        RECT 806.400 700.050 807.450 700.950 ;
        RECT 805.950 697.950 808.050 700.050 ;
        RECT 805.950 695.850 808.050 696.750 ;
        RECT 802.950 691.500 805.050 693.600 ;
        RECT 793.950 688.950 796.050 691.050 ;
        RECT 796.950 688.950 799.050 691.050 ;
        RECT 793.950 685.950 796.050 688.050 ;
        RECT 790.950 658.950 793.050 661.050 ;
        RECT 794.400 660.450 795.450 685.950 ;
        RECT 805.950 670.950 808.050 673.050 ;
        RECT 796.950 668.250 798.750 669.150 ;
        RECT 799.950 667.950 802.050 670.050 ;
        RECT 803.250 668.250 805.050 669.150 ;
        RECT 806.400 667.050 807.450 670.950 ;
        RECT 796.950 664.950 799.050 667.050 ;
        RECT 800.250 665.850 801.750 666.750 ;
        RECT 802.950 666.450 805.050 667.050 ;
        RECT 805.950 666.450 808.050 667.050 ;
        RECT 802.950 665.400 808.050 666.450 ;
        RECT 802.950 664.950 805.050 665.400 ;
        RECT 805.950 664.950 808.050 665.400 ;
        RECT 797.400 664.050 798.450 664.950 ;
        RECT 796.950 661.950 799.050 664.050 ;
        RECT 794.400 659.400 798.450 660.450 ;
        RECT 778.950 655.950 781.050 658.050 ;
        RECT 776.400 653.400 780.450 654.450 ;
        RECT 775.950 649.950 778.050 652.050 ;
        RECT 776.400 622.050 777.450 649.950 ;
        RECT 775.950 619.950 778.050 622.050 ;
        RECT 779.400 598.050 780.450 653.400 ;
        RECT 790.950 631.950 793.050 634.050 ;
        RECT 791.400 631.050 792.450 631.950 ;
        RECT 781.950 629.250 783.750 630.150 ;
        RECT 784.950 628.950 787.050 631.050 ;
        RECT 788.250 629.250 789.750 630.150 ;
        RECT 790.950 628.950 793.050 631.050 ;
        RECT 794.250 629.250 796.050 630.150 ;
        RECT 781.950 625.950 784.050 628.050 ;
        RECT 785.250 626.850 786.750 627.750 ;
        RECT 787.950 625.950 790.050 628.050 ;
        RECT 791.250 626.850 792.750 627.750 ;
        RECT 793.950 625.950 796.050 628.050 ;
        RECT 782.400 625.050 783.450 625.950 ;
        RECT 781.950 622.950 784.050 625.050 ;
        RECT 784.950 622.950 787.050 625.050 ;
        RECT 782.400 601.050 783.450 622.950 ;
        RECT 785.400 601.050 786.450 622.950 ;
        RECT 788.400 622.050 789.450 625.950 ;
        RECT 790.950 622.950 793.050 625.050 ;
        RECT 787.950 619.950 790.050 622.050 ;
        RECT 781.950 598.950 784.050 601.050 ;
        RECT 784.950 598.950 787.050 601.050 ;
        RECT 757.950 595.950 760.050 598.050 ;
        RECT 760.950 595.950 763.050 598.050 ;
        RECT 772.950 595.950 775.050 598.050 ;
        RECT 775.950 596.250 777.750 597.150 ;
        RECT 778.950 595.950 781.050 598.050 ;
        RECT 782.250 596.250 784.050 597.150 ;
        RECT 784.950 595.950 787.050 598.050 ;
        RECT 748.950 574.950 751.050 577.050 ;
        RECT 754.950 556.950 757.050 559.050 ;
        RECT 748.950 553.950 751.050 556.050 ;
        RECT 751.950 554.250 754.050 555.150 ;
        RECT 754.950 554.850 757.050 555.750 ;
        RECT 739.950 550.950 742.050 553.050 ;
        RECT 745.950 550.950 748.050 553.050 ;
        RECT 749.400 552.450 750.450 553.950 ;
        RECT 751.950 552.450 754.050 553.050 ;
        RECT 749.400 551.400 754.050 552.450 ;
        RECT 733.950 547.950 736.050 550.050 ;
        RECT 727.950 529.950 730.050 532.050 ;
        RECT 727.950 527.850 730.050 528.750 ;
        RECT 730.950 527.250 733.050 528.150 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 731.400 523.050 732.450 523.950 ;
        RECT 730.950 520.950 733.050 523.050 ;
        RECT 724.950 496.950 727.050 499.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 722.400 480.450 723.450 490.950 ;
        RECT 728.400 487.050 729.450 490.950 ;
        RECT 727.950 484.950 730.050 487.050 ;
        RECT 724.950 482.250 727.050 483.150 ;
        RECT 727.950 482.850 730.050 483.750 ;
        RECT 724.950 480.450 727.050 481.050 ;
        RECT 722.400 479.400 727.050 480.450 ;
        RECT 724.950 478.950 727.050 479.400 ;
        RECT 721.950 463.950 724.050 466.050 ;
        RECT 718.950 457.950 721.050 460.050 ;
        RECT 722.400 457.050 723.450 463.950 ;
        RECT 725.400 463.050 726.450 478.950 ;
        RECT 724.950 460.950 727.050 463.050 ;
        RECT 721.950 454.950 724.050 457.050 ;
        RECT 725.250 455.250 726.750 456.150 ;
        RECT 727.950 454.950 730.050 457.050 ;
        RECT 730.950 454.950 733.050 457.050 ;
        RECT 718.950 453.450 721.050 454.050 ;
        RECT 716.400 452.400 721.050 453.450 ;
        RECT 722.250 452.850 723.750 453.750 ;
        RECT 716.400 451.050 717.450 452.400 ;
        RECT 718.950 451.950 721.050 452.400 ;
        RECT 724.950 451.950 727.050 454.050 ;
        RECT 728.250 452.850 730.050 453.750 ;
        RECT 715.950 448.950 718.050 451.050 ;
        RECT 718.950 449.850 721.050 450.750 ;
        RECT 727.950 448.950 730.050 451.050 ;
        RECT 718.950 418.950 721.050 421.050 ;
        RECT 719.400 415.050 720.450 418.950 ;
        RECT 724.950 416.250 727.050 417.150 ;
        RECT 715.950 413.250 717.750 414.150 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 722.250 413.250 723.750 414.150 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 715.950 409.950 718.050 412.050 ;
        RECT 719.250 410.850 720.750 411.750 ;
        RECT 721.950 409.950 724.050 412.050 ;
        RECT 716.400 409.050 717.450 409.950 ;
        RECT 715.950 406.950 718.050 409.050 ;
        RECT 712.950 403.950 715.050 406.050 ;
        RECT 703.950 400.950 706.050 403.050 ;
        RECT 700.950 382.950 703.050 385.050 ;
        RECT 700.950 380.850 703.050 381.750 ;
        RECT 694.950 346.950 697.050 349.050 ;
        RECT 679.950 343.950 682.050 346.050 ;
        RECT 676.950 331.950 679.050 334.050 ;
        RECT 658.950 328.950 661.050 331.050 ;
        RECT 676.950 322.950 679.050 325.050 ;
        RECT 664.950 319.950 667.050 322.050 ;
        RECT 658.950 310.950 661.050 313.050 ;
        RECT 659.400 304.050 660.450 310.950 ;
        RECT 661.950 307.950 664.050 310.050 ;
        RECT 665.400 307.050 666.450 319.950 ;
        RECT 673.950 313.950 676.050 316.050 ;
        RECT 667.950 310.950 670.050 313.050 ;
        RECT 668.400 310.050 669.450 310.950 ;
        RECT 667.950 307.950 670.050 310.050 ;
        RECT 671.250 308.250 673.050 309.150 ;
        RECT 674.400 307.050 675.450 313.950 ;
        RECT 677.400 310.050 678.450 322.950 ;
        RECT 676.950 307.950 679.050 310.050 ;
        RECT 661.950 305.850 663.750 306.750 ;
        RECT 664.950 304.950 667.050 307.050 ;
        RECT 668.250 305.850 669.750 306.750 ;
        RECT 670.950 306.450 673.050 307.050 ;
        RECT 673.950 306.450 676.050 307.050 ;
        RECT 670.950 305.400 676.050 306.450 ;
        RECT 670.950 304.950 673.050 305.400 ;
        RECT 673.950 304.950 676.050 305.400 ;
        RECT 658.950 301.950 661.050 304.050 ;
        RECT 664.950 302.850 667.050 303.750 ;
        RECT 652.950 280.950 655.050 283.050 ;
        RECT 670.950 280.950 673.050 283.050 ;
        RECT 664.950 277.950 667.050 280.050 ;
        RECT 634.950 272.250 637.050 273.150 ;
        RECT 619.950 268.950 622.050 271.050 ;
        RECT 634.950 268.950 637.050 271.050 ;
        RECT 638.250 269.250 639.750 270.150 ;
        RECT 640.950 268.950 643.050 271.050 ;
        RECT 644.250 269.250 646.050 270.150 ;
        RECT 655.950 268.950 658.050 271.050 ;
        RECT 616.950 266.250 619.050 267.150 ;
        RECT 619.950 266.850 622.050 267.750 ;
        RECT 616.950 262.950 619.050 265.050 ;
        RECT 635.400 264.450 636.450 268.950 ;
        RECT 665.400 268.050 666.450 277.950 ;
        RECT 671.400 271.050 672.450 280.950 ;
        RECT 676.950 272.250 679.050 273.150 ;
        RECT 667.950 269.250 669.750 270.150 ;
        RECT 670.950 268.950 673.050 271.050 ;
        RECT 674.250 269.250 675.750 270.150 ;
        RECT 676.950 268.950 679.050 271.050 ;
        RECT 637.950 265.950 640.050 268.050 ;
        RECT 641.250 266.850 642.750 267.750 ;
        RECT 643.950 265.950 646.050 268.050 ;
        RECT 655.950 266.850 658.050 267.750 ;
        RECT 664.950 267.450 667.050 268.050 ;
        RECT 667.950 267.450 670.050 268.050 ;
        RECT 658.950 266.250 661.050 267.150 ;
        RECT 664.950 266.400 670.050 267.450 ;
        RECT 671.250 266.850 672.750 267.750 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 667.950 265.950 670.050 266.400 ;
        RECT 673.950 265.950 676.050 268.050 ;
        RECT 635.400 263.400 639.450 264.450 ;
        RECT 614.400 251.400 618.450 252.450 ;
        RECT 613.950 245.400 616.050 247.500 ;
        RECT 610.950 242.250 613.050 243.150 ;
        RECT 610.950 238.950 613.050 241.050 ;
        RECT 611.400 238.050 612.450 238.950 ;
        RECT 610.950 235.950 613.050 238.050 ;
        RECT 614.550 233.400 615.750 245.400 ;
        RECT 613.950 231.300 616.050 233.400 ;
        RECT 610.950 226.950 613.050 229.050 ;
        RECT 614.550 227.700 615.750 231.300 ;
        RECT 607.950 202.950 610.050 205.050 ;
        RECT 608.400 202.050 609.450 202.950 ;
        RECT 605.250 200.250 606.750 201.150 ;
        RECT 607.950 199.950 610.050 202.050 ;
        RECT 611.400 199.050 612.450 226.950 ;
        RECT 613.950 225.600 616.050 227.700 ;
        RECT 601.950 197.850 603.750 198.750 ;
        RECT 604.950 196.950 607.050 199.050 ;
        RECT 608.250 197.850 610.050 198.750 ;
        RECT 610.950 196.950 613.050 199.050 ;
        RECT 589.950 190.950 592.050 193.050 ;
        RECT 589.950 184.950 592.050 187.050 ;
        RECT 583.950 172.950 586.050 175.050 ;
        RECT 583.950 169.950 586.050 172.050 ;
        RECT 584.400 169.050 585.450 169.950 ;
        RECT 590.400 169.050 591.450 184.950 ;
        RECT 604.950 178.950 607.050 181.050 ;
        RECT 598.950 173.400 601.050 175.500 ;
        RECT 577.950 166.950 580.050 169.050 ;
        RECT 581.250 167.250 582.750 168.150 ;
        RECT 583.950 166.950 586.050 169.050 ;
        RECT 587.250 167.250 588.750 168.150 ;
        RECT 589.950 166.950 592.050 169.050 ;
        RECT 577.950 164.850 579.750 165.750 ;
        RECT 580.950 163.950 583.050 166.050 ;
        RECT 584.250 164.850 585.750 165.750 ;
        RECT 586.950 163.950 589.050 166.050 ;
        RECT 590.250 164.850 592.050 165.750 ;
        RECT 587.400 151.050 588.450 163.950 ;
        RECT 599.400 156.600 600.600 173.400 ;
        RECT 605.400 169.050 606.450 178.950 ;
        RECT 610.950 175.950 613.050 178.050 ;
        RECT 611.400 169.050 612.450 175.950 ;
        RECT 617.400 175.050 618.450 251.400 ;
        RECT 634.950 245.400 637.050 247.500 ;
        RECT 622.950 238.950 625.050 241.050 ;
        RECT 628.950 238.950 631.050 241.050 ;
        RECT 622.950 236.850 625.050 237.750 ;
        RECT 628.950 236.850 631.050 237.750 ;
        RECT 635.400 228.600 636.600 245.400 ;
        RECT 634.950 226.500 637.050 228.600 ;
        RECT 619.950 208.950 622.050 211.050 ;
        RECT 620.400 202.050 621.450 208.950 ;
        RECT 619.950 199.950 622.050 202.050 ;
        RECT 625.950 201.450 628.050 202.050 ;
        RECT 623.250 200.250 624.750 201.150 ;
        RECT 625.950 200.400 630.450 201.450 ;
        RECT 625.950 199.950 628.050 200.400 ;
        RECT 619.950 197.850 621.750 198.750 ;
        RECT 622.950 196.950 625.050 199.050 ;
        RECT 626.250 197.850 628.050 198.750 ;
        RECT 629.400 193.050 630.450 200.400 ;
        RECT 638.400 199.050 639.450 263.400 ;
        RECT 658.950 262.950 661.050 265.050 ;
        RECT 652.950 241.950 655.050 244.050 ;
        RECT 653.400 241.050 654.450 241.950 ;
        RECT 652.950 238.950 655.050 241.050 ;
        RECT 656.250 239.250 657.750 240.150 ;
        RECT 658.950 238.950 661.050 241.050 ;
        RECT 652.950 236.850 654.750 237.750 ;
        RECT 655.950 235.950 658.050 238.050 ;
        RECT 659.250 236.850 660.750 237.750 ;
        RECT 661.950 235.950 664.050 238.050 ;
        RECT 649.950 232.950 652.050 235.050 ;
        RECT 650.400 202.050 651.450 232.950 ;
        RECT 656.400 229.050 657.450 235.950 ;
        RECT 665.400 235.050 666.450 265.950 ;
        RECT 667.950 241.950 670.050 244.050 ;
        RECT 661.950 233.850 664.050 234.750 ;
        RECT 664.950 232.950 667.050 235.050 ;
        RECT 655.950 226.950 658.050 229.050 ;
        RECT 661.950 214.950 664.050 217.050 ;
        RECT 652.950 205.950 655.050 208.050 ;
        RECT 647.250 200.250 648.750 201.150 ;
        RECT 649.950 199.950 652.050 202.050 ;
        RECT 637.950 196.950 640.050 199.050 ;
        RECT 643.950 197.850 645.750 198.750 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 650.250 197.850 652.050 198.750 ;
        RECT 628.950 190.950 631.050 193.050 ;
        RECT 616.950 172.950 619.050 175.050 ;
        RECT 619.950 173.400 622.050 175.500 ;
        RECT 604.950 166.950 607.050 169.050 ;
        RECT 610.950 166.950 613.050 169.050 ;
        RECT 604.950 164.850 607.050 165.750 ;
        RECT 610.950 164.850 613.050 165.750 ;
        RECT 620.250 161.400 621.450 173.400 ;
        RECT 622.950 170.250 625.050 171.150 ;
        RECT 629.400 169.050 630.450 190.950 ;
        RECT 622.950 166.950 625.050 169.050 ;
        RECT 628.950 166.950 631.050 169.050 ;
        RECT 637.950 166.950 640.050 169.050 ;
        RECT 643.950 166.950 646.050 169.050 ;
        RECT 647.250 167.250 648.750 168.150 ;
        RECT 649.950 166.950 652.050 169.050 ;
        RECT 619.950 159.300 622.050 161.400 ;
        RECT 598.950 154.500 601.050 156.600 ;
        RECT 620.250 155.700 621.450 159.300 ;
        RECT 619.950 153.600 622.050 155.700 ;
        RECT 586.950 148.950 589.050 151.050 ;
        RECT 629.400 148.050 630.450 166.950 ;
        RECT 638.400 157.050 639.450 166.950 ;
        RECT 640.950 163.950 643.050 166.050 ;
        RECT 644.250 164.850 645.750 165.750 ;
        RECT 646.950 163.950 649.050 166.050 ;
        RECT 650.250 164.850 652.050 165.750 ;
        RECT 640.950 161.850 643.050 162.750 ;
        RECT 643.950 160.950 646.050 163.050 ;
        RECT 637.950 154.950 640.050 157.050 ;
        RECT 628.950 145.950 631.050 148.050 ;
        RECT 553.950 127.950 556.050 130.050 ;
        RECT 556.950 128.250 559.050 129.150 ;
        RECT 574.950 127.950 577.050 130.050 ;
        RECT 589.950 127.950 592.050 130.050 ;
        RECT 595.950 127.950 598.050 130.050 ;
        RECT 535.950 124.950 538.050 127.050 ;
        RECT 547.950 125.250 549.750 126.150 ;
        RECT 550.950 124.950 553.050 127.050 ;
        RECT 554.250 125.250 555.750 126.150 ;
        RECT 556.950 124.950 559.050 127.050 ;
        RECT 571.950 124.950 574.050 127.050 ;
        RECT 535.950 122.850 538.050 123.750 ;
        RECT 538.950 122.250 541.050 123.150 ;
        RECT 547.950 121.950 550.050 124.050 ;
        RECT 551.250 122.850 552.750 123.750 ;
        RECT 553.950 121.950 556.050 124.050 ;
        RECT 568.950 122.250 571.050 123.150 ;
        RECT 571.950 122.850 574.050 123.750 ;
        RECT 554.400 121.050 555.450 121.950 ;
        RECT 538.950 118.950 541.050 121.050 ;
        RECT 553.950 118.950 556.050 121.050 ;
        RECT 568.950 118.950 571.050 121.050 ;
        RECT 554.400 97.050 555.450 118.950 ;
        RECT 569.400 115.050 570.450 118.950 ;
        RECT 568.950 112.950 571.050 115.050 ;
        RECT 565.950 106.950 568.050 109.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 544.950 96.450 547.050 97.050 ;
        RECT 542.400 95.400 547.050 96.450 ;
        RECT 542.400 91.050 543.450 95.400 ;
        RECT 544.950 94.950 547.050 95.400 ;
        RECT 553.950 94.950 556.050 97.050 ;
        RECT 563.400 94.050 564.450 100.950 ;
        RECT 566.400 97.050 567.450 106.950 ;
        RECT 575.400 103.050 576.450 127.950 ;
        RECT 590.400 127.050 591.450 127.950 ;
        RECT 577.950 124.950 580.050 127.050 ;
        RECT 583.950 124.950 586.050 127.050 ;
        RECT 589.950 124.950 592.050 127.050 ;
        RECT 593.250 125.250 595.050 126.150 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 574.950 94.950 577.050 97.050 ;
        RECT 544.950 92.850 547.050 93.750 ;
        RECT 547.950 92.250 550.050 93.150 ;
        RECT 553.950 92.850 556.050 93.750 ;
        RECT 562.950 91.950 565.050 94.050 ;
        RECT 566.400 91.050 567.450 94.950 ;
        RECT 568.950 91.950 571.050 94.050 ;
        RECT 572.250 92.250 574.050 93.150 ;
        RECT 541.950 88.950 544.050 91.050 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 562.950 89.850 564.750 90.750 ;
        RECT 565.950 88.950 568.050 91.050 ;
        RECT 569.250 89.850 570.750 90.750 ;
        RECT 571.950 90.450 574.050 91.050 ;
        RECT 575.400 90.450 576.450 94.950 ;
        RECT 578.400 94.050 579.450 124.950 ;
        RECT 583.950 122.850 586.050 123.750 ;
        RECT 586.950 122.250 589.050 123.150 ;
        RECT 589.950 122.850 591.750 123.750 ;
        RECT 592.950 121.950 595.050 124.050 ;
        RECT 586.950 118.950 589.050 121.050 ;
        RECT 587.400 109.050 588.450 118.950 ;
        RECT 586.950 106.950 589.050 109.050 ;
        RECT 596.400 106.050 597.450 127.950 ;
        RECT 607.950 125.250 609.750 126.150 ;
        RECT 610.950 124.950 613.050 127.050 ;
        RECT 616.950 124.950 619.050 127.050 ;
        RECT 631.950 124.950 634.050 127.050 ;
        RECT 640.950 124.950 643.050 127.050 ;
        RECT 607.950 121.950 610.050 124.050 ;
        RECT 611.250 122.850 613.050 123.750 ;
        RECT 613.950 122.250 616.050 123.150 ;
        RECT 616.950 122.850 619.050 123.750 ;
        RECT 631.950 122.850 634.050 123.750 ;
        RECT 634.950 122.250 637.050 123.150 ;
        RECT 595.950 103.950 598.050 106.050 ;
        RECT 592.950 94.950 595.050 97.050 ;
        RECT 577.950 91.950 580.050 94.050 ;
        RECT 586.950 92.250 588.750 93.150 ;
        RECT 589.950 91.950 592.050 94.050 ;
        RECT 593.400 91.050 594.450 94.950 ;
        RECT 596.400 94.050 597.450 103.950 ;
        RECT 608.400 96.450 609.450 121.950 ;
        RECT 613.950 118.950 616.050 121.050 ;
        RECT 619.950 118.950 622.050 121.050 ;
        RECT 634.950 118.950 637.050 121.050 ;
        RECT 614.400 97.050 615.450 118.950 ;
        RECT 605.400 95.400 609.450 96.450 ;
        RECT 595.950 91.950 598.050 94.050 ;
        RECT 571.950 89.400 576.450 90.450 ;
        RECT 571.950 88.950 574.050 89.400 ;
        RECT 586.950 88.950 589.050 91.050 ;
        RECT 590.250 89.850 591.750 90.750 ;
        RECT 592.950 88.950 595.050 91.050 ;
        RECT 596.250 89.850 598.050 90.750 ;
        RECT 548.400 88.050 549.450 88.950 ;
        RECT 547.950 85.950 550.050 88.050 ;
        RECT 565.950 86.850 568.050 87.750 ;
        RECT 532.950 82.950 535.050 85.050 ;
        RECT 526.950 70.950 529.050 73.050 ;
        RECT 521.400 68.400 525.450 69.450 ;
        RECT 505.950 59.250 508.050 60.150 ;
        RECT 517.950 58.950 520.050 61.050 ;
        RECT 518.400 58.050 519.450 58.950 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 56.250 504.750 57.150 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 511.950 57.450 514.050 58.050 ;
        RECT 509.250 56.250 510.750 57.150 ;
        RECT 511.950 56.400 516.450 57.450 ;
        RECT 511.950 55.950 514.050 56.400 ;
        RECT 500.400 54.450 501.450 55.950 ;
        RECT 506.400 55.050 507.450 55.950 ;
        RECT 502.950 54.450 505.050 55.050 ;
        RECT 500.400 53.400 505.050 54.450 ;
        RECT 502.950 52.950 505.050 53.400 ;
        RECT 505.950 52.950 508.050 55.050 ;
        RECT 508.950 52.950 511.050 55.050 ;
        RECT 512.250 53.850 514.050 54.750 ;
        RECT 503.400 34.050 504.450 52.950 ;
        RECT 509.400 52.050 510.450 52.950 ;
        RECT 508.950 49.950 511.050 52.050 ;
        RECT 502.950 31.950 505.050 34.050 ;
        RECT 505.950 28.950 508.050 31.050 ;
        RECT 496.950 25.950 499.050 28.050 ;
        RECT 497.400 25.050 498.450 25.950 ;
        RECT 496.950 22.950 499.050 25.050 ;
        RECT 500.250 23.250 501.750 24.150 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 506.400 22.050 507.450 28.950 ;
        RECT 515.400 28.050 516.450 56.400 ;
        RECT 517.950 55.950 520.050 58.050 ;
        RECT 518.400 49.050 519.450 55.950 ;
        RECT 517.950 46.950 520.050 49.050 ;
        RECT 521.400 31.050 522.450 68.400 ;
        RECT 527.400 61.050 528.450 70.950 ;
        RECT 587.400 67.050 588.450 88.950 ;
        RECT 592.950 86.850 595.050 87.750 ;
        RECT 605.400 70.050 606.450 95.400 ;
        RECT 613.950 94.950 616.050 97.050 ;
        RECT 607.950 91.950 610.050 94.050 ;
        RECT 610.950 92.250 612.750 93.150 ;
        RECT 613.950 91.950 616.050 94.050 ;
        RECT 617.250 92.250 619.050 93.150 ;
        RECT 608.400 90.450 609.450 91.950 ;
        RECT 610.950 90.450 613.050 91.050 ;
        RECT 608.400 89.400 613.050 90.450 ;
        RECT 614.250 89.850 615.750 90.750 ;
        RECT 616.950 90.450 619.050 91.050 ;
        RECT 620.400 90.450 621.450 118.950 ;
        RECT 635.400 118.050 636.450 118.950 ;
        RECT 634.950 115.950 637.050 118.050 ;
        RECT 634.950 106.950 637.050 109.050 ;
        RECT 625.950 96.450 628.050 97.050 ;
        RECT 623.400 95.400 628.050 96.450 ;
        RECT 623.400 94.050 624.450 95.400 ;
        RECT 625.950 94.950 628.050 95.400 ;
        RECT 629.250 95.250 630.750 96.150 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 635.400 94.050 636.450 106.950 ;
        RECT 637.950 97.950 640.050 100.050 ;
        RECT 622.950 91.950 625.050 94.050 ;
        RECT 625.950 92.850 627.750 93.750 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 632.250 92.850 633.750 93.750 ;
        RECT 634.950 91.950 637.050 94.050 ;
        RECT 610.950 88.950 613.050 89.400 ;
        RECT 616.950 89.400 621.450 90.450 ;
        RECT 616.950 88.950 619.050 89.400 ;
        RECT 604.950 67.950 607.050 70.050 ;
        RECT 586.950 64.950 589.050 67.050 ;
        RECT 620.400 64.050 621.450 89.400 ;
        RECT 625.950 88.950 628.050 91.050 ;
        RECT 622.950 67.950 625.050 70.050 ;
        RECT 610.950 61.950 613.050 64.050 ;
        RECT 613.950 61.950 616.050 64.050 ;
        RECT 619.950 61.950 622.050 64.050 ;
        RECT 526.950 58.950 529.050 61.050 ;
        RECT 523.950 40.950 526.050 43.050 ;
        RECT 520.950 28.950 523.050 31.050 ;
        RECT 514.950 25.950 517.050 28.050 ;
        RECT 524.400 25.050 525.450 40.950 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 521.250 23.250 522.750 24.150 ;
        RECT 523.950 22.950 526.050 25.050 ;
        RECT 527.400 22.050 528.450 58.950 ;
        RECT 611.400 58.050 612.450 61.950 ;
        RECT 529.950 56.250 532.050 57.150 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 608.250 56.250 609.750 57.150 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 529.950 52.950 532.050 55.050 ;
        RECT 533.250 53.250 534.750 54.150 ;
        RECT 535.950 52.950 538.050 55.050 ;
        RECT 539.250 53.250 541.050 54.150 ;
        RECT 541.950 52.950 544.050 55.050 ;
        RECT 550.950 53.250 552.750 54.150 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 559.950 52.950 562.050 55.050 ;
        RECT 574.950 52.950 577.050 55.050 ;
        RECT 583.950 54.450 586.050 55.050 ;
        RECT 580.950 53.250 582.750 54.150 ;
        RECT 583.950 53.400 588.450 54.450 ;
        RECT 583.950 52.950 586.050 53.400 ;
        RECT 532.950 49.950 535.050 52.050 ;
        RECT 536.250 50.850 537.750 51.750 ;
        RECT 538.950 49.950 541.050 52.050 ;
        RECT 539.400 49.050 540.450 49.950 ;
        RECT 538.950 46.950 541.050 49.050 ;
        RECT 542.400 40.050 543.450 52.950 ;
        RECT 550.950 49.950 553.050 52.050 ;
        RECT 554.250 50.850 556.050 51.750 ;
        RECT 556.950 50.250 559.050 51.150 ;
        RECT 559.950 50.850 562.050 51.750 ;
        RECT 574.950 50.850 577.050 51.750 ;
        RECT 580.950 49.950 583.050 52.050 ;
        RECT 584.250 50.850 586.050 51.750 ;
        RECT 541.950 37.950 544.050 40.050 ;
        RECT 551.400 37.050 552.450 49.950 ;
        RECT 556.950 46.950 559.050 49.050 ;
        RECT 581.400 46.050 582.450 49.950 ;
        RECT 580.950 43.950 583.050 46.050 ;
        RECT 550.950 34.950 553.050 37.050 ;
        RECT 571.950 31.950 574.050 34.050 ;
        RECT 572.400 28.050 573.450 31.950 ;
        RECT 541.950 25.950 544.050 28.050 ;
        RECT 571.950 25.950 574.050 28.050 ;
        RECT 542.400 25.050 543.450 25.950 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 545.250 23.250 546.750 24.150 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 569.250 23.250 571.050 24.150 ;
        RECT 571.950 23.850 574.050 24.750 ;
        RECT 574.950 23.250 577.050 24.150 ;
        RECT 493.950 19.950 496.050 22.050 ;
        RECT 496.950 20.850 498.750 21.750 ;
        RECT 499.950 19.950 502.050 22.050 ;
        RECT 503.250 20.850 504.750 21.750 ;
        RECT 505.950 19.950 508.050 22.050 ;
        RECT 517.950 20.850 519.750 21.750 ;
        RECT 520.950 19.950 523.050 22.050 ;
        RECT 524.250 20.850 525.750 21.750 ;
        RECT 526.950 19.950 529.050 22.050 ;
        RECT 541.950 20.850 543.750 21.750 ;
        RECT 544.950 19.950 547.050 22.050 ;
        RECT 548.250 20.850 549.750 21.750 ;
        RECT 550.950 19.950 553.050 22.050 ;
        RECT 505.950 17.850 508.050 18.750 ;
        RECT 521.400 16.050 522.450 19.950 ;
        RECT 554.400 19.050 555.450 22.950 ;
        RECT 581.400 22.050 582.450 43.950 ;
        RECT 587.400 40.050 588.450 53.400 ;
        RECT 589.950 53.250 592.050 54.150 ;
        RECT 589.950 49.950 592.050 52.050 ;
        RECT 589.950 43.950 592.050 46.050 ;
        RECT 583.950 37.950 586.050 40.050 ;
        RECT 586.950 37.950 589.050 40.050 ;
        RECT 584.400 25.050 585.450 37.950 ;
        RECT 586.950 25.950 589.050 28.050 ;
        RECT 590.400 25.050 591.450 43.950 ;
        RECT 602.400 27.450 603.450 55.950 ;
        RECT 604.950 53.850 606.750 54.750 ;
        RECT 607.950 52.950 610.050 55.050 ;
        RECT 611.250 53.850 613.050 54.750 ;
        RECT 608.400 52.050 609.450 52.950 ;
        RECT 607.950 49.950 610.050 52.050 ;
        RECT 608.400 37.050 609.450 49.950 ;
        RECT 607.950 34.950 610.050 37.050 ;
        RECT 614.400 34.050 615.450 61.950 ;
        RECT 623.400 54.450 624.450 67.950 ;
        RECT 626.400 61.050 627.450 88.950 ;
        RECT 629.400 85.050 630.450 91.950 ;
        RECT 634.950 89.850 637.050 90.750 ;
        RECT 628.950 82.950 631.050 85.050 ;
        RECT 638.400 82.050 639.450 97.950 ;
        RECT 637.950 79.950 640.050 82.050 ;
        RECT 637.950 64.950 640.050 67.050 ;
        RECT 625.950 58.950 628.050 61.050 ;
        RECT 625.950 56.250 628.050 57.150 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 632.400 55.050 633.450 55.950 ;
        RECT 625.950 54.450 628.050 55.050 ;
        RECT 623.400 53.400 628.050 54.450 ;
        RECT 625.950 52.950 628.050 53.400 ;
        RECT 629.250 53.250 630.750 54.150 ;
        RECT 631.950 52.950 634.050 55.050 ;
        RECT 635.250 53.250 637.050 54.150 ;
        RECT 628.950 49.950 631.050 52.050 ;
        RECT 632.250 50.850 633.750 51.750 ;
        RECT 634.950 51.450 637.050 52.050 ;
        RECT 638.400 51.450 639.450 64.950 ;
        RECT 641.400 52.050 642.450 124.950 ;
        RECT 634.950 50.400 639.450 51.450 ;
        RECT 634.950 49.950 637.050 50.400 ;
        RECT 640.950 49.950 643.050 52.050 ;
        RECT 616.950 46.950 619.050 49.050 ;
        RECT 617.400 40.050 618.450 46.950 ;
        RECT 629.400 40.050 630.450 49.950 ;
        RECT 644.400 46.050 645.450 160.950 ;
        RECT 647.400 124.050 648.450 163.950 ;
        RECT 653.400 145.050 654.450 205.950 ;
        RECT 662.400 199.050 663.450 214.950 ;
        RECT 661.950 196.950 664.050 199.050 ;
        RECT 658.950 194.250 661.050 195.150 ;
        RECT 661.950 194.850 664.050 195.750 ;
        RECT 658.950 190.950 661.050 193.050 ;
        RECT 658.950 173.400 661.050 175.500 ;
        RECT 655.950 166.950 658.050 169.050 ;
        RECT 656.400 163.050 657.450 166.950 ;
        RECT 655.950 160.950 658.050 163.050 ;
        RECT 659.400 156.600 660.600 173.400 ;
        RECT 664.950 169.950 667.050 172.050 ;
        RECT 665.400 169.050 666.450 169.950 ;
        RECT 664.950 166.950 667.050 169.050 ;
        RECT 664.950 164.850 667.050 165.750 ;
        RECT 658.950 154.500 661.050 156.600 ;
        RECT 652.950 142.950 655.050 145.050 ;
        RECT 661.950 139.950 664.050 142.050 ;
        RECT 649.950 128.250 652.050 129.150 ;
        RECT 655.950 127.950 658.050 130.050 ;
        RECT 656.400 127.050 657.450 127.950 ;
        RECT 649.950 124.950 652.050 127.050 ;
        RECT 653.250 125.250 654.750 126.150 ;
        RECT 655.950 124.950 658.050 127.050 ;
        RECT 659.250 125.250 661.050 126.150 ;
        RECT 646.950 121.950 649.050 124.050 ;
        RECT 652.950 121.950 655.050 124.050 ;
        RECT 656.250 122.850 657.750 123.750 ;
        RECT 658.950 121.950 661.050 124.050 ;
        RECT 659.400 121.050 660.450 121.950 ;
        RECT 658.950 118.950 661.050 121.050 ;
        RECT 655.950 103.950 658.050 106.050 ;
        RECT 649.950 97.950 652.050 100.050 ;
        RECT 650.400 97.050 651.450 97.950 ;
        RECT 656.400 97.050 657.450 103.950 ;
        RECT 662.400 97.050 663.450 139.950 ;
        RECT 668.400 133.050 669.450 241.950 ;
        RECT 677.400 240.450 678.450 268.950 ;
        RECT 680.400 244.050 681.450 343.950 ;
        RECT 682.950 340.950 685.050 343.050 ;
        RECT 694.950 341.250 697.050 342.150 ;
        RECT 700.950 341.250 703.050 342.150 ;
        RECT 682.950 338.850 685.050 339.750 ;
        RECT 700.950 339.450 703.050 340.050 ;
        RECT 704.400 339.450 705.450 400.950 ;
        RECT 712.950 389.400 715.050 391.500 ;
        RECT 706.950 385.950 709.050 388.050 ;
        RECT 707.400 385.050 708.450 385.950 ;
        RECT 706.950 382.950 709.050 385.050 ;
        RECT 706.950 380.850 709.050 381.750 ;
        RECT 713.400 372.600 714.600 389.400 ;
        RECT 724.950 385.950 727.050 388.050 ;
        RECT 712.950 370.500 715.050 372.600 ;
        RECT 721.950 343.950 724.050 346.050 ;
        RECT 712.950 341.250 715.050 342.150 ;
        RECT 718.950 341.250 721.050 342.150 ;
        RECT 685.950 338.250 688.050 339.150 ;
        RECT 700.950 338.400 705.450 339.450 ;
        RECT 700.950 337.950 703.050 338.400 ;
        RECT 712.950 337.950 715.050 340.050 ;
        RECT 718.950 339.450 721.050 340.050 ;
        RECT 722.400 339.450 723.450 343.950 ;
        RECT 716.250 338.250 717.750 339.150 ;
        RECT 718.950 338.400 723.450 339.450 ;
        RECT 718.950 337.950 721.050 338.400 ;
        RECT 685.950 334.950 688.050 337.050 ;
        RECT 686.400 325.050 687.450 334.950 ;
        RECT 685.950 322.950 688.050 325.050 ;
        RECT 694.950 316.950 697.050 319.050 ;
        RECT 695.400 316.050 696.450 316.950 ;
        RECT 685.950 313.950 688.050 316.050 ;
        RECT 694.950 313.950 697.050 316.050 ;
        RECT 682.950 311.250 685.050 312.150 ;
        RECT 685.950 311.850 688.050 312.750 ;
        RECT 688.950 311.250 690.750 312.150 ;
        RECT 691.950 310.950 694.050 313.050 ;
        RECT 695.400 310.050 696.450 313.950 ;
        RECT 682.950 307.950 685.050 310.050 ;
        RECT 688.950 307.950 691.050 310.050 ;
        RECT 692.250 308.850 694.050 309.750 ;
        RECT 694.950 307.950 697.050 310.050 ;
        RECT 688.950 278.400 691.050 280.500 ;
        RECT 685.950 271.950 688.050 274.050 ;
        RECT 679.950 241.950 682.050 244.050 ;
        RECT 677.400 239.400 681.450 240.450 ;
        RECT 680.400 238.050 681.450 239.400 ;
        RECT 676.950 236.250 678.750 237.150 ;
        RECT 679.950 235.950 682.050 238.050 ;
        RECT 683.250 236.250 685.050 237.150 ;
        RECT 676.950 232.950 679.050 235.050 ;
        RECT 680.250 233.850 681.750 234.750 ;
        RECT 676.950 202.950 679.050 205.050 ;
        RECT 677.400 199.050 678.450 202.950 ;
        RECT 682.950 200.250 685.050 201.150 ;
        RECT 670.950 196.950 673.050 199.050 ;
        RECT 673.950 197.250 675.750 198.150 ;
        RECT 676.950 196.950 679.050 199.050 ;
        RECT 680.250 197.250 681.750 198.150 ;
        RECT 682.950 196.950 685.050 199.050 ;
        RECT 671.400 195.450 672.450 196.950 ;
        RECT 673.950 195.450 676.050 196.050 ;
        RECT 671.400 194.400 676.050 195.450 ;
        RECT 677.250 194.850 678.750 195.750 ;
        RECT 673.950 193.950 676.050 194.400 ;
        RECT 679.950 193.950 682.050 196.050 ;
        RECT 680.400 181.050 681.450 193.950 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 670.950 175.950 673.050 178.050 ;
        RECT 671.400 169.050 672.450 175.950 ;
        RECT 679.950 173.400 682.050 175.500 ;
        RECT 670.950 166.950 673.050 169.050 ;
        RECT 670.950 164.850 673.050 165.750 ;
        RECT 680.250 161.400 681.450 173.400 ;
        RECT 682.950 170.250 685.050 171.150 ;
        RECT 682.950 166.950 685.050 169.050 ;
        RECT 682.950 163.950 685.050 166.050 ;
        RECT 679.950 159.300 682.050 161.400 ;
        RECT 680.250 155.700 681.450 159.300 ;
        RECT 679.950 153.600 682.050 155.700 ;
        RECT 670.950 148.950 673.050 151.050 ;
        RECT 667.950 130.950 670.050 133.050 ;
        RECT 668.400 130.050 669.450 130.950 ;
        RECT 667.950 127.950 670.050 130.050 ;
        RECT 667.950 125.250 670.050 126.150 ;
        RECT 667.950 121.950 670.050 124.050 ;
        RECT 668.400 109.050 669.450 121.950 ;
        RECT 667.950 106.950 670.050 109.050 ;
        RECT 671.400 108.450 672.450 148.950 ;
        RECT 673.950 127.950 676.050 130.050 ;
        RECT 673.950 125.850 676.050 126.750 ;
        RECT 676.950 125.250 679.050 126.150 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 683.400 117.450 684.450 163.950 ;
        RECT 686.400 121.050 687.450 271.950 ;
        RECT 689.400 261.600 690.600 278.400 ;
        RECT 701.400 274.050 702.450 337.950 ;
        RECT 713.400 337.050 714.450 337.950 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 713.400 319.050 714.450 334.950 ;
        RECT 716.400 334.050 717.450 334.950 ;
        RECT 715.950 331.950 718.050 334.050 ;
        RECT 712.950 316.950 715.050 319.050 ;
        RECT 706.950 313.950 709.050 316.050 ;
        RECT 703.950 310.950 706.050 313.050 ;
        RECT 706.950 311.850 709.050 312.750 ;
        RECT 721.950 312.450 724.050 313.050 ;
        RECT 709.950 311.250 712.050 312.150 ;
        RECT 719.400 311.400 724.050 312.450 ;
        RECT 700.950 271.950 703.050 274.050 ;
        RECT 694.950 269.250 697.050 270.150 ;
        RECT 700.950 269.250 703.050 270.150 ;
        RECT 694.950 265.950 697.050 268.050 ;
        RECT 700.950 265.950 703.050 268.050 ;
        RECT 701.400 262.050 702.450 265.950 ;
        RECT 688.950 259.500 691.050 261.600 ;
        RECT 700.950 259.950 703.050 262.050 ;
        RECT 704.400 256.050 705.450 310.950 ;
        RECT 719.400 310.050 720.450 311.400 ;
        RECT 721.950 310.950 724.050 311.400 ;
        RECT 709.950 307.950 712.050 310.050 ;
        RECT 718.950 307.950 721.050 310.050 ;
        RECT 721.950 308.850 724.050 309.750 ;
        RECT 709.950 279.300 712.050 281.400 ;
        RECT 710.250 275.700 711.450 279.300 ;
        RECT 709.950 273.600 712.050 275.700 ;
        RECT 710.250 261.600 711.450 273.600 ;
        RECT 712.950 265.950 715.050 268.050 ;
        RECT 712.950 263.850 715.050 264.750 ;
        RECT 709.950 259.500 712.050 261.600 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 688.950 241.950 691.050 244.050 ;
        RECT 689.400 154.050 690.450 241.950 ;
        RECT 704.400 238.050 705.450 253.950 ;
        RECT 712.950 247.950 715.050 250.050 ;
        RECT 713.400 241.050 714.450 247.950 ;
        RECT 725.400 241.050 726.450 385.950 ;
        RECT 728.400 343.050 729.450 448.950 ;
        RECT 731.400 388.050 732.450 454.950 ;
        RECT 734.400 451.050 735.450 547.950 ;
        RECT 740.400 457.050 741.450 550.950 ;
        RECT 742.950 529.950 745.050 532.050 ;
        RECT 743.400 486.450 744.450 529.950 ;
        RECT 749.400 526.050 750.450 551.400 ;
        RECT 751.950 550.950 754.050 551.400 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 745.950 524.250 747.750 525.150 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 752.250 524.250 754.050 525.150 ;
        RECT 755.400 523.050 756.450 526.950 ;
        RECT 745.950 520.950 748.050 523.050 ;
        RECT 749.250 521.850 750.750 522.750 ;
        RECT 751.950 520.950 754.050 523.050 ;
        RECT 754.950 520.950 757.050 523.050 ;
        RECT 746.400 520.050 747.450 520.950 ;
        RECT 745.950 517.950 748.050 520.050 ;
        RECT 751.950 493.950 754.050 496.050 ;
        RECT 745.950 488.250 748.050 489.150 ;
        RECT 752.400 487.050 753.450 493.950 ;
        RECT 745.950 486.450 748.050 487.050 ;
        RECT 743.400 485.400 748.050 486.450 ;
        RECT 745.950 484.950 748.050 485.400 ;
        RECT 749.250 485.250 750.750 486.150 ;
        RECT 751.950 484.950 754.050 487.050 ;
        RECT 755.250 485.250 757.050 486.150 ;
        RECT 748.950 481.950 751.050 484.050 ;
        RECT 752.250 482.850 753.750 483.750 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 755.400 481.050 756.450 481.950 ;
        RECT 754.950 478.950 757.050 481.050 ;
        RECT 758.400 477.450 759.450 595.950 ;
        RECT 761.400 532.050 762.450 595.950 ;
        RECT 775.950 592.950 778.050 595.050 ;
        RECT 779.250 593.850 780.750 594.750 ;
        RECT 781.950 592.950 784.050 595.050 ;
        RECT 776.400 567.450 777.450 592.950 ;
        RECT 782.400 580.050 783.450 592.950 ;
        RECT 781.950 577.950 784.050 580.050 ;
        RECT 781.950 571.950 784.050 574.050 ;
        RECT 776.400 566.400 780.450 567.450 ;
        RECT 779.400 565.050 780.450 566.400 ;
        RECT 778.950 562.950 781.050 565.050 ;
        RECT 775.950 560.250 778.050 561.150 ;
        RECT 778.950 559.950 781.050 562.050 ;
        RECT 766.950 557.250 768.750 558.150 ;
        RECT 769.950 556.950 772.050 559.050 ;
        RECT 775.950 558.450 778.050 559.050 ;
        RECT 779.400 558.450 780.450 559.950 ;
        RECT 773.250 557.250 774.750 558.150 ;
        RECT 775.950 557.400 780.450 558.450 ;
        RECT 775.950 556.950 778.050 557.400 ;
        RECT 766.950 555.450 769.050 556.050 ;
        RECT 764.400 554.400 769.050 555.450 ;
        RECT 770.250 554.850 771.750 555.750 ;
        RECT 772.950 555.450 775.050 556.050 ;
        RECT 775.950 555.450 778.050 556.050 ;
        RECT 764.400 550.050 765.450 554.400 ;
        RECT 766.950 553.950 769.050 554.400 ;
        RECT 772.950 554.400 778.050 555.450 ;
        RECT 772.950 553.950 775.050 554.400 ;
        RECT 775.950 553.950 778.050 554.400 ;
        RECT 775.950 550.950 778.050 553.050 ;
        RECT 763.950 547.950 766.050 550.050 ;
        RECT 764.400 532.050 765.450 547.950 ;
        RECT 760.950 529.950 763.050 532.050 ;
        RECT 763.950 529.950 766.050 532.050 ;
        RECT 769.950 529.950 772.050 532.050 ;
        RECT 760.950 526.950 763.050 529.050 ;
        RECT 764.250 527.850 765.750 528.750 ;
        RECT 766.950 526.950 769.050 529.050 ;
        RECT 760.950 524.850 763.050 525.750 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 766.950 524.850 769.050 525.750 ;
        RECT 764.400 520.050 765.450 523.950 ;
        RECT 763.950 517.950 766.050 520.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 760.950 487.950 763.050 490.050 ;
        RECT 761.400 483.450 762.450 487.950 ;
        RECT 767.400 487.050 768.450 490.950 ;
        RECT 770.400 490.050 771.450 529.950 ;
        RECT 769.950 487.950 772.050 490.050 ;
        RECT 772.950 488.250 775.050 489.150 ;
        RECT 763.950 485.250 765.750 486.150 ;
        RECT 766.950 484.950 769.050 487.050 ;
        RECT 770.250 485.250 771.750 486.150 ;
        RECT 772.950 484.950 775.050 487.050 ;
        RECT 773.400 484.050 774.450 484.950 ;
        RECT 763.950 483.450 766.050 484.050 ;
        RECT 761.400 482.400 766.050 483.450 ;
        RECT 767.250 482.850 768.750 483.750 ;
        RECT 763.950 481.950 766.050 482.400 ;
        RECT 769.950 481.950 772.050 484.050 ;
        RECT 772.950 481.950 775.050 484.050 ;
        RECT 770.400 481.050 771.450 481.950 ;
        RECT 769.950 478.950 772.050 481.050 ;
        RECT 755.400 476.400 759.450 477.450 ;
        RECT 745.950 466.950 748.050 469.050 ;
        RECT 746.400 462.450 747.450 466.950 ;
        RECT 743.400 461.400 747.450 462.450 ;
        RECT 743.400 460.050 744.450 461.400 ;
        RECT 742.950 457.950 745.050 460.050 ;
        RECT 748.950 457.950 751.050 460.050 ;
        RECT 739.950 454.950 742.050 457.050 ;
        RECT 743.250 455.850 744.750 456.750 ;
        RECT 745.950 454.950 748.050 457.050 ;
        RECT 739.950 452.850 742.050 453.750 ;
        RECT 745.950 452.850 748.050 453.750 ;
        RECT 733.950 448.950 736.050 451.050 ;
        RECT 733.950 427.950 736.050 430.050 ;
        RECT 734.400 412.050 735.450 427.950 ;
        RECT 736.950 423.300 739.050 425.400 ;
        RECT 737.550 419.700 738.750 423.300 ;
        RECT 736.950 417.600 739.050 419.700 ;
        RECT 733.950 409.950 736.050 412.050 ;
        RECT 733.950 407.850 736.050 408.750 ;
        RECT 737.550 405.600 738.750 417.600 ;
        RECT 745.950 413.250 748.050 414.150 ;
        RECT 745.950 409.950 748.050 412.050 ;
        RECT 736.950 403.500 739.050 405.600 ;
        RECT 746.400 397.050 747.450 409.950 ;
        RECT 745.950 394.950 748.050 397.050 ;
        RECT 745.950 389.400 748.050 391.500 ;
        RECT 730.950 385.950 733.050 388.050 ;
        RECT 736.950 385.950 739.050 388.050 ;
        RECT 739.950 385.950 742.050 388.050 ;
        RECT 742.950 386.250 745.050 387.150 ;
        RECT 737.400 385.050 738.450 385.950 ;
        RECT 730.950 384.450 733.050 385.050 ;
        RECT 730.950 383.400 735.450 384.450 ;
        RECT 730.950 382.950 733.050 383.400 ;
        RECT 730.950 380.850 733.050 381.750 ;
        RECT 730.950 376.950 733.050 379.050 ;
        RECT 727.950 340.950 730.050 343.050 ;
        RECT 731.400 340.050 732.450 376.950 ;
        RECT 734.400 352.050 735.450 383.400 ;
        RECT 736.950 382.950 739.050 385.050 ;
        RECT 740.400 384.450 741.450 385.950 ;
        RECT 742.950 384.450 745.050 385.050 ;
        RECT 740.400 383.400 745.050 384.450 ;
        RECT 742.950 382.950 745.050 383.400 ;
        RECT 736.950 380.850 739.050 381.750 ;
        RECT 746.550 377.400 747.750 389.400 ;
        RECT 749.400 388.050 750.450 457.950 ;
        RECT 755.400 457.050 756.450 476.400 ;
        RECT 769.950 472.950 772.050 475.050 ;
        RECT 760.950 457.950 763.050 460.050 ;
        RECT 761.400 457.050 762.450 457.950 ;
        RECT 754.950 454.950 757.050 457.050 ;
        RECT 760.950 454.950 763.050 457.050 ;
        RECT 766.950 456.450 769.050 457.050 ;
        RECT 770.400 456.450 771.450 472.950 ;
        RECT 776.400 463.050 777.450 550.950 ;
        RECT 778.950 544.950 781.050 547.050 ;
        RECT 779.400 465.450 780.450 544.950 ;
        RECT 782.400 528.450 783.450 571.950 ;
        RECT 785.400 553.050 786.450 595.950 ;
        RECT 791.400 574.050 792.450 622.950 ;
        RECT 794.400 613.050 795.450 625.950 ;
        RECT 797.400 625.050 798.450 659.400 ;
        RECT 809.400 652.050 810.450 766.950 ;
        RECT 811.950 742.950 814.050 745.050 ;
        RECT 812.400 730.050 813.450 742.950 ;
        RECT 811.950 727.950 814.050 730.050 ;
        RECT 812.400 694.050 813.450 727.950 ;
        RECT 815.400 700.050 816.450 769.950 ;
        RECT 821.400 769.050 822.450 808.950 ;
        RECT 823.950 775.950 826.050 778.050 ;
        RECT 820.950 766.950 823.050 769.050 ;
        RECT 824.400 760.050 825.450 775.950 ;
        RECT 827.400 772.050 828.450 836.400 ;
        RECT 829.950 812.250 831.750 813.150 ;
        RECT 832.950 811.950 835.050 814.050 ;
        RECT 836.250 812.250 838.050 813.150 ;
        RECT 829.950 808.950 832.050 811.050 ;
        RECT 833.250 809.850 834.750 810.750 ;
        RECT 835.950 808.950 838.050 811.050 ;
        RECT 836.400 808.050 837.450 808.950 ;
        RECT 835.950 805.950 838.050 808.050 ;
        RECT 835.950 775.950 838.050 778.050 ;
        RECT 836.400 775.050 837.450 775.950 ;
        RECT 829.950 772.950 832.050 775.050 ;
        RECT 835.950 772.950 838.050 775.050 ;
        RECT 839.250 773.250 841.050 774.150 ;
        RECT 826.950 769.950 829.050 772.050 ;
        RECT 829.950 770.850 832.050 771.750 ;
        RECT 832.950 770.250 835.050 771.150 ;
        RECT 835.950 770.850 837.750 771.750 ;
        RECT 838.950 769.950 841.050 772.050 ;
        RECT 826.950 766.950 829.050 769.050 ;
        RECT 832.950 766.950 835.050 769.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 827.400 733.050 828.450 766.950 ;
        RECT 832.950 763.950 835.050 766.050 ;
        RECT 829.950 742.950 832.050 745.050 ;
        RECT 829.950 740.850 832.050 741.750 ;
        RECT 826.950 730.950 829.050 733.050 ;
        RECT 820.950 703.950 823.050 706.050 ;
        RECT 821.400 703.050 822.450 703.950 ;
        RECT 817.950 701.250 819.750 702.150 ;
        RECT 820.950 700.950 823.050 703.050 ;
        RECT 824.250 701.250 825.750 702.150 ;
        RECT 826.950 700.950 829.050 703.050 ;
        RECT 830.250 701.250 832.050 702.150 ;
        RECT 814.950 697.950 817.050 700.050 ;
        RECT 817.950 697.950 820.050 700.050 ;
        RECT 821.250 698.850 822.750 699.750 ;
        RECT 823.950 697.950 826.050 700.050 ;
        RECT 827.250 698.850 828.750 699.750 ;
        RECT 829.950 697.950 832.050 700.050 ;
        RECT 818.400 696.450 819.450 697.950 ;
        RECT 830.400 697.050 831.450 697.950 ;
        RECT 815.400 695.400 819.450 696.450 ;
        RECT 811.950 691.950 814.050 694.050 ;
        RECT 808.950 649.950 811.050 652.050 ;
        RECT 812.400 637.050 813.450 691.950 ;
        RECT 802.950 634.950 805.050 637.050 ;
        RECT 811.950 634.950 814.050 637.050 ;
        RECT 799.950 631.950 802.050 634.050 ;
        RECT 796.950 622.950 799.050 625.050 ;
        RECT 800.400 619.050 801.450 631.950 ;
        RECT 799.950 616.950 802.050 619.050 ;
        RECT 793.950 610.950 796.050 613.050 ;
        RECT 793.950 596.250 795.750 597.150 ;
        RECT 796.950 595.950 799.050 598.050 ;
        RECT 800.250 596.250 802.050 597.150 ;
        RECT 793.950 592.950 796.050 595.050 ;
        RECT 797.250 593.850 798.750 594.750 ;
        RECT 799.950 592.950 802.050 595.050 ;
        RECT 794.400 577.050 795.450 592.950 ;
        RECT 793.950 574.950 796.050 577.050 ;
        RECT 790.950 571.950 793.050 574.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 790.950 562.950 793.050 565.050 ;
        RECT 791.400 559.050 792.450 562.950 ;
        RECT 790.950 556.950 793.050 559.050 ;
        RECT 787.950 554.250 790.050 555.150 ;
        RECT 790.950 554.850 793.050 555.750 ;
        RECT 784.950 550.950 787.050 553.050 ;
        RECT 787.950 550.950 790.050 553.050 ;
        RECT 788.400 550.050 789.450 550.950 ;
        RECT 787.950 547.950 790.050 550.050 ;
        RECT 784.950 528.450 787.050 529.050 ;
        RECT 782.400 527.400 787.050 528.450 ;
        RECT 782.400 508.050 783.450 527.400 ;
        RECT 784.950 526.950 787.050 527.400 ;
        RECT 788.250 527.250 790.050 528.150 ;
        RECT 784.950 524.850 786.750 525.750 ;
        RECT 787.950 523.950 790.050 526.050 ;
        RECT 788.400 508.050 789.450 523.950 ;
        RECT 794.400 508.050 795.450 568.950 ;
        RECT 796.950 562.950 799.050 565.050 ;
        RECT 797.400 520.050 798.450 562.950 ;
        RECT 803.400 532.050 804.450 634.950 ;
        RECT 805.950 631.950 808.050 634.050 ;
        RECT 809.250 632.250 810.750 633.150 ;
        RECT 811.950 631.950 814.050 634.050 ;
        RECT 805.950 629.850 807.750 630.750 ;
        RECT 808.950 628.950 811.050 631.050 ;
        RECT 812.250 629.850 814.050 630.750 ;
        RECT 815.400 613.050 816.450 695.400 ;
        RECT 829.950 694.950 832.050 697.050 ;
        RECT 817.950 691.950 820.050 694.050 ;
        RECT 829.950 691.950 832.050 694.050 ;
        RECT 818.400 673.050 819.450 691.950 ;
        RECT 817.950 670.950 820.050 673.050 ;
        RECT 823.950 670.950 826.050 673.050 ;
        RECT 817.950 668.850 820.050 669.750 ;
        RECT 823.950 668.850 826.050 669.750 ;
        RECT 830.400 660.450 831.450 691.950 ;
        RECT 833.400 663.450 834.450 763.950 ;
        RECT 839.400 763.050 840.450 769.950 ;
        RECT 842.400 766.050 843.450 838.950 ;
        RECT 845.400 826.050 846.450 841.950 ;
        RECT 844.950 823.950 847.050 826.050 ;
        RECT 845.400 817.050 846.450 823.950 ;
        RECT 844.950 814.950 847.050 817.050 ;
        RECT 841.950 763.950 844.050 766.050 ;
        RECT 838.950 760.950 841.050 763.050 ;
        RECT 845.400 757.050 846.450 814.950 ;
        RECT 844.950 754.950 847.050 757.050 ;
        RECT 835.950 742.950 838.050 745.050 ;
        RECT 844.950 742.950 847.050 745.050 ;
        RECT 845.400 742.050 846.450 742.950 ;
        RECT 835.950 740.850 838.050 741.750 ;
        RECT 844.950 739.950 847.050 742.050 ;
        RECT 841.950 711.300 844.050 713.400 ;
        RECT 842.550 707.700 843.750 711.300 ;
        RECT 835.950 703.950 838.050 706.050 ;
        RECT 841.950 705.600 844.050 707.700 ;
        RECT 836.400 699.450 837.450 703.950 ;
        RECT 838.950 699.450 841.050 700.050 ;
        RECT 836.400 698.400 841.050 699.450 ;
        RECT 836.400 666.450 837.450 698.400 ;
        RECT 838.950 697.950 841.050 698.400 ;
        RECT 838.950 695.850 841.050 696.750 ;
        RECT 842.550 693.600 843.750 705.600 ;
        RECT 845.400 694.050 846.450 739.950 ;
        RECT 848.400 709.050 849.450 848.400 ;
        RECT 850.950 841.950 853.050 844.050 ;
        RECT 850.950 839.850 853.050 840.750 ;
        RECT 854.550 837.600 855.750 849.600 ;
        RECT 857.400 841.050 858.450 889.950 ;
        RECT 863.400 889.050 864.450 892.950 ;
        RECT 862.950 886.950 865.050 889.050 ;
        RECT 859.950 883.950 862.050 886.050 ;
        RECT 862.950 884.850 865.050 885.750 ;
        RECT 868.950 884.850 871.050 885.750 ;
        RECT 856.950 838.950 859.050 841.050 ;
        RECT 853.950 835.500 856.050 837.600 ;
        RECT 853.950 826.950 856.050 829.050 ;
        RECT 850.950 817.950 853.050 820.050 ;
        RECT 851.400 817.050 852.450 817.950 ;
        RECT 850.950 814.950 853.050 817.050 ;
        RECT 850.950 812.850 853.050 813.750 ;
        RECT 854.400 775.050 855.450 826.950 ;
        RECT 856.950 812.850 859.050 813.750 ;
        RECT 853.950 774.450 856.050 775.050 ;
        RECT 853.950 773.400 858.450 774.450 ;
        RECT 853.950 772.950 856.050 773.400 ;
        RECT 853.950 770.850 856.050 771.750 ;
        RECT 850.950 743.250 853.050 744.150 ;
        RECT 850.950 739.950 853.050 742.050 ;
        RECT 847.950 706.950 850.050 709.050 ;
        RECT 851.400 705.450 852.450 739.950 ;
        RECT 857.400 705.450 858.450 773.400 ;
        RECT 848.400 704.400 852.450 705.450 ;
        RECT 854.400 704.400 858.450 705.450 ;
        RECT 848.400 699.450 849.450 704.400 ;
        RECT 850.950 701.250 853.050 702.150 ;
        RECT 850.950 699.450 853.050 700.050 ;
        RECT 848.400 698.400 853.050 699.450 ;
        RECT 841.950 691.500 844.050 693.600 ;
        RECT 844.950 691.950 847.050 694.050 ;
        RECT 848.400 691.050 849.450 698.400 ;
        RECT 850.950 697.950 853.050 698.400 ;
        RECT 847.950 688.950 850.050 691.050 ;
        RECT 838.950 668.250 840.750 669.150 ;
        RECT 841.950 667.950 844.050 670.050 ;
        RECT 845.250 668.250 847.050 669.150 ;
        RECT 838.950 666.450 841.050 667.050 ;
        RECT 836.400 665.400 841.050 666.450 ;
        RECT 842.250 665.850 843.750 666.750 ;
        RECT 838.950 664.950 841.050 665.400 ;
        RECT 844.950 664.950 847.050 667.050 ;
        RECT 833.400 662.400 837.450 663.450 ;
        RECT 830.400 659.400 834.450 660.450 ;
        RECT 829.950 634.950 832.050 637.050 ;
        RECT 826.950 631.950 829.050 634.050 ;
        RECT 823.950 629.250 826.050 630.150 ;
        RECT 823.950 627.450 826.050 628.050 ;
        RECT 827.400 627.450 828.450 631.950 ;
        RECT 830.400 631.050 831.450 634.950 ;
        RECT 829.950 628.950 832.050 631.050 ;
        RECT 820.950 626.250 822.750 627.150 ;
        RECT 823.950 626.400 828.450 627.450 ;
        RECT 829.950 626.850 832.050 627.750 ;
        RECT 823.950 625.950 826.050 626.400 ;
        RECT 820.950 622.950 823.050 625.050 ;
        RECT 821.400 619.050 822.450 622.950 ;
        RECT 820.950 616.950 823.050 619.050 ;
        RECT 820.950 613.950 823.050 616.050 ;
        RECT 814.950 610.950 817.050 613.050 ;
        RECT 808.950 605.400 811.050 607.500 ;
        RECT 805.950 602.250 808.050 603.150 ;
        RECT 805.950 598.950 808.050 601.050 ;
        RECT 806.400 595.050 807.450 598.950 ;
        RECT 805.950 592.950 808.050 595.050 ;
        RECT 809.550 593.400 810.750 605.400 ;
        RECT 817.950 604.950 820.050 607.050 ;
        RECT 818.400 601.050 819.450 604.950 ;
        RECT 817.950 598.950 820.050 601.050 ;
        RECT 817.950 596.850 820.050 597.750 ;
        RECT 808.950 591.300 811.050 593.400 ;
        RECT 809.550 587.700 810.750 591.300 ;
        RECT 808.950 585.600 811.050 587.700 ;
        RECT 814.950 577.950 817.050 580.050 ;
        RECT 808.950 563.250 811.050 564.150 ;
        RECT 815.400 562.050 816.450 577.950 ;
        RECT 805.950 560.250 807.750 561.150 ;
        RECT 808.950 559.950 811.050 562.050 ;
        RECT 812.250 560.250 813.750 561.150 ;
        RECT 814.950 559.950 817.050 562.050 ;
        RECT 805.950 556.950 808.050 559.050 ;
        RECT 809.400 556.050 810.450 559.950 ;
        RECT 811.950 556.950 814.050 559.050 ;
        RECT 815.250 557.850 817.050 558.750 ;
        RECT 808.950 553.950 811.050 556.050 ;
        RECT 812.400 553.050 813.450 556.950 ;
        RECT 811.950 550.950 814.050 553.050 ;
        RECT 817.950 538.950 820.050 541.050 ;
        RECT 802.950 529.950 805.050 532.050 ;
        RECT 814.950 529.950 817.050 532.050 ;
        RECT 808.950 526.950 811.050 529.050 ;
        RECT 811.950 526.950 814.050 529.050 ;
        RECT 799.950 524.250 801.750 525.150 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 806.250 524.250 808.050 525.150 ;
        RECT 803.250 521.850 804.750 522.750 ;
        RECT 805.950 522.450 808.050 523.050 ;
        RECT 809.400 522.450 810.450 526.950 ;
        RECT 805.950 521.400 810.450 522.450 ;
        RECT 805.950 520.950 808.050 521.400 ;
        RECT 796.950 517.950 799.050 520.050 ;
        RECT 802.950 517.950 805.050 520.050 ;
        RECT 799.950 508.950 802.050 511.050 ;
        RECT 781.950 505.950 784.050 508.050 ;
        RECT 787.950 505.950 790.050 508.050 ;
        RECT 793.950 505.950 796.050 508.050 ;
        RECT 796.950 496.950 799.050 499.050 ;
        RECT 781.950 493.950 784.050 496.050 ;
        RECT 787.950 493.950 790.050 496.050 ;
        RECT 782.400 469.050 783.450 493.950 ;
        RECT 788.400 487.050 789.450 493.950 ;
        RECT 793.950 488.250 796.050 489.150 ;
        RECT 784.950 485.250 786.750 486.150 ;
        RECT 787.950 484.950 790.050 487.050 ;
        RECT 791.250 485.250 792.750 486.150 ;
        RECT 793.950 484.950 796.050 487.050 ;
        RECT 784.950 481.950 787.050 484.050 ;
        RECT 788.250 482.850 789.750 483.750 ;
        RECT 790.950 481.950 793.050 484.050 ;
        RECT 785.400 480.450 786.450 481.950 ;
        RECT 785.400 479.400 789.450 480.450 ;
        RECT 785.400 478.050 786.450 479.400 ;
        RECT 784.950 475.950 787.050 478.050 ;
        RECT 781.950 466.950 784.050 469.050 ;
        RECT 779.400 464.400 783.450 465.450 ;
        RECT 775.950 460.950 778.050 463.050 ;
        RECT 766.950 455.400 771.450 456.450 ;
        RECT 766.950 454.950 769.050 455.400 ;
        RECT 751.950 413.250 754.050 414.150 ;
        RECT 751.950 409.950 754.050 412.050 ;
        RECT 755.400 408.450 756.450 454.950 ;
        RECT 760.950 452.850 763.050 453.750 ;
        RECT 766.950 452.850 769.050 453.750 ;
        RECT 760.950 439.950 763.050 442.050 ;
        RECT 757.950 422.400 760.050 424.500 ;
        RECT 752.400 407.400 756.450 408.450 ;
        RECT 748.950 385.950 751.050 388.050 ;
        RECT 745.950 375.300 748.050 377.400 ;
        RECT 746.550 371.700 747.750 375.300 ;
        RECT 745.950 369.600 748.050 371.700 ;
        RECT 733.950 349.950 736.050 352.050 ;
        RECT 742.950 347.250 745.050 348.150 ;
        RECT 736.950 343.950 739.050 346.050 ;
        RECT 740.250 344.250 741.750 345.150 ;
        RECT 742.950 343.950 745.050 346.050 ;
        RECT 746.250 344.250 748.050 345.150 ;
        RECT 748.950 343.950 751.050 346.050 ;
        RECT 736.950 341.850 738.750 342.750 ;
        RECT 739.950 340.950 742.050 343.050 ;
        RECT 730.950 337.950 733.050 340.050 ;
        RECT 730.950 313.950 733.050 316.050 ;
        RECT 733.950 313.950 736.050 316.050 ;
        RECT 731.400 313.050 732.450 313.950 ;
        RECT 730.950 310.950 733.050 313.050 ;
        RECT 727.950 308.250 730.050 309.150 ;
        RECT 730.950 308.850 733.050 309.750 ;
        RECT 727.950 304.950 730.050 307.050 ;
        RECT 730.950 274.950 733.050 277.050 ;
        RECT 731.400 271.050 732.450 274.950 ;
        RECT 734.400 274.050 735.450 313.950 ;
        RECT 733.950 271.950 736.050 274.050 ;
        RECT 736.950 272.250 739.050 273.150 ;
        RECT 727.950 269.250 729.750 270.150 ;
        RECT 730.950 268.950 733.050 271.050 ;
        RECT 734.250 269.250 735.750 270.150 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 727.950 265.950 730.050 268.050 ;
        RECT 731.250 266.850 732.750 267.750 ;
        RECT 733.950 265.950 736.050 268.050 ;
        RECT 734.400 265.050 735.450 265.950 ;
        RECT 733.950 262.950 736.050 265.050 ;
        RECT 733.950 243.450 736.050 244.050 ;
        RECT 731.400 242.400 736.050 243.450 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 716.250 239.250 717.750 240.150 ;
        RECT 718.950 238.950 721.050 241.050 ;
        RECT 724.950 238.950 727.050 241.050 ;
        RECT 694.950 236.250 696.750 237.150 ;
        RECT 697.950 235.950 700.050 238.050 ;
        RECT 701.250 236.250 703.050 237.150 ;
        RECT 703.950 235.950 706.050 238.050 ;
        RECT 712.950 236.850 714.750 237.750 ;
        RECT 715.950 235.950 718.050 238.050 ;
        RECT 719.250 236.850 720.750 237.750 ;
        RECT 721.950 237.450 724.050 238.050 ;
        RECT 721.950 236.400 726.450 237.450 ;
        RECT 721.950 235.950 724.050 236.400 ;
        RECT 698.250 233.850 699.750 234.750 ;
        RECT 700.950 232.950 703.050 235.050 ;
        RECT 718.950 232.950 721.050 235.050 ;
        RECT 721.950 233.850 724.050 234.750 ;
        RECT 701.400 229.050 702.450 232.950 ;
        RECT 700.950 226.950 703.050 229.050 ;
        RECT 701.400 205.050 702.450 226.950 ;
        RECT 700.950 202.950 703.050 205.050 ;
        RECT 701.400 202.050 702.450 202.950 ;
        RECT 698.250 200.250 699.750 201.150 ;
        RECT 700.950 199.950 703.050 202.050 ;
        RECT 694.950 197.850 696.750 198.750 ;
        RECT 697.950 196.950 700.050 199.050 ;
        RECT 701.250 197.850 703.050 198.750 ;
        RECT 703.950 196.950 706.050 199.050 ;
        RECT 715.950 196.950 718.050 199.050 ;
        RECT 694.950 190.950 697.050 193.050 ;
        RECT 695.400 169.050 696.450 190.950 ;
        RECT 704.400 187.050 705.450 196.950 ;
        RECT 712.950 194.250 715.050 195.150 ;
        RECT 715.950 194.850 718.050 195.750 ;
        RECT 712.950 190.950 715.050 193.050 ;
        RECT 703.950 184.950 706.050 187.050 ;
        RECT 706.950 169.950 709.050 172.050 ;
        RECT 707.400 169.050 708.450 169.950 ;
        RECT 694.950 166.950 697.050 169.050 ;
        RECT 700.950 166.950 703.050 169.050 ;
        RECT 704.250 167.250 705.750 168.150 ;
        RECT 706.950 166.950 709.050 169.050 ;
        RECT 710.250 167.250 711.750 168.150 ;
        RECT 712.950 166.950 715.050 169.050 ;
        RECT 700.950 164.850 702.750 165.750 ;
        RECT 703.950 163.950 706.050 166.050 ;
        RECT 707.250 164.850 708.750 165.750 ;
        RECT 709.950 163.950 712.050 166.050 ;
        RECT 713.250 164.850 715.050 165.750 ;
        RECT 704.400 154.050 705.450 163.950 ;
        RECT 688.950 151.950 691.050 154.050 ;
        RECT 703.950 151.950 706.050 154.050 ;
        RECT 710.400 151.050 711.450 163.950 ;
        RECT 709.950 148.950 712.050 151.050 ;
        RECT 688.950 142.950 691.050 145.050 ;
        RECT 685.950 118.950 688.050 121.050 ;
        RECT 683.400 116.400 687.450 117.450 ;
        RECT 671.400 107.400 675.450 108.450 ;
        RECT 670.950 101.400 673.050 103.500 ;
        RECT 664.950 97.950 667.050 100.050 ;
        RECT 649.950 94.950 652.050 97.050 ;
        RECT 653.250 95.250 654.750 96.150 ;
        RECT 655.950 94.950 658.050 97.050 ;
        RECT 659.250 95.250 660.750 96.150 ;
        RECT 661.950 94.950 664.050 97.050 ;
        RECT 649.950 92.850 651.750 93.750 ;
        RECT 652.950 91.950 655.050 94.050 ;
        RECT 656.250 92.850 657.750 93.750 ;
        RECT 658.950 91.950 661.050 94.050 ;
        RECT 662.250 92.850 664.050 93.750 ;
        RECT 653.400 91.050 654.450 91.950 ;
        RECT 652.950 88.950 655.050 91.050 ;
        RECT 646.950 85.950 649.050 88.050 ;
        RECT 647.400 58.050 648.450 85.950 ;
        RECT 665.400 64.050 666.450 97.950 ;
        RECT 667.950 94.950 670.050 97.050 ;
        RECT 652.950 61.950 655.050 64.050 ;
        RECT 658.950 61.950 661.050 64.050 ;
        RECT 664.950 61.950 667.050 64.050 ;
        RECT 653.400 58.050 654.450 61.950 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 650.250 56.250 651.750 57.150 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 646.950 53.850 648.750 54.750 ;
        RECT 649.950 52.950 652.050 55.050 ;
        RECT 653.250 53.850 655.050 54.750 ;
        RECT 646.950 49.950 649.050 52.050 ;
        RECT 643.950 43.950 646.050 46.050 ;
        RECT 616.950 37.950 619.050 40.050 ;
        RECT 628.950 37.950 631.050 40.050 ;
        RECT 613.950 31.950 616.050 34.050 ;
        RECT 604.950 27.450 607.050 28.050 ;
        RECT 602.400 26.400 607.050 27.450 ;
        RECT 604.950 25.950 607.050 26.400 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 587.250 23.850 588.750 24.750 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 604.950 23.850 607.050 24.750 ;
        RECT 607.950 23.250 610.050 24.150 ;
        RECT 565.950 20.850 567.750 21.750 ;
        RECT 568.950 19.950 571.050 22.050 ;
        RECT 574.950 19.950 577.050 22.050 ;
        RECT 580.950 19.950 583.050 22.050 ;
        RECT 583.950 20.850 586.050 21.750 ;
        RECT 589.950 20.850 592.050 21.750 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 617.400 21.450 618.450 37.950 ;
        RECT 622.950 31.950 625.050 34.050 ;
        RECT 623.400 28.050 624.450 31.950 ;
        RECT 622.950 25.950 625.050 28.050 ;
        RECT 619.950 23.250 622.050 24.150 ;
        RECT 622.950 23.850 625.050 24.750 ;
        RECT 625.950 23.250 627.750 24.150 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 619.950 21.450 622.050 22.050 ;
        RECT 617.400 20.400 622.050 21.450 ;
        RECT 619.950 19.950 622.050 20.400 ;
        RECT 625.950 19.950 628.050 22.050 ;
        RECT 629.250 20.850 631.050 21.750 ;
        RECT 575.400 19.050 576.450 19.950 ;
        RECT 608.400 19.050 609.450 19.950 ;
        RECT 526.950 17.850 529.050 18.750 ;
        RECT 550.950 17.850 553.050 18.750 ;
        RECT 553.950 16.950 556.050 19.050 ;
        RECT 574.950 16.950 577.050 19.050 ;
        RECT 607.950 16.950 610.050 19.050 ;
        RECT 641.400 18.450 642.450 22.950 ;
        RECT 647.400 22.050 648.450 49.950 ;
        RECT 650.400 49.050 651.450 52.950 ;
        RECT 649.950 46.950 652.050 49.050 ;
        RECT 652.950 25.950 655.050 28.050 ;
        RECT 643.950 20.250 645.750 21.150 ;
        RECT 646.950 19.950 649.050 22.050 ;
        RECT 650.250 20.250 652.050 21.150 ;
        RECT 643.950 18.450 646.050 19.050 ;
        RECT 641.400 17.400 646.050 18.450 ;
        RECT 647.250 17.850 648.750 18.750 ;
        RECT 649.950 18.450 652.050 19.050 ;
        RECT 653.400 18.450 654.450 25.950 ;
        RECT 659.400 19.050 660.450 61.950 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 665.400 55.050 666.450 55.950 ;
        RECT 668.400 55.050 669.450 94.950 ;
        RECT 671.400 84.600 672.600 101.400 ;
        RECT 674.400 94.050 675.450 107.400 ;
        RECT 676.950 103.950 679.050 106.050 ;
        RECT 682.950 103.950 685.050 106.050 ;
        RECT 677.400 97.050 678.450 103.950 ;
        RECT 683.400 97.050 684.450 103.950 ;
        RECT 676.950 94.950 679.050 97.050 ;
        RECT 682.950 94.950 685.050 97.050 ;
        RECT 673.950 91.950 676.050 94.050 ;
        RECT 676.950 92.850 679.050 93.750 ;
        RECT 682.950 92.850 685.050 93.750 ;
        RECT 670.950 82.500 673.050 84.600 ;
        RECT 670.950 61.950 673.050 64.050 ;
        RECT 671.400 55.050 672.450 61.950 ;
        RECT 664.950 52.950 667.050 55.050 ;
        RECT 667.950 52.950 670.050 55.050 ;
        RECT 670.950 52.950 673.050 55.050 ;
        RECT 674.250 53.250 676.050 54.150 ;
        RECT 676.950 52.950 679.050 55.050 ;
        RECT 664.950 50.850 667.050 51.750 ;
        RECT 667.950 50.250 670.050 51.150 ;
        RECT 670.950 50.850 672.750 51.750 ;
        RECT 673.950 49.950 676.050 52.050 ;
        RECT 667.950 46.950 670.050 49.050 ;
        RECT 664.950 43.950 667.050 46.050 ;
        RECT 665.400 28.050 666.450 43.950 ;
        RECT 677.400 31.050 678.450 52.950 ;
        RECT 686.400 46.050 687.450 116.400 ;
        RECT 689.400 94.050 690.450 142.950 ;
        RECT 694.950 131.250 697.050 132.150 ;
        RECT 719.400 130.050 720.450 232.950 ;
        RECT 725.400 232.050 726.450 236.400 ;
        RECT 731.400 232.050 732.450 242.400 ;
        RECT 733.950 241.950 736.050 242.400 ;
        RECT 733.950 239.850 736.050 240.750 ;
        RECT 736.950 239.250 739.050 240.150 ;
        RECT 736.950 235.950 739.050 238.050 ;
        RECT 740.400 235.050 741.450 340.950 ;
        RECT 743.400 331.050 744.450 343.950 ;
        RECT 745.950 340.950 748.050 343.050 ;
        RECT 742.950 328.950 745.050 331.050 ;
        RECT 745.950 322.950 748.050 325.050 ;
        RECT 742.950 313.950 745.050 316.050 ;
        RECT 746.400 313.050 747.450 322.950 ;
        RECT 742.950 311.850 744.750 312.750 ;
        RECT 745.950 310.950 748.050 313.050 ;
        RECT 745.950 308.850 748.050 309.750 ;
        RECT 749.400 274.050 750.450 343.950 ;
        RECT 752.400 319.050 753.450 407.400 ;
        RECT 758.400 405.600 759.600 422.400 ;
        RECT 757.950 403.500 760.050 405.600 ;
        RECT 761.400 397.050 762.450 439.950 ;
        RECT 754.950 394.950 757.050 397.050 ;
        RECT 757.950 394.950 760.050 397.050 ;
        RECT 760.950 394.950 763.050 397.050 ;
        RECT 755.400 388.050 756.450 394.950 ;
        RECT 754.950 385.950 757.050 388.050 ;
        RECT 755.400 385.050 756.450 385.950 ;
        RECT 754.950 382.950 757.050 385.050 ;
        RECT 754.950 380.850 757.050 381.750 ;
        RECT 754.950 346.950 757.050 349.050 ;
        RECT 751.950 316.950 754.050 319.050 ;
        RECT 751.950 311.250 754.050 312.150 ;
        RECT 755.400 310.050 756.450 346.950 ;
        RECT 758.400 346.050 759.450 394.950 ;
        RECT 766.950 389.400 769.050 391.500 ;
        RECT 760.950 382.950 763.050 385.050 ;
        RECT 760.950 380.850 763.050 381.750 ;
        RECT 767.400 372.600 768.600 389.400 ;
        RECT 770.400 382.050 771.450 455.400 ;
        RECT 772.950 413.250 775.050 414.150 ;
        RECT 772.950 409.950 775.050 412.050 ;
        RECT 769.950 379.950 772.050 382.050 ;
        RECT 766.950 370.500 769.050 372.600 ;
        RECT 763.950 346.950 766.050 349.050 ;
        RECT 764.400 346.050 765.450 346.950 ;
        RECT 757.950 343.950 760.050 346.050 ;
        RECT 761.250 344.250 762.750 345.150 ;
        RECT 763.950 343.950 766.050 346.050 ;
        RECT 757.950 341.850 759.750 342.750 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 764.250 341.850 766.050 342.750 ;
        RECT 761.400 340.050 762.450 340.950 ;
        RECT 760.950 337.950 763.050 340.050 ;
        RECT 770.400 337.050 771.450 379.950 ;
        RECT 776.400 352.050 777.450 460.950 ;
        RECT 782.400 457.050 783.450 464.400 ;
        RECT 788.400 457.050 789.450 479.400 ;
        RECT 781.950 456.450 784.050 457.050 ;
        RECT 781.950 455.400 786.450 456.450 ;
        RECT 781.950 454.950 784.050 455.400 ;
        RECT 781.950 452.850 784.050 453.750 ;
        RECT 778.950 413.250 781.050 414.150 ;
        RECT 785.400 412.050 786.450 455.400 ;
        RECT 787.950 454.950 790.050 457.050 ;
        RECT 787.950 452.850 790.050 453.750 ;
        RECT 797.400 417.450 798.450 496.950 ;
        RECT 800.400 457.050 801.450 508.950 ;
        RECT 803.400 475.050 804.450 517.950 ;
        RECT 806.400 511.050 807.450 520.950 ;
        RECT 805.950 508.950 808.050 511.050 ;
        RECT 805.950 494.400 808.050 496.500 ;
        RECT 806.400 477.600 807.600 494.400 ;
        RECT 812.400 489.450 813.450 526.950 ;
        RECT 809.400 488.400 813.450 489.450 ;
        RECT 805.950 475.500 808.050 477.600 ;
        RECT 802.950 472.950 805.050 475.050 ;
        RECT 805.950 466.950 808.050 469.050 ;
        RECT 802.950 460.950 805.050 463.050 ;
        RECT 803.400 460.050 804.450 460.950 ;
        RECT 802.950 457.950 805.050 460.050 ;
        RECT 806.400 457.050 807.450 466.950 ;
        RECT 799.950 454.950 802.050 457.050 ;
        RECT 803.250 455.850 804.750 456.750 ;
        RECT 805.950 454.950 808.050 457.050 ;
        RECT 799.950 452.850 802.050 453.750 ;
        RECT 805.950 452.850 808.050 453.750 ;
        RECT 797.400 416.400 801.450 417.450 ;
        RECT 790.950 413.250 793.050 414.150 ;
        RECT 796.950 413.250 799.050 414.150 ;
        RECT 778.950 409.950 781.050 412.050 ;
        RECT 784.950 409.950 787.050 412.050 ;
        RECT 790.950 409.950 793.050 412.050 ;
        RECT 796.950 409.950 799.050 412.050 ;
        RECT 779.400 391.050 780.450 409.950 ;
        RECT 797.400 409.050 798.450 409.950 ;
        RECT 796.950 406.950 799.050 409.050 ;
        RECT 778.950 388.950 781.050 391.050 ;
        RECT 781.950 389.400 784.050 391.500 ;
        RECT 778.950 386.250 781.050 387.150 ;
        RECT 778.950 382.950 781.050 385.050 ;
        RECT 775.950 349.950 778.050 352.050 ;
        RECT 779.400 346.050 780.450 382.950 ;
        RECT 782.550 377.400 783.750 389.400 ;
        RECT 787.950 385.950 790.050 388.050 ;
        RECT 788.400 384.450 789.450 385.950 ;
        RECT 790.950 384.450 793.050 385.050 ;
        RECT 788.400 383.400 793.050 384.450 ;
        RECT 781.950 375.300 784.050 377.400 ;
        RECT 782.550 371.700 783.750 375.300 ;
        RECT 781.950 369.600 784.050 371.700 ;
        RECT 775.950 344.250 778.050 345.150 ;
        RECT 778.950 343.950 781.050 346.050 ;
        RECT 772.950 340.950 775.050 343.050 ;
        RECT 775.950 340.950 778.050 343.050 ;
        RECT 779.250 341.250 780.750 342.150 ;
        RECT 781.950 340.950 784.050 343.050 ;
        RECT 785.250 341.250 787.050 342.150 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 760.950 310.950 763.050 313.050 ;
        RECT 751.950 307.950 754.050 310.050 ;
        RECT 754.950 307.950 757.050 310.050 ;
        RECT 748.950 271.950 751.050 274.050 ;
        RECT 748.950 270.450 751.050 271.050 ;
        RECT 752.400 270.450 753.450 307.950 ;
        RECT 755.400 271.050 756.450 307.950 ;
        RECT 748.950 269.400 753.450 270.450 ;
        RECT 748.950 268.950 751.050 269.400 ;
        RECT 754.950 268.950 757.050 271.050 ;
        RECT 758.250 269.250 760.050 270.150 ;
        RECT 748.950 266.850 751.050 267.750 ;
        RECT 751.950 266.250 754.050 267.150 ;
        RECT 754.950 266.850 756.750 267.750 ;
        RECT 757.950 265.950 760.050 268.050 ;
        RECT 751.950 262.950 754.050 265.050 ;
        RECT 761.400 264.450 762.450 310.950 ;
        RECT 758.400 263.400 762.450 264.450 ;
        RECT 754.950 247.950 757.050 250.050 ;
        RECT 751.950 243.450 754.050 244.050 ;
        RECT 749.400 242.400 754.050 243.450 ;
        RECT 745.950 238.950 748.050 241.050 ;
        RECT 739.950 232.950 742.050 235.050 ;
        RECT 724.950 229.950 727.050 232.050 ;
        RECT 730.950 229.950 733.050 232.050 ;
        RECT 736.950 205.950 739.050 208.050 ;
        RECT 742.950 205.950 745.050 208.050 ;
        RECT 737.400 202.050 738.450 205.950 ;
        RECT 730.950 201.450 733.050 202.050 ;
        RECT 728.400 200.400 733.050 201.450 ;
        RECT 728.400 193.050 729.450 200.400 ;
        RECT 730.950 199.950 733.050 200.400 ;
        RECT 734.250 200.250 735.750 201.150 ;
        RECT 736.950 199.950 739.050 202.050 ;
        RECT 730.950 197.850 732.750 198.750 ;
        RECT 733.950 196.950 736.050 199.050 ;
        RECT 737.250 197.850 739.050 198.750 ;
        RECT 743.400 196.050 744.450 205.950 ;
        RECT 742.950 193.950 745.050 196.050 ;
        RECT 727.950 190.950 730.050 193.050 ;
        RECT 739.950 175.950 742.050 178.050 ;
        RECT 736.950 173.400 739.050 175.500 ;
        RECT 727.950 171.450 730.050 172.050 ;
        RECT 727.950 170.400 732.450 171.450 ;
        RECT 727.950 169.950 730.050 170.400 ;
        RECT 721.950 166.950 724.050 169.050 ;
        RECT 724.950 167.250 727.050 168.150 ;
        RECT 727.950 167.850 730.050 168.750 ;
        RECT 731.400 168.450 732.450 170.400 ;
        RECT 733.950 170.250 736.050 171.150 ;
        RECT 733.950 168.450 736.050 169.050 ;
        RECT 731.400 167.400 736.050 168.450 ;
        RECT 733.950 166.950 736.050 167.400 ;
        RECT 722.400 165.450 723.450 166.950 ;
        RECT 724.950 165.450 727.050 166.050 ;
        RECT 722.400 164.400 727.050 165.450 ;
        RECT 724.950 163.950 727.050 164.400 ;
        RECT 725.400 163.050 726.450 163.950 ;
        RECT 724.950 160.950 727.050 163.050 ;
        RECT 737.550 161.400 738.750 173.400 ;
        RECT 740.400 169.050 741.450 175.950 ;
        RECT 746.400 171.450 747.450 238.950 ;
        RECT 749.400 238.050 750.450 242.400 ;
        RECT 751.950 241.950 754.050 242.400 ;
        RECT 755.400 241.050 756.450 247.950 ;
        RECT 751.950 239.850 753.750 240.750 ;
        RECT 754.950 238.950 757.050 241.050 ;
        RECT 748.950 235.950 751.050 238.050 ;
        RECT 754.950 236.850 757.050 237.750 ;
        RECT 758.400 237.450 759.450 263.400 ;
        RECT 760.950 239.250 763.050 240.150 ;
        RECT 760.950 237.450 763.050 238.050 ;
        RECT 758.400 236.400 763.050 237.450 ;
        RECT 760.950 235.950 763.050 236.400 ;
        RECT 764.400 202.050 765.450 334.950 ;
        RECT 769.950 322.950 772.050 325.050 ;
        RECT 770.400 316.050 771.450 322.950 ;
        RECT 773.400 322.050 774.450 340.950 ;
        RECT 776.400 340.050 777.450 340.950 ;
        RECT 775.950 337.950 778.050 340.050 ;
        RECT 778.950 337.950 781.050 340.050 ;
        RECT 782.250 338.850 783.750 339.750 ;
        RECT 784.950 337.950 787.050 340.050 ;
        RECT 785.400 328.050 786.450 337.950 ;
        RECT 788.400 328.050 789.450 383.400 ;
        RECT 790.950 382.950 793.050 383.400 ;
        RECT 796.950 384.450 799.050 385.050 ;
        RECT 800.400 384.450 801.450 416.400 ;
        RECT 809.400 393.450 810.450 488.400 ;
        RECT 811.950 485.250 814.050 486.150 ;
        RECT 811.950 481.950 814.050 484.050 ;
        RECT 812.400 481.050 813.450 481.950 ;
        RECT 811.950 478.950 814.050 481.050 ;
        RECT 811.950 454.950 814.050 457.050 ;
        RECT 812.400 418.050 813.450 454.950 ;
        RECT 811.950 415.950 814.050 418.050 ;
        RECT 811.950 413.250 814.050 414.150 ;
        RECT 811.950 409.950 814.050 412.050 ;
        RECT 815.400 411.450 816.450 529.950 ;
        RECT 818.400 489.450 819.450 538.950 ;
        RECT 821.400 529.050 822.450 613.950 ;
        RECT 829.950 605.400 832.050 607.500 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 823.950 596.850 826.050 597.750 ;
        RECT 830.400 588.600 831.600 605.400 ;
        RECT 829.950 586.500 832.050 588.600 ;
        RECT 833.400 565.050 834.450 659.400 ;
        RECT 832.950 562.950 835.050 565.050 ;
        RECT 832.950 559.950 835.050 562.050 ;
        RECT 833.400 559.050 834.450 559.950 ;
        RECT 832.950 556.950 835.050 559.050 ;
        RECT 829.950 554.250 832.050 555.150 ;
        RECT 832.950 554.850 835.050 555.750 ;
        RECT 829.950 550.950 832.050 553.050 ;
        RECT 823.950 529.950 826.050 532.050 ;
        RECT 824.400 529.050 825.450 529.950 ;
        RECT 820.950 526.950 823.050 529.050 ;
        RECT 823.950 526.950 826.050 529.050 ;
        RECT 827.250 527.250 828.750 528.150 ;
        RECT 829.950 526.950 832.050 529.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 824.250 524.850 825.750 525.750 ;
        RECT 826.950 523.950 829.050 526.050 ;
        RECT 830.250 524.850 832.050 525.750 ;
        RECT 820.950 521.850 823.050 522.750 ;
        RECT 823.950 505.950 826.050 508.050 ;
        RECT 818.400 488.400 822.450 489.450 ;
        RECT 817.950 485.250 820.050 486.150 ;
        RECT 817.950 483.450 820.050 484.050 ;
        RECT 821.400 483.450 822.450 488.400 ;
        RECT 817.950 482.400 822.450 483.450 ;
        RECT 817.950 481.950 820.050 482.400 ;
        RECT 824.400 481.050 825.450 505.950 ;
        RECT 826.950 495.300 829.050 497.400 ;
        RECT 827.250 491.700 828.450 495.300 ;
        RECT 826.950 489.600 829.050 491.700 ;
        RECT 823.950 478.950 826.050 481.050 ;
        RECT 827.250 477.600 828.450 489.600 ;
        RECT 829.950 484.950 832.050 487.050 ;
        RECT 830.400 484.050 831.450 484.950 ;
        RECT 836.400 484.050 837.450 662.400 ;
        RECT 850.950 634.950 853.050 637.050 ;
        RECT 851.400 634.050 852.450 634.950 ;
        RECT 844.950 633.450 847.050 634.050 ;
        RECT 842.400 632.400 847.050 633.450 ;
        RECT 842.400 631.050 843.450 632.400 ;
        RECT 844.950 631.950 847.050 632.400 ;
        RECT 848.250 632.250 849.750 633.150 ;
        RECT 850.950 631.950 853.050 634.050 ;
        RECT 841.950 628.950 844.050 631.050 ;
        RECT 844.950 629.850 846.750 630.750 ;
        RECT 847.950 628.950 850.050 631.050 ;
        RECT 851.250 629.850 853.050 630.750 ;
        RECT 848.400 625.050 849.450 628.950 ;
        RECT 850.950 625.950 853.050 628.050 ;
        RECT 847.950 622.950 850.050 625.050 ;
        RECT 851.400 616.050 852.450 625.950 ;
        RECT 850.950 613.950 853.050 616.050 ;
        RECT 854.400 604.050 855.450 704.400 ;
        RECT 856.950 701.250 859.050 702.150 ;
        RECT 856.950 697.950 859.050 700.050 ;
        RECT 857.400 688.050 858.450 697.950 ;
        RECT 856.950 685.950 859.050 688.050 ;
        RECT 860.400 672.450 861.450 883.950 ;
        RECT 865.950 880.950 868.050 883.050 ;
        RECT 862.950 845.250 865.050 846.150 ;
        RECT 862.950 841.950 865.050 844.050 ;
        RECT 863.400 829.050 864.450 841.950 ;
        RECT 862.950 826.950 865.050 829.050 ;
        RECT 862.950 710.400 865.050 712.500 ;
        RECT 863.400 693.600 864.600 710.400 ;
        RECT 866.400 700.050 867.450 880.950 ;
        RECT 874.950 854.400 877.050 856.500 ;
        RECT 868.950 845.250 871.050 846.150 ;
        RECT 868.950 841.950 871.050 844.050 ;
        RECT 869.400 835.050 870.450 841.950 ;
        RECT 875.400 837.600 876.600 854.400 ;
        RECT 874.950 835.500 877.050 837.600 ;
        RECT 868.950 832.950 871.050 835.050 ;
        RECT 871.950 815.250 873.750 816.150 ;
        RECT 874.950 814.950 877.050 817.050 ;
        RECT 871.950 811.950 874.050 814.050 ;
        RECT 875.250 812.850 877.050 813.750 ;
        RECT 872.400 768.450 873.450 811.950 ;
        RECT 874.950 770.850 877.050 771.750 ;
        RECT 872.400 767.400 876.450 768.450 ;
        RECT 871.950 743.250 874.050 744.150 ;
        RECT 871.950 706.950 874.050 709.050 ;
        RECT 865.950 697.950 868.050 700.050 ;
        RECT 872.400 697.050 873.450 706.950 ;
        RECT 871.950 694.950 874.050 697.050 ;
        RECT 862.950 691.500 865.050 693.600 ;
        RECT 862.950 685.950 865.050 688.050 ;
        RECT 863.400 673.050 864.450 685.950 ;
        RECT 857.400 671.400 861.450 672.450 ;
        RECT 857.400 604.050 858.450 671.400 ;
        RECT 862.950 670.950 865.050 673.050 ;
        RECT 866.250 671.250 867.750 672.150 ;
        RECT 868.950 670.950 871.050 673.050 ;
        RECT 859.950 667.950 862.050 670.050 ;
        RECT 863.250 668.850 864.750 669.750 ;
        RECT 865.950 667.950 868.050 670.050 ;
        RECT 869.250 668.850 871.050 669.750 ;
        RECT 859.950 665.850 862.050 666.750 ;
        RECT 862.950 664.950 865.050 667.050 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 860.400 628.050 861.450 643.950 ;
        RECT 859.950 625.950 862.050 628.050 ;
        RECT 859.950 622.950 862.050 625.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 839.400 541.050 840.450 601.950 ;
        RECT 850.950 598.950 853.050 601.050 ;
        RECT 854.250 599.250 855.750 600.150 ;
        RECT 856.950 598.950 859.050 601.050 ;
        RECT 847.950 595.950 850.050 598.050 ;
        RECT 851.250 596.850 852.750 597.750 ;
        RECT 853.950 595.950 856.050 598.050 ;
        RECT 857.250 596.850 859.050 597.750 ;
        RECT 847.950 593.850 850.050 594.750 ;
        RECT 853.950 592.950 856.050 595.050 ;
        RECT 844.950 561.450 847.050 562.050 ;
        RECT 842.400 560.400 847.050 561.450 ;
        RECT 838.950 538.950 841.050 541.050 ;
        RECT 838.950 533.400 841.050 535.500 ;
        RECT 839.400 516.600 840.600 533.400 ;
        RECT 838.950 514.500 841.050 516.600 ;
        RECT 842.400 511.050 843.450 560.400 ;
        RECT 844.950 559.950 847.050 560.400 ;
        RECT 848.250 560.250 849.750 561.150 ;
        RECT 850.950 559.950 853.050 562.050 ;
        RECT 844.950 557.850 846.750 558.750 ;
        RECT 847.950 556.950 850.050 559.050 ;
        RECT 851.250 557.850 853.050 558.750 ;
        RECT 848.400 553.050 849.450 556.950 ;
        RECT 847.950 550.950 850.050 553.050 ;
        RECT 850.950 538.950 853.050 541.050 ;
        RECT 844.950 529.950 847.050 532.050 ;
        RECT 845.400 529.050 846.450 529.950 ;
        RECT 851.400 529.050 852.450 538.950 ;
        RECT 844.950 526.950 847.050 529.050 ;
        RECT 850.950 526.950 853.050 529.050 ;
        RECT 854.400 526.050 855.450 592.950 ;
        RECT 856.950 589.950 859.050 592.050 ;
        RECT 857.400 559.050 858.450 589.950 ;
        RECT 856.950 556.950 859.050 559.050 ;
        RECT 860.400 540.450 861.450 622.950 ;
        RECT 863.400 622.050 864.450 664.950 ;
        RECT 866.400 646.050 867.450 667.950 ;
        RECT 865.950 643.950 868.050 646.050 ;
        RECT 865.950 629.250 868.050 630.150 ;
        RECT 871.950 629.250 874.050 630.150 ;
        RECT 865.950 625.950 868.050 628.050 ;
        RECT 869.250 626.250 870.750 627.150 ;
        RECT 871.950 625.950 874.050 628.050 ;
        RECT 866.400 625.050 867.450 625.950 ;
        RECT 865.950 622.950 868.050 625.050 ;
        RECT 868.950 622.950 871.050 625.050 ;
        RECT 871.950 622.950 874.050 625.050 ;
        RECT 869.400 622.050 870.450 622.950 ;
        RECT 862.950 619.950 865.050 622.050 ;
        RECT 865.950 619.950 868.050 622.050 ;
        RECT 868.950 619.950 871.050 622.050 ;
        RECT 866.400 604.050 867.450 619.950 ;
        RECT 868.950 616.950 871.050 619.050 ;
        RECT 869.400 604.050 870.450 616.950 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 872.400 601.050 873.450 622.950 ;
        RECT 875.400 601.050 876.450 767.400 ;
        RECT 877.950 701.250 880.050 702.150 ;
        RECT 883.950 701.250 886.050 702.150 ;
        RECT 877.950 697.950 880.050 700.050 ;
        RECT 881.250 698.250 882.750 699.150 ;
        RECT 883.950 697.950 886.050 700.050 ;
        RECT 878.400 697.050 879.450 697.950 ;
        RECT 877.950 694.950 880.050 697.050 ;
        RECT 880.950 694.950 883.050 697.050 ;
        RECT 877.950 631.950 880.050 634.050 ;
        RECT 865.950 600.450 868.050 601.050 ;
        RECT 863.400 599.400 868.050 600.450 ;
        RECT 863.400 598.050 864.450 599.400 ;
        RECT 865.950 598.950 868.050 599.400 ;
        RECT 869.250 599.250 870.750 600.150 ;
        RECT 871.950 598.950 874.050 601.050 ;
        RECT 874.950 598.950 877.050 601.050 ;
        RECT 862.950 595.950 865.050 598.050 ;
        RECT 865.950 596.850 867.750 597.750 ;
        RECT 868.950 595.950 871.050 598.050 ;
        RECT 872.250 596.850 873.750 597.750 ;
        RECT 874.950 595.950 877.050 598.050 ;
        RECT 862.950 592.950 865.050 595.050 ;
        RECT 871.950 592.950 874.050 595.050 ;
        RECT 874.950 593.850 877.050 594.750 ;
        RECT 863.400 562.050 864.450 592.950 ;
        RECT 872.400 565.050 873.450 592.950 ;
        RECT 874.950 589.950 877.050 592.050 ;
        RECT 865.950 562.950 868.050 565.050 ;
        RECT 871.950 562.950 874.050 565.050 ;
        RECT 866.400 562.050 867.450 562.950 ;
        RECT 862.950 559.950 865.050 562.050 ;
        RECT 865.950 559.950 868.050 562.050 ;
        RECT 869.250 560.250 870.750 561.150 ;
        RECT 871.950 559.950 874.050 562.050 ;
        RECT 865.950 557.850 867.750 558.750 ;
        RECT 868.950 556.950 871.050 559.050 ;
        RECT 872.250 557.850 874.050 558.750 ;
        RECT 868.950 553.950 871.050 556.050 ;
        RECT 857.400 539.400 861.450 540.450 ;
        RECT 844.950 524.850 847.050 525.750 ;
        RECT 850.950 524.850 853.050 525.750 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 841.950 508.950 844.050 511.050 ;
        RECT 838.950 487.950 841.050 490.050 ;
        RECT 844.950 489.450 847.050 490.050 ;
        RECT 842.400 488.400 847.050 489.450 ;
        RECT 850.950 489.450 853.050 490.050 ;
        RECT 829.950 481.950 832.050 484.050 ;
        RECT 835.950 481.950 838.050 484.050 ;
        RECT 829.950 479.850 832.050 480.750 ;
        RECT 826.950 475.500 829.050 477.600 ;
        RECT 832.950 475.950 835.050 478.050 ;
        RECT 817.950 466.950 820.050 469.050 ;
        RECT 818.400 453.450 819.450 466.950 ;
        RECT 833.400 466.050 834.450 475.950 ;
        RECT 835.950 466.950 838.050 469.050 ;
        RECT 832.950 463.950 835.050 466.050 ;
        RECT 833.400 460.050 834.450 463.950 ;
        RECT 823.950 459.450 826.050 460.050 ;
        RECT 823.950 458.400 828.450 459.450 ;
        RECT 823.950 457.950 826.050 458.400 ;
        RECT 820.950 455.250 823.050 456.150 ;
        RECT 823.950 455.850 826.050 456.750 ;
        RECT 827.400 454.050 828.450 458.400 ;
        RECT 832.950 457.950 835.050 460.050 ;
        RECT 836.400 457.050 837.450 466.950 ;
        RECT 832.950 455.850 834.750 456.750 ;
        RECT 835.950 454.950 838.050 457.050 ;
        RECT 820.950 453.450 823.050 454.050 ;
        RECT 818.400 452.400 823.050 453.450 ;
        RECT 820.950 451.950 823.050 452.400 ;
        RECT 826.950 451.950 829.050 454.050 ;
        RECT 835.950 452.850 838.050 453.750 ;
        RECT 839.400 453.450 840.450 487.950 ;
        RECT 842.400 487.050 843.450 488.400 ;
        RECT 844.950 487.950 847.050 488.400 ;
        RECT 848.250 488.250 849.750 489.150 ;
        RECT 850.950 488.400 855.450 489.450 ;
        RECT 850.950 487.950 853.050 488.400 ;
        RECT 841.950 484.950 844.050 487.050 ;
        RECT 844.950 485.850 846.750 486.750 ;
        RECT 847.950 484.950 850.050 487.050 ;
        RECT 851.250 485.850 853.050 486.750 ;
        RECT 842.400 469.050 843.450 484.950 ;
        RECT 847.950 478.950 850.050 481.050 ;
        RECT 841.950 466.950 844.050 469.050 ;
        RECT 848.400 456.450 849.450 478.950 ;
        RECT 854.400 478.050 855.450 488.400 ;
        RECT 853.950 475.950 856.050 478.050 ;
        RECT 853.950 461.400 856.050 463.500 ;
        RECT 850.950 458.250 853.050 459.150 ;
        RECT 850.950 456.450 853.050 457.050 ;
        RECT 841.950 455.250 844.050 456.150 ;
        RECT 848.400 455.400 853.050 456.450 ;
        RECT 850.950 454.950 853.050 455.400 ;
        RECT 841.950 453.450 844.050 454.050 ;
        RECT 839.400 452.400 844.050 453.450 ;
        RECT 841.950 451.950 844.050 452.400 ;
        RECT 850.950 451.950 853.050 454.050 ;
        RECT 841.950 427.950 844.050 430.050 ;
        RECT 826.950 422.400 829.050 424.500 ;
        RECT 817.950 413.250 820.050 414.150 ;
        RECT 817.950 411.450 820.050 412.050 ;
        RECT 815.400 410.400 820.050 411.450 ;
        RECT 812.400 397.050 813.450 409.950 ;
        RECT 811.950 394.950 814.050 397.050 ;
        RECT 809.400 392.400 813.450 393.450 ;
        RECT 802.950 389.400 805.050 391.500 ;
        RECT 796.950 383.400 801.450 384.450 ;
        RECT 796.950 382.950 799.050 383.400 ;
        RECT 790.950 380.850 793.050 381.750 ;
        RECT 796.950 380.850 799.050 381.750 ;
        RECT 793.950 350.400 796.050 352.500 ;
        RECT 794.400 333.600 795.600 350.400 ;
        RECT 800.400 349.050 801.450 383.400 ;
        RECT 803.400 372.600 804.600 389.400 ;
        RECT 808.950 388.950 811.050 391.050 ;
        RECT 802.950 370.500 805.050 372.600 ;
        RECT 799.950 346.950 802.050 349.050 ;
        RECT 799.950 341.250 802.050 342.150 ;
        RECT 805.950 341.250 808.050 342.150 ;
        RECT 809.400 340.050 810.450 388.950 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 805.950 337.950 808.050 340.050 ;
        RECT 808.950 337.950 811.050 340.050 ;
        RECT 793.950 331.500 796.050 333.600 ;
        RECT 806.400 328.050 807.450 337.950 ;
        RECT 775.950 325.950 778.050 328.050 ;
        RECT 784.950 325.950 787.050 328.050 ;
        RECT 787.950 325.950 790.050 328.050 ;
        RECT 799.950 325.950 802.050 328.050 ;
        RECT 805.950 325.950 808.050 328.050 ;
        RECT 772.950 319.950 775.050 322.050 ;
        RECT 769.950 313.950 772.050 316.050 ;
        RECT 766.950 310.950 769.050 313.050 ;
        RECT 770.250 311.850 771.750 312.750 ;
        RECT 772.950 310.950 775.050 313.050 ;
        RECT 766.950 308.850 769.050 309.750 ;
        RECT 772.950 308.850 775.050 309.750 ;
        RECT 776.400 273.450 777.450 325.950 ;
        RECT 784.950 319.950 787.050 322.050 ;
        RECT 785.400 313.050 786.450 319.950 ;
        RECT 790.950 313.950 793.050 316.050 ;
        RECT 778.950 310.950 781.050 313.050 ;
        RECT 784.950 310.950 787.050 313.050 ;
        RECT 788.250 311.250 790.050 312.150 ;
        RECT 790.950 311.850 793.050 312.750 ;
        RECT 793.950 311.250 796.050 312.150 ;
        RECT 773.400 272.400 777.450 273.450 ;
        RECT 773.400 271.050 774.450 272.400 ;
        RECT 769.950 268.950 772.050 271.050 ;
        RECT 772.950 268.950 775.050 271.050 ;
        RECT 776.250 269.250 778.050 270.150 ;
        RECT 770.400 211.050 771.450 268.950 ;
        RECT 772.950 266.850 774.750 267.750 ;
        RECT 775.950 265.950 778.050 268.050 ;
        RECT 772.950 247.950 775.050 250.050 ;
        RECT 773.400 241.050 774.450 247.950 ;
        RECT 776.400 247.050 777.450 265.950 ;
        RECT 779.400 256.050 780.450 310.950 ;
        RECT 784.950 308.850 786.750 309.750 ;
        RECT 787.950 307.950 790.050 310.050 ;
        RECT 793.950 307.950 796.050 310.050 ;
        RECT 800.400 298.050 801.450 325.950 ;
        RECT 805.950 322.950 808.050 325.050 ;
        RECT 806.400 316.050 807.450 322.950 ;
        RECT 802.950 313.950 805.050 316.050 ;
        RECT 805.950 313.950 808.050 316.050 ;
        RECT 799.950 295.950 802.050 298.050 ;
        RECT 784.950 271.950 787.050 274.050 ;
        RECT 799.950 272.250 802.050 273.150 ;
        RECT 785.400 268.050 786.450 271.950 ;
        RECT 790.950 269.250 792.750 270.150 ;
        RECT 793.950 268.950 796.050 271.050 ;
        RECT 797.250 269.250 798.750 270.150 ;
        RECT 799.950 268.950 802.050 271.050 ;
        RECT 784.950 265.950 787.050 268.050 ;
        RECT 790.950 265.950 793.050 268.050 ;
        RECT 794.250 266.850 795.750 267.750 ;
        RECT 796.950 265.950 799.050 268.050 ;
        RECT 778.950 253.950 781.050 256.050 ;
        RECT 781.950 253.950 784.050 256.050 ;
        RECT 778.950 250.950 781.050 253.050 ;
        RECT 775.950 244.950 778.050 247.050 ;
        RECT 779.400 241.050 780.450 250.950 ;
        RECT 772.950 238.950 775.050 241.050 ;
        RECT 776.250 239.250 777.750 240.150 ;
        RECT 778.950 238.950 781.050 241.050 ;
        RECT 782.400 238.050 783.450 253.950 ;
        RECT 787.950 244.950 790.050 247.050 ;
        RECT 772.950 236.850 774.750 237.750 ;
        RECT 775.950 235.950 778.050 238.050 ;
        RECT 779.250 236.850 780.750 237.750 ;
        RECT 781.950 235.950 784.050 238.050 ;
        RECT 781.950 233.850 784.050 234.750 ;
        RECT 769.950 208.950 772.050 211.050 ;
        RECT 778.950 202.950 781.050 205.050 ;
        RECT 748.950 200.250 751.050 201.150 ;
        RECT 763.950 199.950 766.050 202.050 ;
        RECT 775.950 200.250 778.050 201.150 ;
        RECT 748.950 196.950 751.050 199.050 ;
        RECT 752.250 197.250 753.750 198.150 ;
        RECT 754.950 196.950 757.050 199.050 ;
        RECT 758.250 197.250 760.050 198.150 ;
        RECT 760.950 196.950 763.050 199.050 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 766.950 197.250 768.750 198.150 ;
        RECT 769.950 196.950 772.050 199.050 ;
        RECT 773.250 197.250 774.750 198.150 ;
        RECT 775.950 196.950 778.050 199.050 ;
        RECT 751.950 193.950 754.050 196.050 ;
        RECT 755.250 194.850 756.750 195.750 ;
        RECT 757.950 193.950 760.050 196.050 ;
        RECT 752.400 187.050 753.450 193.950 ;
        RECT 751.950 184.950 754.050 187.050 ;
        RECT 757.950 173.400 760.050 175.500 ;
        RECT 746.400 170.400 750.450 171.450 ;
        RECT 739.950 166.950 742.050 169.050 ;
        RECT 745.950 166.950 748.050 169.050 ;
        RECT 749.400 166.050 750.450 170.400 ;
        RECT 751.950 169.950 754.050 172.050 ;
        RECT 752.400 169.050 753.450 169.950 ;
        RECT 751.950 166.950 754.050 169.050 ;
        RECT 745.950 164.850 748.050 165.750 ;
        RECT 748.950 163.950 751.050 166.050 ;
        RECT 751.950 164.850 754.050 165.750 ;
        RECT 736.950 159.300 739.050 161.400 ;
        RECT 737.550 155.700 738.750 159.300 ;
        RECT 758.400 156.600 759.600 173.400 ;
        RECT 736.950 153.600 739.050 155.700 ;
        RECT 757.950 154.500 760.050 156.600 ;
        RECT 730.950 145.950 733.050 148.050 ;
        RECT 691.950 128.250 693.750 129.150 ;
        RECT 694.950 127.950 697.050 130.050 ;
        RECT 698.250 128.250 699.750 129.150 ;
        RECT 700.950 127.950 703.050 130.050 ;
        RECT 706.950 127.950 709.050 130.050 ;
        RECT 715.950 127.950 718.050 130.050 ;
        RECT 718.950 127.950 721.050 130.050 ;
        RECT 724.950 127.950 727.050 130.050 ;
        RECT 691.950 124.950 694.050 127.050 ;
        RECT 692.400 118.050 693.450 124.950 ;
        RECT 695.400 124.050 696.450 127.950 ;
        RECT 697.950 124.950 700.050 127.050 ;
        RECT 701.250 125.850 703.050 126.750 ;
        RECT 707.400 124.050 708.450 127.950 ;
        RECT 709.950 126.450 712.050 127.050 ;
        RECT 712.950 126.450 715.050 127.050 ;
        RECT 709.950 125.400 715.050 126.450 ;
        RECT 716.400 126.450 717.450 127.950 ;
        RECT 718.950 126.450 721.050 127.050 ;
        RECT 716.400 125.400 721.050 126.450 ;
        RECT 709.950 124.950 712.050 125.400 ;
        RECT 712.950 124.950 715.050 125.400 ;
        RECT 718.950 124.950 721.050 125.400 ;
        RECT 722.250 125.250 724.050 126.150 ;
        RECT 694.950 121.950 697.050 124.050 ;
        RECT 706.950 121.950 709.050 124.050 ;
        RECT 710.400 120.450 711.450 124.950 ;
        RECT 712.950 122.850 715.050 123.750 ;
        RECT 715.950 122.250 718.050 123.150 ;
        RECT 718.950 122.850 720.750 123.750 ;
        RECT 721.950 121.950 724.050 124.050 ;
        RECT 710.400 119.400 714.450 120.450 ;
        RECT 691.950 115.950 694.050 118.050 ;
        RECT 697.950 112.950 700.050 115.050 ;
        RECT 691.950 101.400 694.050 103.500 ;
        RECT 688.950 91.950 691.050 94.050 ;
        RECT 692.250 89.400 693.450 101.400 ;
        RECT 694.950 98.250 697.050 99.150 ;
        RECT 694.950 96.450 697.050 97.050 ;
        RECT 698.400 96.450 699.450 112.950 ;
        RECT 706.950 99.450 709.050 100.050 ;
        RECT 694.950 95.400 699.450 96.450 ;
        RECT 704.400 98.400 709.050 99.450 ;
        RECT 694.950 94.950 697.050 95.400 ;
        RECT 691.950 87.300 694.050 89.400 ;
        RECT 692.250 83.700 693.450 87.300 ;
        RECT 704.400 85.050 705.450 98.400 ;
        RECT 706.950 97.950 709.050 98.400 ;
        RECT 706.950 95.850 709.050 96.750 ;
        RECT 709.950 95.250 712.050 96.150 ;
        RECT 709.950 93.450 712.050 94.050 ;
        RECT 713.400 93.450 714.450 119.400 ;
        RECT 715.950 118.950 718.050 121.050 ;
        RECT 716.400 118.050 717.450 118.950 ;
        RECT 715.950 115.950 718.050 118.050 ;
        RECT 718.950 94.950 721.050 97.050 ;
        RECT 709.950 92.400 714.450 93.450 ;
        RECT 709.950 91.950 712.050 92.400 ;
        RECT 691.950 81.600 694.050 83.700 ;
        RECT 703.950 82.950 706.050 85.050 ;
        RECT 688.950 56.250 691.050 57.150 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 695.400 55.050 696.450 55.950 ;
        RECT 688.950 52.950 691.050 55.050 ;
        RECT 692.250 53.250 693.750 54.150 ;
        RECT 694.950 52.950 697.050 55.050 ;
        RECT 698.250 53.250 700.050 54.150 ;
        RECT 689.400 52.050 690.450 52.950 ;
        RECT 704.400 52.050 705.450 82.950 ;
        RECT 719.400 55.050 720.450 94.950 ;
        RECT 725.400 94.050 726.450 127.950 ;
        RECT 731.400 102.450 732.450 145.950 ;
        RECT 761.400 142.050 762.450 196.950 ;
        RECT 764.400 160.050 765.450 196.950 ;
        RECT 766.950 193.950 769.050 196.050 ;
        RECT 770.250 194.850 771.750 195.750 ;
        RECT 772.950 193.950 775.050 196.050 ;
        RECT 773.400 193.050 774.450 193.950 ;
        RECT 772.950 190.950 775.050 193.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 773.400 175.050 774.450 178.950 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 769.950 169.950 772.050 172.050 ;
        RECT 766.950 166.950 769.050 169.050 ;
        RECT 763.950 157.950 766.050 160.050 ;
        RECT 760.950 139.950 763.050 142.050 ;
        RECT 736.950 130.950 739.050 133.050 ;
        RECT 737.400 127.050 738.450 130.950 ;
        RECT 742.950 128.250 745.050 129.150 ;
        RECT 763.950 128.250 766.050 129.150 ;
        RECT 733.950 125.250 735.750 126.150 ;
        RECT 736.950 124.950 739.050 127.050 ;
        RECT 740.250 125.250 741.750 126.150 ;
        RECT 742.950 124.950 745.050 127.050 ;
        RECT 754.950 125.250 756.750 126.150 ;
        RECT 757.950 124.950 760.050 127.050 ;
        RECT 761.250 125.250 762.750 126.150 ;
        RECT 763.950 124.950 766.050 127.050 ;
        RECT 733.950 121.950 736.050 124.050 ;
        RECT 737.250 122.850 738.750 123.750 ;
        RECT 739.950 121.950 742.050 124.050 ;
        RECT 754.950 121.950 757.050 124.050 ;
        RECT 758.250 122.850 759.750 123.750 ;
        RECT 760.950 121.950 763.050 124.050 ;
        RECT 734.400 121.050 735.450 121.950 ;
        RECT 755.400 121.050 756.450 121.950 ;
        RECT 733.950 118.950 736.050 121.050 ;
        RECT 754.950 118.950 757.050 121.050 ;
        RECT 767.400 106.050 768.450 166.950 ;
        RECT 770.400 154.050 771.450 169.950 ;
        RECT 773.400 169.050 774.450 172.950 ;
        RECT 779.400 169.050 780.450 202.950 ;
        RECT 781.950 199.950 784.050 202.050 ;
        RECT 784.950 199.950 787.050 202.050 ;
        RECT 782.400 178.050 783.450 199.950 ;
        RECT 781.950 175.950 784.050 178.050 ;
        RECT 785.400 172.050 786.450 199.950 ;
        RECT 788.400 172.050 789.450 244.950 ;
        RECT 796.950 241.950 799.050 244.050 ;
        RECT 797.400 241.050 798.450 241.950 ;
        RECT 800.400 241.050 801.450 268.950 ;
        RECT 803.400 253.050 804.450 313.950 ;
        RECT 805.950 311.850 808.050 312.750 ;
        RECT 808.950 311.250 811.050 312.150 ;
        RECT 808.950 307.950 811.050 310.050 ;
        RECT 812.400 285.450 813.450 392.400 ;
        RECT 815.400 358.050 816.450 410.400 ;
        RECT 817.950 409.950 820.050 410.400 ;
        RECT 827.400 405.600 828.600 422.400 ;
        RECT 832.950 413.250 835.050 414.150 ;
        RECT 838.950 413.250 841.050 414.150 ;
        RECT 832.950 409.950 835.050 412.050 ;
        RECT 838.950 411.450 841.050 412.050 ;
        RECT 842.400 411.450 843.450 427.950 ;
        RECT 847.950 423.300 850.050 425.400 ;
        RECT 848.250 419.700 849.450 423.300 ;
        RECT 847.950 417.600 850.050 419.700 ;
        RECT 838.950 410.400 843.450 411.450 ;
        RECT 838.950 409.950 841.050 410.400 ;
        RECT 826.950 403.500 829.050 405.600 ;
        RECT 839.400 388.050 840.450 409.950 ;
        RECT 848.250 405.600 849.450 417.600 ;
        RECT 851.400 412.050 852.450 451.950 ;
        RECT 854.550 449.400 855.750 461.400 ;
        RECT 853.950 447.300 856.050 449.400 ;
        RECT 854.550 443.700 855.750 447.300 ;
        RECT 853.950 441.600 856.050 443.700 ;
        RECT 850.950 409.950 853.050 412.050 ;
        RECT 850.950 407.850 853.050 408.750 ;
        RECT 847.950 403.500 850.050 405.600 ;
        RECT 853.950 389.400 856.050 391.500 ;
        RECT 838.950 385.950 841.050 388.050 ;
        RECT 844.950 387.450 847.050 388.050 ;
        RECT 844.950 386.400 849.450 387.450 ;
        RECT 844.950 385.950 847.050 386.400 ;
        RECT 823.950 382.950 826.050 385.050 ;
        RECT 829.950 384.450 832.050 385.050 ;
        RECT 827.250 383.250 828.750 384.150 ;
        RECT 829.950 383.400 834.450 384.450 ;
        RECT 829.950 382.950 832.050 383.400 ;
        RECT 833.400 382.050 834.450 383.400 ;
        RECT 841.950 383.250 844.050 384.150 ;
        RECT 844.950 383.850 847.050 384.750 ;
        RECT 848.400 384.450 849.450 386.400 ;
        RECT 850.950 386.250 853.050 387.150 ;
        RECT 850.950 384.450 853.050 385.050 ;
        RECT 848.400 383.400 853.050 384.450 ;
        RECT 820.950 381.450 823.050 382.050 ;
        RECT 818.400 380.400 823.050 381.450 ;
        RECT 824.250 380.850 825.750 381.750 ;
        RECT 818.400 379.050 819.450 380.400 ;
        RECT 820.950 379.950 823.050 380.400 ;
        RECT 826.950 379.950 829.050 382.050 ;
        RECT 830.250 380.850 832.050 381.750 ;
        RECT 832.950 379.950 835.050 382.050 ;
        RECT 841.950 379.950 844.050 382.050 ;
        RECT 817.950 376.950 820.050 379.050 ;
        RECT 820.950 377.850 823.050 378.750 ;
        RECT 814.950 355.950 817.050 358.050 ;
        RECT 820.950 355.950 823.050 358.050 ;
        RECT 814.950 351.300 817.050 353.400 ;
        RECT 815.250 347.700 816.450 351.300 ;
        RECT 814.950 345.600 817.050 347.700 ;
        RECT 815.250 333.600 816.450 345.600 ;
        RECT 817.950 343.950 820.050 346.050 ;
        RECT 818.400 340.050 819.450 343.950 ;
        RECT 817.950 337.950 820.050 340.050 ;
        RECT 817.950 335.850 820.050 336.750 ;
        RECT 814.950 331.500 817.050 333.600 ;
        RECT 817.950 328.950 820.050 331.050 ;
        RECT 814.950 316.950 817.050 319.050 ;
        RECT 809.400 284.400 813.450 285.450 ;
        RECT 802.950 250.950 805.050 253.050 ;
        RECT 805.950 241.950 808.050 244.050 ;
        RECT 806.400 241.050 807.450 241.950 ;
        RECT 796.950 238.950 799.050 241.050 ;
        RECT 799.950 238.950 802.050 241.050 ;
        RECT 802.950 238.950 805.050 241.050 ;
        RECT 805.950 238.950 808.050 241.050 ;
        RECT 796.950 236.850 799.050 237.750 ;
        RECT 799.950 236.250 802.050 237.150 ;
        RECT 799.950 232.950 802.050 235.050 ;
        RECT 799.950 208.950 802.050 211.050 ;
        RECT 790.950 199.950 793.050 202.050 ;
        RECT 794.250 200.250 795.750 201.150 ;
        RECT 796.950 199.950 799.050 202.050 ;
        RECT 790.950 197.850 792.750 198.750 ;
        RECT 793.950 196.950 796.050 199.050 ;
        RECT 797.250 197.850 799.050 198.750 ;
        RECT 796.950 175.950 799.050 178.050 ;
        RECT 784.950 169.950 787.050 172.050 ;
        RECT 787.950 169.950 790.050 172.050 ;
        RECT 772.950 166.950 775.050 169.050 ;
        RECT 776.250 167.250 777.750 168.150 ;
        RECT 778.950 166.950 781.050 169.050 ;
        RECT 782.250 167.250 783.750 168.150 ;
        RECT 784.950 166.950 787.050 169.050 ;
        RECT 787.950 166.950 790.050 169.050 ;
        RECT 790.950 166.950 793.050 169.050 ;
        RECT 772.950 164.850 774.750 165.750 ;
        RECT 775.950 163.950 778.050 166.050 ;
        RECT 779.250 164.850 780.750 165.750 ;
        RECT 781.950 163.950 784.050 166.050 ;
        RECT 785.250 164.850 787.050 165.750 ;
        RECT 776.400 163.050 777.450 163.950 ;
        RECT 782.400 163.050 783.450 163.950 ;
        RECT 775.950 160.950 778.050 163.050 ;
        RECT 781.950 160.950 784.050 163.050 ;
        RECT 772.950 157.950 775.050 160.050 ;
        RECT 769.950 151.950 772.050 154.050 ;
        RECT 770.400 127.050 771.450 151.950 ;
        RECT 769.950 124.950 772.050 127.050 ;
        RECT 766.950 103.950 769.050 106.050 ;
        RECT 731.400 101.400 735.450 102.450 ;
        RECT 757.950 101.400 760.050 103.500 ;
        RECT 767.400 103.050 768.450 103.950 ;
        RECT 734.400 97.050 735.450 101.400 ;
        RECT 748.950 99.450 751.050 100.050 ;
        RECT 748.950 98.400 753.450 99.450 ;
        RECT 748.950 97.950 751.050 98.400 ;
        RECT 727.950 94.950 730.050 97.050 ;
        RECT 733.950 96.450 736.050 97.050 ;
        RECT 731.250 95.250 732.750 96.150 ;
        RECT 733.950 95.400 738.450 96.450 ;
        RECT 733.950 94.950 736.050 95.400 ;
        RECT 724.950 93.450 727.050 94.050 ;
        RECT 722.400 92.400 727.050 93.450 ;
        RECT 728.250 92.850 729.750 93.750 ;
        RECT 722.400 60.450 723.450 92.400 ;
        RECT 724.950 91.950 727.050 92.400 ;
        RECT 730.950 91.950 733.050 94.050 ;
        RECT 734.250 92.850 736.050 93.750 ;
        RECT 724.950 89.850 727.050 90.750 ;
        RECT 731.400 67.050 732.450 91.950 ;
        RECT 730.950 64.950 733.050 67.050 ;
        RECT 737.400 61.050 738.450 95.400 ;
        RECT 745.950 95.250 748.050 96.150 ;
        RECT 748.950 95.850 751.050 96.750 ;
        RECT 752.400 96.450 753.450 98.400 ;
        RECT 754.950 98.250 757.050 99.150 ;
        RECT 754.950 96.450 757.050 97.050 ;
        RECT 752.400 95.400 757.050 96.450 ;
        RECT 754.950 94.950 757.050 95.400 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 758.550 89.400 759.750 101.400 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 757.950 87.300 760.050 89.400 ;
        RECT 758.550 83.700 759.750 87.300 ;
        RECT 757.950 81.600 760.050 83.700 ;
        RECT 757.950 64.950 760.050 67.050 ;
        RECT 722.400 59.400 726.450 60.450 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 709.950 53.250 711.750 54.150 ;
        RECT 712.950 52.950 715.050 55.050 ;
        RECT 718.950 52.950 721.050 55.050 ;
        RECT 722.400 52.050 723.450 55.950 ;
        RECT 688.950 49.950 691.050 52.050 ;
        RECT 691.950 49.950 694.050 52.050 ;
        RECT 695.250 50.850 696.750 51.750 ;
        RECT 697.950 49.950 700.050 52.050 ;
        RECT 703.950 49.950 706.050 52.050 ;
        RECT 709.950 49.950 712.050 52.050 ;
        RECT 713.250 50.850 715.050 51.750 ;
        RECT 715.950 50.250 718.050 51.150 ;
        RECT 718.950 50.850 721.050 51.750 ;
        RECT 721.950 49.950 724.050 52.050 ;
        RECT 692.400 46.050 693.450 49.950 ;
        RECT 698.400 49.050 699.450 49.950 ;
        RECT 697.950 46.950 700.050 49.050 ;
        RECT 715.950 46.950 718.050 49.050 ;
        RECT 685.950 43.950 688.050 46.050 ;
        RECT 691.950 43.950 694.050 46.050 ;
        RECT 685.950 34.950 688.050 37.050 ;
        RECT 703.950 34.950 706.050 37.050 ;
        RECT 676.950 28.950 679.050 31.050 ;
        RECT 661.950 25.950 664.050 28.050 ;
        RECT 664.950 25.950 667.050 28.050 ;
        RECT 662.400 25.050 663.450 25.950 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 665.250 23.850 666.750 24.750 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 677.400 22.050 678.450 28.950 ;
        RECT 686.400 28.050 687.450 34.950 ;
        RECT 685.950 25.950 688.050 28.050 ;
        RECT 704.400 25.050 705.450 34.950 ;
        RECT 725.400 28.050 726.450 59.400 ;
        RECT 736.950 58.950 739.050 61.050 ;
        RECT 751.950 58.950 754.050 61.050 ;
        RECT 752.400 58.050 753.450 58.950 ;
        RECT 758.400 58.050 759.450 64.950 ;
        RECT 736.950 57.450 739.050 58.050 ;
        RECT 734.400 56.400 739.050 57.450 ;
        RECT 727.950 52.950 730.050 55.050 ;
        RECT 730.950 53.250 733.050 54.150 ;
        RECT 728.400 51.450 729.450 52.950 ;
        RECT 730.950 51.450 733.050 52.050 ;
        RECT 728.400 50.400 733.050 51.450 ;
        RECT 730.950 49.950 733.050 50.400 ;
        RECT 734.400 49.050 735.450 56.400 ;
        RECT 736.950 55.950 739.050 56.400 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 755.250 56.250 756.750 57.150 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 736.950 53.850 739.050 54.750 ;
        RECT 739.950 53.250 742.050 54.150 ;
        RECT 751.950 53.850 753.750 54.750 ;
        RECT 754.950 52.950 757.050 55.050 ;
        RECT 758.250 53.850 760.050 54.750 ;
        RECT 739.950 49.950 742.050 52.050 ;
        RECT 755.400 49.050 756.450 52.950 ;
        RECT 733.950 46.950 736.050 49.050 ;
        RECT 754.950 46.950 757.050 49.050 ;
        RECT 730.950 43.950 733.050 46.050 ;
        RECT 724.950 25.950 727.050 28.050 ;
        RECT 682.950 23.250 685.050 24.150 ;
        RECT 685.950 23.850 688.050 24.750 ;
        RECT 691.950 24.450 694.050 25.050 ;
        RECT 688.950 23.250 690.750 24.150 ;
        RECT 691.950 23.400 696.450 24.450 ;
        RECT 691.950 22.950 694.050 23.400 ;
        RECT 661.950 20.850 664.050 21.750 ;
        RECT 667.950 20.850 670.050 21.750 ;
        RECT 676.950 19.950 679.050 22.050 ;
        RECT 682.950 19.950 685.050 22.050 ;
        RECT 688.950 19.950 691.050 22.050 ;
        RECT 692.250 20.850 694.050 21.750 ;
        RECT 689.400 19.050 690.450 19.950 ;
        RECT 695.400 19.050 696.450 23.400 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 707.250 23.250 708.750 24.150 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 724.950 23.850 727.050 24.750 ;
        RECT 727.950 23.250 730.050 24.150 ;
        RECT 703.950 20.850 705.750 21.750 ;
        RECT 706.950 19.950 709.050 22.050 ;
        RECT 710.250 20.850 711.750 21.750 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 727.950 21.450 730.050 22.050 ;
        RECT 731.400 21.450 732.450 43.950 ;
        RECT 757.950 29.400 760.050 31.500 ;
        RECT 764.400 31.050 765.450 100.950 ;
        RECT 767.400 97.050 768.450 100.950 ;
        RECT 766.950 94.950 769.050 97.050 ;
        RECT 766.950 92.850 769.050 93.750 ;
        RECT 770.400 91.050 771.450 124.950 ;
        RECT 773.400 123.450 774.450 157.950 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 779.400 127.050 780.450 133.950 ;
        RECT 784.950 128.250 787.050 129.150 ;
        RECT 775.950 125.250 777.750 126.150 ;
        RECT 778.950 124.950 781.050 127.050 ;
        RECT 782.250 125.250 783.750 126.150 ;
        RECT 784.950 124.950 787.050 127.050 ;
        RECT 775.950 123.450 778.050 124.050 ;
        RECT 773.400 122.400 778.050 123.450 ;
        RECT 779.250 122.850 780.750 123.750 ;
        RECT 775.950 121.950 778.050 122.400 ;
        RECT 781.950 121.950 784.050 124.050 ;
        RECT 772.950 94.950 775.050 97.050 ;
        RECT 776.400 94.050 777.450 121.950 ;
        RECT 778.950 101.400 781.050 103.500 ;
        RECT 772.950 92.850 775.050 93.750 ;
        RECT 775.950 91.950 778.050 94.050 ;
        RECT 769.950 88.950 772.050 91.050 ;
        RECT 779.400 84.600 780.600 101.400 ;
        RECT 782.400 97.050 783.450 121.950 ;
        RECT 781.950 94.950 784.050 97.050 ;
        RECT 778.950 82.500 781.050 84.600 ;
        RECT 778.950 64.950 781.050 67.050 ;
        RECT 766.950 58.950 769.050 61.050 ;
        RECT 767.400 51.450 768.450 58.950 ;
        RECT 769.950 53.250 772.050 54.150 ;
        RECT 775.950 53.250 778.050 54.150 ;
        RECT 769.950 51.450 772.050 52.050 ;
        RECT 767.400 50.400 772.050 51.450 ;
        RECT 775.950 51.450 778.050 52.050 ;
        RECT 779.400 51.450 780.450 64.950 ;
        RECT 769.950 49.950 772.050 50.400 ;
        RECT 773.250 50.250 774.750 51.150 ;
        RECT 775.950 50.400 780.450 51.450 ;
        RECT 775.950 49.950 778.050 50.400 ;
        RECT 772.950 46.950 775.050 49.050 ;
        RECT 785.400 43.050 786.450 124.950 ;
        RECT 784.950 40.950 787.050 43.050 ;
        RECT 745.950 25.950 748.050 28.050 ;
        RECT 746.400 22.050 747.450 25.950 ;
        RECT 727.950 20.400 732.450 21.450 ;
        RECT 727.950 19.950 730.050 20.400 ;
        RECT 742.950 20.250 744.750 21.150 ;
        RECT 745.950 19.950 748.050 22.050 ;
        RECT 749.250 20.250 751.050 21.150 ;
        RECT 751.950 19.950 754.050 22.050 ;
        RECT 643.950 16.950 646.050 17.400 ;
        RECT 649.950 17.400 654.450 18.450 ;
        RECT 649.950 16.950 652.050 17.400 ;
        RECT 658.950 16.950 661.050 19.050 ;
        RECT 688.950 16.950 691.050 19.050 ;
        RECT 694.950 16.950 697.050 19.050 ;
        RECT 712.950 17.850 715.050 18.750 ;
        RECT 742.950 16.950 745.050 19.050 ;
        RECT 746.250 17.850 747.750 18.750 ;
        RECT 748.950 18.450 751.050 19.050 ;
        RECT 752.400 18.450 753.450 19.950 ;
        RECT 748.950 17.400 753.450 18.450 ;
        RECT 748.950 16.950 751.050 17.400 ;
        RECT 484.950 13.950 487.050 16.050 ;
        RECT 520.950 13.950 523.050 16.050 ;
        RECT 743.400 13.050 744.450 16.950 ;
        RECT 151.950 10.950 154.050 13.050 ;
        RECT 280.950 10.950 283.050 13.050 ;
        RECT 388.950 10.950 391.050 13.050 ;
        RECT 742.950 10.950 745.050 13.050 ;
        RECT 758.400 12.600 759.600 29.400 ;
        RECT 763.950 28.950 766.050 31.050 ;
        RECT 769.950 28.950 772.050 31.050 ;
        RECT 778.950 29.400 781.050 31.500 ;
        RECT 763.950 25.950 766.050 28.050 ;
        RECT 764.400 25.050 765.450 25.950 ;
        RECT 770.400 25.050 771.450 28.950 ;
        RECT 763.950 22.950 766.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 763.950 20.850 766.050 21.750 ;
        RECT 769.950 20.850 772.050 21.750 ;
        RECT 779.250 17.400 780.450 29.400 ;
        RECT 781.950 26.250 784.050 27.150 ;
        RECT 781.950 22.950 784.050 25.050 ;
        RECT 782.400 19.050 783.450 22.950 ;
        RECT 788.400 19.050 789.450 166.950 ;
        RECT 791.400 94.050 792.450 166.950 ;
        RECT 793.950 163.950 796.050 166.050 ;
        RECT 794.400 157.050 795.450 163.950 ;
        RECT 793.950 154.950 796.050 157.050 ;
        RECT 793.950 101.400 796.050 103.500 ;
        RECT 790.950 91.950 793.050 94.050 ;
        RECT 794.400 84.600 795.600 101.400 ;
        RECT 793.950 82.500 796.050 84.600 ;
        RECT 793.950 55.950 796.050 58.050 ;
        RECT 794.400 55.050 795.450 55.950 ;
        RECT 793.950 52.950 796.050 55.050 ;
        RECT 790.950 50.250 793.050 51.150 ;
        RECT 793.950 50.850 796.050 51.750 ;
        RECT 790.950 46.950 793.050 49.050 ;
        RECT 797.400 34.050 798.450 175.950 ;
        RECT 800.400 172.050 801.450 208.950 ;
        RECT 803.400 202.050 804.450 238.950 ;
        RECT 805.950 236.850 808.050 237.750 ;
        RECT 802.950 199.950 805.050 202.050 ;
        RECT 803.400 196.050 804.450 199.950 ;
        RECT 802.950 193.950 805.050 196.050 ;
        RECT 802.950 175.950 805.050 178.050 ;
        RECT 799.950 169.950 802.050 172.050 ;
        RECT 803.400 169.050 804.450 175.950 ;
        RECT 809.400 175.050 810.450 284.400 ;
        RECT 811.950 278.400 814.050 280.500 ;
        RECT 812.400 261.600 813.600 278.400 ;
        RECT 811.950 259.500 814.050 261.600 ;
        RECT 811.950 232.950 814.050 235.050 ;
        RECT 812.400 202.050 813.450 232.950 ;
        RECT 815.400 208.050 816.450 316.950 ;
        RECT 818.400 310.050 819.450 328.950 ;
        RECT 821.400 313.050 822.450 355.950 ;
        RECT 829.950 349.950 832.050 352.050 ;
        RECT 823.950 346.950 826.050 349.050 ;
        RECT 824.400 319.050 825.450 346.950 ;
        RECT 830.400 339.450 831.450 349.950 ;
        RECT 835.950 343.950 838.050 346.050 ;
        RECT 836.400 343.050 837.450 343.950 ;
        RECT 848.400 343.050 849.450 383.400 ;
        RECT 850.950 382.950 853.050 383.400 ;
        RECT 854.550 377.400 855.750 389.400 ;
        RECT 853.950 375.300 856.050 377.400 ;
        RECT 854.550 371.700 855.750 375.300 ;
        RECT 853.950 369.600 856.050 371.700 ;
        RECT 857.400 346.050 858.450 539.400 ;
        RECT 859.950 533.400 862.050 535.500 ;
        RECT 860.250 521.400 861.450 533.400 ;
        RECT 862.950 530.250 865.050 531.150 ;
        RECT 865.950 529.950 868.050 532.050 ;
        RECT 862.950 528.450 865.050 529.050 ;
        RECT 866.400 528.450 867.450 529.950 ;
        RECT 862.950 527.400 867.450 528.450 ;
        RECT 862.950 526.950 865.050 527.400 ;
        RECT 869.400 523.050 870.450 553.950 ;
        RECT 871.950 550.950 874.050 553.050 ;
        RECT 859.950 519.300 862.050 521.400 ;
        RECT 868.950 520.950 871.050 523.050 ;
        RECT 860.250 515.700 861.450 519.300 ;
        RECT 859.950 513.600 862.050 515.700 ;
        RECT 859.950 508.950 862.050 511.050 ;
        RECT 860.400 489.450 861.450 508.950 ;
        RECT 862.950 489.450 865.050 490.050 ;
        RECT 860.400 488.400 865.050 489.450 ;
        RECT 860.400 487.050 861.450 488.400 ;
        RECT 862.950 487.950 865.050 488.400 ;
        RECT 866.250 488.250 867.750 489.150 ;
        RECT 868.950 487.950 871.050 490.050 ;
        RECT 859.950 484.950 862.050 487.050 ;
        RECT 862.950 485.850 864.750 486.750 ;
        RECT 865.950 484.950 868.050 487.050 ;
        RECT 869.250 485.850 871.050 486.750 ;
        RECT 866.400 484.050 867.450 484.950 ;
        RECT 865.950 481.950 868.050 484.050 ;
        RECT 865.950 478.950 868.050 481.050 ;
        RECT 862.950 456.450 865.050 457.050 ;
        RECT 860.400 455.400 865.050 456.450 ;
        RECT 860.400 430.050 861.450 455.400 ;
        RECT 862.950 454.950 865.050 455.400 ;
        RECT 862.950 452.850 865.050 453.750 ;
        RECT 866.400 439.050 867.450 478.950 ;
        RECT 868.950 454.950 871.050 457.050 ;
        RECT 868.950 452.850 871.050 453.750 ;
        RECT 865.950 436.950 868.050 439.050 ;
        RECT 859.950 427.950 862.050 430.050 ;
        RECT 859.950 415.950 862.050 418.050 ;
        RECT 860.400 411.450 861.450 415.950 ;
        RECT 862.950 413.250 865.050 414.150 ;
        RECT 868.950 413.250 871.050 414.150 ;
        RECT 862.950 411.450 865.050 412.050 ;
        RECT 860.400 410.400 865.050 411.450 ;
        RECT 862.950 409.950 865.050 410.400 ;
        RECT 866.250 410.250 867.750 411.150 ;
        RECT 868.950 409.950 871.050 412.050 ;
        RECT 865.950 406.950 868.050 409.050 ;
        RECT 862.950 385.950 865.050 388.050 ;
        RECT 863.400 385.050 864.450 385.950 ;
        RECT 862.950 382.950 865.050 385.050 ;
        RECT 868.950 382.950 871.050 385.050 ;
        RECT 862.950 380.850 865.050 381.750 ;
        RECT 868.950 380.850 871.050 381.750 ;
        RECT 856.950 343.950 859.050 346.050 ;
        RECT 862.950 344.250 865.050 345.150 ;
        RECT 865.950 343.950 868.050 346.050 ;
        RECT 832.950 341.250 834.750 342.150 ;
        RECT 835.950 340.950 838.050 343.050 ;
        RECT 839.250 341.250 840.750 342.150 ;
        RECT 841.950 340.950 844.050 343.050 ;
        RECT 845.250 341.250 847.050 342.150 ;
        RECT 847.950 340.950 850.050 343.050 ;
        RECT 850.950 340.950 853.050 343.050 ;
        RECT 853.950 341.250 855.750 342.150 ;
        RECT 856.950 340.950 859.050 343.050 ;
        RECT 860.250 341.250 861.750 342.150 ;
        RECT 862.950 340.950 865.050 343.050 ;
        RECT 832.950 339.450 835.050 340.050 ;
        RECT 830.400 338.400 835.050 339.450 ;
        RECT 836.250 338.850 837.750 339.750 ;
        RECT 823.950 316.950 826.050 319.050 ;
        RECT 824.400 316.050 825.450 316.950 ;
        RECT 823.950 313.950 826.050 316.050 ;
        RECT 820.950 310.950 823.050 313.050 ;
        RECT 823.950 311.850 826.050 312.750 ;
        RECT 826.950 311.250 829.050 312.150 ;
        RECT 817.950 307.950 820.050 310.050 ;
        RECT 820.950 307.950 823.050 310.050 ;
        RECT 826.950 307.950 829.050 310.050 ;
        RECT 817.950 269.250 820.050 270.150 ;
        RECT 817.950 265.950 820.050 268.050 ;
        RECT 821.400 246.450 822.450 307.950 ;
        RECT 826.950 295.950 829.050 298.050 ;
        RECT 827.400 271.050 828.450 295.950 ;
        RECT 823.950 269.250 826.050 270.150 ;
        RECT 826.950 268.950 829.050 271.050 ;
        RECT 823.950 267.450 826.050 268.050 ;
        RECT 827.400 267.450 828.450 268.950 ;
        RECT 823.950 266.400 828.450 267.450 ;
        RECT 823.950 265.950 826.050 266.400 ;
        RECT 824.400 262.050 825.450 265.950 ;
        RECT 826.950 262.950 829.050 265.050 ;
        RECT 823.950 259.950 826.050 262.050 ;
        RECT 823.950 250.950 826.050 253.050 ;
        RECT 818.400 245.400 822.450 246.450 ;
        RECT 818.400 241.050 819.450 245.400 ;
        RECT 820.950 241.950 823.050 244.050 ;
        RECT 824.400 241.050 825.450 250.950 ;
        RECT 817.950 238.950 820.050 241.050 ;
        RECT 821.250 239.850 822.750 240.750 ;
        RECT 823.950 238.950 826.050 241.050 ;
        RECT 817.950 236.850 820.050 237.750 ;
        RECT 823.950 236.850 826.050 237.750 ;
        RECT 814.950 205.950 817.050 208.050 ;
        RECT 817.950 202.950 820.050 205.050 ;
        RECT 811.950 199.950 814.050 202.050 ;
        RECT 812.400 199.050 813.450 199.950 ;
        RECT 818.400 199.050 819.450 202.950 ;
        RECT 811.950 196.950 814.050 199.050 ;
        RECT 817.950 196.950 820.050 199.050 ;
        RECT 821.250 197.250 823.050 198.150 ;
        RECT 823.950 196.950 826.050 199.050 ;
        RECT 811.950 194.850 814.050 195.750 ;
        RECT 814.950 194.250 817.050 195.150 ;
        RECT 817.950 194.850 819.750 195.750 ;
        RECT 820.950 193.950 823.050 196.050 ;
        RECT 814.950 190.950 817.050 193.050 ;
        RECT 815.400 187.050 816.450 190.950 ;
        RECT 814.950 184.950 817.050 187.050 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 808.950 172.950 811.050 175.050 ;
        RECT 811.950 169.950 814.050 172.050 ;
        RECT 802.950 166.950 805.050 169.050 ;
        RECT 806.250 167.250 807.750 168.150 ;
        RECT 808.950 166.950 811.050 169.050 ;
        RECT 799.950 163.950 802.050 166.050 ;
        RECT 803.250 164.850 804.750 165.750 ;
        RECT 805.950 163.950 808.050 166.050 ;
        RECT 809.250 164.850 811.050 165.750 ;
        RECT 799.950 161.850 802.050 162.750 ;
        RECT 802.950 139.950 805.050 142.050 ;
        RECT 803.400 127.050 804.450 139.950 ;
        RECT 806.400 136.050 807.450 163.950 ;
        RECT 805.950 133.950 808.050 136.050 ;
        RECT 802.950 124.950 805.050 127.050 ;
        RECT 799.950 122.250 802.050 123.150 ;
        RECT 802.950 122.850 805.050 123.750 ;
        RECT 799.950 118.950 802.050 121.050 ;
        RECT 800.400 115.050 801.450 118.950 ;
        RECT 799.950 112.950 802.050 115.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 806.400 97.050 807.450 100.950 ;
        RECT 799.950 94.950 802.050 97.050 ;
        RECT 805.950 94.950 808.050 97.050 ;
        RECT 799.950 92.850 802.050 93.750 ;
        RECT 805.950 92.850 808.050 93.750 ;
        RECT 812.400 64.050 813.450 169.950 ;
        RECT 818.400 169.050 819.450 178.950 ;
        RECT 824.400 169.050 825.450 196.950 ;
        RECT 827.400 196.050 828.450 262.950 ;
        RECT 830.400 244.050 831.450 338.400 ;
        RECT 832.950 337.950 835.050 338.400 ;
        RECT 838.950 337.950 841.050 340.050 ;
        RECT 842.250 338.850 843.750 339.750 ;
        RECT 844.950 337.950 847.050 340.050 ;
        RECT 847.950 337.950 850.050 340.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 832.950 279.300 835.050 281.400 ;
        RECT 833.250 275.700 834.450 279.300 ;
        RECT 836.400 277.050 837.450 334.950 ;
        RECT 839.400 316.050 840.450 337.950 ;
        RECT 838.950 313.950 841.050 316.050 ;
        RECT 838.950 310.950 841.050 313.050 ;
        RECT 844.950 312.450 847.050 313.050 ;
        RECT 842.400 311.400 847.050 312.450 ;
        RECT 838.950 308.850 841.050 309.750 ;
        RECT 832.950 273.600 835.050 275.700 ;
        RECT 835.950 274.950 838.050 277.050 ;
        RECT 833.250 261.600 834.450 273.600 ;
        RECT 835.950 267.450 838.050 268.050 ;
        RECT 835.950 266.400 840.450 267.450 ;
        RECT 835.950 265.950 838.050 266.400 ;
        RECT 835.950 263.850 838.050 264.750 ;
        RECT 832.950 259.500 835.050 261.600 ;
        RECT 829.950 241.950 832.050 244.050 ;
        RECT 830.400 229.050 831.450 241.950 ;
        RECT 839.400 241.050 840.450 266.400 ;
        RECT 838.950 238.950 841.050 241.050 ;
        RECT 842.400 240.450 843.450 311.400 ;
        RECT 844.950 310.950 847.050 311.400 ;
        RECT 844.950 308.850 847.050 309.750 ;
        RECT 844.950 304.950 847.050 307.050 ;
        RECT 845.400 265.050 846.450 304.950 ;
        RECT 848.400 280.050 849.450 337.950 ;
        RECT 851.400 337.050 852.450 340.950 ;
        RECT 853.950 337.950 856.050 340.050 ;
        RECT 857.250 338.850 858.750 339.750 ;
        RECT 859.950 337.950 862.050 340.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 854.400 319.050 855.450 337.950 ;
        RECT 863.400 336.450 864.450 340.950 ;
        RECT 860.400 335.400 864.450 336.450 ;
        RECT 853.950 316.950 856.050 319.050 ;
        RECT 850.950 313.950 853.050 316.050 ;
        RECT 851.400 310.050 852.450 313.950 ;
        RECT 854.400 313.050 855.450 316.950 ;
        RECT 856.950 313.950 859.050 316.050 ;
        RECT 853.950 310.950 856.050 313.050 ;
        RECT 850.950 307.950 853.050 310.050 ;
        RECT 847.950 277.950 850.050 280.050 ;
        RECT 847.950 274.950 850.050 277.050 ;
        RECT 844.950 262.950 847.050 265.050 ;
        RECT 842.400 239.400 846.450 240.450 ;
        RECT 835.950 236.250 837.750 237.150 ;
        RECT 838.950 235.950 841.050 238.050 ;
        RECT 842.250 236.250 844.050 237.150 ;
        RECT 835.950 232.950 838.050 235.050 ;
        RECT 839.250 233.850 840.750 234.750 ;
        RECT 841.950 234.450 844.050 235.050 ;
        RECT 845.400 234.450 846.450 239.400 ;
        RECT 841.950 233.400 846.450 234.450 ;
        RECT 841.950 232.950 844.050 233.400 ;
        RECT 829.950 226.950 832.050 229.050 ;
        RECT 832.950 199.950 835.050 202.050 ;
        RECT 833.400 199.050 834.450 199.950 ;
        RECT 832.950 196.950 835.050 199.050 ;
        RECT 838.950 196.950 841.050 199.050 ;
        RECT 842.250 197.250 844.050 198.150 ;
        RECT 826.950 193.950 829.050 196.050 ;
        RECT 832.950 194.850 835.050 195.750 ;
        RECT 835.950 194.250 838.050 195.150 ;
        RECT 838.950 194.850 840.750 195.750 ;
        RECT 841.950 193.950 844.050 196.050 ;
        RECT 835.950 190.950 838.050 193.050 ;
        RECT 835.950 172.950 838.050 175.050 ;
        RECT 817.950 166.950 820.050 169.050 ;
        RECT 821.250 167.250 822.750 168.150 ;
        RECT 823.950 166.950 826.050 169.050 ;
        RECT 827.250 167.250 828.750 168.150 ;
        RECT 829.950 166.950 832.050 169.050 ;
        RECT 817.950 164.850 819.750 165.750 ;
        RECT 820.950 163.950 823.050 166.050 ;
        RECT 824.250 164.850 825.750 165.750 ;
        RECT 826.950 163.950 829.050 166.050 ;
        RECT 830.250 164.850 832.050 165.750 ;
        RECT 821.400 154.050 822.450 163.950 ;
        RECT 827.400 163.050 828.450 163.950 ;
        RECT 826.950 160.950 829.050 163.050 ;
        RECT 820.950 151.950 823.050 154.050 ;
        RECT 832.950 151.950 835.050 154.050 ;
        RECT 826.950 133.950 829.050 136.050 ;
        RECT 820.950 128.250 823.050 129.150 ;
        RECT 827.400 127.050 828.450 133.950 ;
        RECT 833.400 127.050 834.450 151.950 ;
        RECT 820.950 124.950 823.050 127.050 ;
        RECT 824.250 125.250 825.750 126.150 ;
        RECT 826.950 124.950 829.050 127.050 ;
        RECT 830.250 125.250 832.050 126.150 ;
        RECT 832.950 124.950 835.050 127.050 ;
        RECT 821.400 124.050 822.450 124.950 ;
        RECT 820.950 121.950 823.050 124.050 ;
        RECT 823.950 121.950 826.050 124.050 ;
        RECT 827.250 122.850 828.750 123.750 ;
        RECT 829.950 123.450 832.050 124.050 ;
        RECT 833.400 123.450 834.450 124.950 ;
        RECT 829.950 122.400 834.450 123.450 ;
        RECT 829.950 121.950 832.050 122.400 ;
        RECT 836.400 109.050 837.450 172.950 ;
        RECT 845.400 171.450 846.450 233.400 ;
        RECT 848.400 196.050 849.450 274.950 ;
        RECT 854.400 273.450 855.450 310.950 ;
        RECT 857.400 283.050 858.450 313.950 ;
        RECT 860.400 313.050 861.450 335.400 ;
        RECT 862.950 316.950 865.050 319.050 ;
        RECT 863.400 313.050 864.450 316.950 ;
        RECT 866.400 316.050 867.450 343.950 ;
        RECT 872.400 337.050 873.450 550.950 ;
        RECT 875.400 525.450 876.450 589.950 ;
        RECT 878.400 532.050 879.450 631.950 ;
        RECT 881.400 607.050 882.450 694.950 ;
        RECT 884.400 625.050 885.450 697.950 ;
        RECT 883.950 622.950 886.050 625.050 ;
        RECT 880.950 604.950 883.050 607.050 ;
        RECT 880.950 595.950 883.050 598.050 ;
        RECT 881.400 553.050 882.450 595.950 ;
        RECT 880.950 550.950 883.050 553.050 ;
        RECT 877.950 529.950 880.050 532.050 ;
        RECT 877.950 527.850 880.050 528.750 ;
        RECT 880.950 527.250 883.050 528.150 ;
        RECT 875.400 524.400 879.450 525.450 ;
        RECT 874.950 520.950 877.050 523.050 ;
        RECT 875.400 481.050 876.450 520.950 ;
        RECT 874.950 478.950 877.050 481.050 ;
        RECT 874.950 461.400 877.050 463.500 ;
        RECT 875.400 444.600 876.600 461.400 ;
        RECT 874.950 442.500 877.050 444.600 ;
        RECT 874.950 436.950 877.050 439.050 ;
        RECT 875.400 409.050 876.450 436.950 ;
        RECT 874.950 406.950 877.050 409.050 ;
        RECT 874.950 389.400 877.050 391.500 ;
        RECT 875.400 372.600 876.600 389.400 ;
        RECT 874.950 370.500 877.050 372.600 ;
        RECT 874.950 341.250 877.050 342.150 ;
        RECT 874.950 337.950 877.050 340.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 878.400 336.450 879.450 524.400 ;
        RECT 880.950 523.950 883.050 526.050 ;
        RECT 880.950 341.250 883.050 342.150 ;
        RECT 875.400 335.400 879.450 336.450 ;
        RECT 865.950 313.950 868.050 316.050 ;
        RECT 859.950 310.950 862.050 313.050 ;
        RECT 862.950 310.950 865.050 313.050 ;
        RECT 866.250 311.250 867.750 312.150 ;
        RECT 868.950 310.950 871.050 313.050 ;
        RECT 859.950 307.950 862.050 310.050 ;
        RECT 863.250 308.850 864.750 309.750 ;
        RECT 865.950 307.950 868.050 310.050 ;
        RECT 869.250 308.850 871.050 309.750 ;
        RECT 875.400 307.050 876.450 335.400 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 877.950 316.950 880.050 319.050 ;
        RECT 878.400 313.050 879.450 316.950 ;
        RECT 877.950 310.950 880.050 313.050 ;
        RECT 877.950 308.850 880.050 309.750 ;
        RECT 859.950 305.850 862.050 306.750 ;
        RECT 865.950 304.950 868.050 307.050 ;
        RECT 874.950 304.950 877.050 307.050 ;
        RECT 859.950 300.450 862.050 301.050 ;
        RECT 859.950 299.400 864.450 300.450 ;
        RECT 859.950 298.950 862.050 299.400 ;
        RECT 856.950 280.950 859.050 283.050 ;
        RECT 856.950 277.950 859.050 280.050 ;
        RECT 851.400 272.400 855.450 273.450 ;
        RECT 851.400 253.050 852.450 272.400 ;
        RECT 853.950 268.950 856.050 271.050 ;
        RECT 853.950 266.850 856.050 267.750 ;
        RECT 850.950 250.950 853.050 253.050 ;
        RECT 857.400 241.050 858.450 277.950 ;
        RECT 863.400 241.050 864.450 299.400 ;
        RECT 866.400 247.050 867.450 304.950 ;
        RECT 868.950 280.950 871.050 283.050 ;
        RECT 865.950 244.950 868.050 247.050 ;
        RECT 869.400 246.450 870.450 280.950 ;
        RECT 874.950 266.850 877.050 267.750 ;
        RECT 881.400 265.050 882.450 334.950 ;
        RECT 883.950 308.850 886.050 309.750 ;
        RECT 874.950 262.950 877.050 265.050 ;
        RECT 880.950 262.950 883.050 265.050 ;
        RECT 869.400 245.400 873.450 246.450 ;
        RECT 868.950 241.950 871.050 244.050 ;
        RECT 869.400 241.050 870.450 241.950 ;
        RECT 856.950 238.950 859.050 241.050 ;
        RECT 860.250 239.250 861.750 240.150 ;
        RECT 862.950 238.950 865.050 241.050 ;
        RECT 866.250 239.250 867.750 240.150 ;
        RECT 868.950 238.950 871.050 241.050 ;
        RECT 856.950 236.850 858.750 237.750 ;
        RECT 859.950 235.950 862.050 238.050 ;
        RECT 863.250 236.850 864.750 237.750 ;
        RECT 865.950 235.950 868.050 238.050 ;
        RECT 869.250 236.850 871.050 237.750 ;
        RECT 866.400 235.050 867.450 235.950 ;
        RECT 859.950 232.950 862.050 235.050 ;
        RECT 865.950 232.950 868.050 235.050 ;
        RECT 856.950 196.950 859.050 199.050 ;
        RECT 847.950 193.950 850.050 196.050 ;
        RECT 856.950 194.850 859.050 195.750 ;
        RECT 856.950 173.400 859.050 175.500 ;
        RECT 842.400 170.400 846.450 171.450 ;
        RECT 847.950 171.450 850.050 172.050 ;
        RECT 847.950 170.400 852.450 171.450 ;
        RECT 842.400 151.050 843.450 170.400 ;
        RECT 847.950 169.950 850.050 170.400 ;
        RECT 844.950 167.250 847.050 168.150 ;
        RECT 847.950 167.850 850.050 168.750 ;
        RECT 851.400 168.450 852.450 170.400 ;
        RECT 853.950 170.250 856.050 171.150 ;
        RECT 853.950 168.450 856.050 169.050 ;
        RECT 851.400 167.400 856.050 168.450 ;
        RECT 853.950 166.950 856.050 167.400 ;
        RECT 844.950 163.950 847.050 166.050 ;
        RECT 853.950 163.950 856.050 166.050 ;
        RECT 841.950 148.950 844.050 151.050 ;
        RECT 838.950 134.400 841.050 136.500 ;
        RECT 839.400 117.600 840.600 134.400 ;
        RECT 838.950 115.500 841.050 117.600 ;
        RECT 835.950 106.950 838.050 109.050 ;
        RECT 842.400 106.050 843.450 148.950 ;
        RECT 844.950 125.250 847.050 126.150 ;
        RECT 850.950 125.250 853.050 126.150 ;
        RECT 844.950 121.950 847.050 124.050 ;
        RECT 850.950 123.450 853.050 124.050 ;
        RECT 854.400 123.450 855.450 163.950 ;
        RECT 857.550 161.400 858.750 173.400 ;
        RECT 856.950 159.300 859.050 161.400 ;
        RECT 857.550 155.700 858.750 159.300 ;
        RECT 856.950 153.600 859.050 155.700 ;
        RECT 860.400 150.450 861.450 232.950 ;
        RECT 862.950 229.950 865.050 232.050 ;
        RECT 863.400 162.450 864.450 229.950 ;
        RECT 865.950 196.950 868.050 199.050 ;
        RECT 866.400 169.050 867.450 196.950 ;
        RECT 872.400 171.450 873.450 245.400 ;
        RECT 869.400 170.400 873.450 171.450 ;
        RECT 865.950 166.950 868.050 169.050 ;
        RECT 865.950 164.850 868.050 165.750 ;
        RECT 863.400 161.400 867.450 162.450 ;
        RECT 850.950 122.400 855.450 123.450 ;
        RECT 857.400 149.400 861.450 150.450 ;
        RECT 850.950 121.950 853.050 122.400 ;
        RECT 826.950 103.950 829.050 106.050 ;
        RECT 841.950 103.950 844.050 106.050 ;
        RECT 814.950 101.400 817.050 103.500 ;
        RECT 815.250 89.400 816.450 101.400 ;
        RECT 817.950 98.250 820.050 99.150 ;
        RECT 820.950 97.950 823.050 100.050 ;
        RECT 817.950 96.450 820.050 97.050 ;
        RECT 821.400 96.450 822.450 97.950 ;
        RECT 817.950 95.400 822.450 96.450 ;
        RECT 817.950 94.950 820.050 95.400 ;
        RECT 827.400 94.050 828.450 103.950 ;
        RECT 851.400 103.050 852.450 121.950 ;
        RECT 853.950 106.950 856.050 109.050 ;
        RECT 850.950 100.950 853.050 103.050 ;
        RECT 832.950 96.450 835.050 97.050 ;
        RECT 830.400 95.400 835.050 96.450 ;
        RECT 817.950 91.950 820.050 94.050 ;
        RECT 826.950 91.950 829.050 94.050 ;
        RECT 814.950 87.300 817.050 89.400 ;
        RECT 815.250 83.700 816.450 87.300 ;
        RECT 814.950 81.600 817.050 83.700 ;
        RECT 811.950 61.950 814.050 64.050 ;
        RECT 812.400 61.050 813.450 61.950 ;
        RECT 811.950 58.950 814.050 61.050 ;
        RECT 805.950 57.450 808.050 58.050 ;
        RECT 803.400 56.400 808.050 57.450 ;
        RECT 803.400 55.050 804.450 56.400 ;
        RECT 805.950 55.950 808.050 56.400 ;
        RECT 809.250 56.250 810.750 57.150 ;
        RECT 811.950 55.950 814.050 58.050 ;
        RECT 802.950 52.950 805.050 55.050 ;
        RECT 805.950 53.850 807.750 54.750 ;
        RECT 808.950 52.950 811.050 55.050 ;
        RECT 812.250 53.850 814.050 54.750 ;
        RECT 818.400 43.050 819.450 91.950 ;
        RECT 830.400 88.050 831.450 95.400 ;
        RECT 832.950 94.950 835.050 95.400 ;
        RECT 836.250 95.250 837.750 96.150 ;
        RECT 838.950 94.950 841.050 97.050 ;
        RECT 844.950 96.450 847.050 97.050 ;
        RECT 842.250 95.250 843.750 96.150 ;
        RECT 844.950 95.400 849.450 96.450 ;
        RECT 844.950 94.950 847.050 95.400 ;
        RECT 848.400 94.050 849.450 95.400 ;
        RECT 832.950 92.850 834.750 93.750 ;
        RECT 835.950 91.950 838.050 94.050 ;
        RECT 839.250 92.850 840.750 93.750 ;
        RECT 841.950 91.950 844.050 94.050 ;
        RECT 845.250 92.850 847.050 93.750 ;
        RECT 847.950 91.950 850.050 94.050 ;
        RECT 836.400 91.050 837.450 91.950 ;
        RECT 835.950 88.950 838.050 91.050 ;
        RECT 829.950 85.950 832.050 88.050 ;
        RECT 829.950 58.950 832.050 61.050 ;
        RECT 830.400 55.050 831.450 58.950 ;
        RECT 823.950 52.950 826.050 55.050 ;
        RECT 829.950 52.950 832.050 55.050 ;
        RECT 833.250 53.250 835.050 54.150 ;
        RECT 823.950 50.850 826.050 51.750 ;
        RECT 826.950 50.250 829.050 51.150 ;
        RECT 829.950 50.850 831.750 51.750 ;
        RECT 832.950 49.950 835.050 52.050 ;
        RECT 826.950 46.950 829.050 49.050 ;
        RECT 827.400 46.050 828.450 46.950 ;
        RECT 826.950 43.950 829.050 46.050 ;
        RECT 817.950 40.950 820.050 43.050 ;
        RECT 826.950 40.950 829.050 43.050 ;
        RECT 796.950 31.950 799.050 34.050 ;
        RECT 814.950 25.950 817.050 28.050 ;
        RECT 815.400 25.050 816.450 25.950 ;
        RECT 827.400 25.050 828.450 40.950 ;
        RECT 836.400 36.450 837.450 88.950 ;
        RECT 838.950 85.950 841.050 88.050 ;
        RECT 839.400 49.050 840.450 85.950 ;
        RECT 838.950 46.950 841.050 49.050 ;
        RECT 833.400 35.400 837.450 36.450 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 818.250 23.250 819.750 24.150 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 824.250 23.250 825.750 24.150 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 833.400 22.050 834.450 35.400 ;
        RECT 835.950 29.400 838.050 31.500 ;
        RECT 793.950 20.250 795.750 21.150 ;
        RECT 796.950 19.950 799.050 22.050 ;
        RECT 800.250 20.250 802.050 21.150 ;
        RECT 814.950 20.850 816.750 21.750 ;
        RECT 817.950 19.950 820.050 22.050 ;
        RECT 821.250 20.850 822.750 21.750 ;
        RECT 823.950 19.950 826.050 22.050 ;
        RECT 827.250 20.850 829.050 21.750 ;
        RECT 832.950 19.950 835.050 22.050 ;
        RECT 824.400 19.050 825.450 19.950 ;
        RECT 778.950 15.300 781.050 17.400 ;
        RECT 781.950 16.950 784.050 19.050 ;
        RECT 787.950 16.950 790.050 19.050 ;
        RECT 793.950 16.950 796.050 19.050 ;
        RECT 797.250 17.850 798.750 18.750 ;
        RECT 799.950 16.950 802.050 19.050 ;
        RECT 823.950 16.950 826.050 19.050 ;
        RECT 757.950 10.500 760.050 12.600 ;
        RECT 779.250 11.700 780.450 15.300 ;
        RECT 836.400 12.600 837.600 29.400 ;
        RECT 842.400 27.450 843.450 91.950 ;
        RECT 854.400 88.050 855.450 106.950 ;
        RECT 857.400 100.050 858.450 149.400 ;
        RECT 859.950 135.300 862.050 137.400 ;
        RECT 860.250 131.700 861.450 135.300 ;
        RECT 859.950 129.600 862.050 131.700 ;
        RECT 860.250 117.600 861.450 129.600 ;
        RECT 862.950 121.950 865.050 124.050 ;
        RECT 862.950 119.850 865.050 120.750 ;
        RECT 859.950 115.500 862.050 117.600 ;
        RECT 866.400 117.450 867.450 161.400 ;
        RECT 863.400 116.400 867.450 117.450 ;
        RECT 856.950 97.950 859.050 100.050 ;
        RECT 859.950 97.950 862.050 100.050 ;
        RECT 856.950 95.250 859.050 96.150 ;
        RECT 859.950 95.850 862.050 96.750 ;
        RECT 856.950 91.950 859.050 94.050 ;
        RECT 853.950 85.950 856.050 88.050 ;
        RECT 856.950 56.250 859.050 57.150 ;
        RECT 847.950 53.250 849.750 54.150 ;
        RECT 850.950 52.950 853.050 55.050 ;
        RECT 854.250 53.250 855.750 54.150 ;
        RECT 856.950 52.950 859.050 55.050 ;
        RECT 857.400 52.050 858.450 52.950 ;
        RECT 847.950 49.950 850.050 52.050 ;
        RECT 851.250 50.850 852.750 51.750 ;
        RECT 853.950 49.950 856.050 52.050 ;
        RECT 856.950 49.950 859.050 52.050 ;
        RECT 848.400 46.050 849.450 49.950 ;
        RECT 854.400 49.050 855.450 49.950 ;
        RECT 853.950 46.950 856.050 49.050 ;
        RECT 847.950 43.950 850.050 46.050 ;
        RECT 847.950 28.950 850.050 31.050 ;
        RECT 856.950 29.400 859.050 31.500 ;
        RECT 839.400 26.400 843.450 27.450 ;
        RECT 839.400 19.050 840.450 26.400 ;
        RECT 848.400 25.050 849.450 28.950 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 841.950 20.850 844.050 21.750 ;
        RECT 847.950 20.850 850.050 21.750 ;
        RECT 838.950 16.950 841.050 19.050 ;
        RECT 857.250 17.400 858.450 29.400 ;
        RECT 859.950 26.250 862.050 27.150 ;
        RECT 859.950 22.950 862.050 25.050 ;
        RECT 863.400 22.050 864.450 116.400 ;
        RECT 869.400 96.450 870.450 170.400 ;
        RECT 871.950 166.950 874.050 169.050 ;
        RECT 871.950 164.850 874.050 165.750 ;
        RECT 875.400 162.450 876.450 262.950 ;
        RECT 877.950 194.850 880.050 195.750 ;
        RECT 880.950 175.950 883.050 178.050 ;
        RECT 877.950 173.400 880.050 175.500 ;
        RECT 866.400 95.400 870.450 96.450 ;
        RECT 872.400 161.400 876.450 162.450 ;
        RECT 866.400 91.050 867.450 95.400 ;
        RECT 872.400 94.050 873.450 161.400 ;
        RECT 878.400 156.600 879.600 173.400 ;
        RECT 881.400 169.050 882.450 175.950 ;
        RECT 880.950 166.950 883.050 169.050 ;
        RECT 877.950 154.500 880.050 156.600 ;
        RECT 880.950 124.950 883.050 127.050 ;
        RECT 877.950 122.250 880.050 123.150 ;
        RECT 880.950 122.850 883.050 123.750 ;
        RECT 877.950 118.950 880.050 121.050 ;
        RECT 868.950 92.250 870.750 93.150 ;
        RECT 871.950 91.950 874.050 94.050 ;
        RECT 875.250 92.250 877.050 93.150 ;
        RECT 877.950 91.950 880.050 94.050 ;
        RECT 865.950 88.950 868.050 91.050 ;
        RECT 868.950 88.950 871.050 91.050 ;
        RECT 872.250 89.850 873.750 90.750 ;
        RECT 874.950 88.950 877.050 91.050 ;
        RECT 869.400 88.050 870.450 88.950 ;
        RECT 868.950 85.950 871.050 88.050 ;
        RECT 868.950 52.950 871.050 55.050 ;
        RECT 874.950 52.950 877.050 55.050 ;
        RECT 869.400 43.050 870.450 52.950 ;
        RECT 871.950 50.250 874.050 51.150 ;
        RECT 874.950 50.850 877.050 51.750 ;
        RECT 871.950 46.950 874.050 49.050 ;
        RECT 868.950 40.950 871.050 43.050 ;
        RECT 868.950 31.950 871.050 34.050 ;
        RECT 862.950 19.950 865.050 22.050 ;
        RECT 856.950 15.300 859.050 17.400 ;
        RECT 869.400 16.050 870.450 31.950 ;
        RECT 872.400 28.050 873.450 46.950 ;
        RECT 871.950 25.950 874.050 28.050 ;
        RECT 878.400 25.050 879.450 91.950 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 877.950 22.950 880.050 25.050 ;
        RECT 872.400 19.050 873.450 22.950 ;
        RECT 874.950 20.250 876.750 21.150 ;
        RECT 877.950 19.950 880.050 22.050 ;
        RECT 881.250 20.250 883.050 21.150 ;
        RECT 871.950 16.950 874.050 19.050 ;
        RECT 874.950 16.950 877.050 19.050 ;
        RECT 878.250 17.850 879.750 18.750 ;
        RECT 880.950 16.950 883.050 19.050 ;
        RECT 875.400 16.050 876.450 16.950 ;
        RECT 778.950 9.600 781.050 11.700 ;
        RECT 835.950 10.500 838.050 12.600 ;
        RECT 857.250 11.700 858.450 15.300 ;
        RECT 868.950 13.950 871.050 16.050 ;
        RECT 874.950 13.950 877.050 16.050 ;
        RECT 856.950 9.600 859.050 11.700 ;
      LAYER metal3 ;
        RECT 745.950 894.600 748.050 895.050 ;
        RECT 862.950 894.600 865.050 895.050 ;
        RECT 745.950 893.400 865.050 894.600 ;
        RECT 745.950 892.950 748.050 893.400 ;
        RECT 862.950 892.950 865.050 893.400 ;
        RECT 175.950 889.950 178.050 892.050 ;
        RECT 250.950 889.950 253.050 892.050 ;
        RECT 325.950 891.600 328.050 892.050 ;
        RECT 340.950 891.600 343.050 892.050 ;
        RECT 314.400 890.400 343.050 891.600 ;
        RECT 31.950 888.600 34.050 889.050 ;
        RECT 43.950 888.600 46.050 889.050 ;
        RECT 31.950 887.400 46.050 888.600 ;
        RECT 31.950 886.950 34.050 887.400 ;
        RECT 43.950 886.950 46.050 887.400 ;
        RECT 49.950 888.600 52.050 889.050 ;
        RECT 70.950 888.600 73.050 889.050 ;
        RECT 49.950 887.400 73.050 888.600 ;
        RECT 49.950 886.950 52.050 887.400 ;
        RECT 70.950 886.950 73.050 887.400 ;
        RECT 76.950 888.600 79.050 889.050 ;
        RECT 148.950 888.600 151.050 889.050 ;
        RECT 76.950 887.400 151.050 888.600 ;
        RECT 76.950 886.950 79.050 887.400 ;
        RECT 148.950 886.950 151.050 887.400 ;
        RECT 160.950 888.600 163.050 889.050 ;
        RECT 176.400 888.600 177.600 889.950 ;
        RECT 160.950 887.400 177.600 888.600 ;
        RECT 235.950 888.600 238.050 889.050 ;
        RECT 251.400 888.600 252.600 889.950 ;
        RECT 314.400 889.050 315.600 890.400 ;
        RECT 325.950 889.950 328.050 890.400 ;
        RECT 340.950 889.950 343.050 890.400 ;
        RECT 382.950 891.600 385.050 892.050 ;
        RECT 397.950 891.600 400.050 892.050 ;
        RECT 382.950 890.400 400.050 891.600 ;
        RECT 382.950 889.950 385.050 890.400 ;
        RECT 397.950 889.950 400.050 890.400 ;
        RECT 550.950 891.600 553.050 892.050 ;
        RECT 574.950 891.600 577.050 892.050 ;
        RECT 550.950 890.400 577.050 891.600 ;
        RECT 550.950 889.950 553.050 890.400 ;
        RECT 574.950 889.950 577.050 890.400 ;
        RECT 580.950 891.600 583.050 892.050 ;
        RECT 586.950 891.600 589.050 892.050 ;
        RECT 598.950 891.600 601.050 892.050 ;
        RECT 637.950 891.600 640.050 892.050 ;
        RECT 580.950 890.400 585.600 891.600 ;
        RECT 580.950 889.950 583.050 890.400 ;
        RECT 235.950 887.400 252.600 888.600 ;
        RECT 274.950 888.600 277.050 889.050 ;
        RECT 295.950 888.600 298.050 889.050 ;
        RECT 274.950 887.400 298.050 888.600 ;
        RECT 160.950 886.950 163.050 887.400 ;
        RECT 235.950 886.950 238.050 887.400 ;
        RECT 274.950 886.950 277.050 887.400 ;
        RECT 295.950 886.950 298.050 887.400 ;
        RECT 313.950 886.950 316.050 889.050 ;
        RECT 403.950 888.600 406.050 889.050 ;
        RECT 424.950 888.600 427.050 889.050 ;
        RECT 403.950 887.400 427.050 888.600 ;
        RECT 403.950 886.950 406.050 887.400 ;
        RECT 424.950 886.950 427.050 887.400 ;
        RECT 433.950 888.600 436.050 889.050 ;
        RECT 484.950 888.600 487.050 889.050 ;
        RECT 433.950 887.400 487.050 888.600 ;
        RECT 433.950 886.950 436.050 887.400 ;
        RECT 484.950 886.950 487.050 887.400 ;
        RECT 496.950 888.600 499.050 889.050 ;
        RECT 505.950 888.600 508.050 889.050 ;
        RECT 496.950 887.400 508.050 888.600 ;
        RECT 584.400 888.600 585.600 890.400 ;
        RECT 586.950 890.400 601.050 891.600 ;
        RECT 586.950 889.950 589.050 890.400 ;
        RECT 598.950 889.950 601.050 890.400 ;
        RECT 617.400 890.400 640.050 891.600 ;
        RECT 617.400 888.600 618.600 890.400 ;
        RECT 637.950 889.950 640.050 890.400 ;
        RECT 835.950 891.600 838.050 892.050 ;
        RECT 856.950 891.600 859.050 892.050 ;
        RECT 835.950 890.400 859.050 891.600 ;
        RECT 835.950 889.950 838.050 890.400 ;
        RECT 856.950 889.950 859.050 890.400 ;
        RECT 584.400 887.400 618.600 888.600 ;
        RECT 619.950 888.600 622.050 889.050 ;
        RECT 643.950 888.600 646.050 889.050 ;
        RECT 685.950 888.600 688.050 889.050 ;
        RECT 619.950 887.400 642.600 888.600 ;
        RECT 496.950 886.950 499.050 887.400 ;
        RECT 505.950 886.950 508.050 887.400 ;
        RECT 619.950 886.950 622.050 887.400 ;
        RECT 641.400 886.050 642.600 887.400 ;
        RECT 643.950 887.400 688.050 888.600 ;
        RECT 643.950 886.950 646.050 887.400 ;
        RECT 685.950 886.950 688.050 887.400 ;
        RECT 691.950 888.600 694.050 889.050 ;
        RECT 781.950 888.600 784.050 889.050 ;
        RECT 691.950 887.400 784.050 888.600 ;
        RECT 691.950 886.950 694.050 887.400 ;
        RECT 781.950 886.950 784.050 887.400 ;
        RECT 787.950 888.600 790.050 889.050 ;
        RECT 823.950 888.600 826.050 889.050 ;
        RECT 787.950 887.400 826.050 888.600 ;
        RECT 787.950 886.950 790.050 887.400 ;
        RECT 823.950 886.950 826.050 887.400 ;
        RECT 10.950 885.600 13.050 886.050 ;
        RECT 46.950 885.600 49.050 886.050 ;
        RECT 10.950 884.400 49.050 885.600 ;
        RECT 10.950 883.950 13.050 884.400 ;
        RECT 46.950 883.950 49.050 884.400 ;
        RECT 52.950 885.600 55.050 886.050 ;
        RECT 103.950 885.600 106.050 886.050 ;
        RECT 52.950 884.400 106.050 885.600 ;
        RECT 52.950 883.950 55.050 884.400 ;
        RECT 103.950 883.950 106.050 884.400 ;
        RECT 124.950 885.600 127.050 886.050 ;
        RECT 199.950 885.600 202.050 886.050 ;
        RECT 214.950 885.600 217.050 886.050 ;
        RECT 124.950 884.400 198.600 885.600 ;
        RECT 124.950 883.950 127.050 884.400 ;
        RECT 10.950 882.600 13.050 883.050 ;
        RECT 16.950 882.600 19.050 883.050 ;
        RECT 10.950 881.400 19.050 882.600 ;
        RECT 10.950 880.950 13.050 881.400 ;
        RECT 16.950 880.950 19.050 881.400 ;
        RECT 28.950 882.600 31.050 883.050 ;
        RECT 46.950 882.600 49.050 883.050 ;
        RECT 28.950 881.400 49.050 882.600 ;
        RECT 28.950 880.950 31.050 881.400 ;
        RECT 46.950 880.950 49.050 881.400 ;
        RECT 88.950 882.600 91.050 883.050 ;
        RECT 100.950 882.600 103.050 883.050 ;
        RECT 88.950 881.400 103.050 882.600 ;
        RECT 88.950 880.950 91.050 881.400 ;
        RECT 100.950 880.950 103.050 881.400 ;
        RECT 178.950 882.600 181.050 883.050 ;
        RECT 187.950 882.600 190.050 883.050 ;
        RECT 178.950 881.400 190.050 882.600 ;
        RECT 197.400 882.600 198.600 884.400 ;
        RECT 199.950 884.400 217.050 885.600 ;
        RECT 199.950 883.950 202.050 884.400 ;
        RECT 214.950 883.950 217.050 884.400 ;
        RECT 220.950 885.600 223.050 886.050 ;
        RECT 247.950 885.600 250.050 886.050 ;
        RECT 220.950 884.400 250.050 885.600 ;
        RECT 220.950 883.950 223.050 884.400 ;
        RECT 247.950 883.950 250.050 884.400 ;
        RECT 277.950 885.600 280.050 886.050 ;
        RECT 328.950 885.600 331.050 886.050 ;
        RECT 277.950 884.400 331.050 885.600 ;
        RECT 277.950 883.950 280.050 884.400 ;
        RECT 328.950 883.950 331.050 884.400 ;
        RECT 367.950 885.600 370.050 886.050 ;
        RECT 400.950 885.600 403.050 886.050 ;
        RECT 367.950 884.400 403.050 885.600 ;
        RECT 367.950 883.950 370.050 884.400 ;
        RECT 400.950 883.950 403.050 884.400 ;
        RECT 406.950 885.600 409.050 886.050 ;
        RECT 457.950 885.600 460.050 886.050 ;
        RECT 406.950 884.400 460.050 885.600 ;
        RECT 406.950 883.950 409.050 884.400 ;
        RECT 457.950 883.950 460.050 884.400 ;
        RECT 481.950 885.600 484.050 886.050 ;
        RECT 502.950 885.600 505.050 886.050 ;
        RECT 481.950 884.400 505.050 885.600 ;
        RECT 481.950 883.950 484.050 884.400 ;
        RECT 502.950 883.950 505.050 884.400 ;
        RECT 526.950 885.600 529.050 886.050 ;
        RECT 547.950 885.600 550.050 886.050 ;
        RECT 526.950 884.400 550.050 885.600 ;
        RECT 526.950 883.950 529.050 884.400 ;
        RECT 547.950 883.950 550.050 884.400 ;
        RECT 565.950 885.600 568.050 886.050 ;
        RECT 574.950 885.600 577.050 886.050 ;
        RECT 565.950 884.400 577.050 885.600 ;
        RECT 565.950 883.950 568.050 884.400 ;
        RECT 574.950 883.950 577.050 884.400 ;
        RECT 601.950 885.600 604.050 886.050 ;
        RECT 616.950 885.600 619.050 886.050 ;
        RECT 601.950 884.400 619.050 885.600 ;
        RECT 601.950 883.950 604.050 884.400 ;
        RECT 616.950 883.950 619.050 884.400 ;
        RECT 622.950 883.950 625.050 886.050 ;
        RECT 640.950 883.950 643.050 886.050 ;
        RECT 646.950 885.600 649.050 886.050 ;
        RECT 718.950 885.600 721.050 886.050 ;
        RECT 646.950 884.400 721.050 885.600 ;
        RECT 646.950 883.950 649.050 884.400 ;
        RECT 718.950 883.950 721.050 884.400 ;
        RECT 739.950 885.600 742.050 886.050 ;
        RECT 805.950 885.600 808.050 886.050 ;
        RECT 739.950 884.400 808.050 885.600 ;
        RECT 739.950 883.950 742.050 884.400 ;
        RECT 805.950 883.950 808.050 884.400 ;
        RECT 847.950 885.600 850.050 886.050 ;
        RECT 859.950 885.600 862.050 886.050 ;
        RECT 847.950 884.400 862.050 885.600 ;
        RECT 847.950 883.950 850.050 884.400 ;
        RECT 859.950 883.950 862.050 884.400 ;
        RECT 268.950 882.600 271.050 883.050 ;
        RECT 197.400 881.400 271.050 882.600 ;
        RECT 178.950 880.950 181.050 881.400 ;
        RECT 187.950 880.950 190.050 881.400 ;
        RECT 268.950 880.950 271.050 881.400 ;
        RECT 283.950 882.600 286.050 883.050 ;
        RECT 340.950 882.600 343.050 883.050 ;
        RECT 370.950 882.600 373.050 883.050 ;
        RECT 283.950 881.400 373.050 882.600 ;
        RECT 283.950 880.950 286.050 881.400 ;
        RECT 340.950 880.950 343.050 881.400 ;
        RECT 370.950 880.950 373.050 881.400 ;
        RECT 442.950 882.600 445.050 883.050 ;
        RECT 454.950 882.600 457.050 883.050 ;
        RECT 442.950 881.400 457.050 882.600 ;
        RECT 442.950 880.950 445.050 881.400 ;
        RECT 454.950 880.950 457.050 881.400 ;
        RECT 460.950 882.600 463.050 883.050 ;
        RECT 481.950 882.600 484.050 883.050 ;
        RECT 460.950 881.400 484.050 882.600 ;
        RECT 460.950 880.950 463.050 881.400 ;
        RECT 481.950 880.950 484.050 881.400 ;
        RECT 553.950 882.600 556.050 883.050 ;
        RECT 586.950 882.600 589.050 883.050 ;
        RECT 553.950 881.400 589.050 882.600 ;
        RECT 623.400 882.600 624.600 883.950 ;
        RECT 664.950 882.600 667.050 883.050 ;
        RECT 623.400 881.400 667.050 882.600 ;
        RECT 553.950 880.950 556.050 881.400 ;
        RECT 586.950 880.950 589.050 881.400 ;
        RECT 664.950 880.950 667.050 881.400 ;
        RECT 703.950 882.600 706.050 883.050 ;
        RECT 715.950 882.600 718.050 883.050 ;
        RECT 736.950 882.600 739.050 883.050 ;
        RECT 703.950 881.400 739.050 882.600 ;
        RECT 703.950 880.950 706.050 881.400 ;
        RECT 715.950 880.950 718.050 881.400 ;
        RECT 736.950 880.950 739.050 881.400 ;
        RECT 742.950 882.600 745.050 883.050 ;
        RECT 769.950 882.600 772.050 883.050 ;
        RECT 778.950 882.600 781.050 883.050 ;
        RECT 742.950 881.400 781.050 882.600 ;
        RECT 742.950 880.950 745.050 881.400 ;
        RECT 769.950 880.950 772.050 881.400 ;
        RECT 778.950 880.950 781.050 881.400 ;
        RECT 832.950 882.600 835.050 883.050 ;
        RECT 844.950 882.600 847.050 883.050 ;
        RECT 832.950 881.400 847.050 882.600 ;
        RECT 832.950 880.950 835.050 881.400 ;
        RECT 844.950 880.950 847.050 881.400 ;
        RECT 850.950 882.600 853.050 883.050 ;
        RECT 865.950 882.600 868.050 883.050 ;
        RECT 850.950 881.400 868.050 882.600 ;
        RECT 850.950 880.950 853.050 881.400 ;
        RECT 865.950 880.950 868.050 881.400 ;
        RECT 100.950 879.600 103.050 880.050 ;
        RECT 196.950 879.600 199.050 880.050 ;
        RECT 100.950 878.400 199.050 879.600 ;
        RECT 100.950 877.950 103.050 878.400 ;
        RECT 196.950 877.950 199.050 878.400 ;
        RECT 226.950 879.600 229.050 880.050 ;
        RECT 304.950 879.600 307.050 880.050 ;
        RECT 226.950 878.400 307.050 879.600 ;
        RECT 226.950 877.950 229.050 878.400 ;
        RECT 304.950 877.950 307.050 878.400 ;
        RECT 571.950 879.600 574.050 880.050 ;
        RECT 607.950 879.600 610.050 880.050 ;
        RECT 571.950 878.400 610.050 879.600 ;
        RECT 571.950 877.950 574.050 878.400 ;
        RECT 607.950 877.950 610.050 878.400 ;
        RECT 106.950 870.600 109.050 871.050 ;
        RECT 199.950 870.600 202.050 871.050 ;
        RECT 106.950 869.400 202.050 870.600 ;
        RECT 106.950 868.950 109.050 869.400 ;
        RECT 199.950 868.950 202.050 869.400 ;
        RECT 202.950 870.600 205.050 871.050 ;
        RECT 208.950 870.600 211.050 871.050 ;
        RECT 202.950 869.400 211.050 870.600 ;
        RECT 202.950 868.950 205.050 869.400 ;
        RECT 208.950 868.950 211.050 869.400 ;
        RECT 127.950 867.600 130.050 868.050 ;
        RECT 178.950 867.600 181.050 868.050 ;
        RECT 127.950 866.400 181.050 867.600 ;
        RECT 127.950 865.950 130.050 866.400 ;
        RECT 178.950 865.950 181.050 866.400 ;
        RECT 520.950 864.600 523.050 865.050 ;
        RECT 565.950 864.600 568.050 865.050 ;
        RECT 520.950 863.400 568.050 864.600 ;
        RECT 520.950 862.950 523.050 863.400 ;
        RECT 565.950 862.950 568.050 863.400 ;
        RECT 715.950 864.600 718.050 865.050 ;
        RECT 721.950 864.600 724.050 865.050 ;
        RECT 715.950 863.400 724.050 864.600 ;
        RECT 715.950 862.950 718.050 863.400 ;
        RECT 721.950 862.950 724.050 863.400 ;
        RECT 511.950 861.600 514.050 862.050 ;
        RECT 538.950 861.600 541.050 862.050 ;
        RECT 511.950 860.400 541.050 861.600 ;
        RECT 511.950 859.950 514.050 860.400 ;
        RECT 538.950 859.950 541.050 860.400 ;
        RECT 541.950 858.600 544.050 859.050 ;
        RECT 643.950 858.600 646.050 859.050 ;
        RECT 673.950 858.600 676.050 859.050 ;
        RECT 541.950 857.400 676.050 858.600 ;
        RECT 541.950 856.950 544.050 857.400 ;
        RECT 643.950 856.950 646.050 857.400 ;
        RECT 673.950 856.950 676.050 857.400 ;
        RECT 214.950 855.600 217.050 856.050 ;
        RECT 298.950 855.600 301.050 856.050 ;
        RECT 214.950 854.400 301.050 855.600 ;
        RECT 214.950 853.950 217.050 854.400 ;
        RECT 298.950 853.950 301.050 854.400 ;
        RECT 454.950 855.600 457.050 856.050 ;
        RECT 574.950 855.600 577.050 856.050 ;
        RECT 454.950 854.400 577.050 855.600 ;
        RECT 454.950 853.950 457.050 854.400 ;
        RECT 574.950 853.950 577.050 854.400 ;
        RECT 589.950 855.600 592.050 856.050 ;
        RECT 817.950 855.600 820.050 856.050 ;
        RECT 589.950 854.400 820.050 855.600 ;
        RECT 589.950 853.950 592.050 854.400 ;
        RECT 817.950 853.950 820.050 854.400 ;
        RECT 40.950 852.600 43.050 853.050 ;
        RECT 61.950 852.600 64.050 853.050 ;
        RECT 40.950 851.400 64.050 852.600 ;
        RECT 40.950 850.950 43.050 851.400 ;
        RECT 61.950 850.950 64.050 851.400 ;
        RECT 91.950 852.600 94.050 853.050 ;
        RECT 124.950 852.600 127.050 853.050 ;
        RECT 91.950 851.400 127.050 852.600 ;
        RECT 91.950 850.950 94.050 851.400 ;
        RECT 124.950 850.950 127.050 851.400 ;
        RECT 142.950 852.600 145.050 853.050 ;
        RECT 226.950 852.600 229.050 853.050 ;
        RECT 142.950 851.400 229.050 852.600 ;
        RECT 142.950 850.950 145.050 851.400 ;
        RECT 226.950 850.950 229.050 851.400 ;
        RECT 238.950 852.600 241.050 853.050 ;
        RECT 358.950 852.600 361.050 853.050 ;
        RECT 481.950 852.600 484.050 853.050 ;
        RECT 532.950 852.600 535.050 853.050 ;
        RECT 238.950 851.400 535.050 852.600 ;
        RECT 238.950 850.950 241.050 851.400 ;
        RECT 358.950 850.950 361.050 851.400 ;
        RECT 481.950 850.950 484.050 851.400 ;
        RECT 532.950 850.950 535.050 851.400 ;
        RECT 568.950 852.600 571.050 853.050 ;
        RECT 724.950 852.600 727.050 853.050 ;
        RECT 568.950 851.400 727.050 852.600 ;
        RECT 568.950 850.950 571.050 851.400 ;
        RECT 724.950 850.950 727.050 851.400 ;
        RECT 820.950 852.600 823.050 853.050 ;
        RECT 832.950 852.600 835.050 853.050 ;
        RECT 820.950 851.400 835.050 852.600 ;
        RECT 820.950 850.950 823.050 851.400 ;
        RECT 832.950 850.950 835.050 851.400 ;
        RECT 34.950 849.600 37.050 850.050 ;
        RECT 82.950 849.600 85.050 850.050 ;
        RECT 97.950 849.600 100.050 850.050 ;
        RECT 34.950 848.400 63.600 849.600 ;
        RECT 34.950 847.950 37.050 848.400 ;
        RECT 13.950 846.600 16.050 847.050 ;
        RECT 43.950 846.600 46.050 847.050 ;
        RECT 62.400 846.600 63.600 848.400 ;
        RECT 82.950 848.400 100.050 849.600 ;
        RECT 82.950 847.950 85.050 848.400 ;
        RECT 97.950 847.950 100.050 848.400 ;
        RECT 118.950 847.950 121.050 850.050 ;
        RECT 136.950 849.600 139.050 850.050 ;
        RECT 232.950 849.600 235.050 850.050 ;
        RECT 352.950 849.600 355.050 850.050 ;
        RECT 136.950 848.400 355.050 849.600 ;
        RECT 136.950 847.950 139.050 848.400 ;
        RECT 232.950 847.950 235.050 848.400 ;
        RECT 352.950 847.950 355.050 848.400 ;
        RECT 376.950 849.600 379.050 850.050 ;
        RECT 385.950 849.600 388.050 850.050 ;
        RECT 376.950 848.400 388.050 849.600 ;
        RECT 376.950 847.950 379.050 848.400 ;
        RECT 385.950 847.950 388.050 848.400 ;
        RECT 475.950 849.600 478.050 850.050 ;
        RECT 526.950 849.600 529.050 850.050 ;
        RECT 475.950 848.400 529.050 849.600 ;
        RECT 475.950 847.950 478.050 848.400 ;
        RECT 526.950 847.950 529.050 848.400 ;
        RECT 532.950 849.600 535.050 850.050 ;
        RECT 562.950 849.600 565.050 850.050 ;
        RECT 532.950 848.400 565.050 849.600 ;
        RECT 532.950 847.950 535.050 848.400 ;
        RECT 562.950 847.950 565.050 848.400 ;
        RECT 565.950 849.600 568.050 850.050 ;
        RECT 592.950 849.600 595.050 850.050 ;
        RECT 565.950 848.400 595.050 849.600 ;
        RECT 565.950 847.950 568.050 848.400 ;
        RECT 592.950 847.950 595.050 848.400 ;
        RECT 703.950 849.600 706.050 850.050 ;
        RECT 715.950 849.600 718.050 850.050 ;
        RECT 703.950 848.400 718.050 849.600 ;
        RECT 703.950 847.950 706.050 848.400 ;
        RECT 715.950 847.950 718.050 848.400 ;
        RECT 721.950 849.600 724.050 850.050 ;
        RECT 754.950 849.600 757.050 850.050 ;
        RECT 772.950 849.600 775.050 850.050 ;
        RECT 721.950 848.400 775.050 849.600 ;
        RECT 721.950 847.950 724.050 848.400 ;
        RECT 754.950 847.950 757.050 848.400 ;
        RECT 772.950 847.950 775.050 848.400 ;
        RECT 787.950 849.600 790.050 850.050 ;
        RECT 796.950 849.600 799.050 850.050 ;
        RECT 787.950 848.400 799.050 849.600 ;
        RECT 787.950 847.950 790.050 848.400 ;
        RECT 796.950 847.950 799.050 848.400 ;
        RECT 826.950 849.600 829.050 850.050 ;
        RECT 841.950 849.600 844.050 850.050 ;
        RECT 826.950 848.400 844.050 849.600 ;
        RECT 826.950 847.950 829.050 848.400 ;
        RECT 841.950 847.950 844.050 848.400 ;
        RECT 67.950 846.600 70.050 847.050 ;
        RECT 13.950 845.400 30.600 846.600 ;
        RECT 13.950 844.950 16.050 845.400 ;
        RECT 29.400 844.050 30.600 845.400 ;
        RECT 43.950 845.400 60.600 846.600 ;
        RECT 62.400 845.400 70.050 846.600 ;
        RECT 43.950 844.950 46.050 845.400 ;
        RECT 59.400 844.050 60.600 845.400 ;
        RECT 67.950 844.950 70.050 845.400 ;
        RECT 100.950 846.600 103.050 847.050 ;
        RECT 119.400 846.600 120.600 847.950 ;
        RECT 100.950 845.400 120.600 846.600 ;
        RECT 121.950 846.600 124.050 847.050 ;
        RECT 142.950 846.600 145.050 847.050 ;
        RECT 172.950 846.600 175.050 847.050 ;
        RECT 121.950 845.400 145.050 846.600 ;
        RECT 100.950 844.950 103.050 845.400 ;
        RECT 121.950 844.950 124.050 845.400 ;
        RECT 142.950 844.950 145.050 845.400 ;
        RECT 146.400 845.400 175.050 846.600 ;
        RECT 28.950 841.950 31.050 844.050 ;
        RECT 58.950 841.950 61.050 844.050 ;
        RECT 64.950 843.600 67.050 844.050 ;
        RECT 146.400 843.600 147.600 845.400 ;
        RECT 172.950 844.950 175.050 845.400 ;
        RECT 178.950 846.600 181.050 847.050 ;
        RECT 184.950 846.600 187.050 847.050 ;
        RECT 178.950 845.400 187.050 846.600 ;
        RECT 178.950 844.950 181.050 845.400 ;
        RECT 184.950 844.950 187.050 845.400 ;
        RECT 199.950 846.600 202.050 847.050 ;
        RECT 238.950 846.600 241.050 847.050 ;
        RECT 199.950 845.400 241.050 846.600 ;
        RECT 199.950 844.950 202.050 845.400 ;
        RECT 238.950 844.950 241.050 845.400 ;
        RECT 244.950 846.600 247.050 847.050 ;
        RECT 280.950 846.600 283.050 847.050 ;
        RECT 289.950 846.600 292.050 847.050 ;
        RECT 244.950 845.400 292.050 846.600 ;
        RECT 244.950 844.950 247.050 845.400 ;
        RECT 280.950 844.950 283.050 845.400 ;
        RECT 289.950 844.950 292.050 845.400 ;
        RECT 364.950 846.600 367.050 847.050 ;
        RECT 373.950 846.600 376.050 847.050 ;
        RECT 364.950 845.400 376.050 846.600 ;
        RECT 364.950 844.950 367.050 845.400 ;
        RECT 373.950 844.950 376.050 845.400 ;
        RECT 382.950 846.600 385.050 847.050 ;
        RECT 427.950 846.600 430.050 847.050 ;
        RECT 382.950 845.400 430.050 846.600 ;
        RECT 382.950 844.950 385.050 845.400 ;
        RECT 427.950 844.950 430.050 845.400 ;
        RECT 505.950 846.600 508.050 847.050 ;
        RECT 541.950 846.600 544.050 847.050 ;
        RECT 547.950 846.600 550.050 847.050 ;
        RECT 505.950 845.400 525.600 846.600 ;
        RECT 505.950 844.950 508.050 845.400 ;
        RECT 524.400 844.050 525.600 845.400 ;
        RECT 541.950 845.400 550.050 846.600 ;
        RECT 541.950 844.950 544.050 845.400 ;
        RECT 547.950 844.950 550.050 845.400 ;
        RECT 553.950 846.600 556.050 847.050 ;
        RECT 571.950 846.600 574.050 847.050 ;
        RECT 610.950 846.600 613.050 847.050 ;
        RECT 553.950 845.400 574.050 846.600 ;
        RECT 553.950 844.950 556.050 845.400 ;
        RECT 571.950 844.950 574.050 845.400 ;
        RECT 593.400 845.400 613.050 846.600 ;
        RECT 593.400 844.050 594.600 845.400 ;
        RECT 610.950 844.950 613.050 845.400 ;
        RECT 616.950 846.600 619.050 847.050 ;
        RECT 634.950 846.600 637.050 847.050 ;
        RECT 616.950 845.400 637.050 846.600 ;
        RECT 616.950 844.950 619.050 845.400 ;
        RECT 634.950 844.950 637.050 845.400 ;
        RECT 664.950 846.600 667.050 847.050 ;
        RECT 679.950 846.600 682.050 847.050 ;
        RECT 664.950 845.400 682.050 846.600 ;
        RECT 664.950 844.950 667.050 845.400 ;
        RECT 679.950 844.950 682.050 845.400 ;
        RECT 694.950 844.950 697.050 847.050 ;
        RECT 700.950 846.600 703.050 847.050 ;
        RECT 718.950 846.600 721.050 847.050 ;
        RECT 700.950 845.400 721.050 846.600 ;
        RECT 700.950 844.950 703.050 845.400 ;
        RECT 718.950 844.950 721.050 845.400 ;
        RECT 775.950 846.600 778.050 847.050 ;
        RECT 790.950 846.600 793.050 847.050 ;
        RECT 775.950 845.400 793.050 846.600 ;
        RECT 775.950 844.950 778.050 845.400 ;
        RECT 790.950 844.950 793.050 845.400 ;
        RECT 829.950 846.600 832.050 847.050 ;
        RECT 835.950 846.600 838.050 847.050 ;
        RECT 829.950 845.400 838.050 846.600 ;
        RECT 829.950 844.950 832.050 845.400 ;
        RECT 835.950 844.950 838.050 845.400 ;
        RECT 64.950 842.400 147.600 843.600 ;
        RECT 148.950 843.600 151.050 844.050 ;
        RECT 172.950 843.600 175.050 844.050 ;
        RECT 148.950 842.400 175.050 843.600 ;
        RECT 64.950 841.950 67.050 842.400 ;
        RECT 148.950 841.950 151.050 842.400 ;
        RECT 172.950 841.950 175.050 842.400 ;
        RECT 175.950 843.600 178.050 844.050 ;
        RECT 196.950 843.600 199.050 844.050 ;
        RECT 175.950 842.400 199.050 843.600 ;
        RECT 175.950 841.950 178.050 842.400 ;
        RECT 196.950 841.950 199.050 842.400 ;
        RECT 214.950 843.600 217.050 844.050 ;
        RECT 220.950 843.600 223.050 844.050 ;
        RECT 214.950 842.400 223.050 843.600 ;
        RECT 214.950 841.950 217.050 842.400 ;
        RECT 220.950 841.950 223.050 842.400 ;
        RECT 235.950 843.600 238.050 844.050 ;
        RECT 256.950 843.600 259.050 844.050 ;
        RECT 235.950 842.400 259.050 843.600 ;
        RECT 235.950 841.950 238.050 842.400 ;
        RECT 256.950 841.950 259.050 842.400 ;
        RECT 274.950 843.600 277.050 844.050 ;
        RECT 283.950 843.600 286.050 844.050 ;
        RECT 274.950 842.400 286.050 843.600 ;
        RECT 274.950 841.950 277.050 842.400 ;
        RECT 283.950 841.950 286.050 842.400 ;
        RECT 337.950 843.600 340.050 844.050 ;
        RECT 349.950 843.600 352.050 844.050 ;
        RECT 337.950 842.400 352.050 843.600 ;
        RECT 337.950 841.950 340.050 842.400 ;
        RECT 349.950 841.950 352.050 842.400 ;
        RECT 355.950 843.600 358.050 844.050 ;
        RECT 394.950 843.600 397.050 844.050 ;
        RECT 355.950 842.400 397.050 843.600 ;
        RECT 355.950 841.950 358.050 842.400 ;
        RECT 394.950 841.950 397.050 842.400 ;
        RECT 412.950 843.600 415.050 844.050 ;
        RECT 421.950 843.600 424.050 844.050 ;
        RECT 412.950 842.400 424.050 843.600 ;
        RECT 412.950 841.950 415.050 842.400 ;
        RECT 421.950 841.950 424.050 842.400 ;
        RECT 442.950 843.600 445.050 844.050 ;
        RECT 463.950 843.600 466.050 844.050 ;
        RECT 442.950 842.400 466.050 843.600 ;
        RECT 442.950 841.950 445.050 842.400 ;
        RECT 463.950 841.950 466.050 842.400 ;
        RECT 523.950 841.950 526.050 844.050 ;
        RECT 535.950 843.600 538.050 844.050 ;
        RECT 538.950 843.600 541.050 844.050 ;
        RECT 544.950 843.600 547.050 844.050 ;
        RECT 535.950 842.400 547.050 843.600 ;
        RECT 535.950 841.950 538.050 842.400 ;
        RECT 538.950 841.950 541.050 842.400 ;
        RECT 544.950 841.950 547.050 842.400 ;
        RECT 550.950 843.600 553.050 844.050 ;
        RECT 589.950 843.600 592.050 844.050 ;
        RECT 550.950 842.400 592.050 843.600 ;
        RECT 550.950 841.950 553.050 842.400 ;
        RECT 589.950 841.950 592.050 842.400 ;
        RECT 592.950 841.950 595.050 844.050 ;
        RECT 655.950 843.600 658.050 844.050 ;
        RECT 695.400 843.600 696.600 844.950 ;
        RECT 655.950 842.400 696.600 843.600 ;
        RECT 697.950 843.600 700.050 844.050 ;
        RECT 736.950 843.600 739.050 844.050 ;
        RECT 697.950 842.400 739.050 843.600 ;
        RECT 655.950 841.950 658.050 842.400 ;
        RECT 697.950 841.950 700.050 842.400 ;
        RECT 736.950 841.950 739.050 842.400 ;
        RECT 757.950 843.600 760.050 844.050 ;
        RECT 781.950 843.600 784.050 844.050 ;
        RECT 799.950 843.600 802.050 844.050 ;
        RECT 757.950 842.400 802.050 843.600 ;
        RECT 757.950 841.950 760.050 842.400 ;
        RECT 781.950 841.950 784.050 842.400 ;
        RECT 799.950 841.950 802.050 842.400 ;
        RECT 823.950 843.600 826.050 844.050 ;
        RECT 850.950 843.600 853.050 844.050 ;
        RECT 823.950 842.400 853.050 843.600 ;
        RECT 823.950 841.950 826.050 842.400 ;
        RECT 850.950 841.950 853.050 842.400 ;
        RECT 100.950 840.600 103.050 841.050 ;
        RECT 106.950 840.600 109.050 841.050 ;
        RECT 100.950 839.400 109.050 840.600 ;
        RECT 100.950 838.950 103.050 839.400 ;
        RECT 106.950 838.950 109.050 839.400 ;
        RECT 145.950 840.600 148.050 841.050 ;
        RECT 151.950 840.600 154.050 841.050 ;
        RECT 202.950 840.600 205.050 841.050 ;
        RECT 259.950 840.600 262.050 841.050 ;
        RECT 145.950 839.400 262.050 840.600 ;
        RECT 145.950 838.950 148.050 839.400 ;
        RECT 151.950 838.950 154.050 839.400 ;
        RECT 202.950 838.950 205.050 839.400 ;
        RECT 259.950 838.950 262.050 839.400 ;
        RECT 304.950 840.600 307.050 841.050 ;
        RECT 319.950 840.600 322.050 841.050 ;
        RECT 400.950 840.600 403.050 841.050 ;
        RECT 433.950 840.600 436.050 841.050 ;
        RECT 451.950 840.600 454.050 841.050 ;
        RECT 304.950 839.400 454.050 840.600 ;
        RECT 304.950 838.950 307.050 839.400 ;
        RECT 319.950 838.950 322.050 839.400 ;
        RECT 400.950 838.950 403.050 839.400 ;
        RECT 433.950 838.950 436.050 839.400 ;
        RECT 451.950 838.950 454.050 839.400 ;
        RECT 487.950 840.600 490.050 841.050 ;
        RECT 490.950 840.600 493.050 841.050 ;
        RECT 496.950 840.600 499.050 841.050 ;
        RECT 487.950 839.400 499.050 840.600 ;
        RECT 487.950 838.950 490.050 839.400 ;
        RECT 490.950 838.950 493.050 839.400 ;
        RECT 496.950 838.950 499.050 839.400 ;
        RECT 502.950 840.600 505.050 841.050 ;
        RECT 529.950 840.600 532.050 841.050 ;
        RECT 502.950 839.400 532.050 840.600 ;
        RECT 502.950 838.950 505.050 839.400 ;
        RECT 529.950 838.950 532.050 839.400 ;
        RECT 595.950 840.600 598.050 841.050 ;
        RECT 607.950 840.600 610.050 841.050 ;
        RECT 625.950 840.600 628.050 841.050 ;
        RECT 595.950 839.400 628.050 840.600 ;
        RECT 595.950 838.950 598.050 839.400 ;
        RECT 607.950 838.950 610.050 839.400 ;
        RECT 625.950 838.950 628.050 839.400 ;
        RECT 676.950 840.600 679.050 841.050 ;
        RECT 691.950 840.600 694.050 841.050 ;
        RECT 676.950 839.400 694.050 840.600 ;
        RECT 676.950 838.950 679.050 839.400 ;
        RECT 691.950 838.950 694.050 839.400 ;
        RECT 793.950 840.600 796.050 841.050 ;
        RECT 814.950 840.600 817.050 841.050 ;
        RECT 793.950 839.400 817.050 840.600 ;
        RECT 793.950 838.950 796.050 839.400 ;
        RECT 814.950 838.950 817.050 839.400 ;
        RECT 820.950 840.600 823.050 841.050 ;
        RECT 826.950 840.600 829.050 841.050 ;
        RECT 820.950 839.400 829.050 840.600 ;
        RECT 820.950 838.950 823.050 839.400 ;
        RECT 826.950 838.950 829.050 839.400 ;
        RECT 841.950 840.600 844.050 841.050 ;
        RECT 856.950 840.600 859.050 841.050 ;
        RECT 841.950 839.400 859.050 840.600 ;
        RECT 841.950 838.950 844.050 839.400 ;
        RECT 856.950 838.950 859.050 839.400 ;
        RECT 16.950 837.600 19.050 838.050 ;
        RECT 22.950 837.600 25.050 838.050 ;
        RECT 16.950 836.400 25.050 837.600 ;
        RECT 16.950 835.950 19.050 836.400 ;
        RECT 22.950 835.950 25.050 836.400 ;
        RECT 139.950 837.600 142.050 838.050 ;
        RECT 145.950 837.600 148.050 838.050 ;
        RECT 139.950 836.400 148.050 837.600 ;
        RECT 139.950 835.950 142.050 836.400 ;
        RECT 145.950 835.950 148.050 836.400 ;
        RECT 178.950 837.600 181.050 838.050 ;
        RECT 187.950 837.600 190.050 838.050 ;
        RECT 343.950 837.600 346.050 838.050 ;
        RECT 178.950 836.400 346.050 837.600 ;
        RECT 178.950 835.950 181.050 836.400 ;
        RECT 187.950 835.950 190.050 836.400 ;
        RECT 343.950 835.950 346.050 836.400 ;
        RECT 484.950 837.600 487.050 838.050 ;
        RECT 499.950 837.600 502.050 838.050 ;
        RECT 484.950 836.400 502.050 837.600 ;
        RECT 484.950 835.950 487.050 836.400 ;
        RECT 499.950 835.950 502.050 836.400 ;
        RECT 541.950 837.600 544.050 838.050 ;
        RECT 790.950 837.600 793.050 838.050 ;
        RECT 541.950 836.400 793.050 837.600 ;
        RECT 541.950 835.950 544.050 836.400 ;
        RECT 790.950 835.950 793.050 836.400 ;
        RECT 208.950 834.600 211.050 835.050 ;
        RECT 232.950 834.600 235.050 835.050 ;
        RECT 262.950 834.600 265.050 835.050 ;
        RECT 286.950 834.600 289.050 835.050 ;
        RECT 757.950 834.600 760.050 835.050 ;
        RECT 208.950 833.400 760.050 834.600 ;
        RECT 208.950 832.950 211.050 833.400 ;
        RECT 232.950 832.950 235.050 833.400 ;
        RECT 262.950 832.950 265.050 833.400 ;
        RECT 286.950 832.950 289.050 833.400 ;
        RECT 757.950 832.950 760.050 833.400 ;
        RECT 814.950 834.600 817.050 835.050 ;
        RECT 868.950 834.600 871.050 835.050 ;
        RECT 814.950 833.400 871.050 834.600 ;
        RECT 814.950 832.950 817.050 833.400 ;
        RECT 868.950 832.950 871.050 833.400 ;
        RECT 394.950 831.600 397.050 832.050 ;
        RECT 676.950 831.600 679.050 832.050 ;
        RECT 394.950 830.400 679.050 831.600 ;
        RECT 394.950 829.950 397.050 830.400 ;
        RECT 676.950 829.950 679.050 830.400 ;
        RECT 292.950 828.600 295.050 829.050 ;
        RECT 418.950 828.600 421.050 829.050 ;
        RECT 292.950 827.400 421.050 828.600 ;
        RECT 292.950 826.950 295.050 827.400 ;
        RECT 418.950 826.950 421.050 827.400 ;
        RECT 742.950 828.600 745.050 829.050 ;
        RECT 754.950 828.600 757.050 829.050 ;
        RECT 784.950 828.600 787.050 829.050 ;
        RECT 853.950 828.600 856.050 829.050 ;
        RECT 862.950 828.600 865.050 829.050 ;
        RECT 742.950 827.400 865.050 828.600 ;
        RECT 742.950 826.950 745.050 827.400 ;
        RECT 754.950 826.950 757.050 827.400 ;
        RECT 784.950 826.950 787.050 827.400 ;
        RECT 853.950 826.950 856.050 827.400 ;
        RECT 862.950 826.950 865.050 827.400 ;
        RECT 253.950 825.600 256.050 826.050 ;
        RECT 367.950 825.600 370.050 826.050 ;
        RECT 253.950 824.400 370.050 825.600 ;
        RECT 253.950 823.950 256.050 824.400 ;
        RECT 367.950 823.950 370.050 824.400 ;
        RECT 427.950 825.600 430.050 826.050 ;
        RECT 445.950 825.600 448.050 826.050 ;
        RECT 427.950 824.400 448.050 825.600 ;
        RECT 427.950 823.950 430.050 824.400 ;
        RECT 445.950 823.950 448.050 824.400 ;
        RECT 493.950 825.600 496.050 826.050 ;
        RECT 520.950 825.600 523.050 826.050 ;
        RECT 628.950 825.600 631.050 826.050 ;
        RECT 649.950 825.600 652.050 826.050 ;
        RECT 670.950 825.600 673.050 826.050 ;
        RECT 493.950 824.400 673.050 825.600 ;
        RECT 493.950 823.950 496.050 824.400 ;
        RECT 520.950 823.950 523.050 824.400 ;
        RECT 628.950 823.950 631.050 824.400 ;
        RECT 649.950 823.950 652.050 824.400 ;
        RECT 670.950 823.950 673.050 824.400 ;
        RECT 682.950 825.600 685.050 826.050 ;
        RECT 844.950 825.600 847.050 826.050 ;
        RECT 682.950 824.400 847.050 825.600 ;
        RECT 682.950 823.950 685.050 824.400 ;
        RECT 844.950 823.950 847.050 824.400 ;
        RECT 16.950 822.600 19.050 823.050 ;
        RECT 88.950 822.600 91.050 823.050 ;
        RECT 97.950 822.600 100.050 823.050 ;
        RECT 16.950 821.400 100.050 822.600 ;
        RECT 16.950 820.950 19.050 821.400 ;
        RECT 88.950 820.950 91.050 821.400 ;
        RECT 97.950 820.950 100.050 821.400 ;
        RECT 355.950 822.600 358.050 823.050 ;
        RECT 379.950 822.600 382.050 823.050 ;
        RECT 715.950 822.600 718.050 823.050 ;
        RECT 808.950 822.600 811.050 823.050 ;
        RECT 811.950 822.600 814.050 823.050 ;
        RECT 817.950 822.600 820.050 823.050 ;
        RECT 355.950 821.400 718.050 822.600 ;
        RECT 355.950 820.950 358.050 821.400 ;
        RECT 379.950 820.950 382.050 821.400 ;
        RECT 715.950 820.950 718.050 821.400 ;
        RECT 719.400 821.400 798.600 822.600 ;
        RECT 37.950 819.600 40.050 820.050 ;
        RECT 58.950 819.600 61.050 820.050 ;
        RECT 64.950 819.600 67.050 820.050 ;
        RECT 37.950 818.400 67.050 819.600 ;
        RECT 37.950 817.950 40.050 818.400 ;
        RECT 58.950 817.950 61.050 818.400 ;
        RECT 64.950 817.950 67.050 818.400 ;
        RECT 82.950 819.600 85.050 820.050 ;
        RECT 91.950 819.600 94.050 820.050 ;
        RECT 82.950 818.400 94.050 819.600 ;
        RECT 82.950 817.950 85.050 818.400 ;
        RECT 91.950 817.950 94.050 818.400 ;
        RECT 160.950 819.600 163.050 820.050 ;
        RECT 190.950 819.600 193.050 820.050 ;
        RECT 160.950 818.400 193.050 819.600 ;
        RECT 160.950 817.950 163.050 818.400 ;
        RECT 190.950 817.950 193.050 818.400 ;
        RECT 211.950 819.600 214.050 820.050 ;
        RECT 220.950 819.600 223.050 820.050 ;
        RECT 211.950 818.400 223.050 819.600 ;
        RECT 211.950 817.950 214.050 818.400 ;
        RECT 220.950 817.950 223.050 818.400 ;
        RECT 361.950 819.600 364.050 820.050 ;
        RECT 382.950 819.600 385.050 820.050 ;
        RECT 361.950 818.400 385.050 819.600 ;
        RECT 361.950 817.950 364.050 818.400 ;
        RECT 382.950 817.950 385.050 818.400 ;
        RECT 391.950 819.600 394.050 820.050 ;
        RECT 400.950 819.600 403.050 820.050 ;
        RECT 391.950 818.400 403.050 819.600 ;
        RECT 391.950 817.950 394.050 818.400 ;
        RECT 400.950 817.950 403.050 818.400 ;
        RECT 406.950 819.600 409.050 820.050 ;
        RECT 541.950 819.600 544.050 820.050 ;
        RECT 406.950 818.400 544.050 819.600 ;
        RECT 406.950 817.950 409.050 818.400 ;
        RECT 541.950 817.950 544.050 818.400 ;
        RECT 598.950 819.600 601.050 820.050 ;
        RECT 634.950 819.600 637.050 820.050 ;
        RECT 598.950 818.400 637.050 819.600 ;
        RECT 598.950 817.950 601.050 818.400 ;
        RECT 13.950 816.600 16.050 817.050 ;
        RECT 28.950 816.600 31.050 817.050 ;
        RECT 34.950 816.600 37.050 817.050 ;
        RECT 13.950 815.400 37.050 816.600 ;
        RECT 13.950 814.950 16.050 815.400 ;
        RECT 28.950 814.950 31.050 815.400 ;
        RECT 34.950 814.950 37.050 815.400 ;
        RECT 103.950 814.950 106.050 817.050 ;
        RECT 133.950 816.600 136.050 817.050 ;
        RECT 139.950 816.600 142.050 817.050 ;
        RECT 133.950 815.400 142.050 816.600 ;
        RECT 133.950 814.950 136.050 815.400 ;
        RECT 139.950 814.950 142.050 815.400 ;
        RECT 157.950 816.600 160.050 817.050 ;
        RECT 166.950 816.600 169.050 817.050 ;
        RECT 157.950 815.400 169.050 816.600 ;
        RECT 157.950 814.950 160.050 815.400 ;
        RECT 166.950 814.950 169.050 815.400 ;
        RECT 268.950 816.600 271.050 817.050 ;
        RECT 298.950 816.600 301.050 817.050 ;
        RECT 268.950 815.400 301.050 816.600 ;
        RECT 268.950 814.950 271.050 815.400 ;
        RECT 298.950 814.950 301.050 815.400 ;
        RECT 316.950 816.600 319.050 817.050 ;
        RECT 325.950 816.600 328.050 817.050 ;
        RECT 316.950 815.400 328.050 816.600 ;
        RECT 316.950 814.950 319.050 815.400 ;
        RECT 325.950 814.950 328.050 815.400 ;
        RECT 349.950 816.600 352.050 817.050 ;
        RECT 361.950 816.600 364.050 817.050 ;
        RECT 349.950 815.400 364.050 816.600 ;
        RECT 349.950 814.950 352.050 815.400 ;
        RECT 361.950 814.950 364.050 815.400 ;
        RECT 373.950 816.600 376.050 817.050 ;
        RECT 424.950 816.600 427.050 817.050 ;
        RECT 472.950 816.600 475.050 817.050 ;
        RECT 373.950 815.400 423.600 816.600 ;
        RECT 373.950 814.950 376.050 815.400 ;
        RECT 19.950 813.600 22.050 814.050 ;
        RECT 31.950 813.600 34.050 814.050 ;
        RECT 19.950 812.400 34.050 813.600 ;
        RECT 19.950 811.950 22.050 812.400 ;
        RECT 31.950 811.950 34.050 812.400 ;
        RECT 49.950 813.600 52.050 814.050 ;
        RECT 61.950 813.600 64.050 814.050 ;
        RECT 49.950 812.400 64.050 813.600 ;
        RECT 49.950 811.950 52.050 812.400 ;
        RECT 61.950 811.950 64.050 812.400 ;
        RECT 85.950 813.600 88.050 814.050 ;
        RECT 104.400 813.600 105.600 814.950 ;
        RECT 422.400 814.050 423.600 815.400 ;
        RECT 424.950 815.400 475.050 816.600 ;
        RECT 424.950 814.950 427.050 815.400 ;
        RECT 472.950 814.950 475.050 815.400 ;
        RECT 478.950 816.600 481.050 817.050 ;
        RECT 484.950 816.600 487.050 817.050 ;
        RECT 478.950 815.400 487.050 816.600 ;
        RECT 478.950 814.950 481.050 815.400 ;
        RECT 484.950 814.950 487.050 815.400 ;
        RECT 514.950 816.600 517.050 817.050 ;
        RECT 532.950 816.600 535.050 817.050 ;
        RECT 514.950 815.400 535.050 816.600 ;
        RECT 514.950 814.950 517.050 815.400 ;
        RECT 532.950 814.950 535.050 815.400 ;
        RECT 538.950 816.600 541.050 817.050 ;
        RECT 568.950 816.600 571.050 817.050 ;
        RECT 616.950 816.600 619.050 817.050 ;
        RECT 538.950 815.400 619.050 816.600 ;
        RECT 538.950 814.950 541.050 815.400 ;
        RECT 568.950 814.950 571.050 815.400 ;
        RECT 616.950 814.950 619.050 815.400 ;
        RECT 623.400 814.050 624.600 818.400 ;
        RECT 634.950 817.950 637.050 818.400 ;
        RECT 670.950 819.600 673.050 820.050 ;
        RECT 679.950 819.600 682.050 820.050 ;
        RECT 670.950 818.400 682.050 819.600 ;
        RECT 670.950 817.950 673.050 818.400 ;
        RECT 679.950 817.950 682.050 818.400 ;
        RECT 688.950 819.600 691.050 820.050 ;
        RECT 719.400 819.600 720.600 821.400 ;
        RECT 688.950 818.400 720.600 819.600 ;
        RECT 772.950 819.600 775.050 820.050 ;
        RECT 778.950 819.600 781.050 820.050 ;
        RECT 772.950 818.400 781.050 819.600 ;
        RECT 688.950 817.950 691.050 818.400 ;
        RECT 772.950 817.950 775.050 818.400 ;
        RECT 778.950 817.950 781.050 818.400 ;
        RECT 784.950 819.600 787.050 820.050 ;
        RECT 793.950 819.600 796.050 820.050 ;
        RECT 784.950 818.400 796.050 819.600 ;
        RECT 797.400 819.600 798.600 821.400 ;
        RECT 808.950 821.400 820.050 822.600 ;
        RECT 808.950 820.950 811.050 821.400 ;
        RECT 811.950 820.950 814.050 821.400 ;
        RECT 817.950 820.950 820.050 821.400 ;
        RECT 850.950 819.600 853.050 820.050 ;
        RECT 797.400 818.400 853.050 819.600 ;
        RECT 784.950 817.950 787.050 818.400 ;
        RECT 793.950 817.950 796.050 818.400 ;
        RECT 850.950 817.950 853.050 818.400 ;
        RECT 628.950 816.600 631.050 817.050 ;
        RECT 658.950 816.600 661.050 817.050 ;
        RECT 628.950 815.400 661.050 816.600 ;
        RECT 628.950 814.950 631.050 815.400 ;
        RECT 658.950 814.950 661.050 815.400 ;
        RECT 664.950 814.950 667.050 817.050 ;
        RECT 709.950 816.600 712.050 817.050 ;
        RECT 748.950 816.600 751.050 817.050 ;
        RECT 709.950 815.400 751.050 816.600 ;
        RECT 709.950 814.950 712.050 815.400 ;
        RECT 748.950 814.950 751.050 815.400 ;
        RECT 808.950 816.600 811.050 817.050 ;
        RECT 814.950 816.600 817.050 817.050 ;
        RECT 808.950 815.400 817.050 816.600 ;
        RECT 808.950 814.950 811.050 815.400 ;
        RECT 814.950 814.950 817.050 815.400 ;
        RECT 844.950 816.600 847.050 817.050 ;
        RECT 874.950 816.600 877.050 817.050 ;
        RECT 844.950 815.400 877.050 816.600 ;
        RECT 844.950 814.950 847.050 815.400 ;
        RECT 874.950 814.950 877.050 815.400 ;
        RECT 85.950 812.400 105.600 813.600 ;
        RECT 124.950 813.600 127.050 814.050 ;
        RECT 142.950 813.600 145.050 814.050 ;
        RECT 124.950 812.400 145.050 813.600 ;
        RECT 85.950 811.950 88.050 812.400 ;
        RECT 124.950 811.950 127.050 812.400 ;
        RECT 142.950 811.950 145.050 812.400 ;
        RECT 181.950 813.600 184.050 814.050 ;
        RECT 208.950 813.600 211.050 814.050 ;
        RECT 181.950 812.400 211.050 813.600 ;
        RECT 181.950 811.950 184.050 812.400 ;
        RECT 208.950 811.950 211.050 812.400 ;
        RECT 226.950 813.600 229.050 814.050 ;
        RECT 271.950 813.600 274.050 814.050 ;
        RECT 226.950 812.400 274.050 813.600 ;
        RECT 226.950 811.950 229.050 812.400 ;
        RECT 271.950 811.950 274.050 812.400 ;
        RECT 280.950 813.600 283.050 814.050 ;
        RECT 286.950 813.600 289.050 814.050 ;
        RECT 280.950 812.400 289.050 813.600 ;
        RECT 280.950 811.950 283.050 812.400 ;
        RECT 286.950 811.950 289.050 812.400 ;
        RECT 313.950 813.600 316.050 814.050 ;
        RECT 340.950 813.600 343.050 814.050 ;
        RECT 313.950 812.400 343.050 813.600 ;
        RECT 313.950 811.950 316.050 812.400 ;
        RECT 340.950 811.950 343.050 812.400 ;
        RECT 376.950 813.600 379.050 814.050 ;
        RECT 382.950 813.600 385.050 814.050 ;
        RECT 376.950 812.400 385.050 813.600 ;
        RECT 376.950 811.950 379.050 812.400 ;
        RECT 382.950 811.950 385.050 812.400 ;
        RECT 421.950 811.950 424.050 814.050 ;
        RECT 460.950 813.600 463.050 814.050 ;
        RECT 511.950 813.600 514.050 814.050 ;
        RECT 460.950 812.400 514.050 813.600 ;
        RECT 460.950 811.950 463.050 812.400 ;
        RECT 497.400 811.050 498.600 812.400 ;
        RECT 511.950 811.950 514.050 812.400 ;
        RECT 556.950 813.600 559.050 814.050 ;
        RECT 574.950 813.600 577.050 814.050 ;
        RECT 622.950 813.600 625.050 814.050 ;
        RECT 661.950 813.600 664.050 814.050 ;
        RECT 556.950 812.400 573.600 813.600 ;
        RECT 556.950 811.950 559.050 812.400 ;
        RECT 25.950 810.600 28.050 811.050 ;
        RECT 43.950 810.600 46.050 811.050 ;
        RECT 25.950 809.400 46.050 810.600 ;
        RECT 25.950 808.950 28.050 809.400 ;
        RECT 43.950 808.950 46.050 809.400 ;
        RECT 67.950 810.600 70.050 811.050 ;
        RECT 127.950 810.600 130.050 811.050 ;
        RECT 136.950 810.600 139.050 811.050 ;
        RECT 67.950 809.400 139.050 810.600 ;
        RECT 67.950 808.950 70.050 809.400 ;
        RECT 127.950 808.950 130.050 809.400 ;
        RECT 136.950 808.950 139.050 809.400 ;
        RECT 154.950 810.600 157.050 811.050 ;
        RECT 193.950 810.600 196.050 811.050 ;
        RECT 265.950 810.600 268.050 811.050 ;
        RECT 154.950 809.400 268.050 810.600 ;
        RECT 154.950 808.950 157.050 809.400 ;
        RECT 193.950 808.950 196.050 809.400 ;
        RECT 265.950 808.950 268.050 809.400 ;
        RECT 313.950 810.600 316.050 811.050 ;
        RECT 319.950 810.600 322.050 811.050 ;
        RECT 313.950 809.400 322.050 810.600 ;
        RECT 313.950 808.950 316.050 809.400 ;
        RECT 319.950 808.950 322.050 809.400 ;
        RECT 328.950 810.600 331.050 811.050 ;
        RECT 352.950 810.600 355.050 811.050 ;
        RECT 328.950 809.400 355.050 810.600 ;
        RECT 328.950 808.950 331.050 809.400 ;
        RECT 352.950 808.950 355.050 809.400 ;
        RECT 364.950 810.600 367.050 811.050 ;
        RECT 373.950 810.600 376.050 811.050 ;
        RECT 364.950 809.400 376.050 810.600 ;
        RECT 364.950 808.950 367.050 809.400 ;
        RECT 373.950 808.950 376.050 809.400 ;
        RECT 445.950 810.600 448.050 811.050 ;
        RECT 463.950 810.600 466.050 811.050 ;
        RECT 445.950 809.400 466.050 810.600 ;
        RECT 445.950 808.950 448.050 809.400 ;
        RECT 463.950 808.950 466.050 809.400 ;
        RECT 484.950 810.600 487.050 811.050 ;
        RECT 490.950 810.600 493.050 811.050 ;
        RECT 484.950 809.400 493.050 810.600 ;
        RECT 484.950 808.950 487.050 809.400 ;
        RECT 490.950 808.950 493.050 809.400 ;
        RECT 496.950 808.950 499.050 811.050 ;
        RECT 572.400 810.600 573.600 812.400 ;
        RECT 574.950 812.400 615.600 813.600 ;
        RECT 574.950 811.950 577.050 812.400 ;
        RECT 577.950 810.600 580.050 811.050 ;
        RECT 572.400 809.400 580.050 810.600 ;
        RECT 614.400 810.600 615.600 812.400 ;
        RECT 622.950 812.400 664.050 813.600 ;
        RECT 622.950 811.950 625.050 812.400 ;
        RECT 661.950 811.950 664.050 812.400 ;
        RECT 665.400 811.050 666.600 814.950 ;
        RECT 676.950 813.600 679.050 814.050 ;
        RECT 685.950 813.600 688.050 814.050 ;
        RECT 676.950 812.400 688.050 813.600 ;
        RECT 676.950 811.950 679.050 812.400 ;
        RECT 685.950 811.950 688.050 812.400 ;
        RECT 691.950 813.600 694.050 814.050 ;
        RECT 697.950 813.600 700.050 814.050 ;
        RECT 691.950 812.400 700.050 813.600 ;
        RECT 691.950 811.950 694.050 812.400 ;
        RECT 697.950 811.950 700.050 812.400 ;
        RECT 712.950 813.600 715.050 814.050 ;
        RECT 730.950 813.600 733.050 814.050 ;
        RECT 712.950 812.400 733.050 813.600 ;
        RECT 712.950 811.950 715.050 812.400 ;
        RECT 730.950 811.950 733.050 812.400 ;
        RECT 781.950 813.600 784.050 814.050 ;
        RECT 787.950 813.600 790.050 814.050 ;
        RECT 781.950 812.400 790.050 813.600 ;
        RECT 781.950 811.950 784.050 812.400 ;
        RECT 787.950 811.950 790.050 812.400 ;
        RECT 790.950 813.600 793.050 814.050 ;
        RECT 799.950 813.600 802.050 814.050 ;
        RECT 832.950 813.600 835.050 814.050 ;
        RECT 790.950 812.400 835.050 813.600 ;
        RECT 790.950 811.950 793.050 812.400 ;
        RECT 799.950 811.950 802.050 812.400 ;
        RECT 832.950 811.950 835.050 812.400 ;
        RECT 628.950 810.600 631.050 811.050 ;
        RECT 640.950 810.600 643.050 811.050 ;
        RECT 614.400 809.400 643.050 810.600 ;
        RECT 577.950 808.950 580.050 809.400 ;
        RECT 628.950 808.950 631.050 809.400 ;
        RECT 640.950 808.950 643.050 809.400 ;
        RECT 664.950 808.950 667.050 811.050 ;
        RECT 700.950 810.600 703.050 811.050 ;
        RECT 727.950 810.600 730.050 811.050 ;
        RECT 700.950 809.400 730.050 810.600 ;
        RECT 700.950 808.950 703.050 809.400 ;
        RECT 727.950 808.950 730.050 809.400 ;
        RECT 733.950 810.600 736.050 811.050 ;
        RECT 766.950 810.600 769.050 811.050 ;
        RECT 772.950 810.600 775.050 811.050 ;
        RECT 733.950 809.400 775.050 810.600 ;
        RECT 733.950 808.950 736.050 809.400 ;
        RECT 766.950 808.950 769.050 809.400 ;
        RECT 772.950 808.950 775.050 809.400 ;
        RECT 775.950 810.600 778.050 811.050 ;
        RECT 796.950 810.600 799.050 811.050 ;
        RECT 775.950 809.400 799.050 810.600 ;
        RECT 775.950 808.950 778.050 809.400 ;
        RECT 796.950 808.950 799.050 809.400 ;
        RECT 811.950 810.600 814.050 811.050 ;
        RECT 820.950 810.600 823.050 811.050 ;
        RECT 811.950 809.400 823.050 810.600 ;
        RECT 811.950 808.950 814.050 809.400 ;
        RECT 820.950 808.950 823.050 809.400 ;
        RECT 823.950 810.600 826.050 811.050 ;
        RECT 829.950 810.600 832.050 811.050 ;
        RECT 823.950 809.400 832.050 810.600 ;
        RECT 823.950 808.950 826.050 809.400 ;
        RECT 829.950 808.950 832.050 809.400 ;
        RECT 10.950 807.600 13.050 808.050 ;
        RECT 31.950 807.600 34.050 808.050 ;
        RECT 10.950 806.400 34.050 807.600 ;
        RECT 10.950 805.950 13.050 806.400 ;
        RECT 31.950 805.950 34.050 806.400 ;
        RECT 67.950 807.600 70.050 808.050 ;
        RECT 76.950 807.600 79.050 808.050 ;
        RECT 67.950 806.400 79.050 807.600 ;
        RECT 67.950 805.950 70.050 806.400 ;
        RECT 76.950 805.950 79.050 806.400 ;
        RECT 175.950 807.600 178.050 808.050 ;
        RECT 199.950 807.600 202.050 808.050 ;
        RECT 175.950 806.400 202.050 807.600 ;
        RECT 175.950 805.950 178.050 806.400 ;
        RECT 199.950 805.950 202.050 806.400 ;
        RECT 346.950 807.600 349.050 808.050 ;
        RECT 370.950 807.600 373.050 808.050 ;
        RECT 406.950 807.600 409.050 808.050 ;
        RECT 346.950 806.400 409.050 807.600 ;
        RECT 346.950 805.950 349.050 806.400 ;
        RECT 370.950 805.950 373.050 806.400 ;
        RECT 406.950 805.950 409.050 806.400 ;
        RECT 439.950 807.600 442.050 808.050 ;
        RECT 445.950 807.600 448.050 808.050 ;
        RECT 475.950 807.600 478.050 808.050 ;
        RECT 439.950 806.400 478.050 807.600 ;
        RECT 439.950 805.950 442.050 806.400 ;
        RECT 445.950 805.950 448.050 806.400 ;
        RECT 475.950 805.950 478.050 806.400 ;
        RECT 532.950 807.600 535.050 808.050 ;
        RECT 595.950 807.600 598.050 808.050 ;
        RECT 532.950 806.400 598.050 807.600 ;
        RECT 532.950 805.950 535.050 806.400 ;
        RECT 595.950 805.950 598.050 806.400 ;
        RECT 631.950 807.600 634.050 808.050 ;
        RECT 706.950 807.600 709.050 808.050 ;
        RECT 631.950 806.400 709.050 807.600 ;
        RECT 631.950 805.950 634.050 806.400 ;
        RECT 706.950 805.950 709.050 806.400 ;
        RECT 715.950 807.600 718.050 808.050 ;
        RECT 778.950 807.600 781.050 808.050 ;
        RECT 835.950 807.600 838.050 808.050 ;
        RECT 715.950 806.400 838.050 807.600 ;
        RECT 715.950 805.950 718.050 806.400 ;
        RECT 778.950 805.950 781.050 806.400 ;
        RECT 835.950 805.950 838.050 806.400 ;
        RECT 337.950 804.600 340.050 805.050 ;
        RECT 346.950 804.600 349.050 805.050 ;
        RECT 337.950 803.400 349.050 804.600 ;
        RECT 337.950 802.950 340.050 803.400 ;
        RECT 346.950 802.950 349.050 803.400 ;
        RECT 361.950 804.600 364.050 805.050 ;
        RECT 397.950 804.600 400.050 805.050 ;
        RECT 361.950 803.400 400.050 804.600 ;
        RECT 361.950 802.950 364.050 803.400 ;
        RECT 397.950 802.950 400.050 803.400 ;
        RECT 481.950 804.600 484.050 805.050 ;
        RECT 559.950 804.600 562.050 805.050 ;
        RECT 481.950 803.400 562.050 804.600 ;
        RECT 481.950 802.950 484.050 803.400 ;
        RECT 559.950 802.950 562.050 803.400 ;
        RECT 562.950 804.600 565.050 805.050 ;
        RECT 712.950 804.600 715.050 805.050 ;
        RECT 562.950 803.400 715.050 804.600 ;
        RECT 562.950 802.950 565.050 803.400 ;
        RECT 712.950 802.950 715.050 803.400 ;
        RECT 724.950 804.600 727.050 805.050 ;
        RECT 733.950 804.600 736.050 805.050 ;
        RECT 808.950 804.600 811.050 805.050 ;
        RECT 724.950 803.400 811.050 804.600 ;
        RECT 724.950 802.950 727.050 803.400 ;
        RECT 733.950 802.950 736.050 803.400 ;
        RECT 808.950 802.950 811.050 803.400 ;
        RECT 298.950 801.600 301.050 802.050 ;
        RECT 391.950 801.600 394.050 802.050 ;
        RECT 298.950 800.400 394.050 801.600 ;
        RECT 298.950 799.950 301.050 800.400 ;
        RECT 391.950 799.950 394.050 800.400 ;
        RECT 169.950 798.600 172.050 799.050 ;
        RECT 181.950 798.600 184.050 799.050 ;
        RECT 169.950 797.400 184.050 798.600 ;
        RECT 169.950 796.950 172.050 797.400 ;
        RECT 181.950 796.950 184.050 797.400 ;
        RECT 403.950 798.600 406.050 799.050 ;
        RECT 415.950 798.600 418.050 799.050 ;
        RECT 688.950 798.600 691.050 799.050 ;
        RECT 403.950 797.400 691.050 798.600 ;
        RECT 403.950 796.950 406.050 797.400 ;
        RECT 415.950 796.950 418.050 797.400 ;
        RECT 688.950 796.950 691.050 797.400 ;
        RECT 460.950 795.600 463.050 796.050 ;
        RECT 535.950 795.600 538.050 796.050 ;
        RECT 460.950 794.400 538.050 795.600 ;
        RECT 460.950 793.950 463.050 794.400 ;
        RECT 535.950 793.950 538.050 794.400 ;
        RECT 466.950 792.600 469.050 793.050 ;
        RECT 589.950 792.600 592.050 793.050 ;
        RECT 466.950 791.400 592.050 792.600 ;
        RECT 466.950 790.950 469.050 791.400 ;
        RECT 589.950 790.950 592.050 791.400 ;
        RECT 529.950 789.600 532.050 790.050 ;
        RECT 544.950 789.600 547.050 790.050 ;
        RECT 553.950 789.600 556.050 790.050 ;
        RECT 529.950 788.400 556.050 789.600 ;
        RECT 529.950 787.950 532.050 788.400 ;
        RECT 544.950 787.950 547.050 788.400 ;
        RECT 553.950 787.950 556.050 788.400 ;
        RECT 643.950 786.600 646.050 787.050 ;
        RECT 679.950 786.600 682.050 787.050 ;
        RECT 643.950 785.400 682.050 786.600 ;
        RECT 643.950 784.950 646.050 785.400 ;
        RECT 679.950 784.950 682.050 785.400 ;
        RECT 100.950 783.600 103.050 784.050 ;
        RECT 133.950 783.600 136.050 784.050 ;
        RECT 100.950 782.400 136.050 783.600 ;
        RECT 100.950 781.950 103.050 782.400 ;
        RECT 133.950 781.950 136.050 782.400 ;
        RECT 451.950 783.600 454.050 784.050 ;
        RECT 547.950 783.600 550.050 784.050 ;
        RECT 451.950 782.400 550.050 783.600 ;
        RECT 451.950 781.950 454.050 782.400 ;
        RECT 547.950 781.950 550.050 782.400 ;
        RECT 670.950 783.600 673.050 784.050 ;
        RECT 679.950 783.600 682.050 784.050 ;
        RECT 670.950 782.400 682.050 783.600 ;
        RECT 670.950 781.950 673.050 782.400 ;
        RECT 679.950 781.950 682.050 782.400 ;
        RECT 19.950 780.600 22.050 781.050 ;
        RECT 25.950 780.600 28.050 781.050 ;
        RECT 37.950 780.600 40.050 781.050 ;
        RECT 19.950 779.400 40.050 780.600 ;
        RECT 19.950 778.950 22.050 779.400 ;
        RECT 25.950 778.950 28.050 779.400 ;
        RECT 37.950 778.950 40.050 779.400 ;
        RECT 472.950 780.600 475.050 781.050 ;
        RECT 649.950 780.600 652.050 781.050 ;
        RECT 472.950 779.400 652.050 780.600 ;
        RECT 472.950 778.950 475.050 779.400 ;
        RECT 649.950 778.950 652.050 779.400 ;
        RECT 658.950 780.600 661.050 781.050 ;
        RECT 745.950 780.600 748.050 781.050 ;
        RECT 658.950 779.400 748.050 780.600 ;
        RECT 658.950 778.950 661.050 779.400 ;
        RECT 745.950 778.950 748.050 779.400 ;
        RECT 13.950 777.600 16.050 778.050 ;
        RECT 28.950 777.600 31.050 778.050 ;
        RECT 13.950 776.400 31.050 777.600 ;
        RECT 13.950 775.950 16.050 776.400 ;
        RECT 28.950 775.950 31.050 776.400 ;
        RECT 94.950 777.600 97.050 778.050 ;
        RECT 106.950 777.600 109.050 778.050 ;
        RECT 112.950 777.600 115.050 778.050 ;
        RECT 94.950 776.400 115.050 777.600 ;
        RECT 94.950 775.950 97.050 776.400 ;
        RECT 106.950 775.950 109.050 776.400 ;
        RECT 112.950 775.950 115.050 776.400 ;
        RECT 148.950 777.600 151.050 778.050 ;
        RECT 184.950 777.600 187.050 778.050 ;
        RECT 241.950 777.600 244.050 778.050 ;
        RECT 250.950 777.600 253.050 778.050 ;
        RECT 349.950 777.600 352.050 778.050 ;
        RECT 148.950 776.400 352.050 777.600 ;
        RECT 148.950 775.950 151.050 776.400 ;
        RECT 184.950 775.950 187.050 776.400 ;
        RECT 241.950 775.950 244.050 776.400 ;
        RECT 250.950 775.950 253.050 776.400 ;
        RECT 349.950 775.950 352.050 776.400 ;
        RECT 397.950 777.600 400.050 778.050 ;
        RECT 406.950 777.600 409.050 778.050 ;
        RECT 451.950 777.600 454.050 778.050 ;
        RECT 397.950 776.400 454.050 777.600 ;
        RECT 397.950 775.950 400.050 776.400 ;
        RECT 406.950 775.950 409.050 776.400 ;
        RECT 451.950 775.950 454.050 776.400 ;
        RECT 517.950 777.600 520.050 778.050 ;
        RECT 583.950 777.600 586.050 778.050 ;
        RECT 598.950 777.600 601.050 778.050 ;
        RECT 517.950 776.400 543.600 777.600 ;
        RECT 517.950 775.950 520.050 776.400 ;
        RECT 16.950 774.600 19.050 775.050 ;
        RECT 22.950 774.600 25.050 775.050 ;
        RECT 16.950 773.400 25.050 774.600 ;
        RECT 16.950 772.950 19.050 773.400 ;
        RECT 22.950 772.950 25.050 773.400 ;
        RECT 55.950 774.600 58.050 775.050 ;
        RECT 73.950 774.600 76.050 775.050 ;
        RECT 55.950 773.400 76.050 774.600 ;
        RECT 55.950 772.950 58.050 773.400 ;
        RECT 73.950 772.950 76.050 773.400 ;
        RECT 91.950 774.600 94.050 775.050 ;
        RECT 115.950 774.600 118.050 775.050 ;
        RECT 91.950 773.400 118.050 774.600 ;
        RECT 91.950 772.950 94.050 773.400 ;
        RECT 115.950 772.950 118.050 773.400 ;
        RECT 175.950 772.950 178.050 775.050 ;
        RECT 184.950 774.600 187.050 775.050 ;
        RECT 214.950 774.600 217.050 775.050 ;
        RECT 184.950 773.400 217.050 774.600 ;
        RECT 184.950 772.950 187.050 773.400 ;
        RECT 214.950 772.950 217.050 773.400 ;
        RECT 238.950 774.600 241.050 775.050 ;
        RECT 244.950 774.600 247.050 775.050 ;
        RECT 238.950 773.400 247.050 774.600 ;
        RECT 238.950 772.950 241.050 773.400 ;
        RECT 244.950 772.950 247.050 773.400 ;
        RECT 256.950 774.600 259.050 775.050 ;
        RECT 277.950 774.600 280.050 775.050 ;
        RECT 286.950 774.600 289.050 775.050 ;
        RECT 256.950 773.400 276.600 774.600 ;
        RECT 256.950 772.950 259.050 773.400 ;
        RECT 64.950 771.600 67.050 772.050 ;
        RECT 70.950 771.600 73.050 772.050 ;
        RECT 64.950 770.400 73.050 771.600 ;
        RECT 64.950 769.950 67.050 770.400 ;
        RECT 70.950 769.950 73.050 770.400 ;
        RECT 115.950 771.600 118.050 772.050 ;
        RECT 130.950 771.600 133.050 772.050 ;
        RECT 115.950 770.400 133.050 771.600 ;
        RECT 115.950 769.950 118.050 770.400 ;
        RECT 130.950 769.950 133.050 770.400 ;
        RECT 176.400 769.050 177.600 772.950 ;
        RECT 217.950 771.600 220.050 772.050 ;
        RECT 232.950 771.600 235.050 772.050 ;
        RECT 217.950 770.400 235.050 771.600 ;
        RECT 275.400 771.600 276.600 773.400 ;
        RECT 277.950 773.400 289.050 774.600 ;
        RECT 277.950 772.950 280.050 773.400 ;
        RECT 286.950 772.950 289.050 773.400 ;
        RECT 391.950 774.600 394.050 775.050 ;
        RECT 403.950 774.600 406.050 775.050 ;
        RECT 391.950 773.400 406.050 774.600 ;
        RECT 391.950 772.950 394.050 773.400 ;
        RECT 403.950 772.950 406.050 773.400 ;
        RECT 436.950 774.600 439.050 775.050 ;
        RECT 457.950 774.600 460.050 775.050 ;
        RECT 463.950 774.600 466.050 775.050 ;
        RECT 436.950 773.400 450.600 774.600 ;
        RECT 436.950 772.950 439.050 773.400 ;
        RECT 449.400 772.050 450.600 773.400 ;
        RECT 457.950 773.400 466.050 774.600 ;
        RECT 457.950 772.950 460.050 773.400 ;
        RECT 463.950 772.950 466.050 773.400 ;
        RECT 478.950 774.600 481.050 775.050 ;
        RECT 490.950 774.600 493.050 775.050 ;
        RECT 499.950 774.600 502.050 775.050 ;
        RECT 514.950 774.600 517.050 775.050 ;
        RECT 478.950 773.400 493.050 774.600 ;
        RECT 478.950 772.950 481.050 773.400 ;
        RECT 490.950 772.950 493.050 773.400 ;
        RECT 497.400 773.400 517.050 774.600 ;
        RECT 542.400 774.600 543.600 776.400 ;
        RECT 583.950 776.400 601.050 777.600 ;
        RECT 583.950 775.950 586.050 776.400 ;
        RECT 598.950 775.950 601.050 776.400 ;
        RECT 616.950 777.600 619.050 778.050 ;
        RECT 625.950 777.600 628.050 778.050 ;
        RECT 628.950 777.600 631.050 778.050 ;
        RECT 616.950 776.400 631.050 777.600 ;
        RECT 616.950 775.950 619.050 776.400 ;
        RECT 625.950 775.950 628.050 776.400 ;
        RECT 628.950 775.950 631.050 776.400 ;
        RECT 646.950 777.600 649.050 778.050 ;
        RECT 673.950 777.600 676.050 778.050 ;
        RECT 646.950 776.400 676.050 777.600 ;
        RECT 646.950 775.950 649.050 776.400 ;
        RECT 673.950 775.950 676.050 776.400 ;
        RECT 769.950 777.600 772.050 778.050 ;
        RECT 781.950 777.600 784.050 778.050 ;
        RECT 769.950 776.400 784.050 777.600 ;
        RECT 769.950 775.950 772.050 776.400 ;
        RECT 781.950 775.950 784.050 776.400 ;
        RECT 793.950 777.600 796.050 778.050 ;
        RECT 802.950 777.600 805.050 778.050 ;
        RECT 793.950 776.400 805.050 777.600 ;
        RECT 793.950 775.950 796.050 776.400 ;
        RECT 802.950 775.950 805.050 776.400 ;
        RECT 805.950 777.600 808.050 778.050 ;
        RECT 805.950 776.400 816.600 777.600 ;
        RECT 805.950 775.950 808.050 776.400 ;
        RECT 815.400 775.050 816.600 776.400 ;
        RECT 565.950 774.600 568.050 775.050 ;
        RECT 580.950 774.600 583.050 775.050 ;
        RECT 542.400 773.400 583.050 774.600 ;
        RECT 497.400 772.050 498.600 773.400 ;
        RECT 499.950 772.950 502.050 773.400 ;
        RECT 514.950 772.950 517.050 773.400 ;
        RECT 565.950 772.950 568.050 773.400 ;
        RECT 580.950 772.950 583.050 773.400 ;
        RECT 601.950 774.600 604.050 775.050 ;
        RECT 631.950 774.600 634.050 775.050 ;
        RECT 601.950 773.400 634.050 774.600 ;
        RECT 601.950 772.950 604.050 773.400 ;
        RECT 631.950 772.950 634.050 773.400 ;
        RECT 679.950 772.950 682.050 775.050 ;
        RECT 685.950 774.600 688.050 775.050 ;
        RECT 772.950 774.600 775.050 775.050 ;
        RECT 808.950 774.600 811.050 775.050 ;
        RECT 685.950 773.400 811.050 774.600 ;
        RECT 685.950 772.950 688.050 773.400 ;
        RECT 772.950 772.950 775.050 773.400 ;
        RECT 808.950 772.950 811.050 773.400 ;
        RECT 814.950 772.950 817.050 775.050 ;
        RECT 829.950 772.950 832.050 775.050 ;
        RECT 280.950 771.600 283.050 772.050 ;
        RECT 292.950 771.600 295.050 772.050 ;
        RECT 275.400 770.400 295.050 771.600 ;
        RECT 217.950 769.950 220.050 770.400 ;
        RECT 232.950 769.950 235.050 770.400 ;
        RECT 280.950 769.950 283.050 770.400 ;
        RECT 292.950 769.950 295.050 770.400 ;
        RECT 298.950 771.600 301.050 772.050 ;
        RECT 307.950 771.600 310.050 772.050 ;
        RECT 298.950 770.400 310.050 771.600 ;
        RECT 298.950 769.950 301.050 770.400 ;
        RECT 307.950 769.950 310.050 770.400 ;
        RECT 385.950 771.600 388.050 772.050 ;
        RECT 394.950 771.600 397.050 772.050 ;
        RECT 385.950 770.400 397.050 771.600 ;
        RECT 385.950 769.950 388.050 770.400 ;
        RECT 394.950 769.950 397.050 770.400 ;
        RECT 427.950 771.600 430.050 772.050 ;
        RECT 439.950 771.600 442.050 772.050 ;
        RECT 427.950 770.400 442.050 771.600 ;
        RECT 427.950 769.950 430.050 770.400 ;
        RECT 439.950 769.950 442.050 770.400 ;
        RECT 448.950 769.950 451.050 772.050 ;
        RECT 454.950 771.600 457.050 772.050 ;
        RECT 466.950 771.600 469.050 772.050 ;
        RECT 454.950 770.400 469.050 771.600 ;
        RECT 454.950 769.950 457.050 770.400 ;
        RECT 466.950 769.950 469.050 770.400 ;
        RECT 496.950 769.950 499.050 772.050 ;
        RECT 652.950 771.600 655.050 772.050 ;
        RECT 658.950 771.600 661.050 772.050 ;
        RECT 652.950 770.400 661.050 771.600 ;
        RECT 652.950 769.950 655.050 770.400 ;
        RECT 658.950 769.950 661.050 770.400 ;
        RECT 664.950 771.600 667.050 772.050 ;
        RECT 670.950 771.600 673.050 772.050 ;
        RECT 664.950 770.400 673.050 771.600 ;
        RECT 680.400 771.600 681.600 772.950 ;
        RECT 694.950 771.600 697.050 772.050 ;
        RECT 680.400 770.400 697.050 771.600 ;
        RECT 664.950 769.950 667.050 770.400 ;
        RECT 670.950 769.950 673.050 770.400 ;
        RECT 694.950 769.950 697.050 770.400 ;
        RECT 754.950 771.600 757.050 772.050 ;
        RECT 787.950 771.600 790.050 772.050 ;
        RECT 811.950 771.600 814.050 772.050 ;
        RECT 830.400 771.600 831.600 772.950 ;
        RECT 754.950 770.400 771.600 771.600 ;
        RECT 754.950 769.950 757.050 770.400 ;
        RECT 770.400 769.050 771.600 770.400 ;
        RECT 787.950 770.400 795.600 771.600 ;
        RECT 787.950 769.950 790.050 770.400 ;
        RECT 37.950 768.600 40.050 769.050 ;
        RECT 52.950 768.600 55.050 769.050 ;
        RECT 37.950 767.400 55.050 768.600 ;
        RECT 37.950 766.950 40.050 767.400 ;
        RECT 52.950 766.950 55.050 767.400 ;
        RECT 91.950 768.600 94.050 769.050 ;
        RECT 109.950 768.600 112.050 769.050 ;
        RECT 91.950 767.400 112.050 768.600 ;
        RECT 91.950 766.950 94.050 767.400 ;
        RECT 109.950 766.950 112.050 767.400 ;
        RECT 133.950 768.600 136.050 769.050 ;
        RECT 148.950 768.600 151.050 769.050 ;
        RECT 166.950 768.600 169.050 769.050 ;
        RECT 133.950 767.400 169.050 768.600 ;
        RECT 133.950 766.950 136.050 767.400 ;
        RECT 148.950 766.950 151.050 767.400 ;
        RECT 166.950 766.950 169.050 767.400 ;
        RECT 175.950 766.950 178.050 769.050 ;
        RECT 196.950 768.600 199.050 769.050 ;
        RECT 211.950 768.600 214.050 769.050 ;
        RECT 196.950 767.400 214.050 768.600 ;
        RECT 196.950 766.950 199.050 767.400 ;
        RECT 211.950 766.950 214.050 767.400 ;
        RECT 274.950 768.600 277.050 769.050 ;
        RECT 301.950 768.600 304.050 769.050 ;
        RECT 274.950 767.400 304.050 768.600 ;
        RECT 274.950 766.950 277.050 767.400 ;
        RECT 301.950 766.950 304.050 767.400 ;
        RECT 373.950 768.600 376.050 769.050 ;
        RECT 415.950 768.600 418.050 769.050 ;
        RECT 373.950 767.400 418.050 768.600 ;
        RECT 373.950 766.950 376.050 767.400 ;
        RECT 415.950 766.950 418.050 767.400 ;
        RECT 442.950 768.600 445.050 769.050 ;
        RECT 469.950 768.600 472.050 769.050 ;
        RECT 442.950 767.400 472.050 768.600 ;
        RECT 442.950 766.950 445.050 767.400 ;
        RECT 469.950 766.950 472.050 767.400 ;
        RECT 601.950 768.600 604.050 769.050 ;
        RECT 637.950 768.600 640.050 769.050 ;
        RECT 601.950 767.400 640.050 768.600 ;
        RECT 601.950 766.950 604.050 767.400 ;
        RECT 637.950 766.950 640.050 767.400 ;
        RECT 676.950 768.600 679.050 769.050 ;
        RECT 736.950 768.600 739.050 769.050 ;
        RECT 676.950 767.400 739.050 768.600 ;
        RECT 676.950 766.950 679.050 767.400 ;
        RECT 736.950 766.950 739.050 767.400 ;
        RECT 769.950 766.950 772.050 769.050 ;
        RECT 781.950 768.600 784.050 769.050 ;
        RECT 790.950 768.600 793.050 769.050 ;
        RECT 781.950 767.400 793.050 768.600 ;
        RECT 794.400 768.600 795.600 770.400 ;
        RECT 811.950 770.400 831.600 771.600 ;
        RECT 811.950 769.950 814.050 770.400 ;
        RECT 808.950 768.600 811.050 769.050 ;
        RECT 794.400 767.400 811.050 768.600 ;
        RECT 781.950 766.950 784.050 767.400 ;
        RECT 790.950 766.950 793.050 767.400 ;
        RECT 808.950 766.950 811.050 767.400 ;
        RECT 820.950 768.600 823.050 769.050 ;
        RECT 826.950 768.600 829.050 769.050 ;
        RECT 832.950 768.600 835.050 769.050 ;
        RECT 820.950 767.400 835.050 768.600 ;
        RECT 820.950 766.950 823.050 767.400 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 832.950 766.950 835.050 767.400 ;
        RECT 136.950 765.600 139.050 766.050 ;
        RECT 184.950 765.600 187.050 766.050 ;
        RECT 136.950 764.400 187.050 765.600 ;
        RECT 136.950 763.950 139.050 764.400 ;
        RECT 184.950 763.950 187.050 764.400 ;
        RECT 412.950 765.600 415.050 766.050 ;
        RECT 430.950 765.600 433.050 766.050 ;
        RECT 484.950 765.600 487.050 766.050 ;
        RECT 412.950 764.400 487.050 765.600 ;
        RECT 412.950 763.950 415.050 764.400 ;
        RECT 430.950 763.950 433.050 764.400 ;
        RECT 484.950 763.950 487.050 764.400 ;
        RECT 574.950 765.600 577.050 766.050 ;
        RECT 577.950 765.600 580.050 766.050 ;
        RECT 613.950 765.600 616.050 766.050 ;
        RECT 574.950 764.400 616.050 765.600 ;
        RECT 574.950 763.950 577.050 764.400 ;
        RECT 577.950 763.950 580.050 764.400 ;
        RECT 613.950 763.950 616.050 764.400 ;
        RECT 757.950 765.600 760.050 766.050 ;
        RECT 805.950 765.600 808.050 766.050 ;
        RECT 757.950 764.400 808.050 765.600 ;
        RECT 757.950 763.950 760.050 764.400 ;
        RECT 805.950 763.950 808.050 764.400 ;
        RECT 832.950 765.600 835.050 766.050 ;
        RECT 841.950 765.600 844.050 766.050 ;
        RECT 832.950 764.400 844.050 765.600 ;
        RECT 832.950 763.950 835.050 764.400 ;
        RECT 841.950 763.950 844.050 764.400 ;
        RECT 40.950 762.600 43.050 763.050 ;
        RECT 58.950 762.600 61.050 763.050 ;
        RECT 40.950 761.400 61.050 762.600 ;
        RECT 40.950 760.950 43.050 761.400 ;
        RECT 58.950 760.950 61.050 761.400 ;
        RECT 67.950 762.600 70.050 763.050 ;
        RECT 76.950 762.600 79.050 763.050 ;
        RECT 100.950 762.600 103.050 763.050 ;
        RECT 67.950 761.400 103.050 762.600 ;
        RECT 67.950 760.950 70.050 761.400 ;
        RECT 76.950 760.950 79.050 761.400 ;
        RECT 100.950 760.950 103.050 761.400 ;
        RECT 151.950 762.600 154.050 763.050 ;
        RECT 172.950 762.600 175.050 763.050 ;
        RECT 151.950 761.400 175.050 762.600 ;
        RECT 151.950 760.950 154.050 761.400 ;
        RECT 172.950 760.950 175.050 761.400 ;
        RECT 742.950 762.600 745.050 763.050 ;
        RECT 793.950 762.600 796.050 763.050 ;
        RECT 742.950 761.400 796.050 762.600 ;
        RECT 742.950 760.950 745.050 761.400 ;
        RECT 793.950 760.950 796.050 761.400 ;
        RECT 802.950 762.600 805.050 763.050 ;
        RECT 838.950 762.600 841.050 763.050 ;
        RECT 802.950 761.400 841.050 762.600 ;
        RECT 802.950 760.950 805.050 761.400 ;
        RECT 838.950 760.950 841.050 761.400 ;
        RECT 358.950 759.600 361.050 760.050 ;
        RECT 361.950 759.600 364.050 760.050 ;
        RECT 673.950 759.600 676.050 760.050 ;
        RECT 700.950 759.600 703.050 760.050 ;
        RECT 358.950 758.400 703.050 759.600 ;
        RECT 358.950 757.950 361.050 758.400 ;
        RECT 361.950 757.950 364.050 758.400 ;
        RECT 673.950 757.950 676.050 758.400 ;
        RECT 700.950 757.950 703.050 758.400 ;
        RECT 769.950 759.600 772.050 760.050 ;
        RECT 823.950 759.600 826.050 760.050 ;
        RECT 769.950 758.400 826.050 759.600 ;
        RECT 769.950 757.950 772.050 758.400 ;
        RECT 823.950 757.950 826.050 758.400 ;
        RECT 532.950 756.600 535.050 757.050 ;
        RECT 556.950 756.600 559.050 757.050 ;
        RECT 532.950 755.400 559.050 756.600 ;
        RECT 532.950 754.950 535.050 755.400 ;
        RECT 556.950 754.950 559.050 755.400 ;
        RECT 790.950 756.600 793.050 757.050 ;
        RECT 796.950 756.600 799.050 757.050 ;
        RECT 844.950 756.600 847.050 757.050 ;
        RECT 790.950 755.400 847.050 756.600 ;
        RECT 790.950 754.950 793.050 755.400 ;
        RECT 796.950 754.950 799.050 755.400 ;
        RECT 844.950 754.950 847.050 755.400 ;
        RECT 664.950 753.600 667.050 754.050 ;
        RECT 766.950 753.600 769.050 754.050 ;
        RECT 664.950 752.400 769.050 753.600 ;
        RECT 664.950 751.950 667.050 752.400 ;
        RECT 766.950 751.950 769.050 752.400 ;
        RECT 220.950 750.600 223.050 751.050 ;
        RECT 418.950 750.600 421.050 751.050 ;
        RECT 220.950 749.400 421.050 750.600 ;
        RECT 220.950 748.950 223.050 749.400 ;
        RECT 418.950 748.950 421.050 749.400 ;
        RECT 445.950 750.600 448.050 751.050 ;
        RECT 451.950 750.600 454.050 751.050 ;
        RECT 445.950 749.400 454.050 750.600 ;
        RECT 445.950 748.950 448.050 749.400 ;
        RECT 451.950 748.950 454.050 749.400 ;
        RECT 685.950 750.600 688.050 751.050 ;
        RECT 739.950 750.600 742.050 751.050 ;
        RECT 685.950 749.400 742.050 750.600 ;
        RECT 685.950 748.950 688.050 749.400 ;
        RECT 739.950 748.950 742.050 749.400 ;
        RECT 64.950 747.600 67.050 748.050 ;
        RECT 76.950 747.600 79.050 748.050 ;
        RECT 82.950 747.600 85.050 748.050 ;
        RECT 160.950 747.600 163.050 748.050 ;
        RECT 64.950 746.400 163.050 747.600 ;
        RECT 64.950 745.950 67.050 746.400 ;
        RECT 76.950 745.950 79.050 746.400 ;
        RECT 82.950 745.950 85.050 746.400 ;
        RECT 160.950 745.950 163.050 746.400 ;
        RECT 244.950 747.600 247.050 748.050 ;
        RECT 265.950 747.600 268.050 748.050 ;
        RECT 244.950 746.400 268.050 747.600 ;
        RECT 244.950 745.950 247.050 746.400 ;
        RECT 265.950 745.950 268.050 746.400 ;
        RECT 388.950 747.600 391.050 748.050 ;
        RECT 397.950 747.600 400.050 748.050 ;
        RECT 388.950 746.400 400.050 747.600 ;
        RECT 388.950 745.950 391.050 746.400 ;
        RECT 397.950 745.950 400.050 746.400 ;
        RECT 421.950 747.600 424.050 748.050 ;
        RECT 427.950 747.600 430.050 748.050 ;
        RECT 421.950 746.400 430.050 747.600 ;
        RECT 421.950 745.950 424.050 746.400 ;
        RECT 427.950 745.950 430.050 746.400 ;
        RECT 487.950 745.950 490.050 748.050 ;
        RECT 508.950 747.600 511.050 748.050 ;
        RECT 553.950 747.600 556.050 748.050 ;
        RECT 508.950 746.400 556.050 747.600 ;
        RECT 508.950 745.950 511.050 746.400 ;
        RECT 553.950 745.950 556.050 746.400 ;
        RECT 625.950 747.600 628.050 748.050 ;
        RECT 631.950 747.600 634.050 748.050 ;
        RECT 625.950 746.400 634.050 747.600 ;
        RECT 625.950 745.950 628.050 746.400 ;
        RECT 631.950 745.950 634.050 746.400 ;
        RECT 649.950 747.600 652.050 748.050 ;
        RECT 727.950 747.600 730.050 748.050 ;
        RECT 649.950 746.400 730.050 747.600 ;
        RECT 649.950 745.950 652.050 746.400 ;
        RECT 727.950 745.950 730.050 746.400 ;
        RECT 748.950 747.600 751.050 748.050 ;
        RECT 799.950 747.600 802.050 748.050 ;
        RECT 748.950 746.400 802.050 747.600 ;
        RECT 748.950 745.950 751.050 746.400 ;
        RECT 799.950 745.950 802.050 746.400 ;
        RECT 19.950 744.600 22.050 745.050 ;
        RECT 37.950 744.600 40.050 745.050 ;
        RECT 19.950 743.400 40.050 744.600 ;
        RECT 19.950 742.950 22.050 743.400 ;
        RECT 37.950 742.950 40.050 743.400 ;
        RECT 109.950 744.600 112.050 745.050 ;
        RECT 121.950 744.600 124.050 745.050 ;
        RECT 109.950 743.400 124.050 744.600 ;
        RECT 109.950 742.950 112.050 743.400 ;
        RECT 121.950 742.950 124.050 743.400 ;
        RECT 148.950 744.600 151.050 745.050 ;
        RECT 166.950 744.600 169.050 745.050 ;
        RECT 148.950 743.400 169.050 744.600 ;
        RECT 148.950 742.950 151.050 743.400 ;
        RECT 166.950 742.950 169.050 743.400 ;
        RECT 169.950 744.600 172.050 745.050 ;
        RECT 193.950 744.600 196.050 745.050 ;
        RECT 199.950 744.600 202.050 745.050 ;
        RECT 211.950 744.600 214.050 745.050 ;
        RECT 280.950 744.600 283.050 745.050 ;
        RECT 316.950 744.600 319.050 745.050 ;
        RECT 325.950 744.600 328.050 745.050 ;
        RECT 169.950 743.400 214.050 744.600 ;
        RECT 169.950 742.950 172.050 743.400 ;
        RECT 193.950 742.950 196.050 743.400 ;
        RECT 199.950 742.950 202.050 743.400 ;
        RECT 211.950 742.950 214.050 743.400 ;
        RECT 278.400 743.400 328.050 744.600 ;
        RECT 22.950 741.600 25.050 742.050 ;
        RECT 28.950 741.600 31.050 742.050 ;
        RECT 31.950 741.600 34.050 742.050 ;
        RECT 22.950 740.400 34.050 741.600 ;
        RECT 22.950 739.950 25.050 740.400 ;
        RECT 28.950 739.950 31.050 740.400 ;
        RECT 31.950 739.950 34.050 740.400 ;
        RECT 52.950 741.600 55.050 742.050 ;
        RECT 67.950 741.600 70.050 742.050 ;
        RECT 73.950 741.600 76.050 742.050 ;
        RECT 52.950 740.400 76.050 741.600 ;
        RECT 52.950 739.950 55.050 740.400 ;
        RECT 67.950 739.950 70.050 740.400 ;
        RECT 73.950 739.950 76.050 740.400 ;
        RECT 172.950 739.950 175.050 742.050 ;
        RECT 208.950 741.600 211.050 742.050 ;
        RECT 232.950 741.600 235.050 742.050 ;
        RECT 244.950 741.600 247.050 742.050 ;
        RECT 208.950 740.400 213.600 741.600 ;
        RECT 208.950 739.950 211.050 740.400 ;
        RECT 25.950 738.600 28.050 739.050 ;
        RECT 34.950 738.600 37.050 739.050 ;
        RECT 25.950 737.400 37.050 738.600 ;
        RECT 25.950 736.950 28.050 737.400 ;
        RECT 34.950 736.950 37.050 737.400 ;
        RECT 40.950 738.600 43.050 739.050 ;
        RECT 79.950 738.600 82.050 739.050 ;
        RECT 40.950 737.400 82.050 738.600 ;
        RECT 40.950 736.950 43.050 737.400 ;
        RECT 79.950 736.950 82.050 737.400 ;
        RECT 124.950 738.600 127.050 739.050 ;
        RECT 145.950 738.600 148.050 739.050 ;
        RECT 124.950 737.400 148.050 738.600 ;
        RECT 173.400 738.600 174.600 739.950 ;
        RECT 212.400 739.050 213.600 740.400 ;
        RECT 232.950 740.400 247.050 741.600 ;
        RECT 232.950 739.950 235.050 740.400 ;
        RECT 244.950 739.950 247.050 740.400 ;
        RECT 259.950 741.600 262.050 742.050 ;
        RECT 265.950 741.600 268.050 742.050 ;
        RECT 259.950 740.400 268.050 741.600 ;
        RECT 259.950 739.950 262.050 740.400 ;
        RECT 265.950 739.950 268.050 740.400 ;
        RECT 268.950 741.600 271.050 742.050 ;
        RECT 278.400 741.600 279.600 743.400 ;
        RECT 280.950 742.950 283.050 743.400 ;
        RECT 316.950 742.950 319.050 743.400 ;
        RECT 325.950 742.950 328.050 743.400 ;
        RECT 340.950 744.600 343.050 745.050 ;
        RECT 358.950 744.600 361.050 745.050 ;
        RECT 367.950 744.600 370.050 745.050 ;
        RECT 385.950 744.600 388.050 745.050 ;
        RECT 340.950 743.400 388.050 744.600 ;
        RECT 340.950 742.950 343.050 743.400 ;
        RECT 358.950 742.950 361.050 743.400 ;
        RECT 367.950 742.950 370.050 743.400 ;
        RECT 385.950 742.950 388.050 743.400 ;
        RECT 394.950 744.600 397.050 745.050 ;
        RECT 400.950 744.600 403.050 745.050 ;
        RECT 409.950 744.600 412.050 745.050 ;
        RECT 412.950 744.600 415.050 745.050 ;
        RECT 394.950 743.400 415.050 744.600 ;
        RECT 394.950 742.950 397.050 743.400 ;
        RECT 400.950 742.950 403.050 743.400 ;
        RECT 409.950 742.950 412.050 743.400 ;
        RECT 412.950 742.950 415.050 743.400 ;
        RECT 289.950 741.600 292.050 742.050 ;
        RECT 268.950 740.400 279.600 741.600 ;
        RECT 281.400 740.400 292.050 741.600 ;
        RECT 268.950 739.950 271.050 740.400 ;
        RECT 187.950 738.600 190.050 739.050 ;
        RECT 190.950 738.600 193.050 739.050 ;
        RECT 173.400 737.400 193.050 738.600 ;
        RECT 124.950 736.950 127.050 737.400 ;
        RECT 145.950 736.950 148.050 737.400 ;
        RECT 187.950 736.950 190.050 737.400 ;
        RECT 190.950 736.950 193.050 737.400 ;
        RECT 211.950 736.950 214.050 739.050 ;
        RECT 214.950 738.600 217.050 739.050 ;
        RECT 229.950 738.600 232.050 739.050 ;
        RECT 214.950 737.400 232.050 738.600 ;
        RECT 214.950 736.950 217.050 737.400 ;
        RECT 229.950 736.950 232.050 737.400 ;
        RECT 235.950 736.950 238.050 739.050 ;
        RECT 241.950 738.600 244.050 739.050 ;
        RECT 247.950 738.600 250.050 739.050 ;
        RECT 241.950 737.400 250.050 738.600 ;
        RECT 241.950 736.950 244.050 737.400 ;
        RECT 247.950 736.950 250.050 737.400 ;
        RECT 259.950 738.600 262.050 739.050 ;
        RECT 281.400 738.600 282.600 740.400 ;
        RECT 289.950 739.950 292.050 740.400 ;
        RECT 310.950 741.600 313.050 742.050 ;
        RECT 340.950 741.600 343.050 742.050 ;
        RECT 424.950 741.600 427.050 742.050 ;
        RECT 310.950 740.400 343.050 741.600 ;
        RECT 310.950 739.950 313.050 740.400 ;
        RECT 340.950 739.950 343.050 740.400 ;
        RECT 413.400 740.400 427.050 741.600 ;
        RECT 259.950 737.400 282.600 738.600 ;
        RECT 283.950 738.600 286.050 739.050 ;
        RECT 307.950 738.600 310.050 739.050 ;
        RECT 319.950 738.600 322.050 739.050 ;
        RECT 283.950 737.400 322.050 738.600 ;
        RECT 259.950 736.950 262.050 737.400 ;
        RECT 283.950 736.950 286.050 737.400 ;
        RECT 307.950 736.950 310.050 737.400 ;
        RECT 319.950 736.950 322.050 737.400 ;
        RECT 331.950 738.600 334.050 739.050 ;
        RECT 349.950 738.600 352.050 739.050 ;
        RECT 331.950 737.400 352.050 738.600 ;
        RECT 331.950 736.950 334.050 737.400 ;
        RECT 349.950 736.950 352.050 737.400 ;
        RECT 403.950 738.600 406.050 739.050 ;
        RECT 409.950 738.600 412.050 739.050 ;
        RECT 413.400 738.600 414.600 740.400 ;
        RECT 424.950 739.950 427.050 740.400 ;
        RECT 430.950 741.600 433.050 742.050 ;
        RECT 442.950 741.600 445.050 742.050 ;
        RECT 481.950 741.600 484.050 742.050 ;
        RECT 430.950 740.400 484.050 741.600 ;
        RECT 430.950 739.950 433.050 740.400 ;
        RECT 442.950 739.950 445.050 740.400 ;
        RECT 481.950 739.950 484.050 740.400 ;
        RECT 403.950 737.400 414.600 738.600 ;
        RECT 415.950 738.600 418.050 739.050 ;
        RECT 421.950 738.600 424.050 739.050 ;
        RECT 415.950 737.400 424.050 738.600 ;
        RECT 403.950 736.950 406.050 737.400 ;
        RECT 409.950 736.950 412.050 737.400 ;
        RECT 415.950 736.950 418.050 737.400 ;
        RECT 421.950 736.950 424.050 737.400 ;
        RECT 424.950 738.600 427.050 739.050 ;
        RECT 472.950 738.600 475.050 739.050 ;
        RECT 424.950 737.400 475.050 738.600 ;
        RECT 488.400 738.600 489.600 745.950 ;
        RECT 496.950 744.600 499.050 745.050 ;
        RECT 502.950 744.600 505.050 745.050 ;
        RECT 496.950 743.400 505.050 744.600 ;
        RECT 496.950 742.950 499.050 743.400 ;
        RECT 502.950 742.950 505.050 743.400 ;
        RECT 538.950 744.600 541.050 745.050 ;
        RECT 544.950 744.600 547.050 745.050 ;
        RECT 538.950 743.400 547.050 744.600 ;
        RECT 538.950 742.950 541.050 743.400 ;
        RECT 544.950 742.950 547.050 743.400 ;
        RECT 550.950 744.600 553.050 745.050 ;
        RECT 559.950 744.600 562.050 745.050 ;
        RECT 592.950 744.600 595.050 745.050 ;
        RECT 550.950 743.400 595.050 744.600 ;
        RECT 550.950 742.950 553.050 743.400 ;
        RECT 559.950 742.950 562.050 743.400 ;
        RECT 592.950 742.950 595.050 743.400 ;
        RECT 598.950 744.600 601.050 745.050 ;
        RECT 625.950 744.600 628.050 745.050 ;
        RECT 598.950 743.400 628.050 744.600 ;
        RECT 598.950 742.950 601.050 743.400 ;
        RECT 625.950 742.950 628.050 743.400 ;
        RECT 694.950 744.600 697.050 745.050 ;
        RECT 700.950 744.600 703.050 745.050 ;
        RECT 694.950 743.400 703.050 744.600 ;
        RECT 694.950 742.950 697.050 743.400 ;
        RECT 700.950 742.950 703.050 743.400 ;
        RECT 706.950 744.600 709.050 745.050 ;
        RECT 742.950 744.600 745.050 745.050 ;
        RECT 706.950 743.400 745.050 744.600 ;
        RECT 706.950 742.950 709.050 743.400 ;
        RECT 742.950 742.950 745.050 743.400 ;
        RECT 754.950 744.600 757.050 745.050 ;
        RECT 775.950 744.600 778.050 745.050 ;
        RECT 754.950 743.400 778.050 744.600 ;
        RECT 754.950 742.950 757.050 743.400 ;
        RECT 775.950 742.950 778.050 743.400 ;
        RECT 781.950 744.600 784.050 745.050 ;
        RECT 787.950 744.600 790.050 745.050 ;
        RECT 781.950 743.400 790.050 744.600 ;
        RECT 781.950 742.950 784.050 743.400 ;
        RECT 787.950 742.950 790.050 743.400 ;
        RECT 811.950 744.600 814.050 745.050 ;
        RECT 829.950 744.600 832.050 745.050 ;
        RECT 811.950 743.400 832.050 744.600 ;
        RECT 811.950 742.950 814.050 743.400 ;
        RECT 829.950 742.950 832.050 743.400 ;
        RECT 835.950 744.600 838.050 745.050 ;
        RECT 844.950 744.600 847.050 745.050 ;
        RECT 835.950 743.400 847.050 744.600 ;
        RECT 835.950 742.950 838.050 743.400 ;
        RECT 844.950 742.950 847.050 743.400 ;
        RECT 511.950 741.600 514.050 742.050 ;
        RECT 643.950 741.600 646.050 742.050 ;
        RECT 511.950 740.400 646.050 741.600 ;
        RECT 511.950 739.950 514.050 740.400 ;
        RECT 643.950 739.950 646.050 740.400 ;
        RECT 709.950 741.600 712.050 742.050 ;
        RECT 751.950 741.600 754.050 742.050 ;
        RECT 844.950 741.600 847.050 742.050 ;
        RECT 709.950 740.400 847.050 741.600 ;
        RECT 709.950 739.950 712.050 740.400 ;
        RECT 751.950 739.950 754.050 740.400 ;
        RECT 844.950 739.950 847.050 740.400 ;
        RECT 490.950 738.600 493.050 739.050 ;
        RECT 488.400 737.400 493.050 738.600 ;
        RECT 424.950 736.950 427.050 737.400 ;
        RECT 472.950 736.950 475.050 737.400 ;
        RECT 490.950 736.950 493.050 737.400 ;
        RECT 571.950 738.600 574.050 739.050 ;
        RECT 640.950 738.600 643.050 739.050 ;
        RECT 661.950 738.600 664.050 739.050 ;
        RECT 571.950 737.400 664.050 738.600 ;
        RECT 571.950 736.950 574.050 737.400 ;
        RECT 640.950 736.950 643.050 737.400 ;
        RECT 661.950 736.950 664.050 737.400 ;
        RECT 667.950 738.600 670.050 739.050 ;
        RECT 730.950 738.600 733.050 739.050 ;
        RECT 733.950 738.600 736.050 739.050 ;
        RECT 667.950 737.400 736.050 738.600 ;
        RECT 667.950 736.950 670.050 737.400 ;
        RECT 730.950 736.950 733.050 737.400 ;
        RECT 733.950 736.950 736.050 737.400 ;
        RECT 739.950 738.600 742.050 739.050 ;
        RECT 745.950 738.600 748.050 739.050 ;
        RECT 739.950 737.400 748.050 738.600 ;
        RECT 739.950 736.950 742.050 737.400 ;
        RECT 745.950 736.950 748.050 737.400 ;
        RECT 760.950 738.600 763.050 739.050 ;
        RECT 772.950 738.600 775.050 739.050 ;
        RECT 802.950 738.600 805.050 739.050 ;
        RECT 760.950 737.400 805.050 738.600 ;
        RECT 760.950 736.950 763.050 737.400 ;
        RECT 772.950 736.950 775.050 737.400 ;
        RECT 802.950 736.950 805.050 737.400 ;
        RECT 13.950 735.600 16.050 736.050 ;
        RECT 31.950 735.600 34.050 736.050 ;
        RECT 43.950 735.600 46.050 736.050 ;
        RECT 13.950 734.400 46.050 735.600 ;
        RECT 13.950 733.950 16.050 734.400 ;
        RECT 31.950 733.950 34.050 734.400 ;
        RECT 43.950 733.950 46.050 734.400 ;
        RECT 79.950 735.600 82.050 736.050 ;
        RECT 91.950 735.600 94.050 736.050 ;
        RECT 79.950 734.400 94.050 735.600 ;
        RECT 79.950 733.950 82.050 734.400 ;
        RECT 91.950 733.950 94.050 734.400 ;
        RECT 103.950 735.600 106.050 736.050 ;
        RECT 136.950 735.600 139.050 736.050 ;
        RECT 103.950 734.400 139.050 735.600 ;
        RECT 236.400 735.600 237.600 736.950 ;
        RECT 253.950 735.600 256.050 736.050 ;
        RECT 236.400 734.400 256.050 735.600 ;
        RECT 103.950 733.950 106.050 734.400 ;
        RECT 136.950 733.950 139.050 734.400 ;
        RECT 253.950 733.950 256.050 734.400 ;
        RECT 436.950 735.600 439.050 736.050 ;
        RECT 496.950 735.600 499.050 736.050 ;
        RECT 436.950 734.400 499.050 735.600 ;
        RECT 436.950 733.950 439.050 734.400 ;
        RECT 496.950 733.950 499.050 734.400 ;
        RECT 544.950 735.600 547.050 736.050 ;
        RECT 619.950 735.600 622.050 736.050 ;
        RECT 544.950 734.400 622.050 735.600 ;
        RECT 544.950 733.950 547.050 734.400 ;
        RECT 619.950 733.950 622.050 734.400 ;
        RECT 655.950 735.600 658.050 736.050 ;
        RECT 661.950 735.600 664.050 736.050 ;
        RECT 655.950 734.400 664.050 735.600 ;
        RECT 655.950 733.950 658.050 734.400 ;
        RECT 661.950 733.950 664.050 734.400 ;
        RECT 16.950 732.600 19.050 733.050 ;
        RECT 28.950 732.600 31.050 733.050 ;
        RECT 16.950 731.400 31.050 732.600 ;
        RECT 16.950 730.950 19.050 731.400 ;
        RECT 28.950 730.950 31.050 731.400 ;
        RECT 220.950 732.600 223.050 733.050 ;
        RECT 283.950 732.600 286.050 733.050 ;
        RECT 220.950 731.400 286.050 732.600 ;
        RECT 220.950 730.950 223.050 731.400 ;
        RECT 283.950 730.950 286.050 731.400 ;
        RECT 397.950 732.600 400.050 733.050 ;
        RECT 505.950 732.600 508.050 733.050 ;
        RECT 397.950 731.400 508.050 732.600 ;
        RECT 397.950 730.950 400.050 731.400 ;
        RECT 505.950 730.950 508.050 731.400 ;
        RECT 532.950 732.600 535.050 733.050 ;
        RECT 628.950 732.600 631.050 733.050 ;
        RECT 532.950 731.400 631.050 732.600 ;
        RECT 532.950 730.950 535.050 731.400 ;
        RECT 628.950 730.950 631.050 731.400 ;
        RECT 688.950 732.600 691.050 733.050 ;
        RECT 733.950 732.600 736.050 733.050 ;
        RECT 826.950 732.600 829.050 733.050 ;
        RECT 688.950 731.400 829.050 732.600 ;
        RECT 688.950 730.950 691.050 731.400 ;
        RECT 733.950 730.950 736.050 731.400 ;
        RECT 826.950 730.950 829.050 731.400 ;
        RECT 391.950 729.600 394.050 730.050 ;
        RECT 406.950 729.600 409.050 730.050 ;
        RECT 448.950 729.600 451.050 730.050 ;
        RECT 391.950 728.400 451.050 729.600 ;
        RECT 391.950 727.950 394.050 728.400 ;
        RECT 406.950 727.950 409.050 728.400 ;
        RECT 448.950 727.950 451.050 728.400 ;
        RECT 493.950 729.600 496.050 730.050 ;
        RECT 679.950 729.600 682.050 730.050 ;
        RECT 703.950 729.600 706.050 730.050 ;
        RECT 493.950 728.400 706.050 729.600 ;
        RECT 493.950 727.950 496.050 728.400 ;
        RECT 679.950 727.950 682.050 728.400 ;
        RECT 703.950 727.950 706.050 728.400 ;
        RECT 724.950 729.600 727.050 730.050 ;
        RECT 811.950 729.600 814.050 730.050 ;
        RECT 724.950 728.400 814.050 729.600 ;
        RECT 724.950 727.950 727.050 728.400 ;
        RECT 811.950 727.950 814.050 728.400 ;
        RECT 463.950 726.600 466.050 727.050 ;
        RECT 526.950 726.600 529.050 727.050 ;
        RECT 463.950 725.400 529.050 726.600 ;
        RECT 463.950 724.950 466.050 725.400 ;
        RECT 526.950 724.950 529.050 725.400 ;
        RECT 502.950 723.600 505.050 724.050 ;
        RECT 682.950 723.600 685.050 724.050 ;
        RECT 694.950 723.600 697.050 724.050 ;
        RECT 502.950 722.400 697.050 723.600 ;
        RECT 502.950 721.950 505.050 722.400 ;
        RECT 682.950 721.950 685.050 722.400 ;
        RECT 694.950 721.950 697.050 722.400 ;
        RECT 409.950 720.600 412.050 721.050 ;
        RECT 535.950 720.600 538.050 721.050 ;
        RECT 409.950 719.400 538.050 720.600 ;
        RECT 409.950 718.950 412.050 719.400 ;
        RECT 535.950 718.950 538.050 719.400 ;
        RECT 127.950 717.600 130.050 718.050 ;
        RECT 154.950 717.600 157.050 718.050 ;
        RECT 271.950 717.600 274.050 718.050 ;
        RECT 622.950 717.600 625.050 718.050 ;
        RECT 127.950 716.400 625.050 717.600 ;
        RECT 127.950 715.950 130.050 716.400 ;
        RECT 154.950 715.950 157.050 716.400 ;
        RECT 271.950 715.950 274.050 716.400 ;
        RECT 622.950 715.950 625.050 716.400 ;
        RECT 160.950 708.600 163.050 709.050 ;
        RECT 175.950 708.600 178.050 709.050 ;
        RECT 340.950 708.600 343.050 709.050 ;
        RECT 160.950 707.400 343.050 708.600 ;
        RECT 160.950 706.950 163.050 707.400 ;
        RECT 175.950 706.950 178.050 707.400 ;
        RECT 340.950 706.950 343.050 707.400 ;
        RECT 343.950 708.600 346.050 709.050 ;
        RECT 364.950 708.600 367.050 709.050 ;
        RECT 343.950 707.400 367.050 708.600 ;
        RECT 343.950 706.950 346.050 707.400 ;
        RECT 364.950 706.950 367.050 707.400 ;
        RECT 454.950 708.600 457.050 709.050 ;
        RECT 508.950 708.600 511.050 709.050 ;
        RECT 454.950 707.400 511.050 708.600 ;
        RECT 454.950 706.950 457.050 707.400 ;
        RECT 508.950 706.950 511.050 707.400 ;
        RECT 847.950 708.600 850.050 709.050 ;
        RECT 871.950 708.600 874.050 709.050 ;
        RECT 847.950 707.400 874.050 708.600 ;
        RECT 847.950 706.950 850.050 707.400 ;
        RECT 871.950 706.950 874.050 707.400 ;
        RECT 64.950 705.600 67.050 706.050 ;
        RECT 70.950 705.600 73.050 706.050 ;
        RECT 64.950 704.400 73.050 705.600 ;
        RECT 64.950 703.950 67.050 704.400 ;
        RECT 70.950 703.950 73.050 704.400 ;
        RECT 112.950 705.600 115.050 706.050 ;
        RECT 139.950 705.600 142.050 706.050 ;
        RECT 175.950 705.600 178.050 706.050 ;
        RECT 112.950 704.400 120.600 705.600 ;
        RECT 112.950 703.950 115.050 704.400 ;
        RECT 13.950 702.600 16.050 703.050 ;
        RECT 34.950 702.600 37.050 703.050 ;
        RECT 13.950 701.400 37.050 702.600 ;
        RECT 13.950 700.950 16.050 701.400 ;
        RECT 34.950 700.950 37.050 701.400 ;
        RECT 52.950 702.600 55.050 703.050 ;
        RECT 88.950 702.600 91.050 703.050 ;
        RECT 52.950 701.400 91.050 702.600 ;
        RECT 52.950 700.950 55.050 701.400 ;
        RECT 88.950 700.950 91.050 701.400 ;
        RECT 115.950 700.950 118.050 703.050 ;
        RECT 119.400 702.600 120.600 704.400 ;
        RECT 139.950 704.400 178.050 705.600 ;
        RECT 139.950 703.950 142.050 704.400 ;
        RECT 175.950 703.950 178.050 704.400 ;
        RECT 190.950 705.600 193.050 706.050 ;
        RECT 217.950 705.600 220.050 706.050 ;
        RECT 190.950 704.400 220.050 705.600 ;
        RECT 190.950 703.950 193.050 704.400 ;
        RECT 217.950 703.950 220.050 704.400 ;
        RECT 274.950 705.600 277.050 706.050 ;
        RECT 295.950 705.600 298.050 706.050 ;
        RECT 310.950 705.600 313.050 706.050 ;
        RECT 274.950 704.400 313.050 705.600 ;
        RECT 274.950 703.950 277.050 704.400 ;
        RECT 295.950 703.950 298.050 704.400 ;
        RECT 310.950 703.950 313.050 704.400 ;
        RECT 328.950 705.600 331.050 706.050 ;
        RECT 370.950 705.600 373.050 706.050 ;
        RECT 436.950 705.600 439.050 706.050 ;
        RECT 445.950 705.600 448.050 706.050 ;
        RECT 532.950 705.600 535.050 706.050 ;
        RECT 328.950 704.400 396.600 705.600 ;
        RECT 328.950 703.950 331.050 704.400 ;
        RECT 370.950 703.950 373.050 704.400 ;
        RECT 395.400 703.050 396.600 704.400 ;
        RECT 436.950 704.400 535.050 705.600 ;
        RECT 436.950 703.950 439.050 704.400 ;
        RECT 445.950 703.950 448.050 704.400 ;
        RECT 532.950 703.950 535.050 704.400 ;
        RECT 589.950 705.600 592.050 706.050 ;
        RECT 616.950 705.600 619.050 706.050 ;
        RECT 589.950 704.400 619.050 705.600 ;
        RECT 589.950 703.950 592.050 704.400 ;
        RECT 616.950 703.950 619.050 704.400 ;
        RECT 631.950 705.600 634.050 706.050 ;
        RECT 643.950 705.600 646.050 706.050 ;
        RECT 631.950 704.400 646.050 705.600 ;
        RECT 631.950 703.950 634.050 704.400 ;
        RECT 643.950 703.950 646.050 704.400 ;
        RECT 649.950 705.600 652.050 706.050 ;
        RECT 664.950 705.600 667.050 706.050 ;
        RECT 649.950 704.400 667.050 705.600 ;
        RECT 649.950 703.950 652.050 704.400 ;
        RECT 664.950 703.950 667.050 704.400 ;
        RECT 670.950 705.600 673.050 706.050 ;
        RECT 679.950 705.600 682.050 706.050 ;
        RECT 685.950 705.600 688.050 706.050 ;
        RECT 670.950 704.400 688.050 705.600 ;
        RECT 670.950 703.950 673.050 704.400 ;
        RECT 679.950 703.950 682.050 704.400 ;
        RECT 685.950 703.950 688.050 704.400 ;
        RECT 748.950 705.600 751.050 706.050 ;
        RECT 805.950 705.600 808.050 706.050 ;
        RECT 748.950 704.400 808.050 705.600 ;
        RECT 748.950 703.950 751.050 704.400 ;
        RECT 805.950 703.950 808.050 704.400 ;
        RECT 820.950 705.600 823.050 706.050 ;
        RECT 835.950 705.600 838.050 706.050 ;
        RECT 820.950 704.400 838.050 705.600 ;
        RECT 820.950 703.950 823.050 704.400 ;
        RECT 835.950 703.950 838.050 704.400 ;
        RECT 130.950 702.600 133.050 703.050 ;
        RECT 163.950 702.600 166.050 703.050 ;
        RECT 119.400 701.400 166.050 702.600 ;
        RECT 130.950 700.950 133.050 701.400 ;
        RECT 163.950 700.950 166.050 701.400 ;
        RECT 196.950 700.950 199.050 703.050 ;
        RECT 202.950 702.600 205.050 703.050 ;
        RECT 208.950 702.600 211.050 703.050 ;
        RECT 202.950 701.400 211.050 702.600 ;
        RECT 202.950 700.950 205.050 701.400 ;
        RECT 208.950 700.950 211.050 701.400 ;
        RECT 223.950 702.600 226.050 703.050 ;
        RECT 238.950 702.600 241.050 703.050 ;
        RECT 223.950 701.400 241.050 702.600 ;
        RECT 223.950 700.950 226.050 701.400 ;
        RECT 238.950 700.950 241.050 701.400 ;
        RECT 280.950 702.600 283.050 703.050 ;
        RECT 289.950 702.600 292.050 703.050 ;
        RECT 346.950 702.600 349.050 703.050 ;
        RECT 280.950 701.400 349.050 702.600 ;
        RECT 280.950 700.950 283.050 701.400 ;
        RECT 289.950 700.950 292.050 701.400 ;
        RECT 346.950 700.950 349.050 701.400 ;
        RECT 352.950 702.600 355.050 703.050 ;
        RECT 361.950 702.600 364.050 703.050 ;
        RECT 352.950 701.400 364.050 702.600 ;
        RECT 352.950 700.950 355.050 701.400 ;
        RECT 361.950 700.950 364.050 701.400 ;
        RECT 367.950 702.600 370.050 703.050 ;
        RECT 373.950 702.600 376.050 703.050 ;
        RECT 388.950 702.600 391.050 703.050 ;
        RECT 367.950 701.400 391.050 702.600 ;
        RECT 367.950 700.950 370.050 701.400 ;
        RECT 373.950 700.950 376.050 701.400 ;
        RECT 388.950 700.950 391.050 701.400 ;
        RECT 394.950 700.950 397.050 703.050 ;
        RECT 412.950 702.600 415.050 703.050 ;
        RECT 463.950 702.600 466.050 703.050 ;
        RECT 412.950 701.400 466.050 702.600 ;
        RECT 412.950 700.950 415.050 701.400 ;
        RECT 463.950 700.950 466.050 701.400 ;
        RECT 475.950 702.600 478.050 703.050 ;
        RECT 490.950 702.600 493.050 703.050 ;
        RECT 475.950 701.400 493.050 702.600 ;
        RECT 475.950 700.950 478.050 701.400 ;
        RECT 490.950 700.950 493.050 701.400 ;
        RECT 535.950 702.600 538.050 703.050 ;
        RECT 544.950 702.600 547.050 703.050 ;
        RECT 535.950 701.400 547.050 702.600 ;
        RECT 535.950 700.950 538.050 701.400 ;
        RECT 544.950 700.950 547.050 701.400 ;
        RECT 550.950 702.600 553.050 703.050 ;
        RECT 595.950 702.600 598.050 703.050 ;
        RECT 646.950 702.600 649.050 703.050 ;
        RECT 550.950 701.400 567.600 702.600 ;
        RECT 550.950 700.950 553.050 701.400 ;
        RECT 67.950 699.600 70.050 700.050 ;
        RECT 73.950 699.600 76.050 700.050 ;
        RECT 67.950 698.400 76.050 699.600 ;
        RECT 67.950 697.950 70.050 698.400 ;
        RECT 73.950 697.950 76.050 698.400 ;
        RECT 91.950 699.600 94.050 700.050 ;
        RECT 103.950 699.600 106.050 700.050 ;
        RECT 91.950 698.400 106.050 699.600 ;
        RECT 91.950 697.950 94.050 698.400 ;
        RECT 103.950 697.950 106.050 698.400 ;
        RECT 109.950 699.600 112.050 700.050 ;
        RECT 116.400 699.600 117.600 700.950 ;
        RECT 109.950 698.400 117.600 699.600 ;
        RECT 121.950 699.600 124.050 700.050 ;
        RECT 136.950 699.600 139.050 700.050 ;
        RECT 121.950 698.400 139.050 699.600 ;
        RECT 109.950 697.950 112.050 698.400 ;
        RECT 121.950 697.950 124.050 698.400 ;
        RECT 136.950 697.950 139.050 698.400 ;
        RECT 172.950 699.600 175.050 700.050 ;
        RECT 187.950 699.600 190.050 700.050 ;
        RECT 172.950 698.400 190.050 699.600 ;
        RECT 172.950 697.950 175.050 698.400 ;
        RECT 187.950 697.950 190.050 698.400 ;
        RECT 55.950 696.600 58.050 697.050 ;
        RECT 79.950 696.600 82.050 697.050 ;
        RECT 55.950 695.400 82.050 696.600 ;
        RECT 55.950 694.950 58.050 695.400 ;
        RECT 79.950 694.950 82.050 695.400 ;
        RECT 106.950 696.600 109.050 697.050 ;
        RECT 112.950 696.600 115.050 697.050 ;
        RECT 106.950 695.400 115.050 696.600 ;
        RECT 106.950 694.950 109.050 695.400 ;
        RECT 112.950 694.950 115.050 695.400 ;
        RECT 115.950 696.600 118.050 697.050 ;
        RECT 133.950 696.600 136.050 697.050 ;
        RECT 115.950 695.400 136.050 696.600 ;
        RECT 115.950 694.950 118.050 695.400 ;
        RECT 133.950 694.950 136.050 695.400 ;
        RECT 181.950 696.600 184.050 697.050 ;
        RECT 190.950 696.600 193.050 697.050 ;
        RECT 181.950 695.400 193.050 696.600 ;
        RECT 197.400 696.600 198.600 700.950 ;
        RECT 566.400 700.050 567.600 701.400 ;
        RECT 595.950 701.400 649.050 702.600 ;
        RECT 595.950 700.950 598.050 701.400 ;
        RECT 646.950 700.950 649.050 701.400 ;
        RECT 691.950 702.600 694.050 703.050 ;
        RECT 700.950 702.600 703.050 703.050 ;
        RECT 691.950 701.400 703.050 702.600 ;
        RECT 691.950 700.950 694.050 701.400 ;
        RECT 700.950 700.950 703.050 701.400 ;
        RECT 745.950 702.600 748.050 703.050 ;
        RECT 763.950 702.600 766.050 703.050 ;
        RECT 745.950 701.400 766.050 702.600 ;
        RECT 745.950 700.950 748.050 701.400 ;
        RECT 763.950 700.950 766.050 701.400 ;
        RECT 769.950 702.600 772.050 703.050 ;
        RECT 775.950 702.600 778.050 703.050 ;
        RECT 769.950 701.400 778.050 702.600 ;
        RECT 769.950 700.950 772.050 701.400 ;
        RECT 775.950 700.950 778.050 701.400 ;
        RECT 805.950 702.600 808.050 703.050 ;
        RECT 826.950 702.600 829.050 703.050 ;
        RECT 805.950 701.400 829.050 702.600 ;
        RECT 805.950 700.950 808.050 701.400 ;
        RECT 826.950 700.950 829.050 701.400 ;
        RECT 262.950 699.600 265.050 700.050 ;
        RECT 265.950 699.600 268.050 700.050 ;
        RECT 319.950 699.600 322.050 700.050 ;
        RECT 262.950 698.400 322.050 699.600 ;
        RECT 262.950 697.950 265.050 698.400 ;
        RECT 265.950 697.950 268.050 698.400 ;
        RECT 319.950 697.950 322.050 698.400 ;
        RECT 343.950 699.600 346.050 700.050 ;
        RECT 349.950 699.600 352.050 700.050 ;
        RECT 343.950 698.400 352.050 699.600 ;
        RECT 343.950 697.950 346.050 698.400 ;
        RECT 349.950 697.950 352.050 698.400 ;
        RECT 391.950 699.600 394.050 700.050 ;
        RECT 424.950 699.600 427.050 700.050 ;
        RECT 391.950 698.400 427.050 699.600 ;
        RECT 391.950 697.950 394.050 698.400 ;
        RECT 424.950 697.950 427.050 698.400 ;
        RECT 439.950 699.600 442.050 700.050 ;
        RECT 451.950 699.600 454.050 700.050 ;
        RECT 439.950 698.400 454.050 699.600 ;
        RECT 439.950 697.950 442.050 698.400 ;
        RECT 451.950 697.950 454.050 698.400 ;
        RECT 466.950 699.600 469.050 700.050 ;
        RECT 472.950 699.600 475.050 700.050 ;
        RECT 466.950 698.400 475.050 699.600 ;
        RECT 466.950 697.950 469.050 698.400 ;
        RECT 472.950 697.950 475.050 698.400 ;
        RECT 487.950 699.600 490.050 700.050 ;
        RECT 493.950 699.600 496.050 700.050 ;
        RECT 487.950 698.400 496.050 699.600 ;
        RECT 487.950 697.950 490.050 698.400 ;
        RECT 493.950 697.950 496.050 698.400 ;
        RECT 565.950 697.950 568.050 700.050 ;
        RECT 592.950 699.600 595.050 700.050 ;
        RECT 613.950 699.600 616.050 700.050 ;
        RECT 592.950 698.400 616.050 699.600 ;
        RECT 592.950 697.950 595.050 698.400 ;
        RECT 613.950 697.950 616.050 698.400 ;
        RECT 631.950 699.600 634.050 700.050 ;
        RECT 652.950 699.600 655.050 700.050 ;
        RECT 631.950 698.400 655.050 699.600 ;
        RECT 631.950 697.950 634.050 698.400 ;
        RECT 652.950 697.950 655.050 698.400 ;
        RECT 655.950 699.600 658.050 700.050 ;
        RECT 682.950 699.600 685.050 700.050 ;
        RECT 655.950 698.400 685.050 699.600 ;
        RECT 655.950 697.950 658.050 698.400 ;
        RECT 682.950 697.950 685.050 698.400 ;
        RECT 688.950 699.600 691.050 700.050 ;
        RECT 697.950 699.600 700.050 700.050 ;
        RECT 688.950 698.400 700.050 699.600 ;
        RECT 688.950 697.950 691.050 698.400 ;
        RECT 697.950 697.950 700.050 698.400 ;
        RECT 700.950 699.600 703.050 700.050 ;
        RECT 706.950 699.600 709.050 700.050 ;
        RECT 700.950 698.400 709.050 699.600 ;
        RECT 700.950 697.950 703.050 698.400 ;
        RECT 706.950 697.950 709.050 698.400 ;
        RECT 766.950 699.600 769.050 700.050 ;
        RECT 787.950 699.600 790.050 700.050 ;
        RECT 766.950 698.400 790.050 699.600 ;
        RECT 766.950 697.950 769.050 698.400 ;
        RECT 787.950 697.950 790.050 698.400 ;
        RECT 814.950 699.600 817.050 700.050 ;
        RECT 823.950 699.600 826.050 700.050 ;
        RECT 814.950 698.400 826.050 699.600 ;
        RECT 814.950 697.950 817.050 698.400 ;
        RECT 823.950 697.950 826.050 698.400 ;
        RECT 865.950 699.600 868.050 700.050 ;
        RECT 883.950 699.600 886.050 700.050 ;
        RECT 865.950 698.400 886.050 699.600 ;
        RECT 865.950 697.950 868.050 698.400 ;
        RECT 883.950 697.950 886.050 698.400 ;
        RECT 202.950 696.600 205.050 697.050 ;
        RECT 197.400 695.400 205.050 696.600 ;
        RECT 181.950 694.950 184.050 695.400 ;
        RECT 190.950 694.950 193.050 695.400 ;
        RECT 202.950 694.950 205.050 695.400 ;
        RECT 241.950 696.600 244.050 697.050 ;
        RECT 259.950 696.600 262.050 697.050 ;
        RECT 241.950 695.400 262.050 696.600 ;
        RECT 241.950 694.950 244.050 695.400 ;
        RECT 259.950 694.950 262.050 695.400 ;
        RECT 316.950 696.600 319.050 697.050 ;
        RECT 352.950 696.600 355.050 697.050 ;
        RECT 316.950 695.400 355.050 696.600 ;
        RECT 316.950 694.950 319.050 695.400 ;
        RECT 352.950 694.950 355.050 695.400 ;
        RECT 424.950 696.600 427.050 697.050 ;
        RECT 430.950 696.600 433.050 697.050 ;
        RECT 424.950 695.400 433.050 696.600 ;
        RECT 424.950 694.950 427.050 695.400 ;
        RECT 430.950 694.950 433.050 695.400 ;
        RECT 433.950 696.600 436.050 697.050 ;
        RECT 442.950 696.600 445.050 697.050 ;
        RECT 433.950 695.400 445.050 696.600 ;
        RECT 433.950 694.950 436.050 695.400 ;
        RECT 442.950 694.950 445.050 695.400 ;
        RECT 490.950 696.600 493.050 697.050 ;
        RECT 496.950 696.600 499.050 697.050 ;
        RECT 490.950 695.400 499.050 696.600 ;
        RECT 490.950 694.950 493.050 695.400 ;
        RECT 496.950 694.950 499.050 695.400 ;
        RECT 514.950 696.600 517.050 697.050 ;
        RECT 520.950 696.600 523.050 697.050 ;
        RECT 514.950 695.400 523.050 696.600 ;
        RECT 514.950 694.950 517.050 695.400 ;
        RECT 520.950 694.950 523.050 695.400 ;
        RECT 568.950 696.600 571.050 697.050 ;
        RECT 586.950 696.600 589.050 697.050 ;
        RECT 568.950 695.400 589.050 696.600 ;
        RECT 568.950 694.950 571.050 695.400 ;
        RECT 586.950 694.950 589.050 695.400 ;
        RECT 682.950 696.600 685.050 697.050 ;
        RECT 829.950 696.600 832.050 697.050 ;
        RECT 682.950 695.400 832.050 696.600 ;
        RECT 682.950 694.950 685.050 695.400 ;
        RECT 829.950 694.950 832.050 695.400 ;
        RECT 871.950 696.600 874.050 697.050 ;
        RECT 877.950 696.600 880.050 697.050 ;
        RECT 871.950 695.400 880.050 696.600 ;
        RECT 871.950 694.950 874.050 695.400 ;
        RECT 877.950 694.950 880.050 695.400 ;
        RECT 85.950 693.600 88.050 694.050 ;
        RECT 148.950 693.600 151.050 694.050 ;
        RECT 85.950 692.400 151.050 693.600 ;
        RECT 85.950 691.950 88.050 692.400 ;
        RECT 148.950 691.950 151.050 692.400 ;
        RECT 220.950 693.600 223.050 694.050 ;
        RECT 253.950 693.600 256.050 694.050 ;
        RECT 220.950 692.400 256.050 693.600 ;
        RECT 220.950 691.950 223.050 692.400 ;
        RECT 253.950 691.950 256.050 692.400 ;
        RECT 256.950 693.600 259.050 694.050 ;
        RECT 274.950 693.600 277.050 694.050 ;
        RECT 256.950 692.400 277.050 693.600 ;
        RECT 256.950 691.950 259.050 692.400 ;
        RECT 274.950 691.950 277.050 692.400 ;
        RECT 307.950 693.600 310.050 694.050 ;
        RECT 325.950 693.600 328.050 694.050 ;
        RECT 307.950 692.400 328.050 693.600 ;
        RECT 307.950 691.950 310.050 692.400 ;
        RECT 325.950 691.950 328.050 692.400 ;
        RECT 346.950 693.600 349.050 694.050 ;
        RECT 406.950 693.600 409.050 694.050 ;
        RECT 346.950 692.400 409.050 693.600 ;
        RECT 346.950 691.950 349.050 692.400 ;
        RECT 406.950 691.950 409.050 692.400 ;
        RECT 421.950 693.600 424.050 694.050 ;
        RECT 445.950 693.600 448.050 694.050 ;
        RECT 421.950 692.400 448.050 693.600 ;
        RECT 421.950 691.950 424.050 692.400 ;
        RECT 445.950 691.950 448.050 692.400 ;
        RECT 547.950 693.600 550.050 694.050 ;
        RECT 610.950 693.600 613.050 694.050 ;
        RECT 547.950 692.400 613.050 693.600 ;
        RECT 547.950 691.950 550.050 692.400 ;
        RECT 610.950 691.950 613.050 692.400 ;
        RECT 670.950 693.600 673.050 694.050 ;
        RECT 694.950 693.600 697.050 694.050 ;
        RECT 670.950 692.400 697.050 693.600 ;
        RECT 670.950 691.950 673.050 692.400 ;
        RECT 694.950 691.950 697.050 692.400 ;
        RECT 811.950 693.600 814.050 694.050 ;
        RECT 817.950 693.600 820.050 694.050 ;
        RECT 811.950 692.400 820.050 693.600 ;
        RECT 811.950 691.950 814.050 692.400 ;
        RECT 817.950 691.950 820.050 692.400 ;
        RECT 829.950 693.600 832.050 694.050 ;
        RECT 844.950 693.600 847.050 694.050 ;
        RECT 829.950 692.400 847.050 693.600 ;
        RECT 829.950 691.950 832.050 692.400 ;
        RECT 844.950 691.950 847.050 692.400 ;
        RECT 457.950 690.600 460.050 691.050 ;
        RECT 469.950 690.600 472.050 691.050 ;
        RECT 583.950 690.600 586.050 691.050 ;
        RECT 457.950 689.400 586.050 690.600 ;
        RECT 457.950 688.950 460.050 689.400 ;
        RECT 469.950 688.950 472.050 689.400 ;
        RECT 583.950 688.950 586.050 689.400 ;
        RECT 619.950 690.600 622.050 691.050 ;
        RECT 712.950 690.600 715.050 691.050 ;
        RECT 754.950 690.600 757.050 691.050 ;
        RECT 793.950 690.600 796.050 691.050 ;
        RECT 796.950 690.600 799.050 691.050 ;
        RECT 847.950 690.600 850.050 691.050 ;
        RECT 619.950 689.400 850.050 690.600 ;
        RECT 619.950 688.950 622.050 689.400 ;
        RECT 712.950 688.950 715.050 689.400 ;
        RECT 754.950 688.950 757.050 689.400 ;
        RECT 793.950 688.950 796.050 689.400 ;
        RECT 796.950 688.950 799.050 689.400 ;
        RECT 847.950 688.950 850.050 689.400 ;
        RECT 244.950 687.600 247.050 688.050 ;
        RECT 250.950 687.600 253.050 688.050 ;
        RECT 244.950 686.400 253.050 687.600 ;
        RECT 244.950 685.950 247.050 686.400 ;
        RECT 250.950 685.950 253.050 686.400 ;
        RECT 739.950 687.600 742.050 688.050 ;
        RECT 772.950 687.600 775.050 688.050 ;
        RECT 739.950 686.400 775.050 687.600 ;
        RECT 739.950 685.950 742.050 686.400 ;
        RECT 772.950 685.950 775.050 686.400 ;
        RECT 778.950 687.600 781.050 688.050 ;
        RECT 793.950 687.600 796.050 688.050 ;
        RECT 778.950 686.400 796.050 687.600 ;
        RECT 778.950 685.950 781.050 686.400 ;
        RECT 793.950 685.950 796.050 686.400 ;
        RECT 856.950 687.600 859.050 688.050 ;
        RECT 862.950 687.600 865.050 688.050 ;
        RECT 856.950 686.400 865.050 687.600 ;
        RECT 856.950 685.950 859.050 686.400 ;
        RECT 862.950 685.950 865.050 686.400 ;
        RECT 247.950 684.600 250.050 685.050 ;
        RECT 286.950 684.600 289.050 685.050 ;
        RECT 247.950 683.400 289.050 684.600 ;
        RECT 247.950 682.950 250.050 683.400 ;
        RECT 286.950 682.950 289.050 683.400 ;
        RECT 385.950 684.600 388.050 685.050 ;
        RECT 403.950 684.600 406.050 685.050 ;
        RECT 385.950 683.400 406.050 684.600 ;
        RECT 385.950 682.950 388.050 683.400 ;
        RECT 403.950 682.950 406.050 683.400 ;
        RECT 478.950 684.600 481.050 685.050 ;
        RECT 517.950 684.600 520.050 685.050 ;
        RECT 568.950 684.600 571.050 685.050 ;
        RECT 478.950 683.400 571.050 684.600 ;
        RECT 478.950 682.950 481.050 683.400 ;
        RECT 517.950 682.950 520.050 683.400 ;
        RECT 568.950 682.950 571.050 683.400 ;
        RECT 718.950 684.600 721.050 685.050 ;
        RECT 742.950 684.600 745.050 685.050 ;
        RECT 718.950 683.400 745.050 684.600 ;
        RECT 718.950 682.950 721.050 683.400 ;
        RECT 742.950 682.950 745.050 683.400 ;
        RECT 202.950 681.600 205.050 682.050 ;
        RECT 301.950 681.600 304.050 682.050 ;
        RECT 202.950 680.400 304.050 681.600 ;
        RECT 202.950 679.950 205.050 680.400 ;
        RECT 301.950 679.950 304.050 680.400 ;
        RECT 355.950 681.600 358.050 682.050 ;
        RECT 382.950 681.600 385.050 682.050 ;
        RECT 355.950 680.400 385.050 681.600 ;
        RECT 355.950 679.950 358.050 680.400 ;
        RECT 382.950 679.950 385.050 680.400 ;
        RECT 562.950 681.600 565.050 682.050 ;
        RECT 592.950 681.600 595.050 682.050 ;
        RECT 562.950 680.400 595.050 681.600 ;
        RECT 562.950 679.950 565.050 680.400 ;
        RECT 592.950 679.950 595.050 680.400 ;
        RECT 724.950 681.600 727.050 682.050 ;
        RECT 757.950 681.600 760.050 682.050 ;
        RECT 724.950 680.400 760.050 681.600 ;
        RECT 724.950 679.950 727.050 680.400 ;
        RECT 757.950 679.950 760.050 680.400 ;
        RECT 154.950 678.600 157.050 679.050 ;
        RECT 235.950 678.600 238.050 679.050 ;
        RECT 154.950 677.400 238.050 678.600 ;
        RECT 154.950 676.950 157.050 677.400 ;
        RECT 235.950 676.950 238.050 677.400 ;
        RECT 349.950 678.600 352.050 679.050 ;
        RECT 361.950 678.600 364.050 679.050 ;
        RECT 436.950 678.600 439.050 679.050 ;
        RECT 349.950 677.400 439.050 678.600 ;
        RECT 349.950 676.950 352.050 677.400 ;
        RECT 361.950 676.950 364.050 677.400 ;
        RECT 436.950 676.950 439.050 677.400 ;
        RECT 481.950 678.600 484.050 679.050 ;
        RECT 514.950 678.600 517.050 679.050 ;
        RECT 481.950 677.400 517.050 678.600 ;
        RECT 481.950 676.950 484.050 677.400 ;
        RECT 514.950 676.950 517.050 677.400 ;
        RECT 7.950 675.600 10.050 676.050 ;
        RECT 52.950 675.600 55.050 676.050 ;
        RECT 7.950 674.400 55.050 675.600 ;
        RECT 7.950 673.950 10.050 674.400 ;
        RECT 52.950 673.950 55.050 674.400 ;
        RECT 67.950 675.600 70.050 676.050 ;
        RECT 73.950 675.600 76.050 676.050 ;
        RECT 67.950 674.400 76.050 675.600 ;
        RECT 67.950 673.950 70.050 674.400 ;
        RECT 73.950 673.950 76.050 674.400 ;
        RECT 337.950 675.600 340.050 676.050 ;
        RECT 385.950 675.600 388.050 676.050 ;
        RECT 397.950 675.600 400.050 676.050 ;
        RECT 337.950 674.400 400.050 675.600 ;
        RECT 337.950 673.950 340.050 674.400 ;
        RECT 385.950 673.950 388.050 674.400 ;
        RECT 397.950 673.950 400.050 674.400 ;
        RECT 409.950 675.600 412.050 676.050 ;
        RECT 466.950 675.600 469.050 676.050 ;
        RECT 409.950 674.400 469.050 675.600 ;
        RECT 409.950 673.950 412.050 674.400 ;
        RECT 466.950 673.950 469.050 674.400 ;
        RECT 487.950 675.600 490.050 676.050 ;
        RECT 544.950 675.600 547.050 676.050 ;
        RECT 487.950 674.400 547.050 675.600 ;
        RECT 487.950 673.950 490.050 674.400 ;
        RECT 544.950 673.950 547.050 674.400 ;
        RECT 574.950 675.600 577.050 676.050 ;
        RECT 598.950 675.600 601.050 676.050 ;
        RECT 574.950 674.400 601.050 675.600 ;
        RECT 574.950 673.950 577.050 674.400 ;
        RECT 598.950 673.950 601.050 674.400 ;
        RECT 625.950 675.600 628.050 676.050 ;
        RECT 637.950 675.600 640.050 676.050 ;
        RECT 625.950 674.400 640.050 675.600 ;
        RECT 625.950 673.950 628.050 674.400 ;
        RECT 637.950 673.950 640.050 674.400 ;
        RECT 667.950 675.600 670.050 676.050 ;
        RECT 682.950 675.600 685.050 676.050 ;
        RECT 667.950 674.400 685.050 675.600 ;
        RECT 667.950 673.950 670.050 674.400 ;
        RECT 682.950 673.950 685.050 674.400 ;
        RECT 685.950 675.600 688.050 676.050 ;
        RECT 715.950 675.600 718.050 676.050 ;
        RECT 685.950 674.400 718.050 675.600 ;
        RECT 685.950 673.950 688.050 674.400 ;
        RECT 715.950 673.950 718.050 674.400 ;
        RECT 751.950 675.600 754.050 676.050 ;
        RECT 760.950 675.600 763.050 676.050 ;
        RECT 751.950 674.400 763.050 675.600 ;
        RECT 751.950 673.950 754.050 674.400 ;
        RECT 760.950 673.950 763.050 674.400 ;
        RECT 28.950 672.600 31.050 673.050 ;
        RECT 11.400 671.400 31.050 672.600 ;
        RECT 11.400 666.600 12.600 671.400 ;
        RECT 28.950 670.950 31.050 671.400 ;
        RECT 37.950 670.950 40.050 673.050 ;
        RECT 40.950 672.600 43.050 673.050 ;
        RECT 82.950 672.600 85.050 673.050 ;
        RECT 40.950 671.400 85.050 672.600 ;
        RECT 40.950 670.950 43.050 671.400 ;
        RECT 82.950 670.950 85.050 671.400 ;
        RECT 106.950 672.600 109.050 673.050 ;
        RECT 127.950 672.600 130.050 673.050 ;
        RECT 106.950 671.400 130.050 672.600 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 127.950 670.950 130.050 671.400 ;
        RECT 229.950 672.600 232.050 673.050 ;
        RECT 241.950 672.600 244.050 673.050 ;
        RECT 229.950 671.400 244.050 672.600 ;
        RECT 229.950 670.950 232.050 671.400 ;
        RECT 241.950 670.950 244.050 671.400 ;
        RECT 259.950 672.600 262.050 673.050 ;
        RECT 268.950 672.600 271.050 673.050 ;
        RECT 259.950 671.400 271.050 672.600 ;
        RECT 259.950 670.950 262.050 671.400 ;
        RECT 268.950 670.950 271.050 671.400 ;
        RECT 316.950 672.600 319.050 673.050 ;
        RECT 370.950 672.600 373.050 673.050 ;
        RECT 316.950 671.400 373.050 672.600 ;
        RECT 316.950 670.950 319.050 671.400 ;
        RECT 370.950 670.950 373.050 671.400 ;
        RECT 451.950 672.600 454.050 673.050 ;
        RECT 460.950 672.600 463.050 673.050 ;
        RECT 451.950 671.400 463.050 672.600 ;
        RECT 451.950 670.950 454.050 671.400 ;
        RECT 460.950 670.950 463.050 671.400 ;
        RECT 469.950 670.950 472.050 673.050 ;
        RECT 493.950 672.600 496.050 673.050 ;
        RECT 523.950 672.600 526.050 673.050 ;
        RECT 493.950 671.400 526.050 672.600 ;
        RECT 493.950 670.950 496.050 671.400 ;
        RECT 523.950 670.950 526.050 671.400 ;
        RECT 571.950 672.600 574.050 673.050 ;
        RECT 577.950 672.600 580.050 673.050 ;
        RECT 571.950 671.400 580.050 672.600 ;
        RECT 571.950 670.950 574.050 671.400 ;
        RECT 577.950 670.950 580.050 671.400 ;
        RECT 649.950 672.600 652.050 673.050 ;
        RECT 655.950 672.600 658.050 673.050 ;
        RECT 649.950 671.400 658.050 672.600 ;
        RECT 649.950 670.950 652.050 671.400 ;
        RECT 655.950 670.950 658.050 671.400 ;
        RECT 691.950 672.600 694.050 673.050 ;
        RECT 736.950 672.600 739.050 673.050 ;
        RECT 748.950 672.600 751.050 673.050 ;
        RECT 691.950 671.400 751.050 672.600 ;
        RECT 691.950 670.950 694.050 671.400 ;
        RECT 736.950 670.950 739.050 671.400 ;
        RECT 748.950 670.950 751.050 671.400 ;
        RECT 769.950 672.600 772.050 673.050 ;
        RECT 781.950 672.600 784.050 673.050 ;
        RECT 769.950 671.400 784.050 672.600 ;
        RECT 769.950 670.950 772.050 671.400 ;
        RECT 781.950 670.950 784.050 671.400 ;
        RECT 805.950 672.600 808.050 673.050 ;
        RECT 823.950 672.600 826.050 673.050 ;
        RECT 805.950 671.400 826.050 672.600 ;
        RECT 805.950 670.950 808.050 671.400 ;
        RECT 823.950 670.950 826.050 671.400 ;
        RECT 868.950 670.950 871.050 673.050 ;
        RECT 13.950 669.600 16.050 670.050 ;
        RECT 31.950 669.600 34.050 670.050 ;
        RECT 13.950 668.400 34.050 669.600 ;
        RECT 38.400 669.600 39.600 670.950 ;
        RECT 91.950 669.600 94.050 670.050 ;
        RECT 133.950 669.600 136.050 670.050 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 38.400 668.400 48.600 669.600 ;
        RECT 13.950 667.950 16.050 668.400 ;
        RECT 31.950 667.950 34.050 668.400 ;
        RECT 28.950 666.600 31.050 667.050 ;
        RECT 11.400 665.400 31.050 666.600 ;
        RECT 28.950 664.950 31.050 665.400 ;
        RECT 34.950 666.600 37.050 667.050 ;
        RECT 43.950 666.600 46.050 667.050 ;
        RECT 34.950 665.400 46.050 666.600 ;
        RECT 47.400 666.600 48.600 668.400 ;
        RECT 91.950 668.400 111.600 669.600 ;
        RECT 91.950 667.950 94.050 668.400 ;
        RECT 110.400 667.050 111.600 668.400 ;
        RECT 133.950 668.400 163.050 669.600 ;
        RECT 133.950 667.950 136.050 668.400 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 169.950 669.600 172.050 670.050 ;
        RECT 208.950 669.600 211.050 670.050 ;
        RECT 235.950 669.600 238.050 670.050 ;
        RECT 244.950 669.600 247.050 670.050 ;
        RECT 169.950 668.400 189.600 669.600 ;
        RECT 169.950 667.950 172.050 668.400 ;
        RECT 188.400 667.050 189.600 668.400 ;
        RECT 208.950 668.400 222.600 669.600 ;
        RECT 208.950 667.950 211.050 668.400 ;
        RECT 52.950 666.600 55.050 667.050 ;
        RECT 47.400 665.400 55.050 666.600 ;
        RECT 34.950 664.950 37.050 665.400 ;
        RECT 43.950 664.950 46.050 665.400 ;
        RECT 52.950 664.950 55.050 665.400 ;
        RECT 61.950 666.600 64.050 667.050 ;
        RECT 70.950 666.600 73.050 667.050 ;
        RECT 103.950 666.600 106.050 667.050 ;
        RECT 61.950 665.400 106.050 666.600 ;
        RECT 61.950 664.950 64.050 665.400 ;
        RECT 70.950 664.950 73.050 665.400 ;
        RECT 103.950 664.950 106.050 665.400 ;
        RECT 109.950 664.950 112.050 667.050 ;
        RECT 130.950 664.950 133.050 667.050 ;
        RECT 136.950 666.600 139.050 667.050 ;
        RECT 172.950 666.600 175.050 667.050 ;
        RECT 136.950 665.400 175.050 666.600 ;
        RECT 136.950 664.950 139.050 665.400 ;
        RECT 172.950 664.950 175.050 665.400 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 199.950 666.600 202.050 667.050 ;
        RECT 205.950 666.600 208.050 667.050 ;
        RECT 199.950 665.400 208.050 666.600 ;
        RECT 199.950 664.950 202.050 665.400 ;
        RECT 205.950 664.950 208.050 665.400 ;
        RECT 211.950 666.600 214.050 667.050 ;
        RECT 217.950 666.600 220.050 667.050 ;
        RECT 211.950 665.400 220.050 666.600 ;
        RECT 221.400 666.600 222.600 668.400 ;
        RECT 235.950 668.400 247.050 669.600 ;
        RECT 235.950 667.950 238.050 668.400 ;
        RECT 244.950 667.950 247.050 668.400 ;
        RECT 271.950 669.600 274.050 670.050 ;
        RECT 295.950 669.600 298.050 670.050 ;
        RECT 271.950 668.400 298.050 669.600 ;
        RECT 271.950 667.950 274.050 668.400 ;
        RECT 295.950 667.950 298.050 668.400 ;
        RECT 379.950 669.600 382.050 670.050 ;
        RECT 388.950 669.600 391.050 670.050 ;
        RECT 442.950 669.600 445.050 670.050 ;
        RECT 379.950 668.400 445.050 669.600 ;
        RECT 379.950 667.950 382.050 668.400 ;
        RECT 388.950 667.950 391.050 668.400 ;
        RECT 442.950 667.950 445.050 668.400 ;
        RECT 448.950 669.600 451.050 670.050 ;
        RECT 470.400 669.600 471.600 670.950 ;
        RECT 448.950 668.400 471.600 669.600 ;
        RECT 529.950 669.600 532.050 670.050 ;
        RECT 541.950 669.600 544.050 670.050 ;
        RECT 529.950 668.400 544.050 669.600 ;
        RECT 448.950 667.950 451.050 668.400 ;
        RECT 529.950 667.950 532.050 668.400 ;
        RECT 541.950 667.950 544.050 668.400 ;
        RECT 601.950 669.600 604.050 670.050 ;
        RECT 616.950 669.600 619.050 670.050 ;
        RECT 601.950 668.400 619.050 669.600 ;
        RECT 601.950 667.950 604.050 668.400 ;
        RECT 616.950 667.950 619.050 668.400 ;
        RECT 622.950 669.600 625.050 670.050 ;
        RECT 643.950 669.600 646.050 670.050 ;
        RECT 622.950 668.400 646.050 669.600 ;
        RECT 622.950 667.950 625.050 668.400 ;
        RECT 643.950 667.950 646.050 668.400 ;
        RECT 652.950 669.600 655.050 670.050 ;
        RECT 658.950 669.600 661.050 670.050 ;
        RECT 652.950 668.400 661.050 669.600 ;
        RECT 652.950 667.950 655.050 668.400 ;
        RECT 658.950 667.950 661.050 668.400 ;
        RECT 679.950 669.600 682.050 670.050 ;
        RECT 697.950 669.600 700.050 670.050 ;
        RECT 679.950 668.400 700.050 669.600 ;
        RECT 679.950 667.950 682.050 668.400 ;
        RECT 697.950 667.950 700.050 668.400 ;
        RECT 745.950 669.600 748.050 670.050 ;
        RECT 760.950 669.600 763.050 670.050 ;
        RECT 745.950 668.400 763.050 669.600 ;
        RECT 745.950 667.950 748.050 668.400 ;
        RECT 760.950 667.950 763.050 668.400 ;
        RECT 784.950 669.600 787.050 670.050 ;
        RECT 799.950 669.600 802.050 670.050 ;
        RECT 784.950 668.400 802.050 669.600 ;
        RECT 784.950 667.950 787.050 668.400 ;
        RECT 799.950 667.950 802.050 668.400 ;
        RECT 841.950 669.600 844.050 670.050 ;
        RECT 859.950 669.600 862.050 670.050 ;
        RECT 841.950 668.400 862.050 669.600 ;
        RECT 841.950 667.950 844.050 668.400 ;
        RECT 859.950 667.950 862.050 668.400 ;
        RECT 226.950 666.600 229.050 667.050 ;
        RECT 221.400 665.400 229.050 666.600 ;
        RECT 211.950 664.950 214.050 665.400 ;
        RECT 217.950 664.950 220.050 665.400 ;
        RECT 226.950 664.950 229.050 665.400 ;
        RECT 232.950 664.950 235.050 667.050 ;
        RECT 277.950 666.600 280.050 667.050 ;
        RECT 298.950 666.600 301.050 667.050 ;
        RECT 277.950 665.400 301.050 666.600 ;
        RECT 277.950 664.950 280.050 665.400 ;
        RECT 298.950 664.950 301.050 665.400 ;
        RECT 496.950 666.600 499.050 667.050 ;
        RECT 505.950 666.600 508.050 667.050 ;
        RECT 496.950 665.400 508.050 666.600 ;
        RECT 496.950 664.950 499.050 665.400 ;
        RECT 505.950 664.950 508.050 665.400 ;
        RECT 547.950 666.600 550.050 667.050 ;
        RECT 637.950 666.600 640.050 667.050 ;
        RECT 547.950 665.400 640.050 666.600 ;
        RECT 547.950 664.950 550.050 665.400 ;
        RECT 637.950 664.950 640.050 665.400 ;
        RECT 706.950 666.600 709.050 667.050 ;
        RECT 757.950 666.600 760.050 667.050 ;
        RECT 706.950 665.400 760.050 666.600 ;
        RECT 706.950 664.950 709.050 665.400 ;
        RECT 757.950 664.950 760.050 665.400 ;
        RECT 763.950 666.600 766.050 667.050 ;
        RECT 772.950 666.600 775.050 667.050 ;
        RECT 805.950 666.600 808.050 667.050 ;
        RECT 844.950 666.600 847.050 667.050 ;
        RECT 763.950 665.400 847.050 666.600 ;
        RECT 763.950 664.950 766.050 665.400 ;
        RECT 772.950 664.950 775.050 665.400 ;
        RECT 805.950 664.950 808.050 665.400 ;
        RECT 844.950 664.950 847.050 665.400 ;
        RECT 862.950 666.600 865.050 667.050 ;
        RECT 869.400 666.600 870.600 670.950 ;
        RECT 862.950 665.400 870.600 666.600 ;
        RECT 862.950 664.950 865.050 665.400 ;
        RECT 28.950 663.600 31.050 664.050 ;
        RECT 40.950 663.600 43.050 664.050 ;
        RECT 28.950 662.400 43.050 663.600 ;
        RECT 28.950 661.950 31.050 662.400 ;
        RECT 40.950 661.950 43.050 662.400 ;
        RECT 79.950 663.600 82.050 664.050 ;
        RECT 103.950 663.600 106.050 664.050 ;
        RECT 131.400 663.600 132.600 664.950 ;
        RECT 79.950 662.400 132.600 663.600 ;
        RECT 206.400 663.600 207.600 664.950 ;
        RECT 208.950 663.600 211.050 664.050 ;
        RECT 206.400 662.400 211.050 663.600 ;
        RECT 79.950 661.950 82.050 662.400 ;
        RECT 103.950 661.950 106.050 662.400 ;
        RECT 208.950 661.950 211.050 662.400 ;
        RECT 229.950 663.600 232.050 664.050 ;
        RECT 233.400 663.600 234.600 664.950 ;
        RECT 229.950 662.400 234.600 663.600 ;
        RECT 298.950 663.600 301.050 664.050 ;
        RECT 373.950 663.600 376.050 664.050 ;
        RECT 376.950 663.600 379.050 664.050 ;
        RECT 298.950 662.400 379.050 663.600 ;
        RECT 229.950 661.950 232.050 662.400 ;
        RECT 298.950 661.950 301.050 662.400 ;
        RECT 373.950 661.950 376.050 662.400 ;
        RECT 376.950 661.950 379.050 662.400 ;
        RECT 400.950 663.600 403.050 664.050 ;
        RECT 421.950 663.600 424.050 664.050 ;
        RECT 439.950 663.600 442.050 664.050 ;
        RECT 400.950 662.400 442.050 663.600 ;
        RECT 400.950 661.950 403.050 662.400 ;
        RECT 421.950 661.950 424.050 662.400 ;
        RECT 439.950 661.950 442.050 662.400 ;
        RECT 484.950 663.600 487.050 664.050 ;
        RECT 517.950 663.600 520.050 664.050 ;
        RECT 484.950 662.400 520.050 663.600 ;
        RECT 484.950 661.950 487.050 662.400 ;
        RECT 517.950 661.950 520.050 662.400 ;
        RECT 562.950 663.600 565.050 664.050 ;
        RECT 586.950 663.600 589.050 664.050 ;
        RECT 640.950 663.600 643.050 664.050 ;
        RECT 562.950 662.400 643.050 663.600 ;
        RECT 562.950 661.950 565.050 662.400 ;
        RECT 586.950 661.950 589.050 662.400 ;
        RECT 640.950 661.950 643.050 662.400 ;
        RECT 709.950 663.600 712.050 664.050 ;
        RECT 739.950 663.600 742.050 664.050 ;
        RECT 709.950 662.400 742.050 663.600 ;
        RECT 709.950 661.950 712.050 662.400 ;
        RECT 739.950 661.950 742.050 662.400 ;
        RECT 763.950 663.600 766.050 664.050 ;
        RECT 796.950 663.600 799.050 664.050 ;
        RECT 763.950 662.400 799.050 663.600 ;
        RECT 763.950 661.950 766.050 662.400 ;
        RECT 796.950 661.950 799.050 662.400 ;
        RECT 31.950 660.600 34.050 661.050 ;
        RECT 43.950 660.600 46.050 661.050 ;
        RECT 31.950 659.400 46.050 660.600 ;
        RECT 31.950 658.950 34.050 659.400 ;
        RECT 43.950 658.950 46.050 659.400 ;
        RECT 115.950 660.600 118.050 661.050 ;
        RECT 166.950 660.600 169.050 661.050 ;
        RECT 115.950 659.400 169.050 660.600 ;
        RECT 115.950 658.950 118.050 659.400 ;
        RECT 166.950 658.950 169.050 659.400 ;
        RECT 604.950 660.600 607.050 661.050 ;
        RECT 622.950 660.600 625.050 661.050 ;
        RECT 604.950 659.400 625.050 660.600 ;
        RECT 604.950 658.950 607.050 659.400 ;
        RECT 622.950 658.950 625.050 659.400 ;
        RECT 715.950 660.600 718.050 661.050 ;
        RECT 733.950 660.600 736.050 661.050 ;
        RECT 715.950 659.400 736.050 660.600 ;
        RECT 715.950 658.950 718.050 659.400 ;
        RECT 733.950 658.950 736.050 659.400 ;
        RECT 736.950 660.600 739.050 661.050 ;
        RECT 751.950 660.600 754.050 661.050 ;
        RECT 736.950 659.400 754.050 660.600 ;
        RECT 736.950 658.950 739.050 659.400 ;
        RECT 751.950 658.950 754.050 659.400 ;
        RECT 772.950 660.600 775.050 661.050 ;
        RECT 790.950 660.600 793.050 661.050 ;
        RECT 772.950 659.400 793.050 660.600 ;
        RECT 772.950 658.950 775.050 659.400 ;
        RECT 790.950 658.950 793.050 659.400 ;
        RECT 553.950 657.600 556.050 658.050 ;
        RECT 688.950 657.600 691.050 658.050 ;
        RECT 553.950 656.400 691.050 657.600 ;
        RECT 553.950 655.950 556.050 656.400 ;
        RECT 688.950 655.950 691.050 656.400 ;
        RECT 727.950 657.600 730.050 658.050 ;
        RECT 778.950 657.600 781.050 658.050 ;
        RECT 727.950 656.400 781.050 657.600 ;
        RECT 727.950 655.950 730.050 656.400 ;
        RECT 778.950 655.950 781.050 656.400 ;
        RECT 16.950 654.600 19.050 655.050 ;
        RECT 43.950 654.600 46.050 655.050 ;
        RECT 16.950 653.400 46.050 654.600 ;
        RECT 16.950 652.950 19.050 653.400 ;
        RECT 43.950 652.950 46.050 653.400 ;
        RECT 193.950 651.600 196.050 652.050 ;
        RECT 205.950 651.600 208.050 652.050 ;
        RECT 193.950 650.400 208.050 651.600 ;
        RECT 193.950 649.950 196.050 650.400 ;
        RECT 205.950 649.950 208.050 650.400 ;
        RECT 775.950 651.600 778.050 652.050 ;
        RECT 808.950 651.600 811.050 652.050 ;
        RECT 775.950 650.400 811.050 651.600 ;
        RECT 775.950 649.950 778.050 650.400 ;
        RECT 808.950 649.950 811.050 650.400 ;
        RECT 55.950 648.600 58.050 649.050 ;
        RECT 88.950 648.600 91.050 649.050 ;
        RECT 106.950 648.600 109.050 649.050 ;
        RECT 157.950 648.600 160.050 649.050 ;
        RECT 193.950 648.600 196.050 649.050 ;
        RECT 55.950 647.400 196.050 648.600 ;
        RECT 55.950 646.950 58.050 647.400 ;
        RECT 88.950 646.950 91.050 647.400 ;
        RECT 106.950 646.950 109.050 647.400 ;
        RECT 157.950 646.950 160.050 647.400 ;
        RECT 193.950 646.950 196.050 647.400 ;
        RECT 283.950 648.600 286.050 649.050 ;
        RECT 406.950 648.600 409.050 649.050 ;
        RECT 283.950 647.400 409.050 648.600 ;
        RECT 283.950 646.950 286.050 647.400 ;
        RECT 406.950 646.950 409.050 647.400 ;
        RECT 481.950 645.600 484.050 646.050 ;
        RECT 490.950 645.600 493.050 646.050 ;
        RECT 481.950 644.400 493.050 645.600 ;
        RECT 481.950 643.950 484.050 644.400 ;
        RECT 490.950 643.950 493.050 644.400 ;
        RECT 859.950 645.600 862.050 646.050 ;
        RECT 865.950 645.600 868.050 646.050 ;
        RECT 859.950 644.400 868.050 645.600 ;
        RECT 859.950 643.950 862.050 644.400 ;
        RECT 865.950 643.950 868.050 644.400 ;
        RECT 76.950 642.600 79.050 643.050 ;
        RECT 109.950 642.600 112.050 643.050 ;
        RECT 76.950 641.400 112.050 642.600 ;
        RECT 76.950 640.950 79.050 641.400 ;
        RECT 109.950 640.950 112.050 641.400 ;
        RECT 97.950 639.600 100.050 640.050 ;
        RECT 130.950 639.600 133.050 640.050 ;
        RECT 97.950 638.400 133.050 639.600 ;
        RECT 97.950 637.950 100.050 638.400 ;
        RECT 130.950 637.950 133.050 638.400 ;
        RECT 493.950 639.600 496.050 640.050 ;
        RECT 499.950 639.600 502.050 640.050 ;
        RECT 493.950 638.400 502.050 639.600 ;
        RECT 493.950 637.950 496.050 638.400 ;
        RECT 499.950 637.950 502.050 638.400 ;
        RECT 802.950 636.600 805.050 637.050 ;
        RECT 811.950 636.600 814.050 637.050 ;
        RECT 802.950 635.400 814.050 636.600 ;
        RECT 802.950 634.950 805.050 635.400 ;
        RECT 811.950 634.950 814.050 635.400 ;
        RECT 829.950 636.600 832.050 637.050 ;
        RECT 850.950 636.600 853.050 637.050 ;
        RECT 829.950 635.400 853.050 636.600 ;
        RECT 829.950 634.950 832.050 635.400 ;
        RECT 850.950 634.950 853.050 635.400 ;
        RECT 13.950 633.600 16.050 634.050 ;
        RECT 19.950 633.600 22.050 634.050 ;
        RECT 37.950 633.600 40.050 634.050 ;
        RECT 13.950 632.400 40.050 633.600 ;
        RECT 13.950 631.950 16.050 632.400 ;
        RECT 19.950 631.950 22.050 632.400 ;
        RECT 37.950 631.950 40.050 632.400 ;
        RECT 43.950 633.600 46.050 634.050 ;
        RECT 58.950 633.600 61.050 634.050 ;
        RECT 43.950 632.400 61.050 633.600 ;
        RECT 43.950 631.950 46.050 632.400 ;
        RECT 58.950 631.950 61.050 632.400 ;
        RECT 73.950 633.600 76.050 634.050 ;
        RECT 97.950 633.600 100.050 634.050 ;
        RECT 124.950 633.600 127.050 634.050 ;
        RECT 151.950 633.600 154.050 634.050 ;
        RECT 73.950 632.400 154.050 633.600 ;
        RECT 73.950 631.950 76.050 632.400 ;
        RECT 97.950 631.950 100.050 632.400 ;
        RECT 124.950 631.950 127.050 632.400 ;
        RECT 151.950 631.950 154.050 632.400 ;
        RECT 241.950 633.600 244.050 634.050 ;
        RECT 265.950 633.600 268.050 634.050 ;
        RECT 430.950 633.600 433.050 634.050 ;
        RECT 448.950 633.600 451.050 634.050 ;
        RECT 241.950 632.400 264.600 633.600 ;
        RECT 241.950 631.950 244.050 632.400 ;
        RECT 263.400 631.050 264.600 632.400 ;
        RECT 265.950 632.400 285.600 633.600 ;
        RECT 265.950 631.950 268.050 632.400 ;
        RECT 284.400 631.050 285.600 632.400 ;
        RECT 430.950 632.400 451.050 633.600 ;
        RECT 430.950 631.950 433.050 632.400 ;
        RECT 448.950 631.950 451.050 632.400 ;
        RECT 463.950 633.600 466.050 634.050 ;
        RECT 472.950 633.600 475.050 634.050 ;
        RECT 463.950 632.400 475.050 633.600 ;
        RECT 463.950 631.950 466.050 632.400 ;
        RECT 472.950 631.950 475.050 632.400 ;
        RECT 475.950 633.600 478.050 634.050 ;
        RECT 511.950 633.600 514.050 634.050 ;
        RECT 475.950 632.400 514.050 633.600 ;
        RECT 475.950 631.950 478.050 632.400 ;
        RECT 511.950 631.950 514.050 632.400 ;
        RECT 523.950 633.600 526.050 634.050 ;
        RECT 565.950 633.600 568.050 634.050 ;
        RECT 523.950 632.400 568.050 633.600 ;
        RECT 523.950 631.950 526.050 632.400 ;
        RECT 565.950 631.950 568.050 632.400 ;
        RECT 628.950 633.600 631.050 634.050 ;
        RECT 637.950 633.600 640.050 634.050 ;
        RECT 628.950 632.400 640.050 633.600 ;
        RECT 628.950 631.950 631.050 632.400 ;
        RECT 637.950 631.950 640.050 632.400 ;
        RECT 664.950 633.600 667.050 634.050 ;
        RECT 670.950 633.600 673.050 634.050 ;
        RECT 688.950 633.600 691.050 634.050 ;
        RECT 700.950 633.600 703.050 634.050 ;
        RECT 712.950 633.600 715.050 634.050 ;
        RECT 664.950 632.400 691.050 633.600 ;
        RECT 664.950 631.950 667.050 632.400 ;
        RECT 670.950 631.950 673.050 632.400 ;
        RECT 688.950 631.950 691.050 632.400 ;
        RECT 692.400 632.400 715.050 633.600 ;
        RECT 19.950 630.600 22.050 631.050 ;
        RECT 25.950 630.600 28.050 631.050 ;
        RECT 19.950 629.400 28.050 630.600 ;
        RECT 19.950 628.950 22.050 629.400 ;
        RECT 25.950 628.950 28.050 629.400 ;
        RECT 34.950 630.600 37.050 631.050 ;
        RECT 37.950 630.600 40.050 631.050 ;
        RECT 55.950 630.600 58.050 631.050 ;
        RECT 73.950 630.600 76.050 631.050 ;
        RECT 34.950 629.400 76.050 630.600 ;
        RECT 34.950 628.950 37.050 629.400 ;
        RECT 37.950 628.950 40.050 629.400 ;
        RECT 55.950 628.950 58.050 629.400 ;
        RECT 73.950 628.950 76.050 629.400 ;
        RECT 79.950 630.600 82.050 631.050 ;
        RECT 91.950 630.600 94.050 631.050 ;
        RECT 94.950 630.600 97.050 631.050 ;
        RECT 79.950 629.400 97.050 630.600 ;
        RECT 79.950 628.950 82.050 629.400 ;
        RECT 91.950 628.950 94.050 629.400 ;
        RECT 94.950 628.950 97.050 629.400 ;
        RECT 100.950 630.600 103.050 631.050 ;
        RECT 106.950 630.600 109.050 631.050 ;
        RECT 100.950 629.400 109.050 630.600 ;
        RECT 100.950 628.950 103.050 629.400 ;
        RECT 106.950 628.950 109.050 629.400 ;
        RECT 127.950 630.600 130.050 631.050 ;
        RECT 139.950 630.600 142.050 631.050 ;
        RECT 154.950 630.600 157.050 631.050 ;
        RECT 172.950 630.600 175.050 631.050 ;
        RECT 127.950 629.400 153.600 630.600 ;
        RECT 127.950 628.950 130.050 629.400 ;
        RECT 139.950 628.950 142.050 629.400 ;
        RECT 28.950 627.600 31.050 628.050 ;
        RECT 34.950 627.600 37.050 628.050 ;
        RECT 28.950 626.400 37.050 627.600 ;
        RECT 28.950 625.950 31.050 626.400 ;
        RECT 34.950 625.950 37.050 626.400 ;
        RECT 58.950 627.600 61.050 628.050 ;
        RECT 70.950 627.600 73.050 628.050 ;
        RECT 58.950 626.400 73.050 627.600 ;
        RECT 152.400 627.600 153.600 629.400 ;
        RECT 154.950 629.400 175.050 630.600 ;
        RECT 154.950 628.950 157.050 629.400 ;
        RECT 172.950 628.950 175.050 629.400 ;
        RECT 196.950 630.600 199.050 631.050 ;
        RECT 217.950 630.600 220.050 631.050 ;
        RECT 196.950 629.400 220.050 630.600 ;
        RECT 196.950 628.950 199.050 629.400 ;
        RECT 217.950 628.950 220.050 629.400 ;
        RECT 223.950 630.600 226.050 631.050 ;
        RECT 259.950 630.600 262.050 631.050 ;
        RECT 223.950 629.400 262.050 630.600 ;
        RECT 223.950 628.950 226.050 629.400 ;
        RECT 259.950 628.950 262.050 629.400 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 283.950 628.950 286.050 631.050 ;
        RECT 352.950 630.600 355.050 631.050 ;
        RECT 364.950 630.600 367.050 631.050 ;
        RECT 373.950 630.600 376.050 631.050 ;
        RECT 352.950 629.400 357.600 630.600 ;
        RECT 352.950 628.950 355.050 629.400 ;
        RECT 175.950 627.600 178.050 628.050 ;
        RECT 199.950 627.600 202.050 628.050 ;
        RECT 152.400 626.400 202.050 627.600 ;
        RECT 58.950 625.950 61.050 626.400 ;
        RECT 70.950 625.950 73.050 626.400 ;
        RECT 175.950 625.950 178.050 626.400 ;
        RECT 199.950 625.950 202.050 626.400 ;
        RECT 211.950 627.600 214.050 628.050 ;
        RECT 223.950 627.600 226.050 628.050 ;
        RECT 211.950 626.400 226.050 627.600 ;
        RECT 211.950 625.950 214.050 626.400 ;
        RECT 223.950 625.950 226.050 626.400 ;
        RECT 235.950 627.600 238.050 628.050 ;
        RECT 280.950 627.600 283.050 628.050 ;
        RECT 235.950 626.400 283.050 627.600 ;
        RECT 356.400 627.600 357.600 629.400 ;
        RECT 364.950 629.400 376.050 630.600 ;
        RECT 364.950 628.950 367.050 629.400 ;
        RECT 373.950 628.950 376.050 629.400 ;
        RECT 403.950 630.600 406.050 631.050 ;
        RECT 412.950 630.600 415.050 631.050 ;
        RECT 403.950 629.400 415.050 630.600 ;
        RECT 403.950 628.950 406.050 629.400 ;
        RECT 412.950 628.950 415.050 629.400 ;
        RECT 418.950 628.950 421.050 631.050 ;
        RECT 445.950 630.600 448.050 631.050 ;
        RECT 484.950 630.600 487.050 631.050 ;
        RECT 445.950 629.400 487.050 630.600 ;
        RECT 445.950 628.950 448.050 629.400 ;
        RECT 484.950 628.950 487.050 629.400 ;
        RECT 505.950 630.600 508.050 631.050 ;
        RECT 520.950 630.600 523.050 631.050 ;
        RECT 505.950 629.400 523.050 630.600 ;
        RECT 505.950 628.950 508.050 629.400 ;
        RECT 520.950 628.950 523.050 629.400 ;
        RECT 544.950 628.950 547.050 631.050 ;
        RECT 580.950 630.600 583.050 631.050 ;
        RECT 595.950 630.600 598.050 631.050 ;
        RECT 580.950 629.400 598.050 630.600 ;
        RECT 580.950 628.950 583.050 629.400 ;
        RECT 595.950 628.950 598.050 629.400 ;
        RECT 601.950 630.600 604.050 631.050 ;
        RECT 616.950 630.600 619.050 631.050 ;
        RECT 601.950 629.400 619.050 630.600 ;
        RECT 601.950 628.950 604.050 629.400 ;
        RECT 616.950 628.950 619.050 629.400 ;
        RECT 631.950 628.950 634.050 631.050 ;
        RECT 661.950 630.600 664.050 631.050 ;
        RECT 676.950 630.600 679.050 631.050 ;
        RECT 661.950 629.400 679.050 630.600 ;
        RECT 661.950 628.950 664.050 629.400 ;
        RECT 676.950 628.950 679.050 629.400 ;
        RECT 682.950 630.600 685.050 631.050 ;
        RECT 692.400 630.600 693.600 632.400 ;
        RECT 700.950 631.950 703.050 632.400 ;
        RECT 712.950 631.950 715.050 632.400 ;
        RECT 763.950 633.600 766.050 634.050 ;
        RECT 790.950 633.600 793.050 634.050 ;
        RECT 763.950 632.400 793.050 633.600 ;
        RECT 763.950 631.950 766.050 632.400 ;
        RECT 790.950 631.950 793.050 632.400 ;
        RECT 799.950 633.600 802.050 634.050 ;
        RECT 805.950 633.600 808.050 634.050 ;
        RECT 799.950 632.400 808.050 633.600 ;
        RECT 799.950 631.950 802.050 632.400 ;
        RECT 805.950 631.950 808.050 632.400 ;
        RECT 811.950 633.600 814.050 634.050 ;
        RECT 826.950 633.600 829.050 634.050 ;
        RECT 877.950 633.600 880.050 634.050 ;
        RECT 811.950 632.400 880.050 633.600 ;
        RECT 811.950 631.950 814.050 632.400 ;
        RECT 826.950 631.950 829.050 632.400 ;
        RECT 877.950 631.950 880.050 632.400 ;
        RECT 682.950 629.400 693.600 630.600 ;
        RECT 682.950 628.950 685.050 629.400 ;
        RECT 784.950 628.950 787.050 631.050 ;
        RECT 808.950 630.600 811.050 631.050 ;
        RECT 841.950 630.600 844.050 631.050 ;
        RECT 808.950 629.400 844.050 630.600 ;
        RECT 808.950 628.950 811.050 629.400 ;
        RECT 841.950 628.950 844.050 629.400 ;
        RECT 358.950 627.600 361.050 628.050 ;
        RECT 356.400 626.400 361.050 627.600 ;
        RECT 419.400 627.600 420.600 628.950 ;
        RECT 475.950 627.600 478.050 628.050 ;
        RECT 419.400 626.400 478.050 627.600 ;
        RECT 235.950 625.950 238.050 626.400 ;
        RECT 280.950 625.950 283.050 626.400 ;
        RECT 358.950 625.950 361.050 626.400 ;
        RECT 475.950 625.950 478.050 626.400 ;
        RECT 493.950 627.600 496.050 628.050 ;
        RECT 502.950 627.600 505.050 628.050 ;
        RECT 493.950 626.400 505.050 627.600 ;
        RECT 493.950 625.950 496.050 626.400 ;
        RECT 502.950 625.950 505.050 626.400 ;
        RECT 511.950 627.600 514.050 628.050 ;
        RECT 541.950 627.600 544.050 628.050 ;
        RECT 511.950 626.400 544.050 627.600 ;
        RECT 545.400 627.600 546.600 628.950 ;
        RECT 556.950 627.600 559.050 628.050 ;
        RECT 545.400 626.400 559.050 627.600 ;
        RECT 511.950 625.950 514.050 626.400 ;
        RECT 541.950 625.950 544.050 626.400 ;
        RECT 556.950 625.950 559.050 626.400 ;
        RECT 598.950 627.600 601.050 628.050 ;
        RECT 632.400 627.600 633.600 628.950 ;
        RECT 598.950 626.400 633.600 627.600 ;
        RECT 640.950 627.600 643.050 628.050 ;
        RECT 709.950 627.600 712.050 628.050 ;
        RECT 640.950 626.400 712.050 627.600 ;
        RECT 598.950 625.950 601.050 626.400 ;
        RECT 640.950 625.950 643.050 626.400 ;
        RECT 709.950 625.950 712.050 626.400 ;
        RECT 721.950 627.600 724.050 628.050 ;
        RECT 742.950 627.600 745.050 628.050 ;
        RECT 721.950 626.400 745.050 627.600 ;
        RECT 721.950 625.950 724.050 626.400 ;
        RECT 742.950 625.950 745.050 626.400 ;
        RECT 745.950 627.600 748.050 628.050 ;
        RECT 769.950 627.600 772.050 628.050 ;
        RECT 745.950 626.400 772.050 627.600 ;
        RECT 745.950 625.950 748.050 626.400 ;
        RECT 769.950 625.950 772.050 626.400 ;
        RECT 785.400 625.050 786.600 628.950 ;
        RECT 850.950 627.600 853.050 628.050 ;
        RECT 871.950 627.600 874.050 628.050 ;
        RECT 850.950 626.400 874.050 627.600 ;
        RECT 850.950 625.950 853.050 626.400 ;
        RECT 871.950 625.950 874.050 626.400 ;
        RECT 16.950 624.600 19.050 625.050 ;
        RECT 43.950 624.600 46.050 625.050 ;
        RECT 16.950 623.400 46.050 624.600 ;
        RECT 16.950 622.950 19.050 623.400 ;
        RECT 43.950 622.950 46.050 623.400 ;
        RECT 55.950 624.600 58.050 625.050 ;
        RECT 115.950 624.600 118.050 625.050 ;
        RECT 55.950 623.400 118.050 624.600 ;
        RECT 55.950 622.950 58.050 623.400 ;
        RECT 115.950 622.950 118.050 623.400 ;
        RECT 121.950 624.600 124.050 625.050 ;
        RECT 154.950 624.600 157.050 625.050 ;
        RECT 121.950 623.400 157.050 624.600 ;
        RECT 121.950 622.950 124.050 623.400 ;
        RECT 154.950 622.950 157.050 623.400 ;
        RECT 178.950 624.600 181.050 625.050 ;
        RECT 244.950 624.600 247.050 625.050 ;
        RECT 256.950 624.600 259.050 625.050 ;
        RECT 178.950 623.400 259.050 624.600 ;
        RECT 178.950 622.950 181.050 623.400 ;
        RECT 244.950 622.950 247.050 623.400 ;
        RECT 256.950 622.950 259.050 623.400 ;
        RECT 277.950 624.600 280.050 625.050 ;
        RECT 292.950 624.600 295.050 625.050 ;
        RECT 304.950 624.600 307.050 625.050 ;
        RECT 307.950 624.600 310.050 625.050 ;
        RECT 277.950 623.400 310.050 624.600 ;
        RECT 277.950 622.950 280.050 623.400 ;
        RECT 292.950 622.950 295.050 623.400 ;
        RECT 304.950 622.950 307.050 623.400 ;
        RECT 307.950 622.950 310.050 623.400 ;
        RECT 340.950 624.600 343.050 625.050 ;
        RECT 355.950 624.600 358.050 625.050 ;
        RECT 340.950 623.400 358.050 624.600 ;
        RECT 340.950 622.950 343.050 623.400 ;
        RECT 355.950 622.950 358.050 623.400 ;
        RECT 382.950 624.600 385.050 625.050 ;
        RECT 391.950 624.600 394.050 625.050 ;
        RECT 382.950 623.400 394.050 624.600 ;
        RECT 382.950 622.950 385.050 623.400 ;
        RECT 391.950 622.950 394.050 623.400 ;
        RECT 415.950 624.600 418.050 625.050 ;
        RECT 439.950 624.600 442.050 625.050 ;
        RECT 415.950 623.400 442.050 624.600 ;
        RECT 415.950 622.950 418.050 623.400 ;
        RECT 439.950 622.950 442.050 623.400 ;
        RECT 472.950 624.600 475.050 625.050 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 472.950 623.400 502.050 624.600 ;
        RECT 472.950 622.950 475.050 623.400 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 526.950 624.600 529.050 625.050 ;
        RECT 538.950 624.600 541.050 625.050 ;
        RECT 526.950 623.400 541.050 624.600 ;
        RECT 526.950 622.950 529.050 623.400 ;
        RECT 538.950 622.950 541.050 623.400 ;
        RECT 559.950 624.600 562.050 625.050 ;
        RECT 574.950 624.600 577.050 625.050 ;
        RECT 559.950 623.400 577.050 624.600 ;
        RECT 559.950 622.950 562.050 623.400 ;
        RECT 574.950 622.950 577.050 623.400 ;
        RECT 619.950 624.600 622.050 625.050 ;
        RECT 637.950 624.600 640.050 625.050 ;
        RECT 619.950 623.400 640.050 624.600 ;
        RECT 619.950 622.950 622.050 623.400 ;
        RECT 637.950 622.950 640.050 623.400 ;
        RECT 649.950 624.600 652.050 625.050 ;
        RECT 781.950 624.600 784.050 625.050 ;
        RECT 649.950 623.400 784.050 624.600 ;
        RECT 649.950 622.950 652.050 623.400 ;
        RECT 781.950 622.950 784.050 623.400 ;
        RECT 784.950 622.950 787.050 625.050 ;
        RECT 790.950 624.600 793.050 625.050 ;
        RECT 796.950 624.600 799.050 625.050 ;
        RECT 790.950 623.400 799.050 624.600 ;
        RECT 790.950 622.950 793.050 623.400 ;
        RECT 796.950 622.950 799.050 623.400 ;
        RECT 847.950 624.600 850.050 625.050 ;
        RECT 859.950 624.600 862.050 625.050 ;
        RECT 865.950 624.600 868.050 625.050 ;
        RECT 847.950 623.400 868.050 624.600 ;
        RECT 847.950 622.950 850.050 623.400 ;
        RECT 859.950 622.950 862.050 623.400 ;
        RECT 865.950 622.950 868.050 623.400 ;
        RECT 871.950 624.600 874.050 625.050 ;
        RECT 883.950 624.600 886.050 625.050 ;
        RECT 871.950 623.400 886.050 624.600 ;
        RECT 871.950 622.950 874.050 623.400 ;
        RECT 883.950 622.950 886.050 623.400 ;
        RECT 64.950 621.600 67.050 622.050 ;
        RECT 73.950 621.600 76.050 622.050 ;
        RECT 64.950 620.400 76.050 621.600 ;
        RECT 64.950 619.950 67.050 620.400 ;
        RECT 73.950 619.950 76.050 620.400 ;
        RECT 145.950 621.600 148.050 622.050 ;
        RECT 166.950 621.600 169.050 622.050 ;
        RECT 145.950 620.400 169.050 621.600 ;
        RECT 145.950 619.950 148.050 620.400 ;
        RECT 166.950 619.950 169.050 620.400 ;
        RECT 208.950 621.600 211.050 622.050 ;
        RECT 220.950 621.600 223.050 622.050 ;
        RECT 208.950 620.400 223.050 621.600 ;
        RECT 208.950 619.950 211.050 620.400 ;
        RECT 220.950 619.950 223.050 620.400 ;
        RECT 388.950 621.600 391.050 622.050 ;
        RECT 418.950 621.600 421.050 622.050 ;
        RECT 388.950 620.400 421.050 621.600 ;
        RECT 388.950 619.950 391.050 620.400 ;
        RECT 418.950 619.950 421.050 620.400 ;
        RECT 451.950 621.600 454.050 622.050 ;
        RECT 484.950 621.600 487.050 622.050 ;
        RECT 451.950 620.400 487.050 621.600 ;
        RECT 451.950 619.950 454.050 620.400 ;
        RECT 484.950 619.950 487.050 620.400 ;
        RECT 496.950 621.600 499.050 622.050 ;
        RECT 502.950 621.600 505.050 622.050 ;
        RECT 496.950 620.400 505.050 621.600 ;
        RECT 496.950 619.950 499.050 620.400 ;
        RECT 502.950 619.950 505.050 620.400 ;
        RECT 634.950 621.600 637.050 622.050 ;
        RECT 661.950 621.600 664.050 622.050 ;
        RECT 634.950 620.400 664.050 621.600 ;
        RECT 634.950 619.950 637.050 620.400 ;
        RECT 661.950 619.950 664.050 620.400 ;
        RECT 703.950 621.600 706.050 622.050 ;
        RECT 718.950 621.600 721.050 622.050 ;
        RECT 703.950 620.400 721.050 621.600 ;
        RECT 703.950 619.950 706.050 620.400 ;
        RECT 718.950 619.950 721.050 620.400 ;
        RECT 775.950 621.600 778.050 622.050 ;
        RECT 787.950 621.600 790.050 622.050 ;
        RECT 775.950 620.400 790.050 621.600 ;
        RECT 775.950 619.950 778.050 620.400 ;
        RECT 787.950 619.950 790.050 620.400 ;
        RECT 862.950 621.600 865.050 622.050 ;
        RECT 868.950 621.600 871.050 622.050 ;
        RECT 862.950 620.400 871.050 621.600 ;
        RECT 862.950 619.950 865.050 620.400 ;
        RECT 868.950 619.950 871.050 620.400 ;
        RECT 40.950 618.600 43.050 619.050 ;
        RECT 46.950 618.600 49.050 619.050 ;
        RECT 61.950 618.600 64.050 619.050 ;
        RECT 79.950 618.600 82.050 619.050 ;
        RECT 40.950 617.400 82.050 618.600 ;
        RECT 40.950 616.950 43.050 617.400 ;
        RECT 46.950 616.950 49.050 617.400 ;
        RECT 61.950 616.950 64.050 617.400 ;
        RECT 79.950 616.950 82.050 617.400 ;
        RECT 196.950 618.600 199.050 619.050 ;
        RECT 226.950 618.600 229.050 619.050 ;
        RECT 238.950 618.600 241.050 619.050 ;
        RECT 196.950 617.400 241.050 618.600 ;
        RECT 196.950 616.950 199.050 617.400 ;
        RECT 226.950 616.950 229.050 617.400 ;
        RECT 238.950 616.950 241.050 617.400 ;
        RECT 388.950 618.600 391.050 619.050 ;
        RECT 403.950 618.600 406.050 619.050 ;
        RECT 427.950 618.600 430.050 619.050 ;
        RECT 388.950 617.400 430.050 618.600 ;
        RECT 388.950 616.950 391.050 617.400 ;
        RECT 403.950 616.950 406.050 617.400 ;
        RECT 427.950 616.950 430.050 617.400 ;
        RECT 613.950 618.600 616.050 619.050 ;
        RECT 799.950 618.600 802.050 619.050 ;
        RECT 820.950 618.600 823.050 619.050 ;
        RECT 868.950 618.600 871.050 619.050 ;
        RECT 613.950 617.400 871.050 618.600 ;
        RECT 613.950 616.950 616.050 617.400 ;
        RECT 799.950 616.950 802.050 617.400 ;
        RECT 820.950 616.950 823.050 617.400 ;
        RECT 868.950 616.950 871.050 617.400 ;
        RECT 742.950 615.600 745.050 616.050 ;
        RECT 820.950 615.600 823.050 616.050 ;
        RECT 850.950 615.600 853.050 616.050 ;
        RECT 742.950 614.400 853.050 615.600 ;
        RECT 742.950 613.950 745.050 614.400 ;
        RECT 820.950 613.950 823.050 614.400 ;
        RECT 850.950 613.950 853.050 614.400 ;
        RECT 157.950 612.600 160.050 613.050 ;
        RECT 214.950 612.600 217.050 613.050 ;
        RECT 157.950 611.400 217.050 612.600 ;
        RECT 157.950 610.950 160.050 611.400 ;
        RECT 214.950 610.950 217.050 611.400 ;
        RECT 223.950 612.600 226.050 613.050 ;
        RECT 322.950 612.600 325.050 613.050 ;
        RECT 223.950 611.400 325.050 612.600 ;
        RECT 223.950 610.950 226.050 611.400 ;
        RECT 322.950 610.950 325.050 611.400 ;
        RECT 418.950 612.600 421.050 613.050 ;
        RECT 457.950 612.600 460.050 613.050 ;
        RECT 541.950 612.600 544.050 613.050 ;
        RECT 562.950 612.600 565.050 613.050 ;
        RECT 418.950 611.400 565.050 612.600 ;
        RECT 418.950 610.950 421.050 611.400 ;
        RECT 457.950 610.950 460.050 611.400 ;
        RECT 541.950 610.950 544.050 611.400 ;
        RECT 562.950 610.950 565.050 611.400 ;
        RECT 604.950 612.600 607.050 613.050 ;
        RECT 664.950 612.600 667.050 613.050 ;
        RECT 604.950 611.400 667.050 612.600 ;
        RECT 604.950 610.950 607.050 611.400 ;
        RECT 664.950 610.950 667.050 611.400 ;
        RECT 688.950 612.600 691.050 613.050 ;
        RECT 793.950 612.600 796.050 613.050 ;
        RECT 814.950 612.600 817.050 613.050 ;
        RECT 688.950 611.400 817.050 612.600 ;
        RECT 688.950 610.950 691.050 611.400 ;
        RECT 793.950 610.950 796.050 611.400 ;
        RECT 814.950 610.950 817.050 611.400 ;
        RECT 301.950 609.600 304.050 610.050 ;
        RECT 328.950 609.600 331.050 610.050 ;
        RECT 301.950 608.400 331.050 609.600 ;
        RECT 301.950 607.950 304.050 608.400 ;
        RECT 328.950 607.950 331.050 608.400 ;
        RECT 520.950 609.600 523.050 610.050 ;
        RECT 526.950 609.600 529.050 610.050 ;
        RECT 568.950 609.600 571.050 610.050 ;
        RECT 520.950 608.400 571.050 609.600 ;
        RECT 520.950 607.950 523.050 608.400 ;
        RECT 526.950 607.950 529.050 608.400 ;
        RECT 568.950 607.950 571.050 608.400 ;
        RECT 694.950 609.600 697.050 610.050 ;
        RECT 745.950 609.600 748.050 610.050 ;
        RECT 694.950 608.400 748.050 609.600 ;
        RECT 694.950 607.950 697.050 608.400 ;
        RECT 745.950 607.950 748.050 608.400 ;
        RECT 427.950 606.600 430.050 607.050 ;
        RECT 448.950 606.600 451.050 607.050 ;
        RECT 427.950 605.400 451.050 606.600 ;
        RECT 427.950 604.950 430.050 605.400 ;
        RECT 448.950 604.950 451.050 605.400 ;
        RECT 508.950 606.600 511.050 607.050 ;
        RECT 520.950 606.600 523.050 607.050 ;
        RECT 544.950 606.600 547.050 607.050 ;
        RECT 508.950 605.400 547.050 606.600 ;
        RECT 508.950 604.950 511.050 605.400 ;
        RECT 520.950 604.950 523.050 605.400 ;
        RECT 544.950 604.950 547.050 605.400 ;
        RECT 583.950 606.600 586.050 607.050 ;
        RECT 646.950 606.600 649.050 607.050 ;
        RECT 583.950 605.400 649.050 606.600 ;
        RECT 583.950 604.950 586.050 605.400 ;
        RECT 646.950 604.950 649.050 605.400 ;
        RECT 697.950 606.600 700.050 607.050 ;
        RECT 751.950 606.600 754.050 607.050 ;
        RECT 817.950 606.600 820.050 607.050 ;
        RECT 880.950 606.600 883.050 607.050 ;
        RECT 697.950 605.400 820.050 606.600 ;
        RECT 697.950 604.950 700.050 605.400 ;
        RECT 751.950 604.950 754.050 605.400 ;
        RECT 817.950 604.950 820.050 605.400 ;
        RECT 857.400 605.400 883.050 606.600 ;
        RECT 28.950 603.600 31.050 604.050 ;
        RECT 31.950 603.600 34.050 604.050 ;
        RECT 82.950 603.600 85.050 604.050 ;
        RECT 28.950 602.400 85.050 603.600 ;
        RECT 28.950 601.950 31.050 602.400 ;
        RECT 31.950 601.950 34.050 602.400 ;
        RECT 82.950 601.950 85.050 602.400 ;
        RECT 172.950 603.600 175.050 604.050 ;
        RECT 199.950 603.600 202.050 604.050 ;
        RECT 244.950 603.600 247.050 604.050 ;
        RECT 172.950 602.400 247.050 603.600 ;
        RECT 172.950 601.950 175.050 602.400 ;
        RECT 199.950 601.950 202.050 602.400 ;
        RECT 244.950 601.950 247.050 602.400 ;
        RECT 262.950 603.600 265.050 604.050 ;
        RECT 298.950 603.600 301.050 604.050 ;
        RECT 262.950 602.400 301.050 603.600 ;
        RECT 262.950 601.950 265.050 602.400 ;
        RECT 298.950 601.950 301.050 602.400 ;
        RECT 364.950 603.600 367.050 604.050 ;
        RECT 373.950 603.600 376.050 604.050 ;
        RECT 364.950 602.400 376.050 603.600 ;
        RECT 364.950 601.950 367.050 602.400 ;
        RECT 373.950 601.950 376.050 602.400 ;
        RECT 376.950 603.600 379.050 604.050 ;
        RECT 382.950 603.600 385.050 604.050 ;
        RECT 376.950 602.400 385.050 603.600 ;
        RECT 376.950 601.950 379.050 602.400 ;
        RECT 382.950 601.950 385.050 602.400 ;
        RECT 433.950 603.600 436.050 604.050 ;
        RECT 472.950 603.600 475.050 604.050 ;
        RECT 433.950 602.400 475.050 603.600 ;
        RECT 433.950 601.950 436.050 602.400 ;
        RECT 472.950 601.950 475.050 602.400 ;
        RECT 508.950 603.600 511.050 604.050 ;
        RECT 523.950 603.600 526.050 604.050 ;
        RECT 508.950 602.400 526.050 603.600 ;
        RECT 508.950 601.950 511.050 602.400 ;
        RECT 523.950 601.950 526.050 602.400 ;
        RECT 547.950 603.600 550.050 604.050 ;
        RECT 607.950 603.600 610.050 604.050 ;
        RECT 631.950 603.600 634.050 604.050 ;
        RECT 547.950 602.400 634.050 603.600 ;
        RECT 547.950 601.950 550.050 602.400 ;
        RECT 607.950 601.950 610.050 602.400 ;
        RECT 631.950 601.950 634.050 602.400 ;
        RECT 637.950 603.600 640.050 604.050 ;
        RECT 652.950 603.600 655.050 604.050 ;
        RECT 637.950 602.400 655.050 603.600 ;
        RECT 637.950 601.950 640.050 602.400 ;
        RECT 652.950 601.950 655.050 602.400 ;
        RECT 664.950 603.600 667.050 604.050 ;
        RECT 670.950 603.600 673.050 604.050 ;
        RECT 724.950 603.600 727.050 604.050 ;
        RECT 664.950 602.400 673.050 603.600 ;
        RECT 664.950 601.950 667.050 602.400 ;
        RECT 670.950 601.950 673.050 602.400 ;
        RECT 710.400 602.400 727.050 603.600 ;
        RECT 710.400 601.050 711.600 602.400 ;
        RECT 724.950 601.950 727.050 602.400 ;
        RECT 838.950 603.600 841.050 604.050 ;
        RECT 853.950 603.600 856.050 604.050 ;
        RECT 838.950 602.400 856.050 603.600 ;
        RECT 838.950 601.950 841.050 602.400 ;
        RECT 853.950 601.950 856.050 602.400 ;
        RECT 857.400 601.050 858.600 605.400 ;
        RECT 880.950 604.950 883.050 605.400 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 61.950 600.600 64.050 601.050 ;
        RECT 23.400 599.400 64.050 600.600 ;
        RECT 10.950 597.600 13.050 598.050 ;
        RECT 23.400 597.600 24.600 599.400 ;
        RECT 61.950 598.950 64.050 599.400 ;
        RECT 67.950 598.950 70.050 601.050 ;
        RECT 70.950 600.600 73.050 601.050 ;
        RECT 79.950 600.600 82.050 601.050 ;
        RECT 85.950 600.600 88.050 601.050 ;
        RECT 70.950 599.400 88.050 600.600 ;
        RECT 70.950 598.950 73.050 599.400 ;
        RECT 79.950 598.950 82.050 599.400 ;
        RECT 85.950 598.950 88.050 599.400 ;
        RECT 91.950 600.600 94.050 601.050 ;
        RECT 106.950 600.600 109.050 601.050 ;
        RECT 91.950 599.400 109.050 600.600 ;
        RECT 91.950 598.950 94.050 599.400 ;
        RECT 106.950 598.950 109.050 599.400 ;
        RECT 151.950 600.600 154.050 601.050 ;
        RECT 157.950 600.600 160.050 601.050 ;
        RECT 151.950 599.400 160.050 600.600 ;
        RECT 151.950 598.950 154.050 599.400 ;
        RECT 157.950 598.950 160.050 599.400 ;
        RECT 181.950 600.600 184.050 601.050 ;
        RECT 193.950 600.600 196.050 601.050 ;
        RECT 217.950 600.600 220.050 601.050 ;
        RECT 229.950 600.600 232.050 601.050 ;
        RECT 232.950 600.600 235.050 601.050 ;
        RECT 181.950 599.400 220.050 600.600 ;
        RECT 181.950 598.950 184.050 599.400 ;
        RECT 193.950 598.950 196.050 599.400 ;
        RECT 217.950 598.950 220.050 599.400 ;
        RECT 224.400 599.400 235.050 600.600 ;
        RECT 10.950 596.400 24.600 597.600 ;
        RECT 25.950 597.600 28.050 598.050 ;
        RECT 34.950 597.600 37.050 598.050 ;
        RECT 25.950 596.400 37.050 597.600 ;
        RECT 10.950 595.950 13.050 596.400 ;
        RECT 25.950 595.950 28.050 596.400 ;
        RECT 34.950 595.950 37.050 596.400 ;
        RECT 46.950 597.600 49.050 598.050 ;
        RECT 64.950 597.600 67.050 598.050 ;
        RECT 46.950 596.400 67.050 597.600 ;
        RECT 68.400 597.600 69.600 598.950 ;
        RECT 88.950 597.600 91.050 598.050 ;
        RECT 68.400 596.400 91.050 597.600 ;
        RECT 46.950 595.950 49.050 596.400 ;
        RECT 64.950 595.950 67.050 596.400 ;
        RECT 88.950 595.950 91.050 596.400 ;
        RECT 133.950 597.600 136.050 598.050 ;
        RECT 136.950 597.600 139.050 598.050 ;
        RECT 142.950 597.600 145.050 598.050 ;
        RECT 133.950 596.400 145.050 597.600 ;
        RECT 133.950 595.950 136.050 596.400 ;
        RECT 136.950 595.950 139.050 596.400 ;
        RECT 142.950 595.950 145.050 596.400 ;
        RECT 148.950 597.600 151.050 598.050 ;
        RECT 154.950 597.600 157.050 598.050 ;
        RECT 166.950 597.600 169.050 598.050 ;
        RECT 148.950 596.400 169.050 597.600 ;
        RECT 148.950 595.950 151.050 596.400 ;
        RECT 154.950 595.950 157.050 596.400 ;
        RECT 166.950 595.950 169.050 596.400 ;
        RECT 202.950 597.600 205.050 598.050 ;
        RECT 214.950 597.600 217.050 598.050 ;
        RECT 224.400 597.600 225.600 599.400 ;
        RECT 229.950 598.950 232.050 599.400 ;
        RECT 232.950 598.950 235.050 599.400 ;
        RECT 241.950 600.600 244.050 601.050 ;
        RECT 253.950 600.600 256.050 601.050 ;
        RECT 241.950 599.400 256.050 600.600 ;
        RECT 241.950 598.950 244.050 599.400 ;
        RECT 253.950 598.950 256.050 599.400 ;
        RECT 259.950 600.600 262.050 601.050 ;
        RECT 277.950 600.600 280.050 601.050 ;
        RECT 259.950 599.400 280.050 600.600 ;
        RECT 259.950 598.950 262.050 599.400 ;
        RECT 277.950 598.950 280.050 599.400 ;
        RECT 298.950 600.600 301.050 601.050 ;
        RECT 307.950 600.600 310.050 601.050 ;
        RECT 298.950 599.400 310.050 600.600 ;
        RECT 298.950 598.950 301.050 599.400 ;
        RECT 307.950 598.950 310.050 599.400 ;
        RECT 340.950 600.600 343.050 601.050 ;
        RECT 364.950 600.600 367.050 601.050 ;
        RECT 415.950 600.600 418.050 601.050 ;
        RECT 340.950 599.400 367.050 600.600 ;
        RECT 340.950 598.950 343.050 599.400 ;
        RECT 364.950 598.950 367.050 599.400 ;
        RECT 368.400 599.400 418.050 600.600 ;
        RECT 202.950 596.400 225.600 597.600 ;
        RECT 226.950 597.600 229.050 598.050 ;
        RECT 238.950 597.600 241.050 598.050 ;
        RECT 226.950 596.400 241.050 597.600 ;
        RECT 202.950 595.950 205.050 596.400 ;
        RECT 214.950 595.950 217.050 596.400 ;
        RECT 226.950 595.950 229.050 596.400 ;
        RECT 238.950 595.950 241.050 596.400 ;
        RECT 283.950 597.600 286.050 598.050 ;
        RECT 298.950 597.600 301.050 598.050 ;
        RECT 283.950 596.400 301.050 597.600 ;
        RECT 283.950 595.950 286.050 596.400 ;
        RECT 298.950 595.950 301.050 596.400 ;
        RECT 319.950 597.600 322.050 598.050 ;
        RECT 337.950 597.600 340.050 598.050 ;
        RECT 319.950 596.400 340.050 597.600 ;
        RECT 319.950 595.950 322.050 596.400 ;
        RECT 337.950 595.950 340.050 596.400 ;
        RECT 343.950 597.600 346.050 598.050 ;
        RECT 352.950 597.600 355.050 598.050 ;
        RECT 368.400 597.600 369.600 599.400 ;
        RECT 415.950 598.950 418.050 599.400 ;
        RECT 445.950 600.600 448.050 601.050 ;
        RECT 454.950 600.600 457.050 601.050 ;
        RECT 445.950 599.400 457.050 600.600 ;
        RECT 445.950 598.950 448.050 599.400 ;
        RECT 454.950 598.950 457.050 599.400 ;
        RECT 487.950 600.600 490.050 601.050 ;
        RECT 496.950 600.600 499.050 601.050 ;
        RECT 487.950 599.400 499.050 600.600 ;
        RECT 487.950 598.950 490.050 599.400 ;
        RECT 496.950 598.950 499.050 599.400 ;
        RECT 535.950 600.600 538.050 601.050 ;
        RECT 547.950 600.600 550.050 601.050 ;
        RECT 559.950 600.600 562.050 601.050 ;
        RECT 535.950 599.400 562.050 600.600 ;
        RECT 535.950 598.950 538.050 599.400 ;
        RECT 547.950 598.950 550.050 599.400 ;
        RECT 559.950 598.950 562.050 599.400 ;
        RECT 586.950 600.600 589.050 601.050 ;
        RECT 592.950 600.600 595.050 601.050 ;
        RECT 601.950 600.600 604.050 601.050 ;
        RECT 586.950 599.400 591.600 600.600 ;
        RECT 586.950 598.950 589.050 599.400 ;
        RECT 343.950 596.400 355.050 597.600 ;
        RECT 343.950 595.950 346.050 596.400 ;
        RECT 352.950 595.950 355.050 596.400 ;
        RECT 365.400 596.400 369.600 597.600 ;
        RECT 91.950 594.600 94.050 595.050 ;
        RECT 97.950 594.600 100.050 595.050 ;
        RECT 91.950 593.400 100.050 594.600 ;
        RECT 91.950 592.950 94.050 593.400 ;
        RECT 97.950 592.950 100.050 593.400 ;
        RECT 175.950 594.600 178.050 595.050 ;
        RECT 199.950 594.600 202.050 595.050 ;
        RECT 208.950 594.600 211.050 595.050 ;
        RECT 175.950 593.400 211.050 594.600 ;
        RECT 175.950 592.950 178.050 593.400 ;
        RECT 199.950 592.950 202.050 593.400 ;
        RECT 208.950 592.950 211.050 593.400 ;
        RECT 280.950 594.600 283.050 595.050 ;
        RECT 295.950 594.600 298.050 595.050 ;
        RECT 304.950 594.600 307.050 595.050 ;
        RECT 322.950 594.600 325.050 595.050 ;
        RECT 280.950 593.400 325.050 594.600 ;
        RECT 280.950 592.950 283.050 593.400 ;
        RECT 295.950 592.950 298.050 593.400 ;
        RECT 304.950 592.950 307.050 593.400 ;
        RECT 322.950 592.950 325.050 593.400 ;
        RECT 361.950 594.600 364.050 595.050 ;
        RECT 365.400 594.600 366.600 596.400 ;
        RECT 370.950 595.950 373.050 598.050 ;
        RECT 373.950 597.600 376.050 598.050 ;
        RECT 379.950 597.600 382.050 598.050 ;
        RECT 373.950 596.400 382.050 597.600 ;
        RECT 373.950 595.950 376.050 596.400 ;
        RECT 379.950 595.950 382.050 596.400 ;
        RECT 406.950 597.600 409.050 598.050 ;
        RECT 424.950 597.600 427.050 598.050 ;
        RECT 406.950 596.400 427.050 597.600 ;
        RECT 406.950 595.950 409.050 596.400 ;
        RECT 424.950 595.950 427.050 596.400 ;
        RECT 496.950 597.600 499.050 598.050 ;
        RECT 583.950 597.600 586.050 598.050 ;
        RECT 590.400 597.600 591.600 599.400 ;
        RECT 592.950 599.400 604.050 600.600 ;
        RECT 592.950 598.950 595.050 599.400 ;
        RECT 601.950 598.950 604.050 599.400 ;
        RECT 679.950 600.600 682.050 601.050 ;
        RECT 691.950 600.600 694.050 601.050 ;
        RECT 679.950 599.400 694.050 600.600 ;
        RECT 679.950 598.950 682.050 599.400 ;
        RECT 691.950 598.950 694.050 599.400 ;
        RECT 709.950 598.950 712.050 601.050 ;
        RECT 739.950 598.950 742.050 601.050 ;
        RECT 781.950 598.950 784.050 601.050 ;
        RECT 784.950 600.600 787.050 601.050 ;
        RECT 805.950 600.600 808.050 601.050 ;
        RECT 784.950 599.400 808.050 600.600 ;
        RECT 784.950 598.950 787.050 599.400 ;
        RECT 805.950 598.950 808.050 599.400 ;
        RECT 823.950 600.600 826.050 601.050 ;
        RECT 850.950 600.600 853.050 601.050 ;
        RECT 823.950 599.400 853.050 600.600 ;
        RECT 823.950 598.950 826.050 599.400 ;
        RECT 850.950 598.950 853.050 599.400 ;
        RECT 856.950 598.950 859.050 601.050 ;
        RECT 613.950 597.600 616.050 598.050 ;
        RECT 496.950 596.400 588.600 597.600 ;
        RECT 590.400 596.400 616.050 597.600 ;
        RECT 496.950 595.950 499.050 596.400 ;
        RECT 583.950 595.950 586.050 596.400 ;
        RECT 361.950 593.400 366.600 594.600 ;
        RECT 361.950 592.950 364.050 593.400 ;
        RECT 367.950 592.950 370.050 595.050 ;
        RECT 371.400 594.600 372.600 595.950 ;
        RECT 385.950 594.600 388.050 595.050 ;
        RECT 371.400 593.400 388.050 594.600 ;
        RECT 385.950 592.950 388.050 593.400 ;
        RECT 388.950 594.600 391.050 595.050 ;
        RECT 394.950 594.600 397.050 595.050 ;
        RECT 388.950 593.400 397.050 594.600 ;
        RECT 388.950 592.950 391.050 593.400 ;
        RECT 394.950 592.950 397.050 593.400 ;
        RECT 466.950 594.600 469.050 595.050 ;
        RECT 469.950 594.600 472.050 595.050 ;
        RECT 499.950 594.600 502.050 595.050 ;
        RECT 466.950 593.400 502.050 594.600 ;
        RECT 587.400 594.600 588.600 596.400 ;
        RECT 613.950 595.950 616.050 596.400 ;
        RECT 640.950 597.600 643.050 598.050 ;
        RECT 646.950 597.600 649.050 598.050 ;
        RECT 640.950 596.400 649.050 597.600 ;
        RECT 640.950 595.950 643.050 596.400 ;
        RECT 646.950 595.950 649.050 596.400 ;
        RECT 655.950 597.600 658.050 598.050 ;
        RECT 673.950 597.600 676.050 598.050 ;
        RECT 655.950 596.400 676.050 597.600 ;
        RECT 655.950 595.950 658.050 596.400 ;
        RECT 673.950 595.950 676.050 596.400 ;
        RECT 712.950 597.600 715.050 598.050 ;
        RECT 727.950 597.600 730.050 598.050 ;
        RECT 740.400 597.600 741.600 598.950 ;
        RECT 712.950 596.400 741.600 597.600 ;
        RECT 757.950 597.600 760.050 598.050 ;
        RECT 772.950 597.600 775.050 598.050 ;
        RECT 757.950 596.400 775.050 597.600 ;
        RECT 782.400 597.600 783.600 598.950 ;
        RECT 784.950 597.600 787.050 598.050 ;
        RECT 782.400 596.400 787.050 597.600 ;
        RECT 712.950 595.950 715.050 596.400 ;
        RECT 727.950 595.950 730.050 596.400 ;
        RECT 757.950 595.950 760.050 596.400 ;
        RECT 772.950 595.950 775.050 596.400 ;
        RECT 784.950 595.950 787.050 596.400 ;
        RECT 796.950 597.600 799.050 598.050 ;
        RECT 847.950 597.600 850.050 598.050 ;
        RECT 853.950 597.600 856.050 598.050 ;
        RECT 796.950 596.400 850.050 597.600 ;
        RECT 796.950 595.950 799.050 596.400 ;
        RECT 847.950 595.950 850.050 596.400 ;
        RECT 851.400 596.400 856.050 597.600 ;
        RECT 607.950 594.600 610.050 595.050 ;
        RECT 587.400 593.400 610.050 594.600 ;
        RECT 466.950 592.950 469.050 593.400 ;
        RECT 469.950 592.950 472.050 593.400 ;
        RECT 499.950 592.950 502.050 593.400 ;
        RECT 607.950 592.950 610.050 593.400 ;
        RECT 640.950 594.600 643.050 595.050 ;
        RECT 652.950 594.600 655.050 595.050 ;
        RECT 640.950 593.400 655.050 594.600 ;
        RECT 640.950 592.950 643.050 593.400 ;
        RECT 652.950 592.950 655.050 593.400 ;
        RECT 799.950 594.600 802.050 595.050 ;
        RECT 805.950 594.600 808.050 595.050 ;
        RECT 799.950 593.400 808.050 594.600 ;
        RECT 799.950 592.950 802.050 593.400 ;
        RECT 805.950 592.950 808.050 593.400 ;
        RECT 22.950 591.600 25.050 592.050 ;
        RECT 34.950 591.600 37.050 592.050 ;
        RECT 22.950 590.400 37.050 591.600 ;
        RECT 22.950 589.950 25.050 590.400 ;
        RECT 34.950 589.950 37.050 590.400 ;
        RECT 43.950 591.600 46.050 592.050 ;
        RECT 64.950 591.600 67.050 592.050 ;
        RECT 43.950 590.400 67.050 591.600 ;
        RECT 43.950 589.950 46.050 590.400 ;
        RECT 64.950 589.950 67.050 590.400 ;
        RECT 250.950 591.600 253.050 592.050 ;
        RECT 295.950 591.600 298.050 592.050 ;
        RECT 250.950 590.400 298.050 591.600 ;
        RECT 368.400 591.600 369.600 592.950 ;
        RECT 370.950 591.600 373.050 592.050 ;
        RECT 376.950 591.600 379.050 592.050 ;
        RECT 368.400 590.400 379.050 591.600 ;
        RECT 250.950 589.950 253.050 590.400 ;
        RECT 295.950 589.950 298.050 590.400 ;
        RECT 370.950 589.950 373.050 590.400 ;
        RECT 376.950 589.950 379.050 590.400 ;
        RECT 583.950 591.600 586.050 592.050 ;
        RECT 589.950 591.600 592.050 592.050 ;
        RECT 694.950 591.600 697.050 592.050 ;
        RECT 583.950 590.400 697.050 591.600 ;
        RECT 851.400 591.600 852.600 596.400 ;
        RECT 853.950 595.950 856.050 596.400 ;
        RECT 862.950 595.950 865.050 598.050 ;
        RECT 853.950 594.600 856.050 595.050 ;
        RECT 863.400 594.600 864.600 595.950 ;
        RECT 853.950 593.400 864.600 594.600 ;
        RECT 853.950 592.950 856.050 593.400 ;
        RECT 856.950 591.600 859.050 592.050 ;
        RECT 851.400 590.400 859.050 591.600 ;
        RECT 866.400 591.600 867.600 601.950 ;
        RECT 869.400 598.050 870.600 601.950 ;
        RECT 874.950 600.600 877.050 601.050 ;
        RECT 872.400 599.400 877.050 600.600 ;
        RECT 868.950 595.950 871.050 598.050 ;
        RECT 872.400 595.050 873.600 599.400 ;
        RECT 874.950 598.950 877.050 599.400 ;
        RECT 874.950 597.600 877.050 598.050 ;
        RECT 880.950 597.600 883.050 598.050 ;
        RECT 874.950 596.400 883.050 597.600 ;
        RECT 874.950 595.950 877.050 596.400 ;
        RECT 880.950 595.950 883.050 596.400 ;
        RECT 871.950 592.950 874.050 595.050 ;
        RECT 874.950 591.600 877.050 592.050 ;
        RECT 866.400 590.400 877.050 591.600 ;
        RECT 583.950 589.950 586.050 590.400 ;
        RECT 589.950 589.950 592.050 590.400 ;
        RECT 694.950 589.950 697.050 590.400 ;
        RECT 856.950 589.950 859.050 590.400 ;
        RECT 874.950 589.950 877.050 590.400 ;
        RECT 256.950 588.600 259.050 589.050 ;
        RECT 331.950 588.600 334.050 589.050 ;
        RECT 478.950 588.600 481.050 589.050 ;
        RECT 256.950 587.400 481.050 588.600 ;
        RECT 256.950 586.950 259.050 587.400 ;
        RECT 331.950 586.950 334.050 587.400 ;
        RECT 478.950 586.950 481.050 587.400 ;
        RECT 625.950 588.600 628.050 589.050 ;
        RECT 679.950 588.600 682.050 589.050 ;
        RECT 625.950 587.400 682.050 588.600 ;
        RECT 625.950 586.950 628.050 587.400 ;
        RECT 679.950 586.950 682.050 587.400 ;
        RECT 688.950 588.600 691.050 589.050 ;
        RECT 709.950 588.600 712.050 589.050 ;
        RECT 688.950 587.400 712.050 588.600 ;
        RECT 688.950 586.950 691.050 587.400 ;
        RECT 709.950 586.950 712.050 587.400 ;
        RECT 634.950 585.600 637.050 586.050 ;
        RECT 664.950 585.600 667.050 586.050 ;
        RECT 634.950 584.400 667.050 585.600 ;
        RECT 634.950 583.950 637.050 584.400 ;
        RECT 664.950 583.950 667.050 584.400 ;
        RECT 259.950 582.600 262.050 583.050 ;
        RECT 268.950 582.600 271.050 583.050 ;
        RECT 259.950 581.400 271.050 582.600 ;
        RECT 259.950 580.950 262.050 581.400 ;
        RECT 268.950 580.950 271.050 581.400 ;
        RECT 403.950 582.600 406.050 583.050 ;
        RECT 430.950 582.600 433.050 583.050 ;
        RECT 481.950 582.600 484.050 583.050 ;
        RECT 403.950 581.400 484.050 582.600 ;
        RECT 403.950 580.950 406.050 581.400 ;
        RECT 430.950 580.950 433.050 581.400 ;
        RECT 481.950 580.950 484.050 581.400 ;
        RECT 736.950 582.600 739.050 583.050 ;
        RECT 745.950 582.600 748.050 583.050 ;
        RECT 736.950 581.400 748.050 582.600 ;
        RECT 736.950 580.950 739.050 581.400 ;
        RECT 745.950 580.950 748.050 581.400 ;
        RECT 514.950 579.600 517.050 580.050 ;
        RECT 706.950 579.600 709.050 580.050 ;
        RECT 514.950 578.400 709.050 579.600 ;
        RECT 514.950 577.950 517.050 578.400 ;
        RECT 706.950 577.950 709.050 578.400 ;
        RECT 781.950 579.600 784.050 580.050 ;
        RECT 814.950 579.600 817.050 580.050 ;
        RECT 781.950 578.400 817.050 579.600 ;
        RECT 781.950 577.950 784.050 578.400 ;
        RECT 814.950 577.950 817.050 578.400 ;
        RECT 685.950 576.600 688.050 577.050 ;
        RECT 748.950 576.600 751.050 577.050 ;
        RECT 793.950 576.600 796.050 577.050 ;
        RECT 685.950 575.400 796.050 576.600 ;
        RECT 685.950 574.950 688.050 575.400 ;
        RECT 748.950 574.950 751.050 575.400 ;
        RECT 793.950 574.950 796.050 575.400 ;
        RECT 232.950 573.600 235.050 574.050 ;
        RECT 346.950 573.600 349.050 574.050 ;
        RECT 232.950 572.400 349.050 573.600 ;
        RECT 232.950 571.950 235.050 572.400 ;
        RECT 346.950 571.950 349.050 572.400 ;
        RECT 538.950 573.600 541.050 574.050 ;
        RECT 574.950 573.600 577.050 574.050 ;
        RECT 538.950 572.400 577.050 573.600 ;
        RECT 538.950 571.950 541.050 572.400 ;
        RECT 574.950 571.950 577.050 572.400 ;
        RECT 781.950 573.600 784.050 574.050 ;
        RECT 790.950 573.600 793.050 574.050 ;
        RECT 781.950 572.400 793.050 573.600 ;
        RECT 781.950 571.950 784.050 572.400 ;
        RECT 790.950 571.950 793.050 572.400 ;
        RECT 67.950 570.600 70.050 571.050 ;
        RECT 400.950 570.600 403.050 571.050 ;
        RECT 67.950 569.400 403.050 570.600 ;
        RECT 67.950 568.950 70.050 569.400 ;
        RECT 400.950 568.950 403.050 569.400 ;
        RECT 730.950 570.600 733.050 571.050 ;
        RECT 793.950 570.600 796.050 571.050 ;
        RECT 730.950 569.400 796.050 570.600 ;
        RECT 730.950 568.950 733.050 569.400 ;
        RECT 793.950 568.950 796.050 569.400 ;
        RECT 130.950 567.600 133.050 568.050 ;
        RECT 166.950 567.600 169.050 568.050 ;
        RECT 130.950 566.400 169.050 567.600 ;
        RECT 130.950 565.950 133.050 566.400 ;
        RECT 166.950 565.950 169.050 566.400 ;
        RECT 244.950 567.600 247.050 568.050 ;
        RECT 280.950 567.600 283.050 568.050 ;
        RECT 391.950 567.600 394.050 568.050 ;
        RECT 244.950 566.400 394.050 567.600 ;
        RECT 244.950 565.950 247.050 566.400 ;
        RECT 280.950 565.950 283.050 566.400 ;
        RECT 391.950 565.950 394.050 566.400 ;
        RECT 136.950 564.600 139.050 565.050 ;
        RECT 151.950 564.600 154.050 565.050 ;
        RECT 136.950 563.400 154.050 564.600 ;
        RECT 136.950 562.950 139.050 563.400 ;
        RECT 151.950 562.950 154.050 563.400 ;
        RECT 292.950 564.600 295.050 565.050 ;
        RECT 304.950 564.600 307.050 565.050 ;
        RECT 292.950 563.400 307.050 564.600 ;
        RECT 292.950 562.950 295.050 563.400 ;
        RECT 304.950 562.950 307.050 563.400 ;
        RECT 325.950 564.600 328.050 565.050 ;
        RECT 337.950 564.600 340.050 565.050 ;
        RECT 355.950 564.600 358.050 565.050 ;
        RECT 325.950 563.400 358.050 564.600 ;
        RECT 325.950 562.950 328.050 563.400 ;
        RECT 337.950 562.950 340.050 563.400 ;
        RECT 355.950 562.950 358.050 563.400 ;
        RECT 403.950 564.600 406.050 565.050 ;
        RECT 415.950 564.600 418.050 565.050 ;
        RECT 505.950 564.600 508.050 565.050 ;
        RECT 403.950 563.400 508.050 564.600 ;
        RECT 403.950 562.950 406.050 563.400 ;
        RECT 415.950 562.950 418.050 563.400 ;
        RECT 505.950 562.950 508.050 563.400 ;
        RECT 727.950 564.600 730.050 565.050 ;
        RECT 790.950 564.600 793.050 565.050 ;
        RECT 727.950 563.400 793.050 564.600 ;
        RECT 727.950 562.950 730.050 563.400 ;
        RECT 790.950 562.950 793.050 563.400 ;
        RECT 796.950 564.600 799.050 565.050 ;
        RECT 832.950 564.600 835.050 565.050 ;
        RECT 865.950 564.600 868.050 565.050 ;
        RECT 796.950 563.400 868.050 564.600 ;
        RECT 796.950 562.950 799.050 563.400 ;
        RECT 832.950 562.950 835.050 563.400 ;
        RECT 865.950 562.950 868.050 563.400 ;
        RECT 871.950 564.600 874.050 565.050 ;
        RECT 871.950 563.400 876.600 564.600 ;
        RECT 871.950 562.950 874.050 563.400 ;
        RECT 46.950 561.600 49.050 562.050 ;
        RECT 52.950 561.600 55.050 562.050 ;
        RECT 46.950 560.400 55.050 561.600 ;
        RECT 46.950 559.950 49.050 560.400 ;
        RECT 52.950 559.950 55.050 560.400 ;
        RECT 58.950 561.600 61.050 562.050 ;
        RECT 61.950 561.600 64.050 562.050 ;
        RECT 76.950 561.600 79.050 562.050 ;
        RECT 58.950 560.400 79.050 561.600 ;
        RECT 58.950 559.950 61.050 560.400 ;
        RECT 61.950 559.950 64.050 560.400 ;
        RECT 76.950 559.950 79.050 560.400 ;
        RECT 130.950 561.600 133.050 562.050 ;
        RECT 142.950 561.600 145.050 562.050 ;
        RECT 130.950 560.400 145.050 561.600 ;
        RECT 130.950 559.950 133.050 560.400 ;
        RECT 142.950 559.950 145.050 560.400 ;
        RECT 160.950 561.600 163.050 562.050 ;
        RECT 172.950 561.600 175.050 562.050 ;
        RECT 160.950 560.400 175.050 561.600 ;
        RECT 160.950 559.950 163.050 560.400 ;
        RECT 172.950 559.950 175.050 560.400 ;
        RECT 208.950 561.600 211.050 562.050 ;
        RECT 232.950 561.600 235.050 562.050 ;
        RECT 208.950 560.400 235.050 561.600 ;
        RECT 208.950 559.950 211.050 560.400 ;
        RECT 232.950 559.950 235.050 560.400 ;
        RECT 274.950 561.600 277.050 562.050 ;
        RECT 289.950 561.600 292.050 562.050 ;
        RECT 274.950 560.400 292.050 561.600 ;
        RECT 274.950 559.950 277.050 560.400 ;
        RECT 289.950 559.950 292.050 560.400 ;
        RECT 301.950 561.600 304.050 562.050 ;
        RECT 307.950 561.600 310.050 562.050 ;
        RECT 343.950 561.600 346.050 562.050 ;
        RECT 301.950 560.400 310.050 561.600 ;
        RECT 301.950 559.950 304.050 560.400 ;
        RECT 307.950 559.950 310.050 560.400 ;
        RECT 332.400 560.400 346.050 561.600 ;
        RECT 332.400 559.050 333.600 560.400 ;
        RECT 343.950 559.950 346.050 560.400 ;
        RECT 376.950 561.600 379.050 562.050 ;
        RECT 382.950 561.600 385.050 562.050 ;
        RECT 397.950 561.600 400.050 562.050 ;
        RECT 376.950 560.400 400.050 561.600 ;
        RECT 376.950 559.950 379.050 560.400 ;
        RECT 382.950 559.950 385.050 560.400 ;
        RECT 397.950 559.950 400.050 560.400 ;
        RECT 424.950 561.600 427.050 562.050 ;
        RECT 433.950 561.600 436.050 562.050 ;
        RECT 424.950 560.400 436.050 561.600 ;
        RECT 424.950 559.950 427.050 560.400 ;
        RECT 433.950 559.950 436.050 560.400 ;
        RECT 478.950 561.600 481.050 562.050 ;
        RECT 487.950 561.600 490.050 562.050 ;
        RECT 520.950 561.600 523.050 562.050 ;
        RECT 556.950 561.600 559.050 562.050 ;
        RECT 652.950 561.600 655.050 562.050 ;
        RECT 478.950 560.400 523.050 561.600 ;
        RECT 478.950 559.950 481.050 560.400 ;
        RECT 487.950 559.950 490.050 560.400 ;
        RECT 520.950 559.950 523.050 560.400 ;
        RECT 548.400 560.400 559.050 561.600 ;
        RECT 19.950 558.600 22.050 559.050 ;
        RECT 37.950 558.600 40.050 559.050 ;
        RECT 19.950 557.400 40.050 558.600 ;
        RECT 19.950 556.950 22.050 557.400 ;
        RECT 37.950 556.950 40.050 557.400 ;
        RECT 40.950 558.600 43.050 559.050 ;
        RECT 55.950 558.600 58.050 559.050 ;
        RECT 40.950 557.400 58.050 558.600 ;
        RECT 40.950 556.950 43.050 557.400 ;
        RECT 55.950 556.950 58.050 557.400 ;
        RECT 79.950 556.950 82.050 559.050 ;
        RECT 115.950 558.600 118.050 559.050 ;
        RECT 139.950 558.600 142.050 559.050 ;
        RECT 115.950 557.400 142.050 558.600 ;
        RECT 115.950 556.950 118.050 557.400 ;
        RECT 139.950 556.950 142.050 557.400 ;
        RECT 163.950 558.600 166.050 559.050 ;
        RECT 193.950 558.600 196.050 559.050 ;
        RECT 163.950 557.400 196.050 558.600 ;
        RECT 163.950 556.950 166.050 557.400 ;
        RECT 193.950 556.950 196.050 557.400 ;
        RECT 211.950 558.600 214.050 559.050 ;
        RECT 226.950 558.600 229.050 559.050 ;
        RECT 211.950 557.400 229.050 558.600 ;
        RECT 211.950 556.950 214.050 557.400 ;
        RECT 226.950 556.950 229.050 557.400 ;
        RECT 250.950 558.600 253.050 559.050 ;
        RECT 268.950 558.600 271.050 559.050 ;
        RECT 250.950 557.400 271.050 558.600 ;
        RECT 250.950 556.950 253.050 557.400 ;
        RECT 268.950 556.950 271.050 557.400 ;
        RECT 271.950 558.600 274.050 559.050 ;
        RECT 280.950 558.600 283.050 559.050 ;
        RECT 271.950 557.400 283.050 558.600 ;
        RECT 271.950 556.950 274.050 557.400 ;
        RECT 280.950 556.950 283.050 557.400 ;
        RECT 292.950 558.600 295.050 559.050 ;
        RECT 310.950 558.600 313.050 559.050 ;
        RECT 292.950 557.400 313.050 558.600 ;
        RECT 292.950 556.950 295.050 557.400 ;
        RECT 310.950 556.950 313.050 557.400 ;
        RECT 331.950 556.950 334.050 559.050 ;
        RECT 352.950 558.600 355.050 559.050 ;
        RECT 341.400 557.400 355.050 558.600 ;
        RECT 70.950 555.600 73.050 556.050 ;
        RECT 76.950 555.600 79.050 556.050 ;
        RECT 70.950 554.400 79.050 555.600 ;
        RECT 70.950 553.950 73.050 554.400 ;
        RECT 76.950 553.950 79.050 554.400 ;
        RECT 10.950 552.600 13.050 553.050 ;
        RECT 61.950 552.600 64.050 553.050 ;
        RECT 10.950 551.400 64.050 552.600 ;
        RECT 80.400 552.600 81.600 556.950 ;
        RECT 341.400 556.050 342.600 557.400 ;
        RECT 352.950 556.950 355.050 557.400 ;
        RECT 355.950 558.600 358.050 559.050 ;
        RECT 373.950 558.600 376.050 559.050 ;
        RECT 412.950 558.600 415.050 559.050 ;
        RECT 355.950 557.400 415.050 558.600 ;
        RECT 355.950 556.950 358.050 557.400 ;
        RECT 373.950 556.950 376.050 557.400 ;
        RECT 412.950 556.950 415.050 557.400 ;
        RECT 505.950 558.600 508.050 559.050 ;
        RECT 526.950 558.600 529.050 559.050 ;
        RECT 505.950 557.400 529.050 558.600 ;
        RECT 505.950 556.950 508.050 557.400 ;
        RECT 526.950 556.950 529.050 557.400 ;
        RECT 548.400 556.050 549.600 560.400 ;
        RECT 556.950 559.950 559.050 560.400 ;
        RECT 638.400 560.400 655.050 561.600 ;
        RECT 638.400 559.050 639.600 560.400 ;
        RECT 652.950 559.950 655.050 560.400 ;
        RECT 736.950 561.600 739.050 562.050 ;
        RECT 778.950 561.600 781.050 562.050 ;
        RECT 832.950 561.600 835.050 562.050 ;
        RECT 736.950 560.400 835.050 561.600 ;
        RECT 736.950 559.950 739.050 560.400 ;
        RECT 778.950 559.950 781.050 560.400 ;
        RECT 832.950 559.950 835.050 560.400 ;
        RECT 850.950 561.600 853.050 562.050 ;
        RECT 862.950 561.600 865.050 562.050 ;
        RECT 871.950 561.600 874.050 562.050 ;
        RECT 850.950 560.400 874.050 561.600 ;
        RECT 850.950 559.950 853.050 560.400 ;
        RECT 862.950 559.950 865.050 560.400 ;
        RECT 871.950 559.950 874.050 560.400 ;
        RECT 550.950 556.950 553.050 559.050 ;
        RECT 556.950 558.600 559.050 559.050 ;
        RECT 571.950 558.600 574.050 559.050 ;
        RECT 595.950 558.600 598.050 559.050 ;
        RECT 556.950 557.400 598.050 558.600 ;
        RECT 556.950 556.950 559.050 557.400 ;
        RECT 571.950 556.950 574.050 557.400 ;
        RECT 595.950 556.950 598.050 557.400 ;
        RECT 604.950 558.600 607.050 559.050 ;
        RECT 610.950 558.600 613.050 559.050 ;
        RECT 637.950 558.600 640.050 559.050 ;
        RECT 658.950 558.600 661.050 559.050 ;
        RECT 754.950 558.600 757.050 559.050 ;
        RECT 769.950 558.600 772.050 559.050 ;
        RECT 604.950 557.400 613.050 558.600 ;
        RECT 604.950 556.950 607.050 557.400 ;
        RECT 610.950 556.950 613.050 557.400 ;
        RECT 623.400 557.400 640.050 558.600 ;
        RECT 88.950 555.600 91.050 556.050 ;
        RECT 100.950 555.600 103.050 556.050 ;
        RECT 118.950 555.600 121.050 556.050 ;
        RECT 88.950 554.400 121.050 555.600 ;
        RECT 88.950 553.950 91.050 554.400 ;
        RECT 100.950 553.950 103.050 554.400 ;
        RECT 118.950 553.950 121.050 554.400 ;
        RECT 154.950 555.600 157.050 556.050 ;
        RECT 181.950 555.600 184.050 556.050 ;
        RECT 235.950 555.600 238.050 556.050 ;
        RECT 154.950 554.400 238.050 555.600 ;
        RECT 154.950 553.950 157.050 554.400 ;
        RECT 181.950 553.950 184.050 554.400 ;
        RECT 235.950 553.950 238.050 554.400 ;
        RECT 316.950 555.600 319.050 556.050 ;
        RECT 334.950 555.600 337.050 556.050 ;
        RECT 316.950 554.400 337.050 555.600 ;
        RECT 316.950 553.950 319.050 554.400 ;
        RECT 334.950 553.950 337.050 554.400 ;
        RECT 340.950 553.950 343.050 556.050 ;
        RECT 343.950 555.600 346.050 556.050 ;
        RECT 379.950 555.600 382.050 556.050 ;
        RECT 418.950 555.600 421.050 556.050 ;
        RECT 451.950 555.600 454.050 556.050 ;
        RECT 343.950 554.400 454.050 555.600 ;
        RECT 343.950 553.950 346.050 554.400 ;
        RECT 379.950 553.950 382.050 554.400 ;
        RECT 418.950 553.950 421.050 554.400 ;
        RECT 451.950 553.950 454.050 554.400 ;
        RECT 457.950 555.600 460.050 556.050 ;
        RECT 466.950 555.600 469.050 556.050 ;
        RECT 457.950 554.400 469.050 555.600 ;
        RECT 457.950 553.950 460.050 554.400 ;
        RECT 466.950 553.950 469.050 554.400 ;
        RECT 484.950 555.600 487.050 556.050 ;
        RECT 502.950 555.600 505.050 556.050 ;
        RECT 484.950 554.400 505.050 555.600 ;
        RECT 484.950 553.950 487.050 554.400 ;
        RECT 502.950 553.950 505.050 554.400 ;
        RECT 529.950 555.600 532.050 556.050 ;
        RECT 544.950 555.600 547.050 556.050 ;
        RECT 529.950 554.400 547.050 555.600 ;
        RECT 529.950 553.950 532.050 554.400 ;
        RECT 544.950 553.950 547.050 554.400 ;
        RECT 547.950 553.950 550.050 556.050 ;
        RECT 551.400 555.600 552.600 556.950 ;
        RECT 565.950 555.600 568.050 556.050 ;
        RECT 551.400 554.400 568.050 555.600 ;
        RECT 565.950 553.950 568.050 554.400 ;
        RECT 613.950 555.600 616.050 556.050 ;
        RECT 623.400 555.600 624.600 557.400 ;
        RECT 637.950 556.950 640.050 557.400 ;
        RECT 641.400 557.400 661.050 558.600 ;
        RECT 613.950 554.400 624.600 555.600 ;
        RECT 625.950 555.600 628.050 556.050 ;
        RECT 631.950 555.600 634.050 556.050 ;
        RECT 641.400 555.600 642.600 557.400 ;
        RECT 658.950 556.950 661.050 557.400 ;
        RECT 740.400 557.400 772.050 558.600 ;
        RECT 740.400 556.050 741.600 557.400 ;
        RECT 754.950 556.950 757.050 557.400 ;
        RECT 769.950 556.950 772.050 557.400 ;
        RECT 790.950 558.600 793.050 559.050 ;
        RECT 805.950 558.600 808.050 559.050 ;
        RECT 790.950 557.400 808.050 558.600 ;
        RECT 790.950 556.950 793.050 557.400 ;
        RECT 805.950 556.950 808.050 557.400 ;
        RECT 856.950 558.600 859.050 559.050 ;
        RECT 868.950 558.600 871.050 559.050 ;
        RECT 856.950 557.400 871.050 558.600 ;
        RECT 856.950 556.950 859.050 557.400 ;
        RECT 868.950 556.950 871.050 557.400 ;
        RECT 625.950 554.400 642.600 555.600 ;
        RECT 682.950 555.600 685.050 556.050 ;
        RECT 703.950 555.600 706.050 556.050 ;
        RECT 682.950 554.400 706.050 555.600 ;
        RECT 613.950 553.950 616.050 554.400 ;
        RECT 625.950 553.950 628.050 554.400 ;
        RECT 631.950 553.950 634.050 554.400 ;
        RECT 682.950 553.950 685.050 554.400 ;
        RECT 703.950 553.950 706.050 554.400 ;
        RECT 706.950 555.600 709.050 556.050 ;
        RECT 733.950 555.600 736.050 556.050 ;
        RECT 706.950 554.400 736.050 555.600 ;
        RECT 706.950 553.950 709.050 554.400 ;
        RECT 733.950 553.950 736.050 554.400 ;
        RECT 739.950 553.950 742.050 556.050 ;
        RECT 748.950 555.600 751.050 556.050 ;
        RECT 808.950 555.600 811.050 556.050 ;
        RECT 748.950 554.400 811.050 555.600 ;
        RECT 748.950 553.950 751.050 554.400 ;
        RECT 808.950 553.950 811.050 554.400 ;
        RECT 868.950 555.600 871.050 556.050 ;
        RECT 875.400 555.600 876.600 563.400 ;
        RECT 868.950 554.400 876.600 555.600 ;
        RECT 868.950 553.950 871.050 554.400 ;
        RECT 97.950 552.600 100.050 553.050 ;
        RECT 80.400 551.400 100.050 552.600 ;
        RECT 10.950 550.950 13.050 551.400 ;
        RECT 61.950 550.950 64.050 551.400 ;
        RECT 97.950 550.950 100.050 551.400 ;
        RECT 112.950 552.600 115.050 553.050 ;
        RECT 121.950 552.600 124.050 553.050 ;
        RECT 112.950 551.400 124.050 552.600 ;
        RECT 112.950 550.950 115.050 551.400 ;
        RECT 121.950 550.950 124.050 551.400 ;
        RECT 139.950 552.600 142.050 553.050 ;
        RECT 205.950 552.600 208.050 553.050 ;
        RECT 139.950 551.400 208.050 552.600 ;
        RECT 139.950 550.950 142.050 551.400 ;
        RECT 205.950 550.950 208.050 551.400 ;
        RECT 235.950 552.600 238.050 553.050 ;
        RECT 247.950 552.600 250.050 553.050 ;
        RECT 265.950 552.600 268.050 553.050 ;
        RECT 235.950 551.400 268.050 552.600 ;
        RECT 235.950 550.950 238.050 551.400 ;
        RECT 247.950 550.950 250.050 551.400 ;
        RECT 265.950 550.950 268.050 551.400 ;
        RECT 355.950 552.600 358.050 553.050 ;
        RECT 382.950 552.600 385.050 553.050 ;
        RECT 355.950 551.400 385.050 552.600 ;
        RECT 355.950 550.950 358.050 551.400 ;
        RECT 382.950 550.950 385.050 551.400 ;
        RECT 394.950 552.600 397.050 553.050 ;
        RECT 403.950 552.600 406.050 553.050 ;
        RECT 394.950 551.400 406.050 552.600 ;
        RECT 394.950 550.950 397.050 551.400 ;
        RECT 403.950 550.950 406.050 551.400 ;
        RECT 508.950 552.600 511.050 553.050 ;
        RECT 601.950 552.600 604.050 553.050 ;
        RECT 607.950 552.600 610.050 553.050 ;
        RECT 508.950 551.400 610.050 552.600 ;
        RECT 508.950 550.950 511.050 551.400 ;
        RECT 601.950 550.950 604.050 551.400 ;
        RECT 607.950 550.950 610.050 551.400 ;
        RECT 739.950 552.600 742.050 553.050 ;
        RECT 745.950 552.600 748.050 553.050 ;
        RECT 739.950 551.400 748.050 552.600 ;
        RECT 739.950 550.950 742.050 551.400 ;
        RECT 745.950 550.950 748.050 551.400 ;
        RECT 775.950 552.600 778.050 553.050 ;
        RECT 784.950 552.600 787.050 553.050 ;
        RECT 775.950 551.400 787.050 552.600 ;
        RECT 775.950 550.950 778.050 551.400 ;
        RECT 784.950 550.950 787.050 551.400 ;
        RECT 811.950 552.600 814.050 553.050 ;
        RECT 829.950 552.600 832.050 553.050 ;
        RECT 847.950 552.600 850.050 553.050 ;
        RECT 811.950 551.400 850.050 552.600 ;
        RECT 811.950 550.950 814.050 551.400 ;
        RECT 829.950 550.950 832.050 551.400 ;
        RECT 847.950 550.950 850.050 551.400 ;
        RECT 871.950 552.600 874.050 553.050 ;
        RECT 880.950 552.600 883.050 553.050 ;
        RECT 871.950 551.400 883.050 552.600 ;
        RECT 871.950 550.950 874.050 551.400 ;
        RECT 880.950 550.950 883.050 551.400 ;
        RECT 73.950 549.600 76.050 550.050 ;
        RECT 82.950 549.600 85.050 550.050 ;
        RECT 73.950 548.400 85.050 549.600 ;
        RECT 73.950 547.950 76.050 548.400 ;
        RECT 82.950 547.950 85.050 548.400 ;
        RECT 91.950 549.600 94.050 550.050 ;
        RECT 97.950 549.600 100.050 550.050 ;
        RECT 91.950 548.400 100.050 549.600 ;
        RECT 91.950 547.950 94.050 548.400 ;
        RECT 97.950 547.950 100.050 548.400 ;
        RECT 124.950 549.600 127.050 550.050 ;
        RECT 178.950 549.600 181.050 550.050 ;
        RECT 277.950 549.600 280.050 550.050 ;
        RECT 292.950 549.600 295.050 550.050 ;
        RECT 457.950 549.600 460.050 550.050 ;
        RECT 124.950 548.400 181.050 549.600 ;
        RECT 124.950 547.950 127.050 548.400 ;
        RECT 178.950 547.950 181.050 548.400 ;
        RECT 182.400 548.400 460.050 549.600 ;
        RECT 106.950 546.600 109.050 547.050 ;
        RECT 160.950 546.600 163.050 547.050 ;
        RECT 182.400 546.600 183.600 548.400 ;
        RECT 277.950 547.950 280.050 548.400 ;
        RECT 292.950 547.950 295.050 548.400 ;
        RECT 457.950 547.950 460.050 548.400 ;
        RECT 532.950 549.600 535.050 550.050 ;
        RECT 589.950 549.600 592.050 550.050 ;
        RECT 532.950 548.400 592.050 549.600 ;
        RECT 532.950 547.950 535.050 548.400 ;
        RECT 589.950 547.950 592.050 548.400 ;
        RECT 598.950 549.600 601.050 550.050 ;
        RECT 634.950 549.600 637.050 550.050 ;
        RECT 655.950 549.600 658.050 550.050 ;
        RECT 598.950 548.400 658.050 549.600 ;
        RECT 598.950 547.950 601.050 548.400 ;
        RECT 634.950 547.950 637.050 548.400 ;
        RECT 655.950 547.950 658.050 548.400 ;
        RECT 715.950 549.600 718.050 550.050 ;
        RECT 733.950 549.600 736.050 550.050 ;
        RECT 715.950 548.400 736.050 549.600 ;
        RECT 715.950 547.950 718.050 548.400 ;
        RECT 733.950 547.950 736.050 548.400 ;
        RECT 763.950 549.600 766.050 550.050 ;
        RECT 787.950 549.600 790.050 550.050 ;
        RECT 763.950 548.400 790.050 549.600 ;
        RECT 763.950 547.950 766.050 548.400 ;
        RECT 787.950 547.950 790.050 548.400 ;
        RECT 106.950 545.400 183.600 546.600 ;
        RECT 259.950 546.600 262.050 547.050 ;
        RECT 277.950 546.600 280.050 547.050 ;
        RECT 259.950 545.400 280.050 546.600 ;
        RECT 106.950 544.950 109.050 545.400 ;
        RECT 160.950 544.950 163.050 545.400 ;
        RECT 259.950 544.950 262.050 545.400 ;
        RECT 277.950 544.950 280.050 545.400 ;
        RECT 406.950 546.600 409.050 547.050 ;
        RECT 532.950 546.600 535.050 547.050 ;
        RECT 406.950 545.400 535.050 546.600 ;
        RECT 406.950 544.950 409.050 545.400 ;
        RECT 532.950 544.950 535.050 545.400 ;
        RECT 544.950 546.600 547.050 547.050 ;
        RECT 553.950 546.600 556.050 547.050 ;
        RECT 568.950 546.600 571.050 547.050 ;
        RECT 544.950 545.400 571.050 546.600 ;
        RECT 544.950 544.950 547.050 545.400 ;
        RECT 553.950 544.950 556.050 545.400 ;
        RECT 568.950 544.950 571.050 545.400 ;
        RECT 670.950 546.600 673.050 547.050 ;
        RECT 718.950 546.600 721.050 547.050 ;
        RECT 778.950 546.600 781.050 547.050 ;
        RECT 670.950 545.400 781.050 546.600 ;
        RECT 670.950 544.950 673.050 545.400 ;
        RECT 718.950 544.950 721.050 545.400 ;
        RECT 778.950 544.950 781.050 545.400 ;
        RECT 247.950 543.600 250.050 544.050 ;
        RECT 484.950 543.600 487.050 544.050 ;
        RECT 247.950 542.400 487.050 543.600 ;
        RECT 247.950 541.950 250.050 542.400 ;
        RECT 484.950 541.950 487.050 542.400 ;
        RECT 553.950 543.600 556.050 544.050 ;
        RECT 586.950 543.600 589.050 544.050 ;
        RECT 553.950 542.400 589.050 543.600 ;
        RECT 553.950 541.950 556.050 542.400 ;
        RECT 586.950 541.950 589.050 542.400 ;
        RECT 613.950 543.600 616.050 544.050 ;
        RECT 646.950 543.600 649.050 544.050 ;
        RECT 613.950 542.400 649.050 543.600 ;
        RECT 613.950 541.950 616.050 542.400 ;
        RECT 646.950 541.950 649.050 542.400 ;
        RECT 658.950 543.600 661.050 544.050 ;
        RECT 688.950 543.600 691.050 544.050 ;
        RECT 658.950 542.400 691.050 543.600 ;
        RECT 658.950 541.950 661.050 542.400 ;
        RECT 688.950 541.950 691.050 542.400 ;
        RECT 13.950 540.600 16.050 541.050 ;
        RECT 34.950 540.600 37.050 541.050 ;
        RECT 46.950 540.600 49.050 541.050 ;
        RECT 13.950 539.400 49.050 540.600 ;
        RECT 13.950 538.950 16.050 539.400 ;
        RECT 34.950 538.950 37.050 539.400 ;
        RECT 46.950 538.950 49.050 539.400 ;
        RECT 418.950 540.600 421.050 541.050 ;
        RECT 430.950 540.600 433.050 541.050 ;
        RECT 418.950 539.400 433.050 540.600 ;
        RECT 418.950 538.950 421.050 539.400 ;
        RECT 430.950 538.950 433.050 539.400 ;
        RECT 436.950 540.600 439.050 541.050 ;
        RECT 457.950 540.600 460.050 541.050 ;
        RECT 436.950 539.400 460.050 540.600 ;
        RECT 436.950 538.950 439.050 539.400 ;
        RECT 457.950 538.950 460.050 539.400 ;
        RECT 463.950 540.600 466.050 541.050 ;
        RECT 493.950 540.600 496.050 541.050 ;
        RECT 565.950 540.600 568.050 541.050 ;
        RECT 463.950 539.400 568.050 540.600 ;
        RECT 463.950 538.950 466.050 539.400 ;
        RECT 493.950 538.950 496.050 539.400 ;
        RECT 565.950 538.950 568.050 539.400 ;
        RECT 574.950 540.600 577.050 541.050 ;
        RECT 616.950 540.600 619.050 541.050 ;
        RECT 574.950 539.400 619.050 540.600 ;
        RECT 574.950 538.950 577.050 539.400 ;
        RECT 616.950 538.950 619.050 539.400 ;
        RECT 664.950 540.600 667.050 541.050 ;
        RECT 703.950 540.600 706.050 541.050 ;
        RECT 817.950 540.600 820.050 541.050 ;
        RECT 838.950 540.600 841.050 541.050 ;
        RECT 850.950 540.600 853.050 541.050 ;
        RECT 664.950 539.400 853.050 540.600 ;
        RECT 664.950 538.950 667.050 539.400 ;
        RECT 703.950 538.950 706.050 539.400 ;
        RECT 817.950 538.950 820.050 539.400 ;
        RECT 838.950 538.950 841.050 539.400 ;
        RECT 850.950 538.950 853.050 539.400 ;
        RECT 31.950 537.600 34.050 538.050 ;
        RECT 37.950 537.600 40.050 538.050 ;
        RECT 31.950 536.400 40.050 537.600 ;
        RECT 31.950 535.950 34.050 536.400 ;
        RECT 37.950 535.950 40.050 536.400 ;
        RECT 85.950 537.600 88.050 538.050 ;
        RECT 127.950 537.600 130.050 538.050 ;
        RECT 142.950 537.600 145.050 538.050 ;
        RECT 85.950 536.400 145.050 537.600 ;
        RECT 85.950 535.950 88.050 536.400 ;
        RECT 127.950 535.950 130.050 536.400 ;
        RECT 142.950 535.950 145.050 536.400 ;
        RECT 178.950 537.600 181.050 538.050 ;
        RECT 223.950 537.600 226.050 538.050 ;
        RECT 232.950 537.600 235.050 538.050 ;
        RECT 178.950 536.400 235.050 537.600 ;
        RECT 178.950 535.950 181.050 536.400 ;
        RECT 223.950 535.950 226.050 536.400 ;
        RECT 232.950 535.950 235.050 536.400 ;
        RECT 472.950 537.600 475.050 538.050 ;
        RECT 550.950 537.600 553.050 538.050 ;
        RECT 568.950 537.600 571.050 538.050 ;
        RECT 586.950 537.600 589.050 538.050 ;
        RECT 472.950 536.400 589.050 537.600 ;
        RECT 472.950 535.950 475.050 536.400 ;
        RECT 550.950 535.950 553.050 536.400 ;
        RECT 568.950 535.950 571.050 536.400 ;
        RECT 586.950 535.950 589.050 536.400 ;
        RECT 100.950 534.600 103.050 535.050 ;
        RECT 157.950 534.600 160.050 535.050 ;
        RECT 238.950 534.600 241.050 535.050 ;
        RECT 100.950 533.400 241.050 534.600 ;
        RECT 100.950 532.950 103.050 533.400 ;
        RECT 157.950 532.950 160.050 533.400 ;
        RECT 238.950 532.950 241.050 533.400 ;
        RECT 289.950 534.600 292.050 535.050 ;
        RECT 295.950 534.600 298.050 535.050 ;
        RECT 289.950 533.400 298.050 534.600 ;
        RECT 289.950 532.950 292.050 533.400 ;
        RECT 295.950 532.950 298.050 533.400 ;
        RECT 376.950 534.600 379.050 535.050 ;
        RECT 385.950 534.600 388.050 535.050 ;
        RECT 409.950 534.600 412.050 535.050 ;
        RECT 376.950 533.400 412.050 534.600 ;
        RECT 376.950 532.950 379.050 533.400 ;
        RECT 385.950 532.950 388.050 533.400 ;
        RECT 409.950 532.950 412.050 533.400 ;
        RECT 544.950 534.600 547.050 535.050 ;
        RECT 604.950 534.600 607.050 535.050 ;
        RECT 616.950 534.600 619.050 535.050 ;
        RECT 619.950 534.600 622.050 535.050 ;
        RECT 544.950 533.400 622.050 534.600 ;
        RECT 544.950 532.950 547.050 533.400 ;
        RECT 604.950 532.950 607.050 533.400 ;
        RECT 616.950 532.950 619.050 533.400 ;
        RECT 619.950 532.950 622.050 533.400 ;
        RECT 676.950 534.600 679.050 535.050 ;
        RECT 718.950 534.600 721.050 535.050 ;
        RECT 676.950 533.400 721.050 534.600 ;
        RECT 676.950 532.950 679.050 533.400 ;
        RECT 718.950 532.950 721.050 533.400 ;
        RECT 25.950 531.600 28.050 532.050 ;
        RECT 46.950 531.600 49.050 532.050 ;
        RECT 25.950 530.400 49.050 531.600 ;
        RECT 25.950 529.950 28.050 530.400 ;
        RECT 46.950 529.950 49.050 530.400 ;
        RECT 91.950 531.600 94.050 532.050 ;
        RECT 91.950 530.400 117.600 531.600 ;
        RECT 91.950 529.950 94.050 530.400 ;
        RECT 116.400 529.050 117.600 530.400 ;
        RECT 130.950 529.950 133.050 532.050 ;
        RECT 217.950 531.600 220.050 532.050 ;
        RECT 250.950 531.600 253.050 532.050 ;
        RECT 262.950 531.600 265.050 532.050 ;
        RECT 301.950 531.600 304.050 532.050 ;
        RECT 328.950 531.600 331.050 532.050 ;
        RECT 331.950 531.600 334.050 532.050 ;
        RECT 340.950 531.600 343.050 532.050 ;
        RECT 217.950 530.400 304.050 531.600 ;
        RECT 217.950 529.950 220.050 530.400 ;
        RECT 250.950 529.950 253.050 530.400 ;
        RECT 262.950 529.950 265.050 530.400 ;
        RECT 301.950 529.950 304.050 530.400 ;
        RECT 317.400 530.400 343.050 531.600 ;
        RECT 13.950 528.600 16.050 529.050 ;
        RECT 52.950 528.600 55.050 529.050 ;
        RECT 13.950 527.400 55.050 528.600 ;
        RECT 13.950 526.950 16.050 527.400 ;
        RECT 52.950 526.950 55.050 527.400 ;
        RECT 94.950 526.950 97.050 529.050 ;
        RECT 115.950 526.950 118.050 529.050 ;
        RECT 31.950 525.600 34.050 526.050 ;
        RECT 37.950 525.600 40.050 526.050 ;
        RECT 31.950 524.400 40.050 525.600 ;
        RECT 31.950 523.950 34.050 524.400 ;
        RECT 37.950 523.950 40.050 524.400 ;
        RECT 55.950 525.600 58.050 526.050 ;
        RECT 73.950 525.600 76.050 526.050 ;
        RECT 55.950 524.400 76.050 525.600 ;
        RECT 55.950 523.950 58.050 524.400 ;
        RECT 73.950 523.950 76.050 524.400 ;
        RECT 91.950 525.600 94.050 526.050 ;
        RECT 95.400 525.600 96.600 526.950 ;
        RECT 91.950 524.400 96.600 525.600 ;
        RECT 112.950 525.600 115.050 526.050 ;
        RECT 118.950 525.600 121.050 526.050 ;
        RECT 112.950 524.400 121.050 525.600 ;
        RECT 91.950 523.950 94.050 524.400 ;
        RECT 112.950 523.950 115.050 524.400 ;
        RECT 118.950 523.950 121.050 524.400 ;
        RECT 131.400 523.050 132.600 529.950 ;
        RECT 172.950 528.600 175.050 529.050 ;
        RECT 181.950 528.600 184.050 529.050 ;
        RECT 172.950 527.400 184.050 528.600 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 181.950 526.950 184.050 527.400 ;
        RECT 253.950 528.600 256.050 529.050 ;
        RECT 271.950 528.600 274.050 529.050 ;
        RECT 253.950 527.400 274.050 528.600 ;
        RECT 253.950 526.950 256.050 527.400 ;
        RECT 271.950 526.950 274.050 527.400 ;
        RECT 280.950 528.600 283.050 529.050 ;
        RECT 317.400 528.600 318.600 530.400 ;
        RECT 328.950 529.950 331.050 530.400 ;
        RECT 331.950 529.950 334.050 530.400 ;
        RECT 340.950 529.950 343.050 530.400 ;
        RECT 373.950 531.600 376.050 532.050 ;
        RECT 379.950 531.600 382.050 532.050 ;
        RECT 373.950 530.400 382.050 531.600 ;
        RECT 373.950 529.950 376.050 530.400 ;
        RECT 379.950 529.950 382.050 530.400 ;
        RECT 385.950 531.600 388.050 532.050 ;
        RECT 397.950 531.600 400.050 532.050 ;
        RECT 385.950 530.400 400.050 531.600 ;
        RECT 385.950 529.950 388.050 530.400 ;
        RECT 397.950 529.950 400.050 530.400 ;
        RECT 445.950 531.600 448.050 532.050 ;
        RECT 478.950 531.600 481.050 532.050 ;
        RECT 445.950 530.400 481.050 531.600 ;
        RECT 445.950 529.950 448.050 530.400 ;
        RECT 478.950 529.950 481.050 530.400 ;
        RECT 511.950 531.600 514.050 532.050 ;
        RECT 526.950 531.600 529.050 532.050 ;
        RECT 511.950 530.400 529.050 531.600 ;
        RECT 511.950 529.950 514.050 530.400 ;
        RECT 526.950 529.950 529.050 530.400 ;
        RECT 559.950 531.600 562.050 532.050 ;
        RECT 574.950 531.600 577.050 532.050 ;
        RECT 727.950 531.600 730.050 532.050 ;
        RECT 742.950 531.600 745.050 532.050 ;
        RECT 559.950 530.400 577.050 531.600 ;
        RECT 559.950 529.950 562.050 530.400 ;
        RECT 574.950 529.950 577.050 530.400 ;
        RECT 716.400 530.400 745.050 531.600 ;
        RECT 716.400 529.050 717.600 530.400 ;
        RECT 727.950 529.950 730.050 530.400 ;
        RECT 742.950 529.950 745.050 530.400 ;
        RECT 760.950 531.600 763.050 532.050 ;
        RECT 769.950 531.600 772.050 532.050 ;
        RECT 760.950 530.400 772.050 531.600 ;
        RECT 760.950 529.950 763.050 530.400 ;
        RECT 769.950 529.950 772.050 530.400 ;
        RECT 802.950 531.600 805.050 532.050 ;
        RECT 814.950 531.600 817.050 532.050 ;
        RECT 802.950 530.400 817.050 531.600 ;
        RECT 802.950 529.950 805.050 530.400 ;
        RECT 814.950 529.950 817.050 530.400 ;
        RECT 823.950 531.600 826.050 532.050 ;
        RECT 844.950 531.600 847.050 532.050 ;
        RECT 823.950 530.400 847.050 531.600 ;
        RECT 823.950 529.950 826.050 530.400 ;
        RECT 844.950 529.950 847.050 530.400 ;
        RECT 865.950 531.600 868.050 532.050 ;
        RECT 877.950 531.600 880.050 532.050 ;
        RECT 865.950 530.400 880.050 531.600 ;
        RECT 865.950 529.950 868.050 530.400 ;
        RECT 877.950 529.950 880.050 530.400 ;
        RECT 280.950 527.400 318.600 528.600 ;
        RECT 358.950 528.600 361.050 529.050 ;
        RECT 364.950 528.600 367.050 529.050 ;
        RECT 394.950 528.600 397.050 529.050 ;
        RECT 358.950 527.400 397.050 528.600 ;
        RECT 280.950 526.950 283.050 527.400 ;
        RECT 358.950 526.950 361.050 527.400 ;
        RECT 364.950 526.950 367.050 527.400 ;
        RECT 394.950 526.950 397.050 527.400 ;
        RECT 415.950 528.600 418.050 529.050 ;
        RECT 436.950 528.600 439.050 529.050 ;
        RECT 415.950 527.400 439.050 528.600 ;
        RECT 415.950 526.950 418.050 527.400 ;
        RECT 436.950 526.950 439.050 527.400 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 532.950 528.600 535.050 529.050 ;
        RECT 547.950 528.600 550.050 529.050 ;
        RECT 559.950 528.600 562.050 529.050 ;
        RECT 532.950 527.400 546.600 528.600 ;
        RECT 532.950 526.950 535.050 527.400 ;
        RECT 142.950 525.600 145.050 526.050 ;
        RECT 154.950 525.600 157.050 526.050 ;
        RECT 142.950 524.400 157.050 525.600 ;
        RECT 142.950 523.950 145.050 524.400 ;
        RECT 154.950 523.950 157.050 524.400 ;
        RECT 190.950 525.600 193.050 526.050 ;
        RECT 208.950 525.600 211.050 526.050 ;
        RECT 190.950 524.400 211.050 525.600 ;
        RECT 190.950 523.950 193.050 524.400 ;
        RECT 208.950 523.950 211.050 524.400 ;
        RECT 259.950 525.600 262.050 526.050 ;
        RECT 268.950 525.600 271.050 526.050 ;
        RECT 259.950 524.400 271.050 525.600 ;
        RECT 259.950 523.950 262.050 524.400 ;
        RECT 268.950 523.950 271.050 524.400 ;
        RECT 274.950 525.600 277.050 526.050 ;
        RECT 298.950 525.600 301.050 526.050 ;
        RECT 274.950 524.400 301.050 525.600 ;
        RECT 274.950 523.950 277.050 524.400 ;
        RECT 298.950 523.950 301.050 524.400 ;
        RECT 310.950 525.600 313.050 526.050 ;
        RECT 316.950 525.600 319.050 526.050 ;
        RECT 310.950 524.400 319.050 525.600 ;
        RECT 310.950 523.950 313.050 524.400 ;
        RECT 316.950 523.950 319.050 524.400 ;
        RECT 349.950 525.600 352.050 526.050 ;
        RECT 355.950 525.600 358.050 526.050 ;
        RECT 349.950 524.400 358.050 525.600 ;
        RECT 349.950 523.950 352.050 524.400 ;
        RECT 355.950 523.950 358.050 524.400 ;
        RECT 358.950 525.600 361.050 526.050 ;
        RECT 370.950 525.600 373.050 526.050 ;
        RECT 376.950 525.600 379.050 526.050 ;
        RECT 358.950 524.400 379.050 525.600 ;
        RECT 358.950 523.950 361.050 524.400 ;
        RECT 370.950 523.950 373.050 524.400 ;
        RECT 376.950 523.950 379.050 524.400 ;
        RECT 412.950 525.600 415.050 526.050 ;
        RECT 424.950 525.600 427.050 526.050 ;
        RECT 412.950 524.400 427.050 525.600 ;
        RECT 412.950 523.950 415.050 524.400 ;
        RECT 424.950 523.950 427.050 524.400 ;
        RECT 427.950 525.600 430.050 526.050 ;
        RECT 473.400 525.600 474.600 526.950 ;
        RECT 427.950 524.400 474.600 525.600 ;
        RECT 514.950 525.600 517.050 526.050 ;
        RECT 520.950 525.600 523.050 526.050 ;
        RECT 514.950 524.400 523.050 525.600 ;
        RECT 545.400 525.600 546.600 527.400 ;
        RECT 547.950 527.400 562.050 528.600 ;
        RECT 547.950 526.950 550.050 527.400 ;
        RECT 559.950 526.950 562.050 527.400 ;
        RECT 610.950 528.600 613.050 529.050 ;
        RECT 631.950 528.600 634.050 529.050 ;
        RECT 610.950 527.400 634.050 528.600 ;
        RECT 610.950 526.950 613.050 527.400 ;
        RECT 614.400 526.050 615.600 527.400 ;
        RECT 631.950 526.950 634.050 527.400 ;
        RECT 637.950 528.600 640.050 529.050 ;
        RECT 652.950 528.600 655.050 529.050 ;
        RECT 637.950 527.400 655.050 528.600 ;
        RECT 637.950 526.950 640.050 527.400 ;
        RECT 652.950 526.950 655.050 527.400 ;
        RECT 715.950 526.950 718.050 529.050 ;
        RECT 754.950 528.600 757.050 529.050 ;
        RECT 760.950 528.600 763.050 529.050 ;
        RECT 754.950 527.400 763.050 528.600 ;
        RECT 754.950 526.950 757.050 527.400 ;
        RECT 760.950 526.950 763.050 527.400 ;
        RECT 766.950 526.950 769.050 529.050 ;
        RECT 808.950 528.600 811.050 529.050 ;
        RECT 829.950 528.600 832.050 529.050 ;
        RECT 808.950 527.400 832.050 528.600 ;
        RECT 808.950 526.950 811.050 527.400 ;
        RECT 829.950 526.950 832.050 527.400 ;
        RECT 556.950 525.600 559.050 526.050 ;
        RECT 574.950 525.600 577.050 526.050 ;
        RECT 592.950 525.600 595.050 526.050 ;
        RECT 545.400 524.400 595.050 525.600 ;
        RECT 427.950 523.950 430.050 524.400 ;
        RECT 514.950 523.950 517.050 524.400 ;
        RECT 520.950 523.950 523.050 524.400 ;
        RECT 556.950 523.950 559.050 524.400 ;
        RECT 574.950 523.950 577.050 524.400 ;
        RECT 592.950 523.950 595.050 524.400 ;
        RECT 613.950 523.950 616.050 526.050 ;
        RECT 619.950 525.600 622.050 526.050 ;
        RECT 634.950 525.600 637.050 526.050 ;
        RECT 619.950 524.400 637.050 525.600 ;
        RECT 619.950 523.950 622.050 524.400 ;
        RECT 634.950 523.950 637.050 524.400 ;
        RECT 661.950 525.600 664.050 526.050 ;
        RECT 676.950 525.600 679.050 526.050 ;
        RECT 661.950 524.400 679.050 525.600 ;
        RECT 661.950 523.950 664.050 524.400 ;
        RECT 676.950 523.950 679.050 524.400 ;
        RECT 763.950 525.600 766.050 526.050 ;
        RECT 767.400 525.600 768.600 526.950 ;
        RECT 763.950 524.400 768.600 525.600 ;
        RECT 802.950 525.600 805.050 526.050 ;
        RECT 820.950 525.600 823.050 526.050 ;
        RECT 802.950 524.400 823.050 525.600 ;
        RECT 763.950 523.950 766.050 524.400 ;
        RECT 802.950 523.950 805.050 524.400 ;
        RECT 820.950 523.950 823.050 524.400 ;
        RECT 826.950 525.600 829.050 526.050 ;
        RECT 853.950 525.600 856.050 526.050 ;
        RECT 880.950 525.600 883.050 526.050 ;
        RECT 826.950 524.400 883.050 525.600 ;
        RECT 826.950 523.950 829.050 524.400 ;
        RECT 853.950 523.950 856.050 524.400 ;
        RECT 880.950 523.950 883.050 524.400 ;
        RECT 115.950 522.600 118.050 523.050 ;
        RECT 121.950 522.600 124.050 523.050 ;
        RECT 115.950 521.400 124.050 522.600 ;
        RECT 115.950 520.950 118.050 521.400 ;
        RECT 121.950 520.950 124.050 521.400 ;
        RECT 130.950 520.950 133.050 523.050 ;
        RECT 265.950 522.600 268.050 523.050 ;
        RECT 313.950 522.600 316.050 523.050 ;
        RECT 265.950 521.400 316.050 522.600 ;
        RECT 265.950 520.950 268.050 521.400 ;
        RECT 313.950 520.950 316.050 521.400 ;
        RECT 340.950 522.600 343.050 523.050 ;
        RECT 352.950 522.600 355.050 523.050 ;
        RECT 340.950 521.400 355.050 522.600 ;
        RECT 340.950 520.950 343.050 521.400 ;
        RECT 352.950 520.950 355.050 521.400 ;
        RECT 379.950 522.600 382.050 523.050 ;
        RECT 442.950 522.600 445.050 523.050 ;
        RECT 454.950 522.600 457.050 523.050 ;
        RECT 379.950 521.400 457.050 522.600 ;
        RECT 379.950 520.950 382.050 521.400 ;
        RECT 442.950 520.950 445.050 521.400 ;
        RECT 454.950 520.950 457.050 521.400 ;
        RECT 508.950 522.600 511.050 523.050 ;
        RECT 547.950 522.600 550.050 523.050 ;
        RECT 508.950 521.400 550.050 522.600 ;
        RECT 508.950 520.950 511.050 521.400 ;
        RECT 547.950 520.950 550.050 521.400 ;
        RECT 571.950 522.600 574.050 523.050 ;
        RECT 589.950 522.600 592.050 523.050 ;
        RECT 571.950 521.400 592.050 522.600 ;
        RECT 571.950 520.950 574.050 521.400 ;
        RECT 589.950 520.950 592.050 521.400 ;
        RECT 622.950 522.600 625.050 523.050 ;
        RECT 637.950 522.600 640.050 523.050 ;
        RECT 622.950 521.400 640.050 522.600 ;
        RECT 622.950 520.950 625.050 521.400 ;
        RECT 637.950 520.950 640.050 521.400 ;
        RECT 667.950 522.600 670.050 523.050 ;
        RECT 673.950 522.600 676.050 523.050 ;
        RECT 667.950 521.400 676.050 522.600 ;
        RECT 667.950 520.950 670.050 521.400 ;
        RECT 673.950 520.950 676.050 521.400 ;
        RECT 679.950 522.600 682.050 523.050 ;
        RECT 685.950 522.600 688.050 523.050 ;
        RECT 679.950 521.400 688.050 522.600 ;
        RECT 679.950 520.950 682.050 521.400 ;
        RECT 685.950 520.950 688.050 521.400 ;
        RECT 730.950 522.600 733.050 523.050 ;
        RECT 751.950 522.600 754.050 523.050 ;
        RECT 754.950 522.600 757.050 523.050 ;
        RECT 730.950 521.400 757.050 522.600 ;
        RECT 730.950 520.950 733.050 521.400 ;
        RECT 751.950 520.950 754.050 521.400 ;
        RECT 754.950 520.950 757.050 521.400 ;
        RECT 868.950 522.600 871.050 523.050 ;
        RECT 874.950 522.600 877.050 523.050 ;
        RECT 868.950 521.400 877.050 522.600 ;
        RECT 868.950 520.950 871.050 521.400 ;
        RECT 874.950 520.950 877.050 521.400 ;
        RECT 112.950 519.600 115.050 520.050 ;
        RECT 145.950 519.600 148.050 520.050 ;
        RECT 112.950 518.400 148.050 519.600 ;
        RECT 112.950 517.950 115.050 518.400 ;
        RECT 145.950 517.950 148.050 518.400 ;
        RECT 319.950 519.600 322.050 520.050 ;
        RECT 343.950 519.600 346.050 520.050 ;
        RECT 346.950 519.600 349.050 520.050 ;
        RECT 319.950 518.400 349.050 519.600 ;
        RECT 319.950 517.950 322.050 518.400 ;
        RECT 343.950 517.950 346.050 518.400 ;
        RECT 346.950 517.950 349.050 518.400 ;
        RECT 523.950 519.600 526.050 520.050 ;
        RECT 535.950 519.600 538.050 520.050 ;
        RECT 523.950 518.400 538.050 519.600 ;
        RECT 523.950 517.950 526.050 518.400 ;
        RECT 535.950 517.950 538.050 518.400 ;
        RECT 571.950 519.600 574.050 520.050 ;
        RECT 583.950 519.600 586.050 520.050 ;
        RECT 571.950 518.400 586.050 519.600 ;
        RECT 571.950 517.950 574.050 518.400 ;
        RECT 583.950 517.950 586.050 518.400 ;
        RECT 679.950 519.600 682.050 520.050 ;
        RECT 745.950 519.600 748.050 520.050 ;
        RECT 763.950 519.600 766.050 520.050 ;
        RECT 679.950 518.400 766.050 519.600 ;
        RECT 679.950 517.950 682.050 518.400 ;
        RECT 745.950 517.950 748.050 518.400 ;
        RECT 763.950 517.950 766.050 518.400 ;
        RECT 796.950 519.600 799.050 520.050 ;
        RECT 802.950 519.600 805.050 520.050 ;
        RECT 796.950 518.400 805.050 519.600 ;
        RECT 796.950 517.950 799.050 518.400 ;
        RECT 802.950 517.950 805.050 518.400 ;
        RECT 52.950 516.600 55.050 517.050 ;
        RECT 67.950 516.600 70.050 517.050 ;
        RECT 70.950 516.600 73.050 517.050 ;
        RECT 52.950 515.400 73.050 516.600 ;
        RECT 52.950 514.950 55.050 515.400 ;
        RECT 67.950 514.950 70.050 515.400 ;
        RECT 70.950 514.950 73.050 515.400 ;
        RECT 184.950 516.600 187.050 517.050 ;
        RECT 205.950 516.600 208.050 517.050 ;
        RECT 481.950 516.600 484.050 517.050 ;
        RECT 184.950 515.400 484.050 516.600 ;
        RECT 184.950 514.950 187.050 515.400 ;
        RECT 205.950 514.950 208.050 515.400 ;
        RECT 481.950 514.950 484.050 515.400 ;
        RECT 643.950 516.600 646.050 517.050 ;
        RECT 661.950 516.600 664.050 517.050 ;
        RECT 643.950 515.400 664.050 516.600 ;
        RECT 643.950 514.950 646.050 515.400 ;
        RECT 661.950 514.950 664.050 515.400 ;
        RECT 286.950 513.600 289.050 514.050 ;
        RECT 334.950 513.600 337.050 514.050 ;
        RECT 286.950 512.400 337.050 513.600 ;
        RECT 286.950 511.950 289.050 512.400 ;
        RECT 334.950 511.950 337.050 512.400 ;
        RECT 487.950 510.600 490.050 511.050 ;
        RECT 496.950 510.600 499.050 511.050 ;
        RECT 487.950 509.400 499.050 510.600 ;
        RECT 487.950 508.950 490.050 509.400 ;
        RECT 496.950 508.950 499.050 509.400 ;
        RECT 799.950 510.600 802.050 511.050 ;
        RECT 805.950 510.600 808.050 511.050 ;
        RECT 799.950 509.400 808.050 510.600 ;
        RECT 799.950 508.950 802.050 509.400 ;
        RECT 805.950 508.950 808.050 509.400 ;
        RECT 841.950 510.600 844.050 511.050 ;
        RECT 859.950 510.600 862.050 511.050 ;
        RECT 841.950 509.400 862.050 510.600 ;
        RECT 841.950 508.950 844.050 509.400 ;
        RECT 859.950 508.950 862.050 509.400 ;
        RECT 322.950 507.600 325.050 508.050 ;
        RECT 334.950 507.600 337.050 508.050 ;
        RECT 322.950 506.400 337.050 507.600 ;
        RECT 322.950 505.950 325.050 506.400 ;
        RECT 334.950 505.950 337.050 506.400 ;
        RECT 712.950 507.600 715.050 508.050 ;
        RECT 781.950 507.600 784.050 508.050 ;
        RECT 712.950 506.400 784.050 507.600 ;
        RECT 712.950 505.950 715.050 506.400 ;
        RECT 781.950 505.950 784.050 506.400 ;
        RECT 787.950 507.600 790.050 508.050 ;
        RECT 793.950 507.600 796.050 508.050 ;
        RECT 823.950 507.600 826.050 508.050 ;
        RECT 787.950 506.400 826.050 507.600 ;
        RECT 787.950 505.950 790.050 506.400 ;
        RECT 793.950 505.950 796.050 506.400 ;
        RECT 823.950 505.950 826.050 506.400 ;
        RECT 358.950 504.600 361.050 505.050 ;
        RECT 391.950 504.600 394.050 505.050 ;
        RECT 358.950 503.400 394.050 504.600 ;
        RECT 358.950 502.950 361.050 503.400 ;
        RECT 391.950 502.950 394.050 503.400 ;
        RECT 178.950 501.600 181.050 502.050 ;
        RECT 187.950 501.600 190.050 502.050 ;
        RECT 202.950 501.600 205.050 502.050 ;
        RECT 226.950 501.600 229.050 502.050 ;
        RECT 253.950 501.600 256.050 502.050 ;
        RECT 178.950 500.400 256.050 501.600 ;
        RECT 178.950 499.950 181.050 500.400 ;
        RECT 187.950 499.950 190.050 500.400 ;
        RECT 202.950 499.950 205.050 500.400 ;
        RECT 226.950 499.950 229.050 500.400 ;
        RECT 253.950 499.950 256.050 500.400 ;
        RECT 586.950 501.600 589.050 502.050 ;
        RECT 625.950 501.600 628.050 502.050 ;
        RECT 586.950 500.400 628.050 501.600 ;
        RECT 586.950 499.950 589.050 500.400 ;
        RECT 625.950 499.950 628.050 500.400 ;
        RECT 49.950 498.600 52.050 499.050 ;
        RECT 670.950 498.600 673.050 499.050 ;
        RECT 49.950 497.400 673.050 498.600 ;
        RECT 49.950 496.950 52.050 497.400 ;
        RECT 670.950 496.950 673.050 497.400 ;
        RECT 724.950 498.600 727.050 499.050 ;
        RECT 796.950 498.600 799.050 499.050 ;
        RECT 724.950 497.400 799.050 498.600 ;
        RECT 724.950 496.950 727.050 497.400 ;
        RECT 796.950 496.950 799.050 497.400 ;
        RECT 37.950 495.600 40.050 496.050 ;
        RECT 142.950 495.600 145.050 496.050 ;
        RECT 145.950 495.600 148.050 496.050 ;
        RECT 37.950 494.400 148.050 495.600 ;
        RECT 37.950 493.950 40.050 494.400 ;
        RECT 142.950 493.950 145.050 494.400 ;
        RECT 145.950 493.950 148.050 494.400 ;
        RECT 403.950 495.600 406.050 496.050 ;
        RECT 517.950 495.600 520.050 496.050 ;
        RECT 553.950 495.600 556.050 496.050 ;
        RECT 403.950 494.400 556.050 495.600 ;
        RECT 403.950 493.950 406.050 494.400 ;
        RECT 517.950 493.950 520.050 494.400 ;
        RECT 553.950 493.950 556.050 494.400 ;
        RECT 751.950 495.600 754.050 496.050 ;
        RECT 781.950 495.600 784.050 496.050 ;
        RECT 787.950 495.600 790.050 496.050 ;
        RECT 751.950 494.400 790.050 495.600 ;
        RECT 751.950 493.950 754.050 494.400 ;
        RECT 781.950 493.950 784.050 494.400 ;
        RECT 787.950 493.950 790.050 494.400 ;
        RECT 85.950 492.600 88.050 493.050 ;
        RECT 103.950 492.600 106.050 493.050 ;
        RECT 85.950 491.400 106.050 492.600 ;
        RECT 85.950 490.950 88.050 491.400 ;
        RECT 103.950 490.950 106.050 491.400 ;
        RECT 280.950 492.600 283.050 493.050 ;
        RECT 286.950 492.600 289.050 493.050 ;
        RECT 289.950 492.600 292.050 493.050 ;
        RECT 280.950 491.400 292.050 492.600 ;
        RECT 280.950 490.950 283.050 491.400 ;
        RECT 286.950 490.950 289.050 491.400 ;
        RECT 289.950 490.950 292.050 491.400 ;
        RECT 298.950 492.600 301.050 493.050 ;
        RECT 316.950 492.600 319.050 493.050 ;
        RECT 319.950 492.600 322.050 493.050 ;
        RECT 322.950 492.600 325.050 493.050 ;
        RECT 298.950 491.400 325.050 492.600 ;
        RECT 298.950 490.950 301.050 491.400 ;
        RECT 316.950 490.950 319.050 491.400 ;
        RECT 319.950 490.950 322.050 491.400 ;
        RECT 322.950 490.950 325.050 491.400 ;
        RECT 379.950 492.600 382.050 493.050 ;
        RECT 397.950 492.600 400.050 493.050 ;
        RECT 379.950 491.400 400.050 492.600 ;
        RECT 379.950 490.950 382.050 491.400 ;
        RECT 397.950 490.950 400.050 491.400 ;
        RECT 409.950 492.600 412.050 493.050 ;
        RECT 436.950 492.600 439.050 493.050 ;
        RECT 721.950 492.600 724.050 493.050 ;
        RECT 409.950 491.400 724.050 492.600 ;
        RECT 409.950 490.950 412.050 491.400 ;
        RECT 436.950 490.950 439.050 491.400 ;
        RECT 721.950 490.950 724.050 491.400 ;
        RECT 727.950 492.600 730.050 493.050 ;
        RECT 766.950 492.600 769.050 493.050 ;
        RECT 727.950 491.400 769.050 492.600 ;
        RECT 727.950 490.950 730.050 491.400 ;
        RECT 766.950 490.950 769.050 491.400 ;
        RECT 34.950 489.600 37.050 490.050 ;
        RECT 73.950 489.600 76.050 490.050 ;
        RECT 88.950 489.600 91.050 490.050 ;
        RECT 121.950 489.600 124.050 490.050 ;
        RECT 133.950 489.600 136.050 490.050 ;
        RECT 34.950 488.400 76.050 489.600 ;
        RECT 34.950 487.950 37.050 488.400 ;
        RECT 73.950 487.950 76.050 488.400 ;
        RECT 86.400 488.400 136.050 489.600 ;
        RECT 61.950 486.600 64.050 487.050 ;
        RECT 67.950 486.600 70.050 487.050 ;
        RECT 86.400 486.600 87.600 488.400 ;
        RECT 88.950 487.950 91.050 488.400 ;
        RECT 121.950 487.950 124.050 488.400 ;
        RECT 133.950 487.950 136.050 488.400 ;
        RECT 304.950 489.600 307.050 490.050 ;
        RECT 313.950 489.600 316.050 490.050 ;
        RECT 304.950 488.400 316.050 489.600 ;
        RECT 304.950 487.950 307.050 488.400 ;
        RECT 313.950 487.950 316.050 488.400 ;
        RECT 334.950 489.600 337.050 490.050 ;
        RECT 349.950 489.600 352.050 490.050 ;
        RECT 355.950 489.600 358.050 490.050 ;
        RECT 334.950 488.400 352.050 489.600 ;
        RECT 334.950 487.950 337.050 488.400 ;
        RECT 349.950 487.950 352.050 488.400 ;
        RECT 353.400 488.400 358.050 489.600 ;
        RECT 353.400 487.050 354.600 488.400 ;
        RECT 355.950 487.950 358.050 488.400 ;
        RECT 373.950 489.600 376.050 490.050 ;
        RECT 388.950 489.600 391.050 490.050 ;
        RECT 373.950 488.400 391.050 489.600 ;
        RECT 373.950 487.950 376.050 488.400 ;
        RECT 388.950 487.950 391.050 488.400 ;
        RECT 421.950 489.600 424.050 490.050 ;
        RECT 508.950 489.600 511.050 490.050 ;
        RECT 421.950 488.400 511.050 489.600 ;
        RECT 421.950 487.950 424.050 488.400 ;
        RECT 508.950 487.950 511.050 488.400 ;
        RECT 514.950 487.950 517.050 490.050 ;
        RECT 532.950 489.600 535.050 490.050 ;
        RECT 541.950 489.600 544.050 490.050 ;
        RECT 532.950 488.400 544.050 489.600 ;
        RECT 532.950 487.950 535.050 488.400 ;
        RECT 541.950 487.950 544.050 488.400 ;
        RECT 577.950 489.600 580.050 490.050 ;
        RECT 622.950 489.600 625.050 490.050 ;
        RECT 577.950 488.400 625.050 489.600 ;
        RECT 577.950 487.950 580.050 488.400 ;
        RECT 622.950 487.950 625.050 488.400 ;
        RECT 760.950 489.600 763.050 490.050 ;
        RECT 769.950 489.600 772.050 490.050 ;
        RECT 760.950 488.400 772.050 489.600 ;
        RECT 760.950 487.950 763.050 488.400 ;
        RECT 769.950 487.950 772.050 488.400 ;
        RECT 838.950 489.600 841.050 490.050 ;
        RECT 868.950 489.600 871.050 490.050 ;
        RECT 838.950 488.400 871.050 489.600 ;
        RECT 838.950 487.950 841.050 488.400 ;
        RECT 868.950 487.950 871.050 488.400 ;
        RECT 61.950 485.400 70.050 486.600 ;
        RECT 61.950 484.950 64.050 485.400 ;
        RECT 67.950 484.950 70.050 485.400 ;
        RECT 74.400 485.400 87.600 486.600 ;
        RECT 88.950 486.600 91.050 487.050 ;
        RECT 91.950 486.600 94.050 487.050 ;
        RECT 94.950 486.600 97.050 487.050 ;
        RECT 88.950 485.400 97.050 486.600 ;
        RECT 70.950 483.600 73.050 484.050 ;
        RECT 74.400 483.600 75.600 485.400 ;
        RECT 88.950 484.950 91.050 485.400 ;
        RECT 91.950 484.950 94.050 485.400 ;
        RECT 94.950 484.950 97.050 485.400 ;
        RECT 148.950 486.600 151.050 487.050 ;
        RECT 163.950 486.600 166.050 487.050 ;
        RECT 148.950 485.400 166.050 486.600 ;
        RECT 148.950 484.950 151.050 485.400 ;
        RECT 163.950 484.950 166.050 485.400 ;
        RECT 184.950 486.600 187.050 487.050 ;
        RECT 217.950 486.600 220.050 487.050 ;
        RECT 184.950 485.400 220.050 486.600 ;
        RECT 184.950 484.950 187.050 485.400 ;
        RECT 217.950 484.950 220.050 485.400 ;
        RECT 223.950 486.600 226.050 487.050 ;
        RECT 259.950 486.600 262.050 487.050 ;
        RECT 223.950 485.400 262.050 486.600 ;
        RECT 223.950 484.950 226.050 485.400 ;
        RECT 259.950 484.950 262.050 485.400 ;
        RECT 286.950 486.600 289.050 487.050 ;
        RECT 301.950 486.600 304.050 487.050 ;
        RECT 286.950 485.400 304.050 486.600 ;
        RECT 286.950 484.950 289.050 485.400 ;
        RECT 301.950 484.950 304.050 485.400 ;
        RECT 352.950 484.950 355.050 487.050 ;
        RECT 376.950 486.600 379.050 487.050 ;
        RECT 403.950 486.600 406.050 487.050 ;
        RECT 376.950 485.400 406.050 486.600 ;
        RECT 376.950 484.950 379.050 485.400 ;
        RECT 403.950 484.950 406.050 485.400 ;
        RECT 412.950 486.600 415.050 487.050 ;
        RECT 430.950 486.600 433.050 487.050 ;
        RECT 412.950 485.400 433.050 486.600 ;
        RECT 412.950 484.950 415.050 485.400 ;
        RECT 430.950 484.950 433.050 485.400 ;
        RECT 475.950 486.600 478.050 487.050 ;
        RECT 490.950 486.600 493.050 487.050 ;
        RECT 475.950 485.400 493.050 486.600 ;
        RECT 475.950 484.950 478.050 485.400 ;
        RECT 490.950 484.950 493.050 485.400 ;
        RECT 496.950 486.600 499.050 487.050 ;
        RECT 502.950 486.600 505.050 487.050 ;
        RECT 496.950 485.400 505.050 486.600 ;
        RECT 515.400 486.600 516.600 487.950 ;
        RECT 538.950 486.600 541.050 487.050 ;
        RECT 515.400 485.400 541.050 486.600 ;
        RECT 496.950 484.950 499.050 485.400 ;
        RECT 502.950 484.950 505.050 485.400 ;
        RECT 538.950 484.950 541.050 485.400 ;
        RECT 562.950 486.600 565.050 487.050 ;
        RECT 604.950 486.600 607.050 487.050 ;
        RECT 562.950 485.400 607.050 486.600 ;
        RECT 562.950 484.950 565.050 485.400 ;
        RECT 604.950 484.950 607.050 485.400 ;
        RECT 613.950 486.600 616.050 487.050 ;
        RECT 631.950 486.600 634.050 487.050 ;
        RECT 613.950 485.400 634.050 486.600 ;
        RECT 613.950 484.950 616.050 485.400 ;
        RECT 631.950 484.950 634.050 485.400 ;
        RECT 658.950 486.600 661.050 487.050 ;
        RECT 670.950 486.600 673.050 487.050 ;
        RECT 658.950 485.400 673.050 486.600 ;
        RECT 658.950 484.950 661.050 485.400 ;
        RECT 670.950 484.950 673.050 485.400 ;
        RECT 676.950 486.600 679.050 487.050 ;
        RECT 688.950 486.600 691.050 487.050 ;
        RECT 703.950 486.600 706.050 487.050 ;
        RECT 727.950 486.600 730.050 487.050 ;
        RECT 676.950 485.400 702.600 486.600 ;
        RECT 676.950 484.950 679.050 485.400 ;
        RECT 688.950 484.950 691.050 485.400 ;
        RECT 701.400 484.050 702.600 485.400 ;
        RECT 703.950 485.400 730.050 486.600 ;
        RECT 703.950 484.950 706.050 485.400 ;
        RECT 727.950 484.950 730.050 485.400 ;
        RECT 793.950 486.600 796.050 487.050 ;
        RECT 829.950 486.600 832.050 487.050 ;
        RECT 841.950 486.600 844.050 487.050 ;
        RECT 793.950 485.400 844.050 486.600 ;
        RECT 793.950 484.950 796.050 485.400 ;
        RECT 829.950 484.950 832.050 485.400 ;
        RECT 841.950 484.950 844.050 485.400 ;
        RECT 847.950 486.600 850.050 487.050 ;
        RECT 859.950 486.600 862.050 487.050 ;
        RECT 847.950 485.400 862.050 486.600 ;
        RECT 847.950 484.950 850.050 485.400 ;
        RECT 859.950 484.950 862.050 485.400 ;
        RECT 70.950 482.400 75.600 483.600 ;
        RECT 76.950 483.600 79.050 484.050 ;
        RECT 100.950 483.600 103.050 484.050 ;
        RECT 109.950 483.600 112.050 484.050 ;
        RECT 76.950 482.400 112.050 483.600 ;
        RECT 70.950 481.950 73.050 482.400 ;
        RECT 76.950 481.950 79.050 482.400 ;
        RECT 100.950 481.950 103.050 482.400 ;
        RECT 109.950 481.950 112.050 482.400 ;
        RECT 124.950 483.600 127.050 484.050 ;
        RECT 130.950 483.600 133.050 484.050 ;
        RECT 124.950 482.400 133.050 483.600 ;
        RECT 124.950 481.950 127.050 482.400 ;
        RECT 130.950 481.950 133.050 482.400 ;
        RECT 268.950 483.600 271.050 484.050 ;
        RECT 277.950 483.600 280.050 484.050 ;
        RECT 295.950 483.600 298.050 484.050 ;
        RECT 268.950 482.400 298.050 483.600 ;
        RECT 268.950 481.950 271.050 482.400 ;
        RECT 277.950 481.950 280.050 482.400 ;
        RECT 295.950 481.950 298.050 482.400 ;
        RECT 382.950 483.600 385.050 484.050 ;
        RECT 391.950 483.600 394.050 484.050 ;
        RECT 382.950 482.400 394.050 483.600 ;
        RECT 382.950 481.950 385.050 482.400 ;
        RECT 391.950 481.950 394.050 482.400 ;
        RECT 400.950 483.600 403.050 484.050 ;
        RECT 412.950 483.600 415.050 484.050 ;
        RECT 400.950 482.400 415.050 483.600 ;
        RECT 400.950 481.950 403.050 482.400 ;
        RECT 412.950 481.950 415.050 482.400 ;
        RECT 427.950 483.600 430.050 484.050 ;
        RECT 433.950 483.600 436.050 484.050 ;
        RECT 427.950 482.400 436.050 483.600 ;
        RECT 427.950 481.950 430.050 482.400 ;
        RECT 433.950 481.950 436.050 482.400 ;
        RECT 439.950 483.600 442.050 484.050 ;
        RECT 448.950 483.600 451.050 484.050 ;
        RECT 439.950 482.400 451.050 483.600 ;
        RECT 439.950 481.950 442.050 482.400 ;
        RECT 448.950 481.950 451.050 482.400 ;
        RECT 460.950 483.600 463.050 484.050 ;
        RECT 466.950 483.600 469.050 484.050 ;
        RECT 460.950 482.400 469.050 483.600 ;
        RECT 460.950 481.950 463.050 482.400 ;
        RECT 466.950 481.950 469.050 482.400 ;
        RECT 487.950 483.600 490.050 484.050 ;
        RECT 493.950 483.600 496.050 484.050 ;
        RECT 487.950 482.400 496.050 483.600 ;
        RECT 487.950 481.950 490.050 482.400 ;
        RECT 493.950 481.950 496.050 482.400 ;
        RECT 514.950 483.600 517.050 484.050 ;
        RECT 523.950 483.600 526.050 484.050 ;
        RECT 514.950 482.400 526.050 483.600 ;
        RECT 514.950 481.950 517.050 482.400 ;
        RECT 523.950 481.950 526.050 482.400 ;
        RECT 535.950 483.600 538.050 484.050 ;
        RECT 544.950 483.600 547.050 484.050 ;
        RECT 535.950 482.400 547.050 483.600 ;
        RECT 535.950 481.950 538.050 482.400 ;
        RECT 544.950 481.950 547.050 482.400 ;
        RECT 547.950 483.600 550.050 484.050 ;
        RECT 556.950 483.600 559.050 484.050 ;
        RECT 547.950 482.400 559.050 483.600 ;
        RECT 547.950 481.950 550.050 482.400 ;
        RECT 556.950 481.950 559.050 482.400 ;
        RECT 559.950 483.600 562.050 484.050 ;
        RECT 571.950 483.600 574.050 484.050 ;
        RECT 559.950 482.400 574.050 483.600 ;
        RECT 559.950 481.950 562.050 482.400 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 601.950 483.600 604.050 484.050 ;
        RECT 622.950 483.600 625.050 484.050 ;
        RECT 601.950 482.400 625.050 483.600 ;
        RECT 601.950 481.950 604.050 482.400 ;
        RECT 622.950 481.950 625.050 482.400 ;
        RECT 640.950 483.600 643.050 484.050 ;
        RECT 667.950 483.600 670.050 484.050 ;
        RECT 640.950 482.400 670.050 483.600 ;
        RECT 640.950 481.950 643.050 482.400 ;
        RECT 667.950 481.950 670.050 482.400 ;
        RECT 700.950 481.950 703.050 484.050 ;
        RECT 709.950 483.600 712.050 484.050 ;
        RECT 748.950 483.600 751.050 484.050 ;
        RECT 709.950 482.400 751.050 483.600 ;
        RECT 709.950 481.950 712.050 482.400 ;
        RECT 748.950 481.950 751.050 482.400 ;
        RECT 772.950 483.600 775.050 484.050 ;
        RECT 790.950 483.600 793.050 484.050 ;
        RECT 772.950 482.400 793.050 483.600 ;
        RECT 772.950 481.950 775.050 482.400 ;
        RECT 790.950 481.950 793.050 482.400 ;
        RECT 835.950 483.600 838.050 484.050 ;
        RECT 865.950 483.600 868.050 484.050 ;
        RECT 835.950 482.400 868.050 483.600 ;
        RECT 835.950 481.950 838.050 482.400 ;
        RECT 865.950 481.950 868.050 482.400 ;
        RECT 64.950 480.600 67.050 481.050 ;
        RECT 100.950 480.600 103.050 481.050 ;
        RECT 64.950 479.400 103.050 480.600 ;
        RECT 64.950 478.950 67.050 479.400 ;
        RECT 100.950 478.950 103.050 479.400 ;
        RECT 106.950 480.600 109.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 106.950 479.400 121.050 480.600 ;
        RECT 106.950 478.950 109.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 163.950 480.600 166.050 481.050 ;
        RECT 190.950 480.600 193.050 481.050 ;
        RECT 163.950 479.400 193.050 480.600 ;
        RECT 163.950 478.950 166.050 479.400 ;
        RECT 190.950 478.950 193.050 479.400 ;
        RECT 262.950 480.600 265.050 481.050 ;
        RECT 271.950 480.600 274.050 481.050 ;
        RECT 262.950 479.400 274.050 480.600 ;
        RECT 262.950 478.950 265.050 479.400 ;
        RECT 271.950 478.950 274.050 479.400 ;
        RECT 361.950 480.600 364.050 481.050 ;
        RECT 400.950 480.600 403.050 481.050 ;
        RECT 361.950 479.400 403.050 480.600 ;
        RECT 361.950 478.950 364.050 479.400 ;
        RECT 400.950 478.950 403.050 479.400 ;
        RECT 406.950 480.600 409.050 481.050 ;
        RECT 433.950 480.600 436.050 481.050 ;
        RECT 406.950 479.400 436.050 480.600 ;
        RECT 406.950 478.950 409.050 479.400 ;
        RECT 433.950 478.950 436.050 479.400 ;
        RECT 454.950 480.600 457.050 481.050 ;
        RECT 463.950 480.600 466.050 481.050 ;
        RECT 454.950 479.400 466.050 480.600 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 463.950 478.950 466.050 479.400 ;
        RECT 472.950 480.600 475.050 481.050 ;
        RECT 493.950 480.600 496.050 481.050 ;
        RECT 472.950 479.400 496.050 480.600 ;
        RECT 472.950 478.950 475.050 479.400 ;
        RECT 493.950 478.950 496.050 479.400 ;
        RECT 499.950 480.600 502.050 481.050 ;
        RECT 514.950 480.600 517.050 481.050 ;
        RECT 520.950 480.600 523.050 481.050 ;
        RECT 499.950 479.400 523.050 480.600 ;
        RECT 499.950 478.950 502.050 479.400 ;
        RECT 514.950 478.950 517.050 479.400 ;
        RECT 520.950 478.950 523.050 479.400 ;
        RECT 577.950 480.600 580.050 481.050 ;
        RECT 583.950 480.600 586.050 481.050 ;
        RECT 610.950 480.600 613.050 481.050 ;
        RECT 577.950 479.400 613.050 480.600 ;
        RECT 577.950 478.950 580.050 479.400 ;
        RECT 583.950 478.950 586.050 479.400 ;
        RECT 610.950 478.950 613.050 479.400 ;
        RECT 634.950 480.600 637.050 481.050 ;
        RECT 664.950 480.600 667.050 481.050 ;
        RECT 634.950 479.400 667.050 480.600 ;
        RECT 634.950 478.950 637.050 479.400 ;
        RECT 664.950 478.950 667.050 479.400 ;
        RECT 697.950 480.600 700.050 481.050 ;
        RECT 706.950 480.600 709.050 481.050 ;
        RECT 697.950 479.400 709.050 480.600 ;
        RECT 697.950 478.950 700.050 479.400 ;
        RECT 706.950 478.950 709.050 479.400 ;
        RECT 754.950 480.600 757.050 481.050 ;
        RECT 769.950 480.600 772.050 481.050 ;
        RECT 811.950 480.600 814.050 481.050 ;
        RECT 754.950 479.400 768.600 480.600 ;
        RECT 754.950 478.950 757.050 479.400 ;
        RECT 91.950 477.600 94.050 478.050 ;
        RECT 115.950 477.600 118.050 478.050 ;
        RECT 121.950 477.600 124.050 478.050 ;
        RECT 91.950 476.400 124.050 477.600 ;
        RECT 91.950 475.950 94.050 476.400 ;
        RECT 115.950 475.950 118.050 476.400 ;
        RECT 121.950 475.950 124.050 476.400 ;
        RECT 151.950 477.600 154.050 478.050 ;
        RECT 154.950 477.600 157.050 478.050 ;
        RECT 172.950 477.600 175.050 478.050 ;
        RECT 184.950 477.600 187.050 478.050 ;
        RECT 151.950 476.400 187.050 477.600 ;
        RECT 151.950 475.950 154.050 476.400 ;
        RECT 154.950 475.950 157.050 476.400 ;
        RECT 172.950 475.950 175.050 476.400 ;
        RECT 184.950 475.950 187.050 476.400 ;
        RECT 196.950 477.600 199.050 478.050 ;
        RECT 214.950 477.600 217.050 478.050 ;
        RECT 196.950 476.400 217.050 477.600 ;
        RECT 196.950 475.950 199.050 476.400 ;
        RECT 214.950 475.950 217.050 476.400 ;
        RECT 370.950 477.600 373.050 478.050 ;
        RECT 445.950 477.600 448.050 478.050 ;
        RECT 370.950 476.400 448.050 477.600 ;
        RECT 370.950 475.950 373.050 476.400 ;
        RECT 445.950 475.950 448.050 476.400 ;
        RECT 463.950 477.600 466.050 478.050 ;
        RECT 526.950 477.600 529.050 478.050 ;
        RECT 463.950 476.400 529.050 477.600 ;
        RECT 463.950 475.950 466.050 476.400 ;
        RECT 526.950 475.950 529.050 476.400 ;
        RECT 598.950 477.600 601.050 478.050 ;
        RECT 658.950 477.600 661.050 478.050 ;
        RECT 598.950 476.400 661.050 477.600 ;
        RECT 598.950 475.950 601.050 476.400 ;
        RECT 658.950 475.950 661.050 476.400 ;
        RECT 664.950 477.600 667.050 478.050 ;
        RECT 682.950 477.600 685.050 478.050 ;
        RECT 664.950 476.400 685.050 477.600 ;
        RECT 767.400 477.600 768.600 479.400 ;
        RECT 769.950 479.400 814.050 480.600 ;
        RECT 769.950 478.950 772.050 479.400 ;
        RECT 811.950 478.950 814.050 479.400 ;
        RECT 823.950 480.600 826.050 481.050 ;
        RECT 847.950 480.600 850.050 481.050 ;
        RECT 823.950 479.400 850.050 480.600 ;
        RECT 823.950 478.950 826.050 479.400 ;
        RECT 847.950 478.950 850.050 479.400 ;
        RECT 865.950 480.600 868.050 481.050 ;
        RECT 874.950 480.600 877.050 481.050 ;
        RECT 865.950 479.400 877.050 480.600 ;
        RECT 865.950 478.950 868.050 479.400 ;
        RECT 874.950 478.950 877.050 479.400 ;
        RECT 784.950 477.600 787.050 478.050 ;
        RECT 767.400 476.400 787.050 477.600 ;
        RECT 664.950 475.950 667.050 476.400 ;
        RECT 682.950 475.950 685.050 476.400 ;
        RECT 784.950 475.950 787.050 476.400 ;
        RECT 832.950 477.600 835.050 478.050 ;
        RECT 853.950 477.600 856.050 478.050 ;
        RECT 832.950 476.400 856.050 477.600 ;
        RECT 832.950 475.950 835.050 476.400 ;
        RECT 853.950 475.950 856.050 476.400 ;
        RECT 16.950 474.600 19.050 475.050 ;
        RECT 34.950 474.600 37.050 475.050 ;
        RECT 16.950 473.400 37.050 474.600 ;
        RECT 16.950 472.950 19.050 473.400 ;
        RECT 34.950 472.950 37.050 473.400 ;
        RECT 43.950 474.600 46.050 475.050 ;
        RECT 58.950 474.600 61.050 475.050 ;
        RECT 43.950 473.400 61.050 474.600 ;
        RECT 43.950 472.950 46.050 473.400 ;
        RECT 58.950 472.950 61.050 473.400 ;
        RECT 91.950 474.600 94.050 475.050 ;
        RECT 112.950 474.600 115.050 475.050 ;
        RECT 91.950 473.400 115.050 474.600 ;
        RECT 91.950 472.950 94.050 473.400 ;
        RECT 112.950 472.950 115.050 473.400 ;
        RECT 508.950 474.600 511.050 475.050 ;
        RECT 523.950 474.600 526.050 475.050 ;
        RECT 508.950 473.400 526.050 474.600 ;
        RECT 508.950 472.950 511.050 473.400 ;
        RECT 523.950 472.950 526.050 473.400 ;
        RECT 580.950 474.600 583.050 475.050 ;
        RECT 655.950 474.600 658.050 475.050 ;
        RECT 580.950 473.400 658.050 474.600 ;
        RECT 580.950 472.950 583.050 473.400 ;
        RECT 655.950 472.950 658.050 473.400 ;
        RECT 769.950 474.600 772.050 475.050 ;
        RECT 802.950 474.600 805.050 475.050 ;
        RECT 769.950 473.400 805.050 474.600 ;
        RECT 769.950 472.950 772.050 473.400 ;
        RECT 802.950 472.950 805.050 473.400 ;
        RECT 10.950 471.600 13.050 472.050 ;
        RECT 31.950 471.600 34.050 472.050 ;
        RECT 10.950 470.400 34.050 471.600 ;
        RECT 10.950 469.950 13.050 470.400 ;
        RECT 31.950 469.950 34.050 470.400 ;
        RECT 43.950 471.600 46.050 472.050 ;
        RECT 127.950 471.600 130.050 472.050 ;
        RECT 43.950 470.400 130.050 471.600 ;
        RECT 43.950 469.950 46.050 470.400 ;
        RECT 127.950 469.950 130.050 470.400 ;
        RECT 355.950 471.600 358.050 472.050 ;
        RECT 364.950 471.600 367.050 472.050 ;
        RECT 355.950 470.400 367.050 471.600 ;
        RECT 355.950 469.950 358.050 470.400 ;
        RECT 364.950 469.950 367.050 470.400 ;
        RECT 418.950 471.600 421.050 472.050 ;
        RECT 502.950 471.600 505.050 472.050 ;
        RECT 418.950 470.400 505.050 471.600 ;
        RECT 418.950 469.950 421.050 470.400 ;
        RECT 502.950 469.950 505.050 470.400 ;
        RECT 19.950 468.600 22.050 469.050 ;
        RECT 37.950 468.600 40.050 469.050 ;
        RECT 46.950 468.600 49.050 469.050 ;
        RECT 19.950 467.400 49.050 468.600 ;
        RECT 19.950 466.950 22.050 467.400 ;
        RECT 37.950 466.950 40.050 467.400 ;
        RECT 46.950 466.950 49.050 467.400 ;
        RECT 358.950 468.600 361.050 469.050 ;
        RECT 364.950 468.600 367.050 469.050 ;
        RECT 358.950 467.400 367.050 468.600 ;
        RECT 358.950 466.950 361.050 467.400 ;
        RECT 364.950 466.950 367.050 467.400 ;
        RECT 490.950 468.600 493.050 469.050 ;
        RECT 547.950 468.600 550.050 469.050 ;
        RECT 490.950 467.400 550.050 468.600 ;
        RECT 490.950 466.950 493.050 467.400 ;
        RECT 547.950 466.950 550.050 467.400 ;
        RECT 595.950 468.600 598.050 469.050 ;
        RECT 673.950 468.600 676.050 469.050 ;
        RECT 745.950 468.600 748.050 469.050 ;
        RECT 595.950 467.400 748.050 468.600 ;
        RECT 595.950 466.950 598.050 467.400 ;
        RECT 673.950 466.950 676.050 467.400 ;
        RECT 745.950 466.950 748.050 467.400 ;
        RECT 781.950 468.600 784.050 469.050 ;
        RECT 805.950 468.600 808.050 469.050 ;
        RECT 817.950 468.600 820.050 469.050 ;
        RECT 781.950 467.400 820.050 468.600 ;
        RECT 781.950 466.950 784.050 467.400 ;
        RECT 805.950 466.950 808.050 467.400 ;
        RECT 817.950 466.950 820.050 467.400 ;
        RECT 835.950 468.600 838.050 469.050 ;
        RECT 841.950 468.600 844.050 469.050 ;
        RECT 835.950 467.400 844.050 468.600 ;
        RECT 835.950 466.950 838.050 467.400 ;
        RECT 841.950 466.950 844.050 467.400 ;
        RECT 82.950 465.600 85.050 466.050 ;
        RECT 103.950 465.600 106.050 466.050 ;
        RECT 82.950 464.400 106.050 465.600 ;
        RECT 82.950 463.950 85.050 464.400 ;
        RECT 103.950 463.950 106.050 464.400 ;
        RECT 481.950 465.600 484.050 466.050 ;
        RECT 595.950 465.600 598.050 466.050 ;
        RECT 481.950 464.400 598.050 465.600 ;
        RECT 481.950 463.950 484.050 464.400 ;
        RECT 595.950 463.950 598.050 464.400 ;
        RECT 613.950 465.600 616.050 466.050 ;
        RECT 700.950 465.600 703.050 466.050 ;
        RECT 613.950 464.400 703.050 465.600 ;
        RECT 613.950 463.950 616.050 464.400 ;
        RECT 700.950 463.950 703.050 464.400 ;
        RECT 721.950 465.600 724.050 466.050 ;
        RECT 832.950 465.600 835.050 466.050 ;
        RECT 721.950 464.400 835.050 465.600 ;
        RECT 721.950 463.950 724.050 464.400 ;
        RECT 832.950 463.950 835.050 464.400 ;
        RECT 7.950 462.600 10.050 463.050 ;
        RECT 13.950 462.600 16.050 463.050 ;
        RECT 7.950 461.400 16.050 462.600 ;
        RECT 7.950 460.950 10.050 461.400 ;
        RECT 13.950 460.950 16.050 461.400 ;
        RECT 31.950 462.600 34.050 463.050 ;
        RECT 61.950 462.600 64.050 463.050 ;
        RECT 31.950 461.400 64.050 462.600 ;
        RECT 31.950 460.950 34.050 461.400 ;
        RECT 61.950 460.950 64.050 461.400 ;
        RECT 166.950 462.600 169.050 463.050 ;
        RECT 202.950 462.600 205.050 463.050 ;
        RECT 166.950 461.400 205.050 462.600 ;
        RECT 166.950 460.950 169.050 461.400 ;
        RECT 202.950 460.950 205.050 461.400 ;
        RECT 262.950 462.600 265.050 463.050 ;
        RECT 313.950 462.600 316.050 463.050 ;
        RECT 262.950 461.400 316.050 462.600 ;
        RECT 262.950 460.950 265.050 461.400 ;
        RECT 313.950 460.950 316.050 461.400 ;
        RECT 337.950 462.600 340.050 463.050 ;
        RECT 349.950 462.600 352.050 463.050 ;
        RECT 337.950 461.400 352.050 462.600 ;
        RECT 337.950 460.950 340.050 461.400 ;
        RECT 349.950 460.950 352.050 461.400 ;
        RECT 484.950 462.600 487.050 463.050 ;
        RECT 502.950 462.600 505.050 463.050 ;
        RECT 568.950 462.600 571.050 463.050 ;
        RECT 619.950 462.600 622.050 463.050 ;
        RECT 673.950 462.600 676.050 463.050 ;
        RECT 484.950 461.400 501.600 462.600 ;
        RECT 484.950 460.950 487.050 461.400 ;
        RECT 13.950 459.600 16.050 460.050 ;
        RECT 22.950 459.600 25.050 460.050 ;
        RECT 13.950 458.400 25.050 459.600 ;
        RECT 13.950 457.950 16.050 458.400 ;
        RECT 22.950 457.950 25.050 458.400 ;
        RECT 46.950 459.600 49.050 460.050 ;
        RECT 76.950 459.600 79.050 460.050 ;
        RECT 163.950 459.600 166.050 460.050 ;
        RECT 46.950 458.400 166.050 459.600 ;
        RECT 46.950 457.950 49.050 458.400 ;
        RECT 76.950 457.950 79.050 458.400 ;
        RECT 163.950 457.950 166.050 458.400 ;
        RECT 193.950 459.600 196.050 460.050 ;
        RECT 196.950 459.600 199.050 460.050 ;
        RECT 208.950 459.600 211.050 460.050 ;
        RECT 193.950 458.400 211.050 459.600 ;
        RECT 193.950 457.950 196.050 458.400 ;
        RECT 196.950 457.950 199.050 458.400 ;
        RECT 208.950 457.950 211.050 458.400 ;
        RECT 238.950 459.600 241.050 460.050 ;
        RECT 283.950 459.600 286.050 460.050 ;
        RECT 238.950 458.400 286.050 459.600 ;
        RECT 238.950 457.950 241.050 458.400 ;
        RECT 283.950 457.950 286.050 458.400 ;
        RECT 307.950 459.600 310.050 460.050 ;
        RECT 319.950 459.600 322.050 460.050 ;
        RECT 418.950 459.600 421.050 460.050 ;
        RECT 307.950 458.400 421.050 459.600 ;
        RECT 307.950 457.950 310.050 458.400 ;
        RECT 319.950 457.950 322.050 458.400 ;
        RECT 418.950 457.950 421.050 458.400 ;
        RECT 430.950 459.600 433.050 460.050 ;
        RECT 439.950 459.600 442.050 460.050 ;
        RECT 430.950 458.400 442.050 459.600 ;
        RECT 430.950 457.950 433.050 458.400 ;
        RECT 439.950 457.950 442.050 458.400 ;
        RECT 451.950 459.600 454.050 460.050 ;
        RECT 466.950 459.600 469.050 460.050 ;
        RECT 451.950 458.400 469.050 459.600 ;
        RECT 500.400 459.600 501.600 461.400 ;
        RECT 502.950 461.400 676.050 462.600 ;
        RECT 502.950 460.950 505.050 461.400 ;
        RECT 568.950 460.950 571.050 461.400 ;
        RECT 619.950 460.950 622.050 461.400 ;
        RECT 673.950 460.950 676.050 461.400 ;
        RECT 724.950 462.600 727.050 463.050 ;
        RECT 775.950 462.600 778.050 463.050 ;
        RECT 802.950 462.600 805.050 463.050 ;
        RECT 724.950 461.400 805.050 462.600 ;
        RECT 724.950 460.950 727.050 461.400 ;
        RECT 775.950 460.950 778.050 461.400 ;
        RECT 802.950 460.950 805.050 461.400 ;
        RECT 529.950 459.600 532.050 460.050 ;
        RECT 565.950 459.600 568.050 460.050 ;
        RECT 500.400 458.400 568.050 459.600 ;
        RECT 451.950 457.950 454.050 458.400 ;
        RECT 466.950 457.950 469.050 458.400 ;
        RECT 529.950 457.950 532.050 458.400 ;
        RECT 565.950 457.950 568.050 458.400 ;
        RECT 592.950 459.600 595.050 460.050 ;
        RECT 682.950 459.600 685.050 460.050 ;
        RECT 592.950 458.400 685.050 459.600 ;
        RECT 592.950 457.950 595.050 458.400 ;
        RECT 682.950 457.950 685.050 458.400 ;
        RECT 718.950 459.600 721.050 460.050 ;
        RECT 748.950 459.600 751.050 460.050 ;
        RECT 760.950 459.600 763.050 460.050 ;
        RECT 718.950 458.400 763.050 459.600 ;
        RECT 718.950 457.950 721.050 458.400 ;
        RECT 748.950 457.950 751.050 458.400 ;
        RECT 760.950 457.950 763.050 458.400 ;
        RECT 40.950 456.600 43.050 457.050 ;
        RECT 11.400 455.400 43.050 456.600 ;
        RECT 11.400 454.050 12.600 455.400 ;
        RECT 40.950 454.950 43.050 455.400 ;
        RECT 82.950 456.600 85.050 457.050 ;
        RECT 112.950 456.600 115.050 457.050 ;
        RECT 82.950 455.400 115.050 456.600 ;
        RECT 82.950 454.950 85.050 455.400 ;
        RECT 112.950 454.950 115.050 455.400 ;
        RECT 160.950 456.600 163.050 457.050 ;
        RECT 166.950 456.600 169.050 457.050 ;
        RECT 169.950 456.600 172.050 457.050 ;
        RECT 160.950 455.400 172.050 456.600 ;
        RECT 160.950 454.950 163.050 455.400 ;
        RECT 166.950 454.950 169.050 455.400 ;
        RECT 169.950 454.950 172.050 455.400 ;
        RECT 178.950 456.600 181.050 457.050 ;
        RECT 187.950 456.600 190.050 457.050 ;
        RECT 178.950 455.400 190.050 456.600 ;
        RECT 178.950 454.950 181.050 455.400 ;
        RECT 187.950 454.950 190.050 455.400 ;
        RECT 283.950 456.600 286.050 457.050 ;
        RECT 292.950 456.600 295.050 457.050 ;
        RECT 283.950 455.400 295.050 456.600 ;
        RECT 283.950 454.950 286.050 455.400 ;
        RECT 292.950 454.950 295.050 455.400 ;
        RECT 313.950 456.600 316.050 457.050 ;
        RECT 319.950 456.600 322.050 457.050 ;
        RECT 313.950 455.400 322.050 456.600 ;
        RECT 313.950 454.950 316.050 455.400 ;
        RECT 319.950 454.950 322.050 455.400 ;
        RECT 328.950 456.600 331.050 457.050 ;
        RECT 334.950 456.600 337.050 457.050 ;
        RECT 346.950 456.600 349.050 457.050 ;
        RECT 376.950 456.600 379.050 457.050 ;
        RECT 328.950 455.400 345.600 456.600 ;
        RECT 328.950 454.950 331.050 455.400 ;
        RECT 334.950 454.950 337.050 455.400 ;
        RECT 10.950 451.950 13.050 454.050 ;
        RECT 16.950 453.600 19.050 454.050 ;
        RECT 22.950 453.600 25.050 454.050 ;
        RECT 55.950 453.600 58.050 454.050 ;
        RECT 70.950 453.600 73.050 454.050 ;
        RECT 16.950 452.400 73.050 453.600 ;
        RECT 16.950 451.950 19.050 452.400 ;
        RECT 22.950 451.950 25.050 452.400 ;
        RECT 55.950 451.950 58.050 452.400 ;
        RECT 70.950 451.950 73.050 452.400 ;
        RECT 115.950 453.600 118.050 454.050 ;
        RECT 130.950 453.600 133.050 454.050 ;
        RECT 115.950 452.400 133.050 453.600 ;
        RECT 115.950 451.950 118.050 452.400 ;
        RECT 130.950 451.950 133.050 452.400 ;
        RECT 205.950 453.600 208.050 454.050 ;
        RECT 211.950 453.600 214.050 454.050 ;
        RECT 205.950 452.400 214.050 453.600 ;
        RECT 205.950 451.950 208.050 452.400 ;
        RECT 211.950 451.950 214.050 452.400 ;
        RECT 217.950 453.600 220.050 454.050 ;
        RECT 232.950 453.600 235.050 454.050 ;
        RECT 217.950 452.400 235.050 453.600 ;
        RECT 217.950 451.950 220.050 452.400 ;
        RECT 232.950 451.950 235.050 452.400 ;
        RECT 292.950 453.600 295.050 454.050 ;
        RECT 301.950 453.600 304.050 454.050 ;
        RECT 292.950 452.400 304.050 453.600 ;
        RECT 292.950 451.950 295.050 452.400 ;
        RECT 301.950 451.950 304.050 452.400 ;
        RECT 316.950 453.600 319.050 454.050 ;
        RECT 331.950 453.600 334.050 454.050 ;
        RECT 316.950 452.400 334.050 453.600 ;
        RECT 344.400 453.600 345.600 455.400 ;
        RECT 346.950 455.400 379.050 456.600 ;
        RECT 346.950 454.950 349.050 455.400 ;
        RECT 376.950 454.950 379.050 455.400 ;
        RECT 430.950 456.600 433.050 457.050 ;
        RECT 472.950 456.600 475.050 457.050 ;
        RECT 478.950 456.600 481.050 457.050 ;
        RECT 430.950 455.400 468.600 456.600 ;
        RECT 430.950 454.950 433.050 455.400 ;
        RECT 358.950 453.600 361.050 454.050 ;
        RECT 344.400 452.400 361.050 453.600 ;
        RECT 316.950 451.950 319.050 452.400 ;
        RECT 331.950 451.950 334.050 452.400 ;
        RECT 358.950 451.950 361.050 452.400 ;
        RECT 373.950 453.600 376.050 454.050 ;
        RECT 388.950 453.600 391.050 454.050 ;
        RECT 400.950 453.600 403.050 454.050 ;
        RECT 373.950 452.400 403.050 453.600 ;
        RECT 373.950 451.950 376.050 452.400 ;
        RECT 388.950 451.950 391.050 452.400 ;
        RECT 400.950 451.950 403.050 452.400 ;
        RECT 406.950 453.600 409.050 454.050 ;
        RECT 424.950 453.600 427.050 454.050 ;
        RECT 406.950 452.400 427.050 453.600 ;
        RECT 406.950 451.950 409.050 452.400 ;
        RECT 424.950 451.950 427.050 452.400 ;
        RECT 445.950 453.600 448.050 454.050 ;
        RECT 463.950 453.600 466.050 454.050 ;
        RECT 445.950 452.400 466.050 453.600 ;
        RECT 467.400 453.600 468.600 455.400 ;
        RECT 472.950 455.400 481.050 456.600 ;
        RECT 472.950 454.950 475.050 455.400 ;
        RECT 478.950 454.950 481.050 455.400 ;
        RECT 499.950 456.600 502.050 457.050 ;
        RECT 511.950 456.600 514.050 457.050 ;
        RECT 499.950 455.400 514.050 456.600 ;
        RECT 499.950 454.950 502.050 455.400 ;
        RECT 511.950 454.950 514.050 455.400 ;
        RECT 514.950 456.600 517.050 457.050 ;
        RECT 544.950 456.600 547.050 457.050 ;
        RECT 514.950 455.400 547.050 456.600 ;
        RECT 514.950 454.950 517.050 455.400 ;
        RECT 544.950 454.950 547.050 455.400 ;
        RECT 553.950 456.600 556.050 457.050 ;
        RECT 601.950 456.600 604.050 457.050 ;
        RECT 553.950 455.400 604.050 456.600 ;
        RECT 553.950 454.950 556.050 455.400 ;
        RECT 601.950 454.950 604.050 455.400 ;
        RECT 604.950 456.600 607.050 457.050 ;
        RECT 646.950 456.600 649.050 457.050 ;
        RECT 604.950 455.400 649.050 456.600 ;
        RECT 604.950 454.950 607.050 455.400 ;
        RECT 646.950 454.950 649.050 455.400 ;
        RECT 655.950 456.600 658.050 457.050 ;
        RECT 661.950 456.600 664.050 457.050 ;
        RECT 691.950 456.600 694.050 457.050 ;
        RECT 727.950 456.600 730.050 457.050 ;
        RECT 655.950 455.400 660.600 456.600 ;
        RECT 655.950 454.950 658.050 455.400 ;
        RECT 469.950 453.600 472.050 454.050 ;
        RECT 467.400 452.400 472.050 453.600 ;
        RECT 445.950 451.950 448.050 452.400 ;
        RECT 463.950 451.950 466.050 452.400 ;
        RECT 469.950 451.950 472.050 452.400 ;
        RECT 487.950 451.950 490.050 454.050 ;
        RECT 529.950 453.600 532.050 454.050 ;
        RECT 541.950 453.600 544.050 454.050 ;
        RECT 529.950 452.400 544.050 453.600 ;
        RECT 529.950 451.950 532.050 452.400 ;
        RECT 541.950 451.950 544.050 452.400 ;
        RECT 550.950 453.600 553.050 454.050 ;
        RECT 568.950 453.600 571.050 454.050 ;
        RECT 550.950 452.400 571.050 453.600 ;
        RECT 550.950 451.950 553.050 452.400 ;
        RECT 568.950 451.950 571.050 452.400 ;
        RECT 571.950 453.600 574.050 454.050 ;
        RECT 598.950 453.600 601.050 454.050 ;
        RECT 571.950 452.400 601.050 453.600 ;
        RECT 571.950 451.950 574.050 452.400 ;
        RECT 598.950 451.950 601.050 452.400 ;
        RECT 604.950 453.600 607.050 454.050 ;
        RECT 610.950 453.600 613.050 454.050 ;
        RECT 652.950 453.600 655.050 454.050 ;
        RECT 659.400 453.600 660.600 455.400 ;
        RECT 661.950 455.400 730.050 456.600 ;
        RECT 661.950 454.950 664.050 455.400 ;
        RECT 691.950 454.950 694.050 455.400 ;
        RECT 727.950 454.950 730.050 455.400 ;
        RECT 730.950 456.600 733.050 457.050 ;
        RECT 739.950 456.600 742.050 457.050 ;
        RECT 730.950 455.400 742.050 456.600 ;
        RECT 730.950 454.950 733.050 455.400 ;
        RECT 739.950 454.950 742.050 455.400 ;
        RECT 745.950 456.600 748.050 457.050 ;
        RECT 754.950 456.600 757.050 457.050 ;
        RECT 745.950 455.400 757.050 456.600 ;
        RECT 745.950 454.950 748.050 455.400 ;
        RECT 754.950 454.950 757.050 455.400 ;
        RECT 787.950 456.600 790.050 457.050 ;
        RECT 799.950 456.600 802.050 457.050 ;
        RECT 811.950 456.600 814.050 457.050 ;
        RECT 868.950 456.600 871.050 457.050 ;
        RECT 787.950 455.400 814.050 456.600 ;
        RECT 787.950 454.950 790.050 455.400 ;
        RECT 799.950 454.950 802.050 455.400 ;
        RECT 811.950 454.950 814.050 455.400 ;
        RECT 857.400 455.400 871.050 456.600 ;
        RECT 676.950 453.600 679.050 454.050 ;
        RECT 604.950 452.400 655.050 453.600 ;
        RECT 604.950 451.950 607.050 452.400 ;
        RECT 610.950 451.950 613.050 452.400 ;
        RECT 652.950 451.950 655.050 452.400 ;
        RECT 656.400 452.400 679.050 453.600 ;
        RECT 64.950 450.600 67.050 451.050 ;
        RECT 85.950 450.600 88.050 451.050 ;
        RECT 94.950 450.600 97.050 451.050 ;
        RECT 64.950 449.400 97.050 450.600 ;
        RECT 64.950 448.950 67.050 449.400 ;
        RECT 85.950 448.950 88.050 449.400 ;
        RECT 94.950 448.950 97.050 449.400 ;
        RECT 109.950 450.600 112.050 451.050 ;
        RECT 133.950 450.600 136.050 451.050 ;
        RECT 139.950 450.600 142.050 451.050 ;
        RECT 109.950 449.400 142.050 450.600 ;
        RECT 109.950 448.950 112.050 449.400 ;
        RECT 133.950 448.950 136.050 449.400 ;
        RECT 139.950 448.950 142.050 449.400 ;
        RECT 172.950 450.600 175.050 451.050 ;
        RECT 178.950 450.600 181.050 451.050 ;
        RECT 172.950 449.400 181.050 450.600 ;
        RECT 172.950 448.950 175.050 449.400 ;
        RECT 178.950 448.950 181.050 449.400 ;
        RECT 211.950 450.600 214.050 451.050 ;
        RECT 235.950 450.600 238.050 451.050 ;
        RECT 244.950 450.600 247.050 451.050 ;
        RECT 211.950 449.400 247.050 450.600 ;
        RECT 211.950 448.950 214.050 449.400 ;
        RECT 235.950 448.950 238.050 449.400 ;
        RECT 244.950 448.950 247.050 449.400 ;
        RECT 289.950 450.600 292.050 451.050 ;
        RECT 298.950 450.600 301.050 451.050 ;
        RECT 337.950 450.600 340.050 451.050 ;
        RECT 289.950 449.400 340.050 450.600 ;
        RECT 289.950 448.950 292.050 449.400 ;
        RECT 298.950 448.950 301.050 449.400 ;
        RECT 337.950 448.950 340.050 449.400 ;
        RECT 394.950 450.600 397.050 451.050 ;
        RECT 403.950 450.600 406.050 451.050 ;
        RECT 394.950 449.400 406.050 450.600 ;
        RECT 394.950 448.950 397.050 449.400 ;
        RECT 403.950 448.950 406.050 449.400 ;
        RECT 412.950 450.600 415.050 451.050 ;
        RECT 448.950 450.600 451.050 451.050 ;
        RECT 478.950 450.600 481.050 451.050 ;
        RECT 412.950 449.400 481.050 450.600 ;
        RECT 412.950 448.950 415.050 449.400 ;
        RECT 448.950 448.950 451.050 449.400 ;
        RECT 478.950 448.950 481.050 449.400 ;
        RECT 460.950 447.600 463.050 448.050 ;
        RECT 488.400 447.600 489.600 451.950 ;
        RECT 511.950 450.600 514.050 451.050 ;
        RECT 535.950 450.600 538.050 451.050 ;
        RECT 511.950 449.400 538.050 450.600 ;
        RECT 511.950 448.950 514.050 449.400 ;
        RECT 535.950 448.950 538.050 449.400 ;
        RECT 538.950 450.600 541.050 451.050 ;
        RECT 553.950 450.600 556.050 451.050 ;
        RECT 538.950 449.400 556.050 450.600 ;
        RECT 538.950 448.950 541.050 449.400 ;
        RECT 553.950 448.950 556.050 449.400 ;
        RECT 640.950 450.600 643.050 451.050 ;
        RECT 656.400 450.600 657.600 452.400 ;
        RECT 676.950 451.950 679.050 452.400 ;
        RECT 700.950 453.600 703.050 454.050 ;
        RECT 724.950 453.600 727.050 454.050 ;
        RECT 700.950 452.400 727.050 453.600 ;
        RECT 700.950 451.950 703.050 452.400 ;
        RECT 724.950 451.950 727.050 452.400 ;
        RECT 826.950 453.600 829.050 454.050 ;
        RECT 850.950 453.600 853.050 454.050 ;
        RECT 857.400 453.600 858.600 455.400 ;
        RECT 868.950 454.950 871.050 455.400 ;
        RECT 826.950 452.400 858.600 453.600 ;
        RECT 826.950 451.950 829.050 452.400 ;
        RECT 850.950 451.950 853.050 452.400 ;
        RECT 697.950 450.600 700.050 451.050 ;
        RECT 640.950 449.400 657.600 450.600 ;
        RECT 665.400 449.400 700.050 450.600 ;
        RECT 640.950 448.950 643.050 449.400 ;
        RECT 460.950 446.400 489.600 447.600 ;
        RECT 505.950 447.600 508.050 448.050 ;
        RECT 514.950 447.600 517.050 448.050 ;
        RECT 505.950 446.400 517.050 447.600 ;
        RECT 460.950 445.950 463.050 446.400 ;
        RECT 505.950 445.950 508.050 446.400 ;
        RECT 514.950 445.950 517.050 446.400 ;
        RECT 574.950 447.600 577.050 448.050 ;
        RECT 619.950 447.600 622.050 448.050 ;
        RECT 574.950 446.400 622.050 447.600 ;
        RECT 574.950 445.950 577.050 446.400 ;
        RECT 619.950 445.950 622.050 446.400 ;
        RECT 646.950 447.600 649.050 448.050 ;
        RECT 665.400 447.600 666.600 449.400 ;
        RECT 697.950 448.950 700.050 449.400 ;
        RECT 703.950 450.600 706.050 451.050 ;
        RECT 715.950 450.600 718.050 451.050 ;
        RECT 703.950 449.400 718.050 450.600 ;
        RECT 703.950 448.950 706.050 449.400 ;
        RECT 715.950 448.950 718.050 449.400 ;
        RECT 727.950 450.600 730.050 451.050 ;
        RECT 733.950 450.600 736.050 451.050 ;
        RECT 727.950 449.400 736.050 450.600 ;
        RECT 727.950 448.950 730.050 449.400 ;
        RECT 733.950 448.950 736.050 449.400 ;
        RECT 646.950 446.400 666.600 447.600 ;
        RECT 646.950 445.950 649.050 446.400 ;
        RECT 79.950 444.600 82.050 445.050 ;
        RECT 91.950 444.600 94.050 445.050 ;
        RECT 79.950 443.400 94.050 444.600 ;
        RECT 79.950 442.950 82.050 443.400 ;
        RECT 91.950 442.950 94.050 443.400 ;
        RECT 127.950 444.600 130.050 445.050 ;
        RECT 136.950 444.600 139.050 445.050 ;
        RECT 127.950 443.400 139.050 444.600 ;
        RECT 127.950 442.950 130.050 443.400 ;
        RECT 136.950 442.950 139.050 443.400 ;
        RECT 280.950 444.600 283.050 445.050 ;
        RECT 322.950 444.600 325.050 445.050 ;
        RECT 280.950 443.400 325.050 444.600 ;
        RECT 280.950 442.950 283.050 443.400 ;
        RECT 322.950 442.950 325.050 443.400 ;
        RECT 343.950 444.600 346.050 445.050 ;
        RECT 352.950 444.600 355.050 445.050 ;
        RECT 412.950 444.600 415.050 445.050 ;
        RECT 343.950 443.400 415.050 444.600 ;
        RECT 343.950 442.950 346.050 443.400 ;
        RECT 352.950 442.950 355.050 443.400 ;
        RECT 412.950 442.950 415.050 443.400 ;
        RECT 457.950 444.600 460.050 445.050 ;
        RECT 505.950 444.600 508.050 445.050 ;
        RECT 457.950 443.400 508.050 444.600 ;
        RECT 457.950 442.950 460.050 443.400 ;
        RECT 505.950 442.950 508.050 443.400 ;
        RECT 574.950 444.600 577.050 445.050 ;
        RECT 589.950 444.600 592.050 445.050 ;
        RECT 574.950 443.400 592.050 444.600 ;
        RECT 574.950 442.950 577.050 443.400 ;
        RECT 589.950 442.950 592.050 443.400 ;
        RECT 352.950 441.600 355.050 442.050 ;
        RECT 367.950 441.600 370.050 442.050 ;
        RECT 352.950 440.400 370.050 441.600 ;
        RECT 352.950 439.950 355.050 440.400 ;
        RECT 367.950 439.950 370.050 440.400 ;
        RECT 595.950 441.600 598.050 442.050 ;
        RECT 601.950 441.600 604.050 442.050 ;
        RECT 658.950 441.600 661.050 442.050 ;
        RECT 595.950 440.400 661.050 441.600 ;
        RECT 595.950 439.950 598.050 440.400 ;
        RECT 601.950 439.950 604.050 440.400 ;
        RECT 658.950 439.950 661.050 440.400 ;
        RECT 685.950 441.600 688.050 442.050 ;
        RECT 760.950 441.600 763.050 442.050 ;
        RECT 685.950 440.400 763.050 441.600 ;
        RECT 685.950 439.950 688.050 440.400 ;
        RECT 760.950 439.950 763.050 440.400 ;
        RECT 442.950 438.600 445.050 439.050 ;
        RECT 454.950 438.600 457.050 439.050 ;
        RECT 442.950 437.400 457.050 438.600 ;
        RECT 442.950 436.950 445.050 437.400 ;
        RECT 454.950 436.950 457.050 437.400 ;
        RECT 865.950 438.600 868.050 439.050 ;
        RECT 874.950 438.600 877.050 439.050 ;
        RECT 865.950 437.400 877.050 438.600 ;
        RECT 865.950 436.950 868.050 437.400 ;
        RECT 874.950 436.950 877.050 437.400 ;
        RECT 304.950 429.600 307.050 430.050 ;
        RECT 511.950 429.600 514.050 430.050 ;
        RECT 304.950 428.400 514.050 429.600 ;
        RECT 304.950 427.950 307.050 428.400 ;
        RECT 511.950 427.950 514.050 428.400 ;
        RECT 577.950 429.600 580.050 430.050 ;
        RECT 733.950 429.600 736.050 430.050 ;
        RECT 577.950 428.400 736.050 429.600 ;
        RECT 577.950 427.950 580.050 428.400 ;
        RECT 733.950 427.950 736.050 428.400 ;
        RECT 841.950 429.600 844.050 430.050 ;
        RECT 859.950 429.600 862.050 430.050 ;
        RECT 841.950 428.400 862.050 429.600 ;
        RECT 841.950 427.950 844.050 428.400 ;
        RECT 859.950 427.950 862.050 428.400 ;
        RECT 517.950 426.600 520.050 427.050 ;
        RECT 598.950 426.600 601.050 427.050 ;
        RECT 625.950 426.600 628.050 427.050 ;
        RECT 517.950 425.400 628.050 426.600 ;
        RECT 517.950 424.950 520.050 425.400 ;
        RECT 598.950 424.950 601.050 425.400 ;
        RECT 625.950 424.950 628.050 425.400 ;
        RECT 628.950 426.600 631.050 427.050 ;
        RECT 694.950 426.600 697.050 427.050 ;
        RECT 628.950 425.400 697.050 426.600 ;
        RECT 628.950 424.950 631.050 425.400 ;
        RECT 694.950 424.950 697.050 425.400 ;
        RECT 172.950 423.600 175.050 424.050 ;
        RECT 181.950 423.600 184.050 424.050 ;
        RECT 172.950 422.400 184.050 423.600 ;
        RECT 172.950 421.950 175.050 422.400 ;
        RECT 181.950 421.950 184.050 422.400 ;
        RECT 253.950 423.600 256.050 424.050 ;
        RECT 304.950 423.600 307.050 424.050 ;
        RECT 253.950 422.400 307.050 423.600 ;
        RECT 253.950 421.950 256.050 422.400 ;
        RECT 304.950 421.950 307.050 422.400 ;
        RECT 364.950 423.600 367.050 424.050 ;
        RECT 442.950 423.600 445.050 424.050 ;
        RECT 364.950 422.400 445.050 423.600 ;
        RECT 364.950 421.950 367.050 422.400 ;
        RECT 442.950 421.950 445.050 422.400 ;
        RECT 460.950 423.600 463.050 424.050 ;
        RECT 589.950 423.600 592.050 424.050 ;
        RECT 616.950 423.600 619.050 424.050 ;
        RECT 460.950 422.400 619.050 423.600 ;
        RECT 460.950 421.950 463.050 422.400 ;
        RECT 589.950 421.950 592.050 422.400 ;
        RECT 616.950 421.950 619.050 422.400 ;
        RECT 619.950 423.600 622.050 424.050 ;
        RECT 634.950 423.600 637.050 424.050 ;
        RECT 682.950 423.600 685.050 424.050 ;
        RECT 619.950 422.400 685.050 423.600 ;
        RECT 619.950 421.950 622.050 422.400 ;
        RECT 634.950 421.950 637.050 422.400 ;
        RECT 682.950 421.950 685.050 422.400 ;
        RECT 271.950 420.600 274.050 421.050 ;
        RECT 271.950 419.400 279.600 420.600 ;
        RECT 271.950 418.950 274.050 419.400 ;
        RECT 199.950 417.600 202.050 418.050 ;
        RECT 205.950 417.600 208.050 418.050 ;
        RECT 199.950 416.400 208.050 417.600 ;
        RECT 199.950 415.950 202.050 416.400 ;
        RECT 205.950 415.950 208.050 416.400 ;
        RECT 217.950 417.600 220.050 418.050 ;
        RECT 232.950 417.600 235.050 418.050 ;
        RECT 217.950 416.400 235.050 417.600 ;
        RECT 217.950 415.950 220.050 416.400 ;
        RECT 232.950 415.950 235.050 416.400 ;
        RECT 250.950 415.950 253.050 418.050 ;
        RECT 262.950 417.600 265.050 418.050 ;
        RECT 268.950 417.600 271.050 418.050 ;
        RECT 274.950 417.600 277.050 418.050 ;
        RECT 262.950 416.400 271.050 417.600 ;
        RECT 262.950 415.950 265.050 416.400 ;
        RECT 268.950 415.950 271.050 416.400 ;
        RECT 272.400 416.400 277.050 417.600 ;
        RECT 7.950 414.600 10.050 415.050 ;
        RECT 16.950 414.600 19.050 415.050 ;
        RECT 52.950 414.600 55.050 415.050 ;
        RECT 7.950 413.400 55.050 414.600 ;
        RECT 7.950 412.950 10.050 413.400 ;
        RECT 16.950 412.950 19.050 413.400 ;
        RECT 52.950 412.950 55.050 413.400 ;
        RECT 76.950 414.600 79.050 415.050 ;
        RECT 91.950 414.600 94.050 415.050 ;
        RECT 76.950 413.400 94.050 414.600 ;
        RECT 76.950 412.950 79.050 413.400 ;
        RECT 91.950 412.950 94.050 413.400 ;
        RECT 115.950 414.600 118.050 415.050 ;
        RECT 130.950 414.600 133.050 415.050 ;
        RECT 115.950 413.400 133.050 414.600 ;
        RECT 115.950 412.950 118.050 413.400 ;
        RECT 130.950 412.950 133.050 413.400 ;
        RECT 169.950 414.600 172.050 415.050 ;
        RECT 184.950 414.600 187.050 415.050 ;
        RECT 169.950 413.400 187.050 414.600 ;
        RECT 169.950 412.950 172.050 413.400 ;
        RECT 184.950 412.950 187.050 413.400 ;
        RECT 208.950 414.600 211.050 415.050 ;
        RECT 247.950 414.600 250.050 415.050 ;
        RECT 208.950 413.400 250.050 414.600 ;
        RECT 208.950 412.950 211.050 413.400 ;
        RECT 247.950 412.950 250.050 413.400 ;
        RECT 251.400 412.050 252.600 415.950 ;
        RECT 268.950 414.600 271.050 415.050 ;
        RECT 272.400 414.600 273.600 416.400 ;
        RECT 274.950 415.950 277.050 416.400 ;
        RECT 268.950 413.400 273.600 414.600 ;
        RECT 278.400 414.600 279.600 419.400 ;
        RECT 292.950 418.950 295.050 421.050 ;
        RECT 310.950 420.600 313.050 421.050 ;
        RECT 296.400 419.400 313.050 420.600 ;
        RECT 293.400 415.050 294.600 418.950 ;
        RECT 296.400 418.050 297.600 419.400 ;
        RECT 310.950 418.950 313.050 419.400 ;
        RECT 358.950 420.600 361.050 421.050 ;
        RECT 373.950 420.600 376.050 421.050 ;
        RECT 385.950 420.600 388.050 421.050 ;
        RECT 409.950 420.600 412.050 421.050 ;
        RECT 358.950 419.400 376.050 420.600 ;
        RECT 358.950 418.950 361.050 419.400 ;
        RECT 373.950 418.950 376.050 419.400 ;
        RECT 377.400 419.400 388.050 420.600 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 307.950 417.600 310.050 418.050 ;
        RECT 319.950 417.600 322.050 418.050 ;
        RECT 307.950 416.400 322.050 417.600 ;
        RECT 307.950 415.950 310.050 416.400 ;
        RECT 319.950 415.950 322.050 416.400 ;
        RECT 325.950 417.600 328.050 418.050 ;
        RECT 337.950 417.600 340.050 418.050 ;
        RECT 377.400 417.600 378.600 419.400 ;
        RECT 385.950 418.950 388.050 419.400 ;
        RECT 389.400 419.400 412.050 420.600 ;
        RECT 325.950 416.400 340.050 417.600 ;
        RECT 325.950 415.950 328.050 416.400 ;
        RECT 337.950 415.950 340.050 416.400 ;
        RECT 341.400 416.400 378.600 417.600 ;
        RECT 379.950 417.600 382.050 418.050 ;
        RECT 389.400 417.600 390.600 419.400 ;
        RECT 409.950 418.950 412.050 419.400 ;
        RECT 484.950 420.600 487.050 421.050 ;
        RECT 526.950 420.600 529.050 421.050 ;
        RECT 544.950 420.600 547.050 421.050 ;
        RECT 547.950 420.600 550.050 421.050 ;
        RECT 484.950 419.400 550.050 420.600 ;
        RECT 484.950 418.950 487.050 419.400 ;
        RECT 526.950 418.950 529.050 419.400 ;
        RECT 544.950 418.950 547.050 419.400 ;
        RECT 547.950 418.950 550.050 419.400 ;
        RECT 613.950 420.600 616.050 421.050 ;
        RECT 631.950 420.600 634.050 421.050 ;
        RECT 718.950 420.600 721.050 421.050 ;
        RECT 613.950 419.400 721.050 420.600 ;
        RECT 613.950 418.950 616.050 419.400 ;
        RECT 631.950 418.950 634.050 419.400 ;
        RECT 718.950 418.950 721.050 419.400 ;
        RECT 379.950 416.400 390.600 417.600 ;
        RECT 397.950 417.600 400.050 418.050 ;
        RECT 409.950 417.600 412.050 418.050 ;
        RECT 415.950 417.600 418.050 418.050 ;
        RECT 397.950 416.400 418.050 417.600 ;
        RECT 286.950 414.600 289.050 415.050 ;
        RECT 278.400 413.400 289.050 414.600 ;
        RECT 268.950 412.950 271.050 413.400 ;
        RECT 286.950 412.950 289.050 413.400 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 301.950 414.600 304.050 415.050 ;
        RECT 313.950 414.600 316.050 415.050 ;
        RECT 341.400 414.600 342.600 416.400 ;
        RECT 379.950 415.950 382.050 416.400 ;
        RECT 397.950 415.950 400.050 416.400 ;
        RECT 409.950 415.950 412.050 416.400 ;
        RECT 415.950 415.950 418.050 416.400 ;
        RECT 445.950 417.600 448.050 418.050 ;
        RECT 481.950 417.600 484.050 418.050 ;
        RECT 445.950 416.400 484.050 417.600 ;
        RECT 445.950 415.950 448.050 416.400 ;
        RECT 481.950 415.950 484.050 416.400 ;
        RECT 526.950 417.600 529.050 418.050 ;
        RECT 565.950 417.600 568.050 418.050 ;
        RECT 580.950 417.600 583.050 418.050 ;
        RECT 586.950 417.600 589.050 418.050 ;
        RECT 631.950 417.600 634.050 418.050 ;
        RECT 526.950 416.400 564.600 417.600 ;
        RECT 526.950 415.950 529.050 416.400 ;
        RECT 301.950 413.400 316.050 414.600 ;
        RECT 301.950 412.950 304.050 413.400 ;
        RECT 313.950 412.950 316.050 413.400 ;
        RECT 317.400 413.400 342.600 414.600 ;
        RECT 343.950 414.600 346.050 415.050 ;
        RECT 361.950 414.600 364.050 415.050 ;
        RECT 343.950 413.400 364.050 414.600 ;
        RECT 13.950 411.600 16.050 412.050 ;
        RECT 34.950 411.600 37.050 412.050 ;
        RECT 13.950 410.400 37.050 411.600 ;
        RECT 13.950 409.950 16.050 410.400 ;
        RECT 34.950 409.950 37.050 410.400 ;
        RECT 52.950 411.600 55.050 412.050 ;
        RECT 61.950 411.600 64.050 412.050 ;
        RECT 88.950 411.600 91.050 412.050 ;
        RECT 52.950 410.400 91.050 411.600 ;
        RECT 52.950 409.950 55.050 410.400 ;
        RECT 61.950 409.950 64.050 410.400 ;
        RECT 88.950 409.950 91.050 410.400 ;
        RECT 100.950 411.600 103.050 412.050 ;
        RECT 112.950 411.600 115.050 412.050 ;
        RECT 100.950 410.400 115.050 411.600 ;
        RECT 100.950 409.950 103.050 410.400 ;
        RECT 112.950 409.950 115.050 410.400 ;
        RECT 187.950 411.600 190.050 412.050 ;
        RECT 223.950 411.600 226.050 412.050 ;
        RECT 187.950 410.400 226.050 411.600 ;
        RECT 187.950 409.950 190.050 410.400 ;
        RECT 223.950 409.950 226.050 410.400 ;
        RECT 250.950 409.950 253.050 412.050 ;
        RECT 256.950 411.600 259.050 412.050 ;
        RECT 265.950 411.600 268.050 412.050 ;
        RECT 256.950 410.400 268.050 411.600 ;
        RECT 256.950 409.950 259.050 410.400 ;
        RECT 265.950 409.950 268.050 410.400 ;
        RECT 280.950 411.600 283.050 412.050 ;
        RECT 289.950 411.600 292.050 412.050 ;
        RECT 280.950 410.400 292.050 411.600 ;
        RECT 280.950 409.950 283.050 410.400 ;
        RECT 289.950 409.950 292.050 410.400 ;
        RECT 310.950 411.600 313.050 412.050 ;
        RECT 317.400 411.600 318.600 413.400 ;
        RECT 343.950 412.950 346.050 413.400 ;
        RECT 361.950 412.950 364.050 413.400 ;
        RECT 382.950 414.600 385.050 415.050 ;
        RECT 418.950 414.600 421.050 415.050 ;
        RECT 382.950 413.400 421.050 414.600 ;
        RECT 382.950 412.950 385.050 413.400 ;
        RECT 418.950 412.950 421.050 413.400 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 469.950 414.600 472.050 415.050 ;
        RECT 446.400 413.400 472.050 414.600 ;
        RECT 310.950 410.400 318.600 411.600 ;
        RECT 349.950 411.600 352.050 412.050 ;
        RECT 376.950 411.600 379.050 412.050 ;
        RECT 349.950 410.400 379.050 411.600 ;
        RECT 310.950 409.950 313.050 410.400 ;
        RECT 349.950 409.950 352.050 410.400 ;
        RECT 376.950 409.950 379.050 410.400 ;
        RECT 409.950 411.600 412.050 412.050 ;
        RECT 437.400 411.600 438.600 412.950 ;
        RECT 409.950 410.400 438.600 411.600 ;
        RECT 409.950 409.950 412.050 410.400 ;
        RECT 446.400 409.050 447.600 413.400 ;
        RECT 469.950 412.950 472.050 413.400 ;
        RECT 511.950 414.600 514.050 415.050 ;
        RECT 526.950 414.600 529.050 415.050 ;
        RECT 511.950 413.400 529.050 414.600 ;
        RECT 511.950 412.950 514.050 413.400 ;
        RECT 526.950 412.950 529.050 413.400 ;
        RECT 541.950 414.600 544.050 415.050 ;
        RECT 559.950 414.600 562.050 415.050 ;
        RECT 541.950 413.400 562.050 414.600 ;
        RECT 563.400 414.600 564.600 416.400 ;
        RECT 565.950 416.400 589.050 417.600 ;
        RECT 565.950 415.950 568.050 416.400 ;
        RECT 580.950 415.950 583.050 416.400 ;
        RECT 586.950 415.950 589.050 416.400 ;
        RECT 599.400 416.400 634.050 417.600 ;
        RECT 599.400 414.600 600.600 416.400 ;
        RECT 631.950 415.950 634.050 416.400 ;
        RECT 664.950 415.950 667.050 418.050 ;
        RECT 673.950 417.600 676.050 418.050 ;
        RECT 688.950 417.600 691.050 418.050 ;
        RECT 673.950 416.400 691.050 417.600 ;
        RECT 673.950 415.950 676.050 416.400 ;
        RECT 688.950 415.950 691.050 416.400 ;
        RECT 811.950 417.600 814.050 418.050 ;
        RECT 859.950 417.600 862.050 418.050 ;
        RECT 811.950 416.400 862.050 417.600 ;
        RECT 811.950 415.950 814.050 416.400 ;
        RECT 859.950 415.950 862.050 416.400 ;
        RECT 563.400 413.400 600.600 414.600 ;
        RECT 601.950 414.600 604.050 415.050 ;
        RECT 607.950 414.600 610.050 415.050 ;
        RECT 601.950 413.400 610.050 414.600 ;
        RECT 541.950 412.950 544.050 413.400 ;
        RECT 559.950 412.950 562.050 413.400 ;
        RECT 601.950 412.950 604.050 413.400 ;
        RECT 607.950 412.950 610.050 413.400 ;
        RECT 628.950 414.600 631.050 415.050 ;
        RECT 637.950 414.600 640.050 415.050 ;
        RECT 628.950 413.400 640.050 414.600 ;
        RECT 628.950 412.950 631.050 413.400 ;
        RECT 637.950 412.950 640.050 413.400 ;
        RECT 646.950 414.600 649.050 415.050 ;
        RECT 652.950 414.600 655.050 415.050 ;
        RECT 646.950 413.400 655.050 414.600 ;
        RECT 646.950 412.950 649.050 413.400 ;
        RECT 652.950 412.950 655.050 413.400 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 665.400 414.600 666.600 415.950 ;
        RECT 685.950 414.600 688.050 415.050 ;
        RECT 665.400 413.400 688.050 414.600 ;
        RECT 685.950 412.950 688.050 413.400 ;
        RECT 703.950 414.600 706.050 415.050 ;
        RECT 724.950 414.600 727.050 415.050 ;
        RECT 703.950 413.400 727.050 414.600 ;
        RECT 703.950 412.950 706.050 413.400 ;
        RECT 724.950 412.950 727.050 413.400 ;
        RECT 451.950 411.600 454.050 412.050 ;
        RECT 463.950 411.600 466.050 412.050 ;
        RECT 451.950 410.400 466.050 411.600 ;
        RECT 451.950 409.950 454.050 410.400 ;
        RECT 463.950 409.950 466.050 410.400 ;
        RECT 466.950 411.600 469.050 412.050 ;
        RECT 478.950 411.600 481.050 412.050 ;
        RECT 487.950 411.600 490.050 412.050 ;
        RECT 466.950 410.400 490.050 411.600 ;
        RECT 466.950 409.950 469.050 410.400 ;
        RECT 478.950 409.950 481.050 410.400 ;
        RECT 487.950 409.950 490.050 410.400 ;
        RECT 520.950 411.600 523.050 412.050 ;
        RECT 556.950 411.600 559.050 412.050 ;
        RECT 520.950 410.400 559.050 411.600 ;
        RECT 520.950 409.950 523.050 410.400 ;
        RECT 556.950 409.950 559.050 410.400 ;
        RECT 574.950 411.600 577.050 412.050 ;
        RECT 586.950 411.600 589.050 412.050 ;
        RECT 574.950 410.400 589.050 411.600 ;
        RECT 574.950 409.950 577.050 410.400 ;
        RECT 586.950 409.950 589.050 410.400 ;
        RECT 616.950 411.600 619.050 412.050 ;
        RECT 662.400 411.600 663.600 412.950 ;
        RECT 616.950 410.400 663.600 411.600 ;
        RECT 664.950 411.600 667.050 412.050 ;
        RECT 673.950 411.600 676.050 412.050 ;
        RECT 664.950 410.400 676.050 411.600 ;
        RECT 616.950 409.950 619.050 410.400 ;
        RECT 664.950 409.950 667.050 410.400 ;
        RECT 673.950 409.950 676.050 410.400 ;
        RECT 721.950 411.600 724.050 412.050 ;
        RECT 751.950 411.600 754.050 412.050 ;
        RECT 721.950 410.400 754.050 411.600 ;
        RECT 721.950 409.950 724.050 410.400 ;
        RECT 751.950 409.950 754.050 410.400 ;
        RECT 772.950 411.600 775.050 412.050 ;
        RECT 784.950 411.600 787.050 412.050 ;
        RECT 790.950 411.600 793.050 412.050 ;
        RECT 772.950 410.400 793.050 411.600 ;
        RECT 772.950 409.950 775.050 410.400 ;
        RECT 784.950 409.950 787.050 410.400 ;
        RECT 790.950 409.950 793.050 410.400 ;
        RECT 796.950 411.600 799.050 412.050 ;
        RECT 832.950 411.600 835.050 412.050 ;
        RECT 796.950 410.400 835.050 411.600 ;
        RECT 796.950 409.950 799.050 410.400 ;
        RECT 832.950 409.950 835.050 410.400 ;
        RECT 850.950 411.600 853.050 412.050 ;
        RECT 868.950 411.600 871.050 412.050 ;
        RECT 850.950 410.400 871.050 411.600 ;
        RECT 850.950 409.950 853.050 410.400 ;
        RECT 868.950 409.950 871.050 410.400 ;
        RECT 22.950 408.600 25.050 409.050 ;
        RECT 40.950 408.600 43.050 409.050 ;
        RECT 46.950 408.600 49.050 409.050 ;
        RECT 22.950 407.400 49.050 408.600 ;
        RECT 22.950 406.950 25.050 407.400 ;
        RECT 40.950 406.950 43.050 407.400 ;
        RECT 46.950 406.950 49.050 407.400 ;
        RECT 82.950 408.600 85.050 409.050 ;
        RECT 103.950 408.600 106.050 409.050 ;
        RECT 82.950 407.400 106.050 408.600 ;
        RECT 82.950 406.950 85.050 407.400 ;
        RECT 103.950 406.950 106.050 407.400 ;
        RECT 148.950 408.600 151.050 409.050 ;
        RECT 181.950 408.600 184.050 409.050 ;
        RECT 193.950 408.600 196.050 409.050 ;
        RECT 148.950 407.400 196.050 408.600 ;
        RECT 148.950 406.950 151.050 407.400 ;
        RECT 181.950 406.950 184.050 407.400 ;
        RECT 193.950 406.950 196.050 407.400 ;
        RECT 214.950 408.600 217.050 409.050 ;
        RECT 256.950 408.600 259.050 409.050 ;
        RECT 214.950 407.400 259.050 408.600 ;
        RECT 214.950 406.950 217.050 407.400 ;
        RECT 256.950 406.950 259.050 407.400 ;
        RECT 262.950 408.600 265.050 409.050 ;
        RECT 277.950 408.600 280.050 409.050 ;
        RECT 262.950 407.400 280.050 408.600 ;
        RECT 262.950 406.950 265.050 407.400 ;
        RECT 277.950 406.950 280.050 407.400 ;
        RECT 298.950 408.600 301.050 409.050 ;
        RECT 334.950 408.600 337.050 409.050 ;
        RECT 298.950 407.400 337.050 408.600 ;
        RECT 298.950 406.950 301.050 407.400 ;
        RECT 334.950 406.950 337.050 407.400 ;
        RECT 376.950 408.600 379.050 409.050 ;
        RECT 391.950 408.600 394.050 409.050 ;
        RECT 376.950 407.400 394.050 408.600 ;
        RECT 376.950 406.950 379.050 407.400 ;
        RECT 391.950 406.950 394.050 407.400 ;
        RECT 445.950 406.950 448.050 409.050 ;
        RECT 514.950 408.600 517.050 409.050 ;
        RECT 583.950 408.600 586.050 409.050 ;
        RECT 514.950 407.400 586.050 408.600 ;
        RECT 514.950 406.950 517.050 407.400 ;
        RECT 583.950 406.950 586.050 407.400 ;
        RECT 682.950 408.600 685.050 409.050 ;
        RECT 709.950 408.600 712.050 409.050 ;
        RECT 715.950 408.600 718.050 409.050 ;
        RECT 796.950 408.600 799.050 409.050 ;
        RECT 682.950 407.400 799.050 408.600 ;
        RECT 682.950 406.950 685.050 407.400 ;
        RECT 709.950 406.950 712.050 407.400 ;
        RECT 715.950 406.950 718.050 407.400 ;
        RECT 796.950 406.950 799.050 407.400 ;
        RECT 865.950 408.600 868.050 409.050 ;
        RECT 874.950 408.600 877.050 409.050 ;
        RECT 865.950 407.400 877.050 408.600 ;
        RECT 865.950 406.950 868.050 407.400 ;
        RECT 874.950 406.950 877.050 407.400 ;
        RECT 55.950 405.600 58.050 406.050 ;
        RECT 67.950 405.600 70.050 406.050 ;
        RECT 85.950 405.600 88.050 406.050 ;
        RECT 145.950 405.600 148.050 406.050 ;
        RECT 55.950 404.400 148.050 405.600 ;
        RECT 55.950 403.950 58.050 404.400 ;
        RECT 67.950 403.950 70.050 404.400 ;
        RECT 85.950 403.950 88.050 404.400 ;
        RECT 145.950 403.950 148.050 404.400 ;
        RECT 268.950 405.600 271.050 406.050 ;
        RECT 301.950 405.600 304.050 406.050 ;
        RECT 268.950 404.400 304.050 405.600 ;
        RECT 268.950 403.950 271.050 404.400 ;
        RECT 301.950 403.950 304.050 404.400 ;
        RECT 340.950 405.600 343.050 406.050 ;
        RECT 400.950 405.600 403.050 406.050 ;
        RECT 340.950 404.400 403.050 405.600 ;
        RECT 340.950 403.950 343.050 404.400 ;
        RECT 400.950 403.950 403.050 404.400 ;
        RECT 406.950 405.600 409.050 406.050 ;
        RECT 448.950 405.600 451.050 406.050 ;
        RECT 406.950 404.400 451.050 405.600 ;
        RECT 406.950 403.950 409.050 404.400 ;
        RECT 448.950 403.950 451.050 404.400 ;
        RECT 508.950 405.600 511.050 406.050 ;
        RECT 523.950 405.600 526.050 406.050 ;
        RECT 508.950 404.400 526.050 405.600 ;
        RECT 508.950 403.950 511.050 404.400 ;
        RECT 523.950 403.950 526.050 404.400 ;
        RECT 613.950 405.600 616.050 406.050 ;
        RECT 712.950 405.600 715.050 406.050 ;
        RECT 613.950 404.400 715.050 405.600 ;
        RECT 613.950 403.950 616.050 404.400 ;
        RECT 712.950 403.950 715.050 404.400 ;
        RECT 85.950 402.600 88.050 403.050 ;
        RECT 97.950 402.600 100.050 403.050 ;
        RECT 85.950 401.400 100.050 402.600 ;
        RECT 85.950 400.950 88.050 401.400 ;
        RECT 97.950 400.950 100.050 401.400 ;
        RECT 133.950 402.600 136.050 403.050 ;
        RECT 151.950 402.600 154.050 403.050 ;
        RECT 199.950 402.600 202.050 403.050 ;
        RECT 133.950 401.400 202.050 402.600 ;
        RECT 133.950 400.950 136.050 401.400 ;
        RECT 151.950 400.950 154.050 401.400 ;
        RECT 199.950 400.950 202.050 401.400 ;
        RECT 229.950 402.600 232.050 403.050 ;
        RECT 271.950 402.600 274.050 403.050 ;
        RECT 229.950 401.400 274.050 402.600 ;
        RECT 229.950 400.950 232.050 401.400 ;
        RECT 271.950 400.950 274.050 401.400 ;
        RECT 424.950 402.600 427.050 403.050 ;
        RECT 472.950 402.600 475.050 403.050 ;
        RECT 610.950 402.600 613.050 403.050 ;
        RECT 424.950 401.400 613.050 402.600 ;
        RECT 424.950 400.950 427.050 401.400 ;
        RECT 472.950 400.950 475.050 401.400 ;
        RECT 610.950 400.950 613.050 401.400 ;
        RECT 658.950 402.600 661.050 403.050 ;
        RECT 691.950 402.600 694.050 403.050 ;
        RECT 703.950 402.600 706.050 403.050 ;
        RECT 658.950 401.400 706.050 402.600 ;
        RECT 658.950 400.950 661.050 401.400 ;
        RECT 691.950 400.950 694.050 401.400 ;
        RECT 703.950 400.950 706.050 401.400 ;
        RECT 529.950 399.600 532.050 400.050 ;
        RECT 532.950 399.600 535.050 400.050 ;
        RECT 619.950 399.600 622.050 400.050 ;
        RECT 643.950 399.600 646.050 400.050 ;
        RECT 529.950 398.400 646.050 399.600 ;
        RECT 529.950 397.950 532.050 398.400 ;
        RECT 532.950 397.950 535.050 398.400 ;
        RECT 619.950 397.950 622.050 398.400 ;
        RECT 643.950 397.950 646.050 398.400 ;
        RECT 448.950 396.600 451.050 397.050 ;
        RECT 562.950 396.600 565.050 397.050 ;
        RECT 448.950 395.400 565.050 396.600 ;
        RECT 448.950 394.950 451.050 395.400 ;
        RECT 562.950 394.950 565.050 395.400 ;
        RECT 604.950 396.600 607.050 397.050 ;
        RECT 610.950 396.600 613.050 397.050 ;
        RECT 667.950 396.600 670.050 397.050 ;
        RECT 604.950 395.400 670.050 396.600 ;
        RECT 604.950 394.950 607.050 395.400 ;
        RECT 610.950 394.950 613.050 395.400 ;
        RECT 667.950 394.950 670.050 395.400 ;
        RECT 745.950 396.600 748.050 397.050 ;
        RECT 754.950 396.600 757.050 397.050 ;
        RECT 745.950 395.400 757.050 396.600 ;
        RECT 745.950 394.950 748.050 395.400 ;
        RECT 754.950 394.950 757.050 395.400 ;
        RECT 757.950 396.600 760.050 397.050 ;
        RECT 760.950 396.600 763.050 397.050 ;
        RECT 811.950 396.600 814.050 397.050 ;
        RECT 757.950 395.400 814.050 396.600 ;
        RECT 757.950 394.950 760.050 395.400 ;
        RECT 760.950 394.950 763.050 395.400 ;
        RECT 811.950 394.950 814.050 395.400 ;
        RECT 70.950 393.600 73.050 394.050 ;
        RECT 109.950 393.600 112.050 394.050 ;
        RECT 70.950 392.400 112.050 393.600 ;
        RECT 70.950 391.950 73.050 392.400 ;
        RECT 109.950 391.950 112.050 392.400 ;
        RECT 118.950 393.600 121.050 394.050 ;
        RECT 124.950 393.600 127.050 394.050 ;
        RECT 175.950 393.600 178.050 394.050 ;
        RECT 214.950 393.600 217.050 394.050 ;
        RECT 118.950 392.400 217.050 393.600 ;
        RECT 118.950 391.950 121.050 392.400 ;
        RECT 124.950 391.950 127.050 392.400 ;
        RECT 175.950 391.950 178.050 392.400 ;
        RECT 214.950 391.950 217.050 392.400 ;
        RECT 508.950 393.600 511.050 394.050 ;
        RECT 535.950 393.600 538.050 394.050 ;
        RECT 562.950 393.600 565.050 394.050 ;
        RECT 568.950 393.600 571.050 394.050 ;
        RECT 589.950 393.600 592.050 394.050 ;
        RECT 592.950 393.600 595.050 394.050 ;
        RECT 616.950 393.600 619.050 394.050 ;
        RECT 622.950 393.600 625.050 394.050 ;
        RECT 508.950 392.400 625.050 393.600 ;
        RECT 508.950 391.950 511.050 392.400 ;
        RECT 535.950 391.950 538.050 392.400 ;
        RECT 562.950 391.950 565.050 392.400 ;
        RECT 568.950 391.950 571.050 392.400 ;
        RECT 589.950 391.950 592.050 392.400 ;
        RECT 592.950 391.950 595.050 392.400 ;
        RECT 616.950 391.950 619.050 392.400 ;
        RECT 622.950 391.950 625.050 392.400 ;
        RECT 73.950 390.600 76.050 391.050 ;
        RECT 106.950 390.600 109.050 391.050 ;
        RECT 73.950 389.400 109.050 390.600 ;
        RECT 73.950 388.950 76.050 389.400 ;
        RECT 106.950 388.950 109.050 389.400 ;
        RECT 274.950 390.600 277.050 391.050 ;
        RECT 487.950 390.600 490.050 391.050 ;
        RECT 274.950 389.400 490.050 390.600 ;
        RECT 274.950 388.950 277.050 389.400 ;
        RECT 487.950 388.950 490.050 389.400 ;
        RECT 490.950 390.600 493.050 391.050 ;
        RECT 502.950 390.600 505.050 391.050 ;
        RECT 490.950 389.400 505.050 390.600 ;
        RECT 490.950 388.950 493.050 389.400 ;
        RECT 502.950 388.950 505.050 389.400 ;
        RECT 556.950 390.600 559.050 391.050 ;
        RECT 574.950 390.600 577.050 391.050 ;
        RECT 625.950 390.600 628.050 391.050 ;
        RECT 556.950 389.400 628.050 390.600 ;
        RECT 556.950 388.950 559.050 389.400 ;
        RECT 574.950 388.950 577.050 389.400 ;
        RECT 625.950 388.950 628.050 389.400 ;
        RECT 664.950 390.600 667.050 391.050 ;
        RECT 682.950 390.600 685.050 391.050 ;
        RECT 664.950 389.400 685.050 390.600 ;
        RECT 664.950 388.950 667.050 389.400 ;
        RECT 682.950 388.950 685.050 389.400 ;
        RECT 778.950 390.600 781.050 391.050 ;
        RECT 808.950 390.600 811.050 391.050 ;
        RECT 778.950 389.400 811.050 390.600 ;
        RECT 778.950 388.950 781.050 389.400 ;
        RECT 808.950 388.950 811.050 389.400 ;
        RECT 34.950 387.600 37.050 388.050 ;
        RECT 64.950 387.600 67.050 388.050 ;
        RECT 34.950 386.400 67.050 387.600 ;
        RECT 34.950 385.950 37.050 386.400 ;
        RECT 64.950 385.950 67.050 386.400 ;
        RECT 76.950 387.600 79.050 388.050 ;
        RECT 103.950 387.600 106.050 388.050 ;
        RECT 76.950 386.400 106.050 387.600 ;
        RECT 76.950 385.950 79.050 386.400 ;
        RECT 103.950 385.950 106.050 386.400 ;
        RECT 136.950 387.600 139.050 388.050 ;
        RECT 163.950 387.600 166.050 388.050 ;
        RECT 136.950 386.400 166.050 387.600 ;
        RECT 136.950 385.950 139.050 386.400 ;
        RECT 163.950 385.950 166.050 386.400 ;
        RECT 253.950 387.600 256.050 388.050 ;
        RECT 319.950 387.600 322.050 388.050 ;
        RECT 253.950 386.400 322.050 387.600 ;
        RECT 253.950 385.950 256.050 386.400 ;
        RECT 319.950 385.950 322.050 386.400 ;
        RECT 406.950 387.600 409.050 388.050 ;
        RECT 418.950 387.600 421.050 388.050 ;
        RECT 406.950 386.400 421.050 387.600 ;
        RECT 406.950 385.950 409.050 386.400 ;
        RECT 418.950 385.950 421.050 386.400 ;
        RECT 421.950 387.600 424.050 388.050 ;
        RECT 427.950 387.600 430.050 388.050 ;
        RECT 421.950 386.400 430.050 387.600 ;
        RECT 421.950 385.950 424.050 386.400 ;
        RECT 427.950 385.950 430.050 386.400 ;
        RECT 460.950 387.600 463.050 388.050 ;
        RECT 484.950 387.600 487.050 388.050 ;
        RECT 460.950 386.400 487.050 387.600 ;
        RECT 460.950 385.950 463.050 386.400 ;
        RECT 484.950 385.950 487.050 386.400 ;
        RECT 499.950 387.600 502.050 388.050 ;
        RECT 526.950 387.600 529.050 388.050 ;
        RECT 499.950 386.400 529.050 387.600 ;
        RECT 499.950 385.950 502.050 386.400 ;
        RECT 526.950 385.950 529.050 386.400 ;
        RECT 577.950 387.600 580.050 388.050 ;
        RECT 583.950 387.600 586.050 388.050 ;
        RECT 577.950 386.400 586.050 387.600 ;
        RECT 577.950 385.950 580.050 386.400 ;
        RECT 583.950 385.950 586.050 386.400 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 676.950 387.600 679.050 388.050 ;
        RECT 706.950 387.600 709.050 388.050 ;
        RECT 676.950 386.400 709.050 387.600 ;
        RECT 676.950 385.950 679.050 386.400 ;
        RECT 706.950 385.950 709.050 386.400 ;
        RECT 724.950 387.600 727.050 388.050 ;
        RECT 730.950 387.600 733.050 388.050 ;
        RECT 724.950 386.400 733.050 387.600 ;
        RECT 724.950 385.950 727.050 386.400 ;
        RECT 730.950 385.950 733.050 386.400 ;
        RECT 736.950 387.600 739.050 388.050 ;
        RECT 739.950 387.600 742.050 388.050 ;
        RECT 748.950 387.600 751.050 388.050 ;
        RECT 736.950 386.400 751.050 387.600 ;
        RECT 736.950 385.950 739.050 386.400 ;
        RECT 739.950 385.950 742.050 386.400 ;
        RECT 748.950 385.950 751.050 386.400 ;
        RECT 754.950 387.600 757.050 388.050 ;
        RECT 787.950 387.600 790.050 388.050 ;
        RECT 838.950 387.600 841.050 388.050 ;
        RECT 862.950 387.600 865.050 388.050 ;
        RECT 754.950 386.400 865.050 387.600 ;
        RECT 754.950 385.950 757.050 386.400 ;
        RECT 787.950 385.950 790.050 386.400 ;
        RECT 838.950 385.950 841.050 386.400 ;
        RECT 862.950 385.950 865.050 386.400 ;
        RECT 88.950 384.600 91.050 385.050 ;
        RECT 74.400 383.400 91.050 384.600 ;
        RECT 74.400 382.050 75.600 383.400 ;
        RECT 88.950 382.950 91.050 383.400 ;
        RECT 97.950 384.600 100.050 385.050 ;
        RECT 145.950 384.600 148.050 385.050 ;
        RECT 97.950 383.400 148.050 384.600 ;
        RECT 97.950 382.950 100.050 383.400 ;
        RECT 145.950 382.950 148.050 383.400 ;
        RECT 190.950 384.600 193.050 385.050 ;
        RECT 220.950 384.600 223.050 385.050 ;
        RECT 190.950 383.400 223.050 384.600 ;
        RECT 190.950 382.950 193.050 383.400 ;
        RECT 220.950 382.950 223.050 383.400 ;
        RECT 223.950 384.600 226.050 385.050 ;
        RECT 229.950 384.600 232.050 385.050 ;
        RECT 223.950 383.400 232.050 384.600 ;
        RECT 223.950 382.950 226.050 383.400 ;
        RECT 229.950 382.950 232.050 383.400 ;
        RECT 262.950 384.600 265.050 385.050 ;
        RECT 271.950 384.600 274.050 385.050 ;
        RECT 262.950 383.400 274.050 384.600 ;
        RECT 262.950 382.950 265.050 383.400 ;
        RECT 271.950 382.950 274.050 383.400 ;
        RECT 280.950 384.600 283.050 385.050 ;
        RECT 286.950 384.600 289.050 385.050 ;
        RECT 280.950 383.400 289.050 384.600 ;
        RECT 280.950 382.950 283.050 383.400 ;
        RECT 286.950 382.950 289.050 383.400 ;
        RECT 337.950 384.600 340.050 385.050 ;
        RECT 358.950 384.600 361.050 385.050 ;
        RECT 337.950 383.400 361.050 384.600 ;
        RECT 337.950 382.950 340.050 383.400 ;
        RECT 358.950 382.950 361.050 383.400 ;
        RECT 367.950 384.600 370.050 385.050 ;
        RECT 451.950 384.600 454.050 385.050 ;
        RECT 367.950 383.400 454.050 384.600 ;
        RECT 367.950 382.950 370.050 383.400 ;
        RECT 451.950 382.950 454.050 383.400 ;
        RECT 595.950 384.600 598.050 385.050 ;
        RECT 616.950 384.600 619.050 385.050 ;
        RECT 595.950 383.400 619.050 384.600 ;
        RECT 595.950 382.950 598.050 383.400 ;
        RECT 616.950 382.950 619.050 383.400 ;
        RECT 625.950 384.600 628.050 385.050 ;
        RECT 641.400 384.600 642.600 385.950 ;
        RECT 688.950 384.600 691.050 385.050 ;
        RECT 625.950 383.400 691.050 384.600 ;
        RECT 625.950 382.950 628.050 383.400 ;
        RECT 688.950 382.950 691.050 383.400 ;
        RECT 700.950 384.600 703.050 385.050 ;
        RECT 754.950 384.600 757.050 385.050 ;
        RECT 700.950 383.400 757.050 384.600 ;
        RECT 700.950 382.950 703.050 383.400 ;
        RECT 754.950 382.950 757.050 383.400 ;
        RECT 760.950 384.600 763.050 385.050 ;
        RECT 778.950 384.600 781.050 385.050 ;
        RECT 760.950 383.400 781.050 384.600 ;
        RECT 760.950 382.950 763.050 383.400 ;
        RECT 778.950 382.950 781.050 383.400 ;
        RECT 823.950 384.600 826.050 385.050 ;
        RECT 868.950 384.600 871.050 385.050 ;
        RECT 823.950 383.400 871.050 384.600 ;
        RECT 823.950 382.950 826.050 383.400 ;
        RECT 868.950 382.950 871.050 383.400 ;
        RECT 49.950 381.600 52.050 382.050 ;
        RECT 67.950 381.600 70.050 382.050 ;
        RECT 49.950 380.400 70.050 381.600 ;
        RECT 49.950 379.950 52.050 380.400 ;
        RECT 67.950 379.950 70.050 380.400 ;
        RECT 73.950 379.950 76.050 382.050 ;
        RECT 109.950 381.600 112.050 382.050 ;
        RECT 187.950 381.600 190.050 382.050 ;
        RECT 109.950 380.400 190.050 381.600 ;
        RECT 109.950 379.950 112.050 380.400 ;
        RECT 187.950 379.950 190.050 380.400 ;
        RECT 193.950 381.600 196.050 382.050 ;
        RECT 208.950 381.600 211.050 382.050 ;
        RECT 193.950 380.400 211.050 381.600 ;
        RECT 193.950 379.950 196.050 380.400 ;
        RECT 208.950 379.950 211.050 380.400 ;
        RECT 298.950 381.600 301.050 382.050 ;
        RECT 322.950 381.600 325.050 382.050 ;
        RECT 298.950 380.400 325.050 381.600 ;
        RECT 298.950 379.950 301.050 380.400 ;
        RECT 322.950 379.950 325.050 380.400 ;
        RECT 337.950 381.600 340.050 382.050 ;
        RECT 343.950 381.600 346.050 382.050 ;
        RECT 355.950 381.600 358.050 382.050 ;
        RECT 379.950 381.600 382.050 382.050 ;
        RECT 409.950 381.600 412.050 382.050 ;
        RECT 424.950 381.600 427.050 382.050 ;
        RECT 337.950 380.400 358.050 381.600 ;
        RECT 337.950 379.950 340.050 380.400 ;
        RECT 343.950 379.950 346.050 380.400 ;
        RECT 355.950 379.950 358.050 380.400 ;
        RECT 359.400 380.400 427.050 381.600 ;
        RECT 31.950 378.600 34.050 379.050 ;
        RECT 46.950 378.600 49.050 379.050 ;
        RECT 70.950 378.600 73.050 379.050 ;
        RECT 82.950 378.600 85.050 379.050 ;
        RECT 31.950 377.400 85.050 378.600 ;
        RECT 31.950 376.950 34.050 377.400 ;
        RECT 46.950 376.950 49.050 377.400 ;
        RECT 70.950 376.950 73.050 377.400 ;
        RECT 82.950 376.950 85.050 377.400 ;
        RECT 100.950 378.600 103.050 379.050 ;
        RECT 103.950 378.600 106.050 379.050 ;
        RECT 133.950 378.600 136.050 379.050 ;
        RECT 148.950 378.600 151.050 379.050 ;
        RECT 100.950 377.400 151.050 378.600 ;
        RECT 100.950 376.950 103.050 377.400 ;
        RECT 103.950 376.950 106.050 377.400 ;
        RECT 133.950 376.950 136.050 377.400 ;
        RECT 148.950 376.950 151.050 377.400 ;
        RECT 202.950 378.600 205.050 379.050 ;
        RECT 211.950 378.600 214.050 379.050 ;
        RECT 256.950 378.600 259.050 379.050 ;
        RECT 262.950 378.600 265.050 379.050 ;
        RECT 202.950 377.400 265.050 378.600 ;
        RECT 202.950 376.950 205.050 377.400 ;
        RECT 211.950 376.950 214.050 377.400 ;
        RECT 256.950 376.950 259.050 377.400 ;
        RECT 262.950 376.950 265.050 377.400 ;
        RECT 265.950 378.600 268.050 379.050 ;
        RECT 277.950 378.600 280.050 379.050 ;
        RECT 265.950 377.400 280.050 378.600 ;
        RECT 265.950 376.950 268.050 377.400 ;
        RECT 277.950 376.950 280.050 377.400 ;
        RECT 286.950 378.600 289.050 379.050 ;
        RECT 301.950 378.600 304.050 379.050 ;
        RECT 286.950 377.400 304.050 378.600 ;
        RECT 286.950 376.950 289.050 377.400 ;
        RECT 301.950 376.950 304.050 377.400 ;
        RECT 307.950 378.600 310.050 379.050 ;
        RECT 316.950 378.600 319.050 379.050 ;
        RECT 307.950 377.400 319.050 378.600 ;
        RECT 307.950 376.950 310.050 377.400 ;
        RECT 316.950 376.950 319.050 377.400 ;
        RECT 334.950 378.600 337.050 379.050 ;
        RECT 340.950 378.600 343.050 379.050 ;
        RECT 359.400 378.600 360.600 380.400 ;
        RECT 379.950 379.950 382.050 380.400 ;
        RECT 409.950 379.950 412.050 380.400 ;
        RECT 424.950 379.950 427.050 380.400 ;
        RECT 439.950 381.600 442.050 382.050 ;
        RECT 577.950 381.600 580.050 382.050 ;
        RECT 439.950 380.400 580.050 381.600 ;
        RECT 439.950 379.950 442.050 380.400 ;
        RECT 577.950 379.950 580.050 380.400 ;
        RECT 580.950 381.600 583.050 382.050 ;
        RECT 637.950 381.600 640.050 382.050 ;
        RECT 580.950 380.400 640.050 381.600 ;
        RECT 580.950 379.950 583.050 380.400 ;
        RECT 637.950 379.950 640.050 380.400 ;
        RECT 658.950 381.600 661.050 382.050 ;
        RECT 673.950 381.600 676.050 382.050 ;
        RECT 658.950 380.400 676.050 381.600 ;
        RECT 658.950 379.950 661.050 380.400 ;
        RECT 673.950 379.950 676.050 380.400 ;
        RECT 769.950 381.600 772.050 382.050 ;
        RECT 826.950 381.600 829.050 382.050 ;
        RECT 769.950 380.400 829.050 381.600 ;
        RECT 769.950 379.950 772.050 380.400 ;
        RECT 826.950 379.950 829.050 380.400 ;
        RECT 832.950 381.600 835.050 382.050 ;
        RECT 841.950 381.600 844.050 382.050 ;
        RECT 832.950 380.400 844.050 381.600 ;
        RECT 832.950 379.950 835.050 380.400 ;
        RECT 841.950 379.950 844.050 380.400 ;
        RECT 334.950 377.400 360.600 378.600 ;
        RECT 370.950 378.600 373.050 379.050 ;
        RECT 463.950 378.600 466.050 379.050 ;
        RECT 370.950 377.400 466.050 378.600 ;
        RECT 334.950 376.950 337.050 377.400 ;
        RECT 340.950 376.950 343.050 377.400 ;
        RECT 370.950 376.950 373.050 377.400 ;
        RECT 463.950 376.950 466.050 377.400 ;
        RECT 589.950 378.600 592.050 379.050 ;
        RECT 598.950 378.600 601.050 379.050 ;
        RECT 589.950 377.400 601.050 378.600 ;
        RECT 589.950 376.950 592.050 377.400 ;
        RECT 598.950 376.950 601.050 377.400 ;
        RECT 604.950 378.600 607.050 379.050 ;
        RECT 625.950 378.600 628.050 379.050 ;
        RECT 604.950 377.400 628.050 378.600 ;
        RECT 604.950 376.950 607.050 377.400 ;
        RECT 625.950 376.950 628.050 377.400 ;
        RECT 637.950 378.600 640.050 379.050 ;
        RECT 679.950 378.600 682.050 379.050 ;
        RECT 637.950 377.400 682.050 378.600 ;
        RECT 637.950 376.950 640.050 377.400 ;
        RECT 679.950 376.950 682.050 377.400 ;
        RECT 730.950 378.600 733.050 379.050 ;
        RECT 817.950 378.600 820.050 379.050 ;
        RECT 730.950 377.400 820.050 378.600 ;
        RECT 730.950 376.950 733.050 377.400 ;
        RECT 817.950 376.950 820.050 377.400 ;
        RECT 46.950 375.600 49.050 376.050 ;
        RECT 139.950 375.600 142.050 376.050 ;
        RECT 676.950 375.600 679.050 376.050 ;
        RECT 46.950 374.400 679.050 375.600 ;
        RECT 46.950 373.950 49.050 374.400 ;
        RECT 139.950 373.950 142.050 374.400 ;
        RECT 676.950 373.950 679.050 374.400 ;
        RECT 13.950 372.600 16.050 373.050 ;
        RECT 112.950 372.600 115.050 373.050 ;
        RECT 13.950 371.400 115.050 372.600 ;
        RECT 13.950 370.950 16.050 371.400 ;
        RECT 112.950 370.950 115.050 371.400 ;
        RECT 148.950 372.600 151.050 373.050 ;
        RECT 166.950 372.600 169.050 373.050 ;
        RECT 202.950 372.600 205.050 373.050 ;
        RECT 217.950 372.600 220.050 373.050 ;
        RECT 250.950 372.600 253.050 373.050 ;
        RECT 148.950 371.400 253.050 372.600 ;
        RECT 148.950 370.950 151.050 371.400 ;
        RECT 166.950 370.950 169.050 371.400 ;
        RECT 202.950 370.950 205.050 371.400 ;
        RECT 217.950 370.950 220.050 371.400 ;
        RECT 250.950 370.950 253.050 371.400 ;
        RECT 322.950 372.600 325.050 373.050 ;
        RECT 328.950 372.600 331.050 373.050 ;
        RECT 322.950 371.400 331.050 372.600 ;
        RECT 322.950 370.950 325.050 371.400 ;
        RECT 328.950 370.950 331.050 371.400 ;
        RECT 394.950 372.600 397.050 373.050 ;
        RECT 550.950 372.600 553.050 373.050 ;
        RECT 394.950 371.400 553.050 372.600 ;
        RECT 394.950 370.950 397.050 371.400 ;
        RECT 550.950 370.950 553.050 371.400 ;
        RECT 28.950 369.600 31.050 370.050 ;
        RECT 37.950 369.600 40.050 370.050 ;
        RECT 28.950 368.400 40.050 369.600 ;
        RECT 28.950 367.950 31.050 368.400 ;
        RECT 37.950 367.950 40.050 368.400 ;
        RECT 142.950 369.600 145.050 370.050 ;
        RECT 211.950 369.600 214.050 370.050 ;
        RECT 142.950 368.400 214.050 369.600 ;
        RECT 142.950 367.950 145.050 368.400 ;
        RECT 211.950 367.950 214.050 368.400 ;
        RECT 334.950 369.600 337.050 370.050 ;
        RECT 421.950 369.600 424.050 370.050 ;
        RECT 454.950 369.600 457.050 370.050 ;
        RECT 334.950 368.400 457.050 369.600 ;
        RECT 334.950 367.950 337.050 368.400 ;
        RECT 421.950 367.950 424.050 368.400 ;
        RECT 454.950 367.950 457.050 368.400 ;
        RECT 310.950 366.600 313.050 367.050 ;
        RECT 361.950 366.600 364.050 367.050 ;
        RECT 385.950 366.600 388.050 367.050 ;
        RECT 310.950 365.400 388.050 366.600 ;
        RECT 310.950 364.950 313.050 365.400 ;
        RECT 361.950 364.950 364.050 365.400 ;
        RECT 385.950 364.950 388.050 365.400 ;
        RECT 412.950 366.600 415.050 367.050 ;
        RECT 430.950 366.600 433.050 367.050 ;
        RECT 412.950 365.400 433.050 366.600 ;
        RECT 412.950 364.950 415.050 365.400 ;
        RECT 430.950 364.950 433.050 365.400 ;
        RECT 442.950 366.600 445.050 367.050 ;
        RECT 475.950 366.600 478.050 367.050 ;
        RECT 442.950 365.400 478.050 366.600 ;
        RECT 442.950 364.950 445.050 365.400 ;
        RECT 475.950 364.950 478.050 365.400 ;
        RECT 181.950 363.600 184.050 364.050 ;
        RECT 205.950 363.600 208.050 364.050 ;
        RECT 214.950 363.600 217.050 364.050 ;
        RECT 226.950 363.600 229.050 364.050 ;
        RECT 268.950 363.600 271.050 364.050 ;
        RECT 295.950 363.600 298.050 364.050 ;
        RECT 181.950 362.400 298.050 363.600 ;
        RECT 181.950 361.950 184.050 362.400 ;
        RECT 205.950 361.950 208.050 362.400 ;
        RECT 214.950 361.950 217.050 362.400 ;
        RECT 226.950 361.950 229.050 362.400 ;
        RECT 268.950 361.950 271.050 362.400 ;
        RECT 295.950 361.950 298.050 362.400 ;
        RECT 304.950 360.600 307.050 361.050 ;
        RECT 358.950 360.600 361.050 361.050 ;
        RECT 304.950 359.400 361.050 360.600 ;
        RECT 304.950 358.950 307.050 359.400 ;
        RECT 358.950 358.950 361.050 359.400 ;
        RECT 457.950 360.600 460.050 361.050 ;
        RECT 469.950 360.600 472.050 361.050 ;
        RECT 457.950 359.400 472.050 360.600 ;
        RECT 457.950 358.950 460.050 359.400 ;
        RECT 469.950 358.950 472.050 359.400 ;
        RECT 235.950 357.600 238.050 358.050 ;
        RECT 448.950 357.600 451.050 358.050 ;
        RECT 235.950 356.400 451.050 357.600 ;
        RECT 235.950 355.950 238.050 356.400 ;
        RECT 448.950 355.950 451.050 356.400 ;
        RECT 814.950 357.600 817.050 358.050 ;
        RECT 820.950 357.600 823.050 358.050 ;
        RECT 814.950 356.400 823.050 357.600 ;
        RECT 814.950 355.950 817.050 356.400 ;
        RECT 820.950 355.950 823.050 356.400 ;
        RECT 352.950 354.600 355.050 355.050 ;
        RECT 394.950 354.600 397.050 355.050 ;
        RECT 352.950 353.400 397.050 354.600 ;
        RECT 352.950 352.950 355.050 353.400 ;
        RECT 394.950 352.950 397.050 353.400 ;
        RECT 103.950 351.600 106.050 352.050 ;
        RECT 169.950 351.600 172.050 352.050 ;
        RECT 103.950 350.400 172.050 351.600 ;
        RECT 103.950 349.950 106.050 350.400 ;
        RECT 169.950 349.950 172.050 350.400 ;
        RECT 223.950 351.600 226.050 352.050 ;
        RECT 424.950 351.600 427.050 352.050 ;
        RECT 523.950 351.600 526.050 352.050 ;
        RECT 556.950 351.600 559.050 352.050 ;
        RECT 223.950 350.400 427.050 351.600 ;
        RECT 223.950 349.950 226.050 350.400 ;
        RECT 424.950 349.950 427.050 350.400 ;
        RECT 497.400 350.400 559.050 351.600 ;
        RECT 55.950 348.600 58.050 349.050 ;
        RECT 67.950 348.600 70.050 349.050 ;
        RECT 55.950 347.400 70.050 348.600 ;
        RECT 55.950 346.950 58.050 347.400 ;
        RECT 67.950 346.950 70.050 347.400 ;
        RECT 91.950 348.600 94.050 349.050 ;
        RECT 133.950 348.600 136.050 349.050 ;
        RECT 91.950 347.400 136.050 348.600 ;
        RECT 91.950 346.950 94.050 347.400 ;
        RECT 133.950 346.950 136.050 347.400 ;
        RECT 136.950 348.600 139.050 349.050 ;
        RECT 229.950 348.600 232.050 349.050 ;
        RECT 136.950 347.400 232.050 348.600 ;
        RECT 136.950 346.950 139.050 347.400 ;
        RECT 229.950 346.950 232.050 347.400 ;
        RECT 259.950 348.600 262.050 349.050 ;
        RECT 346.950 348.600 349.050 349.050 ;
        RECT 349.950 348.600 352.050 349.050 ;
        RECT 259.950 347.400 352.050 348.600 ;
        RECT 259.950 346.950 262.050 347.400 ;
        RECT 346.950 346.950 349.050 347.400 ;
        RECT 349.950 346.950 352.050 347.400 ;
        RECT 385.950 348.600 388.050 349.050 ;
        RECT 472.950 348.600 475.050 349.050 ;
        RECT 497.400 348.600 498.600 350.400 ;
        RECT 523.950 349.950 526.050 350.400 ;
        RECT 556.950 349.950 559.050 350.400 ;
        RECT 592.950 351.600 595.050 352.050 ;
        RECT 733.950 351.600 736.050 352.050 ;
        RECT 592.950 350.400 736.050 351.600 ;
        RECT 592.950 349.950 595.050 350.400 ;
        RECT 733.950 349.950 736.050 350.400 ;
        RECT 775.950 351.600 778.050 352.050 ;
        RECT 829.950 351.600 832.050 352.050 ;
        RECT 775.950 350.400 832.050 351.600 ;
        RECT 775.950 349.950 778.050 350.400 ;
        RECT 829.950 349.950 832.050 350.400 ;
        RECT 385.950 347.400 498.600 348.600 ;
        RECT 499.950 348.600 502.050 349.050 ;
        RECT 511.950 348.600 514.050 349.050 ;
        RECT 499.950 347.400 514.050 348.600 ;
        RECT 385.950 346.950 388.050 347.400 ;
        RECT 472.950 346.950 475.050 347.400 ;
        RECT 499.950 346.950 502.050 347.400 ;
        RECT 511.950 346.950 514.050 347.400 ;
        RECT 580.950 348.600 583.050 349.050 ;
        RECT 634.950 348.600 637.050 349.050 ;
        RECT 580.950 347.400 637.050 348.600 ;
        RECT 580.950 346.950 583.050 347.400 ;
        RECT 634.950 346.950 637.050 347.400 ;
        RECT 694.950 348.600 697.050 349.050 ;
        RECT 754.950 348.600 757.050 349.050 ;
        RECT 694.950 347.400 757.050 348.600 ;
        RECT 694.950 346.950 697.050 347.400 ;
        RECT 754.950 346.950 757.050 347.400 ;
        RECT 763.950 348.600 766.050 349.050 ;
        RECT 799.950 348.600 802.050 349.050 ;
        RECT 823.950 348.600 826.050 349.050 ;
        RECT 763.950 347.400 798.600 348.600 ;
        RECT 763.950 346.950 766.050 347.400 ;
        RECT 40.950 345.600 43.050 346.050 ;
        RECT 73.950 345.600 76.050 346.050 ;
        RECT 40.950 344.400 76.050 345.600 ;
        RECT 40.950 343.950 43.050 344.400 ;
        RECT 73.950 343.950 76.050 344.400 ;
        RECT 109.950 345.600 112.050 346.050 ;
        RECT 154.950 345.600 157.050 346.050 ;
        RECT 109.950 344.400 157.050 345.600 ;
        RECT 109.950 343.950 112.050 344.400 ;
        RECT 154.950 343.950 157.050 344.400 ;
        RECT 169.950 345.600 172.050 346.050 ;
        RECT 175.950 345.600 178.050 346.050 ;
        RECT 169.950 344.400 178.050 345.600 ;
        RECT 169.950 343.950 172.050 344.400 ;
        RECT 175.950 343.950 178.050 344.400 ;
        RECT 250.950 345.600 253.050 346.050 ;
        RECT 259.950 345.600 262.050 346.050 ;
        RECT 250.950 344.400 262.050 345.600 ;
        RECT 250.950 343.950 253.050 344.400 ;
        RECT 259.950 343.950 262.050 344.400 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 367.950 345.600 370.050 346.050 ;
        RECT 373.950 345.600 376.050 346.050 ;
        RECT 355.950 344.400 376.050 345.600 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 367.950 343.950 370.050 344.400 ;
        RECT 373.950 343.950 376.050 344.400 ;
        RECT 433.950 345.600 436.050 346.050 ;
        RECT 454.950 345.600 457.050 346.050 ;
        RECT 493.950 345.600 496.050 346.050 ;
        RECT 625.950 345.600 628.050 346.050 ;
        RECT 640.950 345.600 643.050 346.050 ;
        RECT 433.950 344.400 438.600 345.600 ;
        RECT 433.950 343.950 436.050 344.400 ;
        RECT 19.950 342.600 22.050 343.050 ;
        RECT 34.950 342.600 37.050 343.050 ;
        RECT 49.950 342.600 52.050 343.050 ;
        RECT 55.950 342.600 58.050 343.050 ;
        RECT 19.950 341.400 58.050 342.600 ;
        RECT 19.950 340.950 22.050 341.400 ;
        RECT 34.950 340.950 37.050 341.400 ;
        RECT 49.950 340.950 52.050 341.400 ;
        RECT 55.950 340.950 58.050 341.400 ;
        RECT 94.950 340.950 97.050 343.050 ;
        RECT 112.950 342.600 115.050 343.050 ;
        RECT 118.950 342.600 121.050 343.050 ;
        RECT 112.950 341.400 121.050 342.600 ;
        RECT 112.950 340.950 115.050 341.400 ;
        RECT 118.950 340.950 121.050 341.400 ;
        RECT 124.950 342.600 127.050 343.050 ;
        RECT 136.950 342.600 139.050 343.050 ;
        RECT 163.950 342.600 166.050 343.050 ;
        RECT 124.950 341.400 139.050 342.600 ;
        RECT 124.950 340.950 127.050 341.400 ;
        RECT 136.950 340.950 139.050 341.400 ;
        RECT 158.400 341.400 166.050 342.600 ;
        RECT 79.950 339.600 82.050 340.050 ;
        RECT 88.950 339.600 91.050 340.050 ;
        RECT 79.950 338.400 91.050 339.600 ;
        RECT 79.950 337.950 82.050 338.400 ;
        RECT 88.950 337.950 91.050 338.400 ;
        RECT 82.950 336.600 85.050 337.050 ;
        RECT 95.400 336.600 96.600 340.950 ;
        RECT 97.950 339.600 100.050 340.050 ;
        RECT 109.950 339.600 112.050 340.050 ;
        RECT 97.950 338.400 112.050 339.600 ;
        RECT 97.950 337.950 100.050 338.400 ;
        RECT 109.950 337.950 112.050 338.400 ;
        RECT 121.950 339.600 124.050 340.050 ;
        RECT 127.950 339.600 130.050 340.050 ;
        RECT 121.950 338.400 130.050 339.600 ;
        RECT 121.950 337.950 124.050 338.400 ;
        RECT 127.950 337.950 130.050 338.400 ;
        RECT 142.950 336.600 145.050 337.050 ;
        RECT 82.950 335.400 145.050 336.600 ;
        RECT 158.400 336.600 159.600 341.400 ;
        RECT 163.950 340.950 166.050 341.400 ;
        RECT 184.950 342.600 187.050 343.050 ;
        RECT 214.950 342.600 217.050 343.050 ;
        RECT 184.950 341.400 217.050 342.600 ;
        RECT 184.950 340.950 187.050 341.400 ;
        RECT 214.950 340.950 217.050 341.400 ;
        RECT 229.950 342.600 232.050 343.050 ;
        RECT 262.950 342.600 265.050 343.050 ;
        RECT 229.950 341.400 265.050 342.600 ;
        RECT 229.950 340.950 232.050 341.400 ;
        RECT 262.950 340.950 265.050 341.400 ;
        RECT 289.950 340.950 292.050 343.050 ;
        RECT 304.950 342.600 307.050 343.050 ;
        RECT 328.950 342.600 331.050 343.050 ;
        RECT 352.950 342.600 355.050 343.050 ;
        RECT 361.950 342.600 364.050 343.050 ;
        RECT 304.950 341.400 364.050 342.600 ;
        RECT 304.950 340.950 307.050 341.400 ;
        RECT 328.950 340.950 331.050 341.400 ;
        RECT 352.950 340.950 355.050 341.400 ;
        RECT 361.950 340.950 364.050 341.400 ;
        RECT 379.950 342.600 382.050 343.050 ;
        RECT 400.950 342.600 403.050 343.050 ;
        RECT 379.950 341.400 403.050 342.600 ;
        RECT 379.950 340.950 382.050 341.400 ;
        RECT 400.950 340.950 403.050 341.400 ;
        RECT 406.950 340.950 409.050 343.050 ;
        RECT 160.950 339.600 163.050 340.050 ;
        RECT 196.950 339.600 199.050 340.050 ;
        RECT 160.950 338.400 199.050 339.600 ;
        RECT 160.950 337.950 163.050 338.400 ;
        RECT 196.950 337.950 199.050 338.400 ;
        RECT 226.950 339.600 229.050 340.050 ;
        RECT 290.400 339.600 291.600 340.950 ;
        RECT 313.950 339.600 316.050 340.050 ;
        RECT 337.950 339.600 340.050 340.050 ;
        RECT 340.950 339.600 343.050 340.050 ;
        RECT 226.950 338.400 303.600 339.600 ;
        RECT 226.950 337.950 229.050 338.400 ;
        RECT 298.950 336.600 301.050 337.050 ;
        RECT 158.400 335.400 301.050 336.600 ;
        RECT 302.400 336.600 303.600 338.400 ;
        RECT 313.950 338.400 343.050 339.600 ;
        RECT 313.950 337.950 316.050 338.400 ;
        RECT 337.950 337.950 340.050 338.400 ;
        RECT 340.950 337.950 343.050 338.400 ;
        RECT 346.950 339.600 349.050 340.050 ;
        RECT 376.950 339.600 379.050 340.050 ;
        RECT 346.950 338.400 379.050 339.600 ;
        RECT 346.950 337.950 349.050 338.400 ;
        RECT 376.950 337.950 379.050 338.400 ;
        RECT 325.950 336.600 328.050 337.050 ;
        RECT 302.400 335.400 328.050 336.600 ;
        RECT 82.950 334.950 85.050 335.400 ;
        RECT 142.950 334.950 145.050 335.400 ;
        RECT 298.950 334.950 301.050 335.400 ;
        RECT 325.950 334.950 328.050 335.400 ;
        RECT 58.950 333.600 61.050 334.050 ;
        RECT 115.950 333.600 118.050 334.050 ;
        RECT 58.950 332.400 118.050 333.600 ;
        RECT 58.950 331.950 61.050 332.400 ;
        RECT 115.950 331.950 118.050 332.400 ;
        RECT 151.950 333.600 154.050 334.050 ;
        RECT 172.950 333.600 175.050 334.050 ;
        RECT 151.950 332.400 175.050 333.600 ;
        RECT 151.950 331.950 154.050 332.400 ;
        RECT 172.950 331.950 175.050 332.400 ;
        RECT 178.950 333.600 181.050 334.050 ;
        RECT 217.950 333.600 220.050 334.050 ;
        RECT 178.950 332.400 220.050 333.600 ;
        RECT 178.950 331.950 181.050 332.400 ;
        RECT 217.950 331.950 220.050 332.400 ;
        RECT 268.950 333.600 271.050 334.050 ;
        RECT 277.950 333.600 280.050 334.050 ;
        RECT 379.950 333.600 382.050 334.050 ;
        RECT 268.950 332.400 382.050 333.600 ;
        RECT 407.400 333.600 408.600 340.950 ;
        RECT 437.400 340.050 438.600 344.400 ;
        RECT 454.950 344.400 643.050 345.600 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 493.950 343.950 496.050 344.400 ;
        RECT 625.950 343.950 628.050 344.400 ;
        RECT 640.950 343.950 643.050 344.400 ;
        RECT 652.950 345.600 655.050 346.050 ;
        RECT 679.950 345.600 682.050 346.050 ;
        RECT 652.950 344.400 682.050 345.600 ;
        RECT 652.950 343.950 655.050 344.400 ;
        RECT 679.950 343.950 682.050 344.400 ;
        RECT 721.950 345.600 724.050 346.050 ;
        RECT 736.950 345.600 739.050 346.050 ;
        RECT 721.950 344.400 739.050 345.600 ;
        RECT 721.950 343.950 724.050 344.400 ;
        RECT 736.950 343.950 739.050 344.400 ;
        RECT 748.950 345.600 751.050 346.050 ;
        RECT 757.950 345.600 760.050 346.050 ;
        RECT 778.950 345.600 781.050 346.050 ;
        RECT 748.950 344.400 760.050 345.600 ;
        RECT 748.950 343.950 751.050 344.400 ;
        RECT 757.950 343.950 760.050 344.400 ;
        RECT 770.400 344.400 781.050 345.600 ;
        RECT 797.400 345.600 798.600 347.400 ;
        RECT 799.950 347.400 826.050 348.600 ;
        RECT 799.950 346.950 802.050 347.400 ;
        RECT 823.950 346.950 826.050 347.400 ;
        RECT 817.950 345.600 820.050 346.050 ;
        RECT 835.950 345.600 838.050 346.050 ;
        RECT 797.400 344.400 838.050 345.600 ;
        RECT 457.950 342.600 460.050 343.050 ;
        RECT 490.950 342.600 493.050 343.050 ;
        RECT 457.950 341.400 493.050 342.600 ;
        RECT 457.950 340.950 460.050 341.400 ;
        RECT 490.950 340.950 493.050 341.400 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 553.950 342.600 556.050 343.050 ;
        RECT 559.950 342.600 562.050 343.050 ;
        RECT 553.950 341.400 562.050 342.600 ;
        RECT 553.950 340.950 556.050 341.400 ;
        RECT 559.950 340.950 562.050 341.400 ;
        RECT 574.950 342.600 577.050 343.050 ;
        RECT 586.950 342.600 589.050 343.050 ;
        RECT 592.950 342.600 595.050 343.050 ;
        RECT 574.950 341.400 595.050 342.600 ;
        RECT 574.950 340.950 577.050 341.400 ;
        RECT 586.950 340.950 589.050 341.400 ;
        RECT 592.950 340.950 595.050 341.400 ;
        RECT 661.950 342.600 664.050 343.050 ;
        RECT 682.950 342.600 685.050 343.050 ;
        RECT 661.950 341.400 685.050 342.600 ;
        RECT 661.950 340.950 664.050 341.400 ;
        RECT 682.950 340.950 685.050 341.400 ;
        RECT 727.950 342.600 730.050 343.050 ;
        RECT 739.950 342.600 742.050 343.050 ;
        RECT 727.950 341.400 742.050 342.600 ;
        RECT 727.950 340.950 730.050 341.400 ;
        RECT 739.950 340.950 742.050 341.400 ;
        RECT 745.950 342.600 748.050 343.050 ;
        RECT 770.400 342.600 771.600 344.400 ;
        RECT 778.950 343.950 781.050 344.400 ;
        RECT 817.950 343.950 820.050 344.400 ;
        RECT 835.950 343.950 838.050 344.400 ;
        RECT 856.950 345.600 859.050 346.050 ;
        RECT 865.950 345.600 868.050 346.050 ;
        RECT 856.950 344.400 868.050 345.600 ;
        RECT 856.950 343.950 859.050 344.400 ;
        RECT 865.950 343.950 868.050 344.400 ;
        RECT 745.950 341.400 771.600 342.600 ;
        RECT 772.950 342.600 775.050 343.050 ;
        RECT 781.950 342.600 784.050 343.050 ;
        RECT 772.950 341.400 784.050 342.600 ;
        RECT 745.950 340.950 748.050 341.400 ;
        RECT 772.950 340.950 775.050 341.400 ;
        RECT 781.950 340.950 784.050 341.400 ;
        RECT 841.950 342.600 844.050 343.050 ;
        RECT 847.950 342.600 850.050 343.050 ;
        RECT 841.950 341.400 850.050 342.600 ;
        RECT 841.950 340.950 844.050 341.400 ;
        RECT 847.950 340.950 850.050 341.400 ;
        RECT 850.950 342.600 853.050 343.050 ;
        RECT 856.950 342.600 859.050 343.050 ;
        RECT 850.950 341.400 859.050 342.600 ;
        RECT 850.950 340.950 853.050 341.400 ;
        RECT 856.950 340.950 859.050 341.400 ;
        RECT 436.950 337.950 439.050 340.050 ;
        RECT 445.950 339.600 448.050 340.050 ;
        RECT 460.950 339.600 463.050 340.050 ;
        RECT 445.950 338.400 463.050 339.600 ;
        RECT 445.950 337.950 448.050 338.400 ;
        RECT 460.950 337.950 463.050 338.400 ;
        RECT 466.950 339.600 469.050 340.050 ;
        RECT 478.950 339.600 481.050 340.050 ;
        RECT 514.950 339.600 517.050 340.050 ;
        RECT 530.400 339.600 531.600 340.950 ;
        RECT 466.950 338.400 531.600 339.600 ;
        RECT 544.950 339.600 547.050 340.050 ;
        RECT 577.950 339.600 580.050 340.050 ;
        RECT 595.950 339.600 598.050 340.050 ;
        RECT 544.950 338.400 598.050 339.600 ;
        RECT 466.950 337.950 469.050 338.400 ;
        RECT 478.950 337.950 481.050 338.400 ;
        RECT 514.950 337.950 517.050 338.400 ;
        RECT 544.950 337.950 547.050 338.400 ;
        RECT 577.950 337.950 580.050 338.400 ;
        RECT 595.950 337.950 598.050 338.400 ;
        RECT 634.950 339.600 637.050 340.050 ;
        RECT 649.950 339.600 652.050 340.050 ;
        RECT 634.950 338.400 652.050 339.600 ;
        RECT 634.950 337.950 637.050 338.400 ;
        RECT 649.950 337.950 652.050 338.400 ;
        RECT 664.950 339.600 667.050 340.050 ;
        RECT 730.950 339.600 733.050 340.050 ;
        RECT 664.950 338.400 733.050 339.600 ;
        RECT 664.950 337.950 667.050 338.400 ;
        RECT 730.950 337.950 733.050 338.400 ;
        RECT 760.950 339.600 763.050 340.050 ;
        RECT 775.950 339.600 778.050 340.050 ;
        RECT 760.950 338.400 778.050 339.600 ;
        RECT 760.950 337.950 763.050 338.400 ;
        RECT 775.950 337.950 778.050 338.400 ;
        RECT 778.950 339.600 781.050 340.050 ;
        RECT 799.950 339.600 802.050 340.050 ;
        RECT 778.950 338.400 802.050 339.600 ;
        RECT 778.950 337.950 781.050 338.400 ;
        RECT 799.950 337.950 802.050 338.400 ;
        RECT 808.950 339.600 811.050 340.050 ;
        RECT 844.950 339.600 847.050 340.050 ;
        RECT 847.950 339.600 850.050 340.050 ;
        RECT 808.950 338.400 850.050 339.600 ;
        RECT 808.950 337.950 811.050 338.400 ;
        RECT 844.950 337.950 847.050 338.400 ;
        RECT 847.950 337.950 850.050 338.400 ;
        RECT 859.950 339.600 862.050 340.050 ;
        RECT 874.950 339.600 877.050 340.050 ;
        RECT 859.950 338.400 877.050 339.600 ;
        RECT 859.950 337.950 862.050 338.400 ;
        RECT 874.950 337.950 877.050 338.400 ;
        RECT 415.950 336.600 418.050 337.050 ;
        RECT 604.950 336.600 607.050 337.050 ;
        RECT 415.950 335.400 607.050 336.600 ;
        RECT 415.950 334.950 418.050 335.400 ;
        RECT 604.950 334.950 607.050 335.400 ;
        RECT 607.950 336.600 610.050 337.050 ;
        RECT 712.950 336.600 715.050 337.050 ;
        RECT 607.950 335.400 715.050 336.600 ;
        RECT 607.950 334.950 610.050 335.400 ;
        RECT 712.950 334.950 715.050 335.400 ;
        RECT 763.950 336.600 766.050 337.050 ;
        RECT 769.950 336.600 772.050 337.050 ;
        RECT 763.950 335.400 772.050 336.600 ;
        RECT 763.950 334.950 766.050 335.400 ;
        RECT 769.950 334.950 772.050 335.400 ;
        RECT 835.950 336.600 838.050 337.050 ;
        RECT 850.950 336.600 853.050 337.050 ;
        RECT 835.950 335.400 853.050 336.600 ;
        RECT 835.950 334.950 838.050 335.400 ;
        RECT 850.950 334.950 853.050 335.400 ;
        RECT 871.950 336.600 874.050 337.050 ;
        RECT 880.950 336.600 883.050 337.050 ;
        RECT 871.950 335.400 883.050 336.600 ;
        RECT 871.950 334.950 874.050 335.400 ;
        RECT 880.950 334.950 883.050 335.400 ;
        RECT 415.950 333.600 418.050 334.050 ;
        RECT 407.400 332.400 418.050 333.600 ;
        RECT 268.950 331.950 271.050 332.400 ;
        RECT 277.950 331.950 280.050 332.400 ;
        RECT 379.950 331.950 382.050 332.400 ;
        RECT 415.950 331.950 418.050 332.400 ;
        RECT 676.950 333.600 679.050 334.050 ;
        RECT 715.950 333.600 718.050 334.050 ;
        RECT 676.950 332.400 718.050 333.600 ;
        RECT 676.950 331.950 679.050 332.400 ;
        RECT 715.950 331.950 718.050 332.400 ;
        RECT 52.950 330.600 55.050 331.050 ;
        RECT 85.950 330.600 88.050 331.050 ;
        RECT 52.950 329.400 88.050 330.600 ;
        RECT 52.950 328.950 55.050 329.400 ;
        RECT 85.950 328.950 88.050 329.400 ;
        RECT 196.950 330.600 199.050 331.050 ;
        RECT 319.950 330.600 322.050 331.050 ;
        RECT 418.950 330.600 421.050 331.050 ;
        RECT 445.950 330.600 448.050 331.050 ;
        RECT 196.950 329.400 448.050 330.600 ;
        RECT 196.950 328.950 199.050 329.400 ;
        RECT 319.950 328.950 322.050 329.400 ;
        RECT 418.950 328.950 421.050 329.400 ;
        RECT 445.950 328.950 448.050 329.400 ;
        RECT 484.950 330.600 487.050 331.050 ;
        RECT 496.950 330.600 499.050 331.050 ;
        RECT 484.950 329.400 499.050 330.600 ;
        RECT 484.950 328.950 487.050 329.400 ;
        RECT 496.950 328.950 499.050 329.400 ;
        RECT 646.950 330.600 649.050 331.050 ;
        RECT 658.950 330.600 661.050 331.050 ;
        RECT 646.950 329.400 661.050 330.600 ;
        RECT 646.950 328.950 649.050 329.400 ;
        RECT 658.950 328.950 661.050 329.400 ;
        RECT 742.950 330.600 745.050 331.050 ;
        RECT 817.950 330.600 820.050 331.050 ;
        RECT 742.950 329.400 820.050 330.600 ;
        RECT 742.950 328.950 745.050 329.400 ;
        RECT 817.950 328.950 820.050 329.400 ;
        RECT 64.950 327.600 67.050 328.050 ;
        RECT 148.950 327.600 151.050 328.050 ;
        RECT 64.950 326.400 151.050 327.600 ;
        RECT 64.950 325.950 67.050 326.400 ;
        RECT 148.950 325.950 151.050 326.400 ;
        RECT 298.950 327.600 301.050 328.050 ;
        RECT 517.950 327.600 520.050 328.050 ;
        RECT 298.950 326.400 520.050 327.600 ;
        RECT 298.950 325.950 301.050 326.400 ;
        RECT 517.950 325.950 520.050 326.400 ;
        RECT 583.950 327.600 586.050 328.050 ;
        RECT 775.950 327.600 778.050 328.050 ;
        RECT 784.950 327.600 787.050 328.050 ;
        RECT 583.950 326.400 787.050 327.600 ;
        RECT 583.950 325.950 586.050 326.400 ;
        RECT 775.950 325.950 778.050 326.400 ;
        RECT 784.950 325.950 787.050 326.400 ;
        RECT 787.950 327.600 790.050 328.050 ;
        RECT 799.950 327.600 802.050 328.050 ;
        RECT 805.950 327.600 808.050 328.050 ;
        RECT 787.950 326.400 808.050 327.600 ;
        RECT 787.950 325.950 790.050 326.400 ;
        RECT 799.950 325.950 802.050 326.400 ;
        RECT 805.950 325.950 808.050 326.400 ;
        RECT 256.950 324.600 259.050 325.050 ;
        RECT 301.950 324.600 304.050 325.050 ;
        RECT 256.950 323.400 304.050 324.600 ;
        RECT 256.950 322.950 259.050 323.400 ;
        RECT 301.950 322.950 304.050 323.400 ;
        RECT 373.950 324.600 376.050 325.050 ;
        RECT 382.950 324.600 385.050 325.050 ;
        RECT 373.950 323.400 385.050 324.600 ;
        RECT 373.950 322.950 376.050 323.400 ;
        RECT 382.950 322.950 385.050 323.400 ;
        RECT 514.950 324.600 517.050 325.050 ;
        RECT 610.950 324.600 613.050 325.050 ;
        RECT 514.950 323.400 613.050 324.600 ;
        RECT 514.950 322.950 517.050 323.400 ;
        RECT 610.950 322.950 613.050 323.400 ;
        RECT 628.950 324.600 631.050 325.050 ;
        RECT 676.950 324.600 679.050 325.050 ;
        RECT 685.950 324.600 688.050 325.050 ;
        RECT 745.950 324.600 748.050 325.050 ;
        RECT 628.950 323.400 748.050 324.600 ;
        RECT 628.950 322.950 631.050 323.400 ;
        RECT 676.950 322.950 679.050 323.400 ;
        RECT 685.950 322.950 688.050 323.400 ;
        RECT 745.950 322.950 748.050 323.400 ;
        RECT 769.950 324.600 772.050 325.050 ;
        RECT 805.950 324.600 808.050 325.050 ;
        RECT 769.950 323.400 808.050 324.600 ;
        RECT 769.950 322.950 772.050 323.400 ;
        RECT 805.950 322.950 808.050 323.400 ;
        RECT 175.950 321.600 178.050 322.050 ;
        RECT 196.950 321.600 199.050 322.050 ;
        RECT 175.950 320.400 199.050 321.600 ;
        RECT 175.950 319.950 178.050 320.400 ;
        RECT 196.950 319.950 199.050 320.400 ;
        RECT 244.950 321.600 247.050 322.050 ;
        RECT 265.950 321.600 268.050 322.050 ;
        RECT 244.950 320.400 268.050 321.600 ;
        RECT 244.950 319.950 247.050 320.400 ;
        RECT 265.950 319.950 268.050 320.400 ;
        RECT 286.950 321.600 289.050 322.050 ;
        RECT 307.950 321.600 310.050 322.050 ;
        RECT 286.950 320.400 310.050 321.600 ;
        RECT 286.950 319.950 289.050 320.400 ;
        RECT 307.950 319.950 310.050 320.400 ;
        RECT 403.950 321.600 406.050 322.050 ;
        RECT 442.950 321.600 445.050 322.050 ;
        RECT 403.950 320.400 445.050 321.600 ;
        RECT 403.950 319.950 406.050 320.400 ;
        RECT 442.950 319.950 445.050 320.400 ;
        RECT 502.950 321.600 505.050 322.050 ;
        RECT 643.950 321.600 646.050 322.050 ;
        RECT 664.950 321.600 667.050 322.050 ;
        RECT 502.950 320.400 667.050 321.600 ;
        RECT 502.950 319.950 505.050 320.400 ;
        RECT 643.950 319.950 646.050 320.400 ;
        RECT 664.950 319.950 667.050 320.400 ;
        RECT 772.950 321.600 775.050 322.050 ;
        RECT 784.950 321.600 787.050 322.050 ;
        RECT 772.950 320.400 787.050 321.600 ;
        RECT 772.950 319.950 775.050 320.400 ;
        RECT 784.950 319.950 787.050 320.400 ;
        RECT 34.950 318.600 37.050 319.050 ;
        RECT 43.950 318.600 46.050 319.050 ;
        RECT 64.950 318.600 67.050 319.050 ;
        RECT 34.950 317.400 67.050 318.600 ;
        RECT 34.950 316.950 37.050 317.400 ;
        RECT 43.950 316.950 46.050 317.400 ;
        RECT 64.950 316.950 67.050 317.400 ;
        RECT 106.950 318.600 109.050 319.050 ;
        RECT 124.950 318.600 127.050 319.050 ;
        RECT 106.950 317.400 127.050 318.600 ;
        RECT 106.950 316.950 109.050 317.400 ;
        RECT 124.950 316.950 127.050 317.400 ;
        RECT 148.950 318.600 151.050 319.050 ;
        RECT 334.950 318.600 337.050 319.050 ;
        RECT 148.950 317.400 337.050 318.600 ;
        RECT 148.950 316.950 151.050 317.400 ;
        RECT 334.950 316.950 337.050 317.400 ;
        RECT 337.950 318.600 340.050 319.050 ;
        RECT 430.950 318.600 433.050 319.050 ;
        RECT 337.950 317.400 433.050 318.600 ;
        RECT 337.950 316.950 340.050 317.400 ;
        RECT 430.950 316.950 433.050 317.400 ;
        RECT 439.950 318.600 442.050 319.050 ;
        RECT 490.950 318.600 493.050 319.050 ;
        RECT 508.950 318.600 511.050 319.050 ;
        RECT 439.950 317.400 511.050 318.600 ;
        RECT 439.950 316.950 442.050 317.400 ;
        RECT 490.950 316.950 493.050 317.400 ;
        RECT 508.950 316.950 511.050 317.400 ;
        RECT 541.950 318.600 544.050 319.050 ;
        RECT 625.950 318.600 628.050 319.050 ;
        RECT 541.950 317.400 628.050 318.600 ;
        RECT 541.950 316.950 544.050 317.400 ;
        RECT 625.950 316.950 628.050 317.400 ;
        RECT 649.950 318.600 652.050 319.050 ;
        RECT 694.950 318.600 697.050 319.050 ;
        RECT 649.950 317.400 697.050 318.600 ;
        RECT 649.950 316.950 652.050 317.400 ;
        RECT 694.950 316.950 697.050 317.400 ;
        RECT 712.950 318.600 715.050 319.050 ;
        RECT 751.950 318.600 754.050 319.050 ;
        RECT 853.950 318.600 856.050 319.050 ;
        RECT 712.950 317.400 856.050 318.600 ;
        RECT 712.950 316.950 715.050 317.400 ;
        RECT 751.950 316.950 754.050 317.400 ;
        RECT 853.950 316.950 856.050 317.400 ;
        RECT 862.950 318.600 865.050 319.050 ;
        RECT 877.950 318.600 880.050 319.050 ;
        RECT 862.950 317.400 880.050 318.600 ;
        RECT 862.950 316.950 865.050 317.400 ;
        RECT 877.950 316.950 880.050 317.400 ;
        RECT 37.950 315.600 40.050 316.050 ;
        RECT 46.950 315.600 49.050 316.050 ;
        RECT 58.950 315.600 61.050 316.050 ;
        RECT 37.950 314.400 61.050 315.600 ;
        RECT 37.950 313.950 40.050 314.400 ;
        RECT 46.950 313.950 49.050 314.400 ;
        RECT 58.950 313.950 61.050 314.400 ;
        RECT 67.950 315.600 70.050 316.050 ;
        RECT 73.950 315.600 76.050 316.050 ;
        RECT 67.950 314.400 76.050 315.600 ;
        RECT 67.950 313.950 70.050 314.400 ;
        RECT 73.950 313.950 76.050 314.400 ;
        RECT 88.950 315.600 91.050 316.050 ;
        RECT 100.950 315.600 103.050 316.050 ;
        RECT 106.950 315.600 109.050 316.050 ;
        RECT 88.950 314.400 99.600 315.600 ;
        RECT 88.950 313.950 91.050 314.400 ;
        RECT 55.950 312.600 58.050 313.050 ;
        RECT 85.950 312.600 88.050 313.050 ;
        RECT 55.950 311.400 88.050 312.600 ;
        RECT 55.950 310.950 58.050 311.400 ;
        RECT 85.950 310.950 88.050 311.400 ;
        RECT 91.950 310.950 94.050 313.050 ;
        RECT 98.400 312.600 99.600 314.400 ;
        RECT 100.950 314.400 109.050 315.600 ;
        RECT 100.950 313.950 103.050 314.400 ;
        RECT 106.950 313.950 109.050 314.400 ;
        RECT 133.950 315.600 136.050 316.050 ;
        RECT 166.950 315.600 169.050 316.050 ;
        RECT 133.950 314.400 169.050 315.600 ;
        RECT 133.950 313.950 136.050 314.400 ;
        RECT 166.950 313.950 169.050 314.400 ;
        RECT 262.950 315.600 265.050 316.050 ;
        RECT 295.950 315.600 298.050 316.050 ;
        RECT 262.950 314.400 298.050 315.600 ;
        RECT 262.950 313.950 265.050 314.400 ;
        RECT 295.950 313.950 298.050 314.400 ;
        RECT 322.950 315.600 325.050 316.050 ;
        RECT 340.950 315.600 343.050 316.050 ;
        RECT 322.950 314.400 343.050 315.600 ;
        RECT 322.950 313.950 325.050 314.400 ;
        RECT 340.950 313.950 343.050 314.400 ;
        RECT 499.950 315.600 502.050 316.050 ;
        RECT 511.950 315.600 514.050 316.050 ;
        RECT 499.950 314.400 514.050 315.600 ;
        RECT 499.950 313.950 502.050 314.400 ;
        RECT 511.950 313.950 514.050 314.400 ;
        RECT 565.950 313.950 568.050 316.050 ;
        RECT 601.950 315.600 604.050 316.050 ;
        RECT 613.950 315.600 616.050 316.050 ;
        RECT 601.950 314.400 616.050 315.600 ;
        RECT 601.950 313.950 604.050 314.400 ;
        RECT 613.950 313.950 616.050 314.400 ;
        RECT 673.950 315.600 676.050 316.050 ;
        RECT 685.950 315.600 688.050 316.050 ;
        RECT 673.950 314.400 688.050 315.600 ;
        RECT 673.950 313.950 676.050 314.400 ;
        RECT 685.950 313.950 688.050 314.400 ;
        RECT 694.950 315.600 697.050 316.050 ;
        RECT 706.950 315.600 709.050 316.050 ;
        RECT 694.950 314.400 709.050 315.600 ;
        RECT 694.950 313.950 697.050 314.400 ;
        RECT 706.950 313.950 709.050 314.400 ;
        RECT 730.950 315.600 733.050 316.050 ;
        RECT 733.950 315.600 736.050 316.050 ;
        RECT 742.950 315.600 745.050 316.050 ;
        RECT 730.950 314.400 745.050 315.600 ;
        RECT 730.950 313.950 733.050 314.400 ;
        RECT 733.950 313.950 736.050 314.400 ;
        RECT 742.950 313.950 745.050 314.400 ;
        RECT 790.950 315.600 793.050 316.050 ;
        RECT 802.950 315.600 805.050 316.050 ;
        RECT 790.950 314.400 805.050 315.600 ;
        RECT 790.950 313.950 793.050 314.400 ;
        RECT 802.950 313.950 805.050 314.400 ;
        RECT 838.950 315.600 841.050 316.050 ;
        RECT 850.950 315.600 853.050 316.050 ;
        RECT 838.950 314.400 853.050 315.600 ;
        RECT 838.950 313.950 841.050 314.400 ;
        RECT 850.950 313.950 853.050 314.400 ;
        RECT 856.950 315.600 859.050 316.050 ;
        RECT 865.950 315.600 868.050 316.050 ;
        RECT 856.950 314.400 868.050 315.600 ;
        RECT 856.950 313.950 859.050 314.400 ;
        RECT 865.950 313.950 868.050 314.400 ;
        RECT 130.950 312.600 133.050 313.050 ;
        RECT 169.950 312.600 172.050 313.050 ;
        RECT 98.400 311.400 111.600 312.600 ;
        RECT 16.950 309.600 19.050 310.050 ;
        RECT 67.950 309.600 70.050 310.050 ;
        RECT 76.950 309.600 79.050 310.050 ;
        RECT 16.950 308.400 33.600 309.600 ;
        RECT 16.950 307.950 19.050 308.400 ;
        RECT 32.400 307.050 33.600 308.400 ;
        RECT 67.950 308.400 79.050 309.600 ;
        RECT 92.400 309.600 93.600 310.950 ;
        RECT 110.400 310.050 111.600 311.400 ;
        RECT 130.950 311.400 172.050 312.600 ;
        RECT 130.950 310.950 133.050 311.400 ;
        RECT 169.950 310.950 172.050 311.400 ;
        RECT 178.950 312.600 181.050 313.050 ;
        RECT 187.950 312.600 190.050 313.050 ;
        RECT 178.950 311.400 190.050 312.600 ;
        RECT 178.950 310.950 181.050 311.400 ;
        RECT 187.950 310.950 190.050 311.400 ;
        RECT 211.950 312.600 214.050 313.050 ;
        RECT 226.950 312.600 229.050 313.050 ;
        RECT 247.950 312.600 250.050 313.050 ;
        RECT 211.950 311.400 250.050 312.600 ;
        RECT 211.950 310.950 214.050 311.400 ;
        RECT 226.950 310.950 229.050 311.400 ;
        RECT 247.950 310.950 250.050 311.400 ;
        RECT 271.950 312.600 274.050 313.050 ;
        RECT 325.950 312.600 328.050 313.050 ;
        RECT 328.950 312.600 331.050 313.050 ;
        RECT 271.950 311.400 331.050 312.600 ;
        RECT 271.950 310.950 274.050 311.400 ;
        RECT 103.950 309.600 106.050 310.050 ;
        RECT 92.400 308.400 106.050 309.600 ;
        RECT 67.950 307.950 70.050 308.400 ;
        RECT 76.950 307.950 79.050 308.400 ;
        RECT 103.950 307.950 106.050 308.400 ;
        RECT 109.950 307.950 112.050 310.050 ;
        RECT 136.950 309.600 139.050 310.050 ;
        RECT 145.950 309.600 148.050 310.050 ;
        RECT 136.950 308.400 148.050 309.600 ;
        RECT 136.950 307.950 139.050 308.400 ;
        RECT 145.950 307.950 148.050 308.400 ;
        RECT 151.950 309.600 154.050 310.050 ;
        RECT 211.950 309.600 214.050 310.050 ;
        RECT 151.950 308.400 214.050 309.600 ;
        RECT 151.950 307.950 154.050 308.400 ;
        RECT 211.950 307.950 214.050 308.400 ;
        RECT 223.950 309.600 226.050 310.050 ;
        RECT 232.950 309.600 235.050 310.050 ;
        RECT 223.950 308.400 235.050 309.600 ;
        RECT 223.950 307.950 226.050 308.400 ;
        RECT 232.950 307.950 235.050 308.400 ;
        RECT 244.950 309.600 247.050 310.050 ;
        RECT 272.400 309.600 273.600 310.950 ;
        RECT 293.400 310.050 294.600 311.400 ;
        RECT 325.950 310.950 328.050 311.400 ;
        RECT 328.950 310.950 331.050 311.400 ;
        RECT 382.950 312.600 385.050 313.050 ;
        RECT 388.950 312.600 391.050 313.050 ;
        RECT 382.950 311.400 391.050 312.600 ;
        RECT 382.950 310.950 385.050 311.400 ;
        RECT 388.950 310.950 391.050 311.400 ;
        RECT 394.950 312.600 397.050 313.050 ;
        RECT 427.950 312.600 430.050 313.050 ;
        RECT 394.950 311.400 430.050 312.600 ;
        RECT 394.950 310.950 397.050 311.400 ;
        RECT 427.950 310.950 430.050 311.400 ;
        RECT 451.950 312.600 454.050 313.050 ;
        RECT 469.950 312.600 472.050 313.050 ;
        RECT 517.950 312.600 520.050 313.050 ;
        RECT 451.950 311.400 520.050 312.600 ;
        RECT 451.950 310.950 454.050 311.400 ;
        RECT 469.950 310.950 472.050 311.400 ;
        RECT 517.950 310.950 520.050 311.400 ;
        RECT 526.950 312.600 529.050 313.050 ;
        RECT 532.950 312.600 535.050 313.050 ;
        RECT 526.950 311.400 535.050 312.600 ;
        RECT 526.950 310.950 529.050 311.400 ;
        RECT 532.950 310.950 535.050 311.400 ;
        RECT 566.400 310.050 567.600 313.950 ;
        RECT 568.950 312.600 571.050 313.050 ;
        RECT 586.950 312.600 589.050 313.050 ;
        RECT 568.950 311.400 589.050 312.600 ;
        RECT 568.950 310.950 571.050 311.400 ;
        RECT 586.950 310.950 589.050 311.400 ;
        RECT 595.950 312.600 598.050 313.050 ;
        RECT 619.950 312.600 622.050 313.050 ;
        RECT 595.950 311.400 622.050 312.600 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 619.950 310.950 622.050 311.400 ;
        RECT 658.950 312.600 661.050 313.050 ;
        RECT 667.950 312.600 670.050 313.050 ;
        RECT 658.950 311.400 670.050 312.600 ;
        RECT 658.950 310.950 661.050 311.400 ;
        RECT 667.950 310.950 670.050 311.400 ;
        RECT 691.950 312.600 694.050 313.050 ;
        RECT 703.950 312.600 706.050 313.050 ;
        RECT 691.950 311.400 706.050 312.600 ;
        RECT 691.950 310.950 694.050 311.400 ;
        RECT 703.950 310.950 706.050 311.400 ;
        RECT 760.950 312.600 763.050 313.050 ;
        RECT 766.950 312.600 769.050 313.050 ;
        RECT 760.950 311.400 769.050 312.600 ;
        RECT 760.950 310.950 763.050 311.400 ;
        RECT 766.950 310.950 769.050 311.400 ;
        RECT 772.950 312.600 775.050 313.050 ;
        RECT 778.950 312.600 781.050 313.050 ;
        RECT 772.950 311.400 781.050 312.600 ;
        RECT 772.950 310.950 775.050 311.400 ;
        RECT 778.950 310.950 781.050 311.400 ;
        RECT 820.950 312.600 823.050 313.050 ;
        RECT 838.950 312.600 841.050 313.050 ;
        RECT 820.950 311.400 841.050 312.600 ;
        RECT 820.950 310.950 823.050 311.400 ;
        RECT 838.950 310.950 841.050 311.400 ;
        RECT 853.950 312.600 856.050 313.050 ;
        RECT 868.950 312.600 871.050 313.050 ;
        RECT 853.950 311.400 871.050 312.600 ;
        RECT 853.950 310.950 856.050 311.400 ;
        RECT 868.950 310.950 871.050 311.400 ;
        RECT 244.950 308.400 273.600 309.600 ;
        RECT 244.950 307.950 247.050 308.400 ;
        RECT 280.950 307.950 283.050 310.050 ;
        RECT 292.950 307.950 295.050 310.050 ;
        RECT 343.950 309.600 346.050 310.050 ;
        RECT 397.950 309.600 400.050 310.050 ;
        RECT 343.950 308.400 400.050 309.600 ;
        RECT 343.950 307.950 346.050 308.400 ;
        RECT 397.950 307.950 400.050 308.400 ;
        RECT 421.950 309.600 424.050 310.050 ;
        RECT 472.950 309.600 475.050 310.050 ;
        RECT 421.950 308.400 475.050 309.600 ;
        RECT 421.950 307.950 424.050 308.400 ;
        RECT 472.950 307.950 475.050 308.400 ;
        RECT 478.950 309.600 481.050 310.050 ;
        RECT 493.950 309.600 496.050 310.050 ;
        RECT 478.950 308.400 496.050 309.600 ;
        RECT 478.950 307.950 481.050 308.400 ;
        RECT 493.950 307.950 496.050 308.400 ;
        RECT 523.950 309.600 526.050 310.050 ;
        RECT 538.950 309.600 541.050 310.050 ;
        RECT 523.950 308.400 541.050 309.600 ;
        RECT 523.950 307.950 526.050 308.400 ;
        RECT 538.950 307.950 541.050 308.400 ;
        RECT 565.950 307.950 568.050 310.050 ;
        RECT 571.950 309.600 574.050 310.050 ;
        RECT 583.950 309.600 586.050 310.050 ;
        RECT 571.950 308.400 586.050 309.600 ;
        RECT 571.950 307.950 574.050 308.400 ;
        RECT 583.950 307.950 586.050 308.400 ;
        RECT 607.950 309.600 610.050 310.050 ;
        RECT 628.950 309.600 631.050 310.050 ;
        RECT 607.950 308.400 631.050 309.600 ;
        RECT 607.950 307.950 610.050 308.400 ;
        RECT 628.950 307.950 631.050 308.400 ;
        RECT 646.950 309.600 649.050 310.050 ;
        RECT 661.950 309.600 664.050 310.050 ;
        RECT 646.950 308.400 664.050 309.600 ;
        RECT 646.950 307.950 649.050 308.400 ;
        RECT 661.950 307.950 664.050 308.400 ;
        RECT 676.950 309.600 679.050 310.050 ;
        RECT 682.950 309.600 685.050 310.050 ;
        RECT 676.950 308.400 685.050 309.600 ;
        RECT 676.950 307.950 679.050 308.400 ;
        RECT 682.950 307.950 685.050 308.400 ;
        RECT 688.950 309.600 691.050 310.050 ;
        RECT 694.950 309.600 697.050 310.050 ;
        RECT 688.950 308.400 697.050 309.600 ;
        RECT 688.950 307.950 691.050 308.400 ;
        RECT 694.950 307.950 697.050 308.400 ;
        RECT 709.950 309.600 712.050 310.050 ;
        RECT 718.950 309.600 721.050 310.050 ;
        RECT 709.950 308.400 721.050 309.600 ;
        RECT 709.950 307.950 712.050 308.400 ;
        RECT 718.950 307.950 721.050 308.400 ;
        RECT 754.950 309.600 757.050 310.050 ;
        RECT 787.950 309.600 790.050 310.050 ;
        RECT 754.950 308.400 790.050 309.600 ;
        RECT 754.950 307.950 757.050 308.400 ;
        RECT 787.950 307.950 790.050 308.400 ;
        RECT 793.950 309.600 796.050 310.050 ;
        RECT 808.950 309.600 811.050 310.050 ;
        RECT 793.950 308.400 811.050 309.600 ;
        RECT 793.950 307.950 796.050 308.400 ;
        RECT 808.950 307.950 811.050 308.400 ;
        RECT 817.950 309.600 820.050 310.050 ;
        RECT 820.950 309.600 823.050 310.050 ;
        RECT 826.950 309.600 829.050 310.050 ;
        RECT 817.950 308.400 829.050 309.600 ;
        RECT 817.950 307.950 820.050 308.400 ;
        RECT 820.950 307.950 823.050 308.400 ;
        RECT 826.950 307.950 829.050 308.400 ;
        RECT 850.950 309.600 853.050 310.050 ;
        RECT 859.950 309.600 862.050 310.050 ;
        RECT 865.950 309.600 868.050 310.050 ;
        RECT 850.950 308.400 862.050 309.600 ;
        RECT 850.950 307.950 853.050 308.400 ;
        RECT 859.950 307.950 862.050 308.400 ;
        RECT 863.400 308.400 868.050 309.600 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 100.950 306.600 103.050 307.050 ;
        RECT 127.950 306.600 130.050 307.050 ;
        RECT 100.950 305.400 130.050 306.600 ;
        RECT 100.950 304.950 103.050 305.400 ;
        RECT 127.950 304.950 130.050 305.400 ;
        RECT 193.950 306.600 196.050 307.050 ;
        RECT 208.950 306.600 211.050 307.050 ;
        RECT 193.950 305.400 211.050 306.600 ;
        RECT 193.950 304.950 196.050 305.400 ;
        RECT 208.950 304.950 211.050 305.400 ;
        RECT 256.950 306.600 259.050 307.050 ;
        RECT 274.950 306.600 277.050 307.050 ;
        RECT 256.950 305.400 277.050 306.600 ;
        RECT 256.950 304.950 259.050 305.400 ;
        RECT 274.950 304.950 277.050 305.400 ;
        RECT 277.950 306.600 280.050 307.050 ;
        RECT 281.400 306.600 282.600 307.950 ;
        RECT 277.950 305.400 282.600 306.600 ;
        RECT 364.950 306.600 367.050 307.050 ;
        RECT 379.950 306.600 382.050 307.050 ;
        RECT 364.950 305.400 382.050 306.600 ;
        RECT 277.950 304.950 280.050 305.400 ;
        RECT 364.950 304.950 367.050 305.400 ;
        RECT 379.950 304.950 382.050 305.400 ;
        RECT 388.950 306.600 391.050 307.050 ;
        RECT 394.950 306.600 397.050 307.050 ;
        RECT 388.950 305.400 397.050 306.600 ;
        RECT 388.950 304.950 391.050 305.400 ;
        RECT 394.950 304.950 397.050 305.400 ;
        RECT 433.950 306.600 436.050 307.050 ;
        RECT 469.950 306.600 472.050 307.050 ;
        RECT 490.950 306.600 493.050 307.050 ;
        RECT 505.950 306.600 508.050 307.050 ;
        RECT 433.950 305.400 508.050 306.600 ;
        RECT 433.950 304.950 436.050 305.400 ;
        RECT 469.950 304.950 472.050 305.400 ;
        RECT 490.950 304.950 493.050 305.400 ;
        RECT 505.950 304.950 508.050 305.400 ;
        RECT 517.950 306.600 520.050 307.050 ;
        RECT 529.950 306.600 532.050 307.050 ;
        RECT 556.950 306.600 559.050 307.050 ;
        RECT 517.950 305.400 559.050 306.600 ;
        RECT 517.950 304.950 520.050 305.400 ;
        RECT 529.950 304.950 532.050 305.400 ;
        RECT 556.950 304.950 559.050 305.400 ;
        RECT 619.950 306.600 622.050 307.050 ;
        RECT 622.950 306.600 625.050 307.050 ;
        RECT 646.950 306.600 649.050 307.050 ;
        RECT 619.950 305.400 649.050 306.600 ;
        RECT 619.950 304.950 622.050 305.400 ;
        RECT 622.950 304.950 625.050 305.400 ;
        RECT 646.950 304.950 649.050 305.400 ;
        RECT 673.950 306.600 676.050 307.050 ;
        RECT 727.950 306.600 730.050 307.050 ;
        RECT 673.950 305.400 730.050 306.600 ;
        RECT 673.950 304.950 676.050 305.400 ;
        RECT 727.950 304.950 730.050 305.400 ;
        RECT 844.950 306.600 847.050 307.050 ;
        RECT 863.400 306.600 864.600 308.400 ;
        RECT 865.950 307.950 868.050 308.400 ;
        RECT 844.950 305.400 864.600 306.600 ;
        RECT 865.950 306.600 868.050 307.050 ;
        RECT 874.950 306.600 877.050 307.050 ;
        RECT 865.950 305.400 877.050 306.600 ;
        RECT 844.950 304.950 847.050 305.400 ;
        RECT 865.950 304.950 868.050 305.400 ;
        RECT 874.950 304.950 877.050 305.400 ;
        RECT 13.950 303.600 16.050 304.050 ;
        RECT 55.950 303.600 58.050 304.050 ;
        RECT 13.950 302.400 58.050 303.600 ;
        RECT 13.950 301.950 16.050 302.400 ;
        RECT 55.950 301.950 58.050 302.400 ;
        RECT 133.950 303.600 136.050 304.050 ;
        RECT 187.950 303.600 190.050 304.050 ;
        RECT 133.950 302.400 190.050 303.600 ;
        RECT 133.950 301.950 136.050 302.400 ;
        RECT 187.950 301.950 190.050 302.400 ;
        RECT 232.950 303.600 235.050 304.050 ;
        RECT 238.950 303.600 241.050 304.050 ;
        RECT 232.950 302.400 241.050 303.600 ;
        RECT 232.950 301.950 235.050 302.400 ;
        RECT 238.950 301.950 241.050 302.400 ;
        RECT 340.950 303.600 343.050 304.050 ;
        RECT 358.950 303.600 361.050 304.050 ;
        RECT 340.950 302.400 361.050 303.600 ;
        RECT 340.950 301.950 343.050 302.400 ;
        RECT 358.950 301.950 361.050 302.400 ;
        RECT 394.950 303.600 397.050 304.050 ;
        RECT 403.950 303.600 406.050 304.050 ;
        RECT 394.950 302.400 406.050 303.600 ;
        RECT 394.950 301.950 397.050 302.400 ;
        RECT 403.950 301.950 406.050 302.400 ;
        RECT 475.950 303.600 478.050 304.050 ;
        RECT 538.950 303.600 541.050 304.050 ;
        RECT 562.950 303.600 565.050 304.050 ;
        RECT 475.950 302.400 565.050 303.600 ;
        RECT 475.950 301.950 478.050 302.400 ;
        RECT 538.950 301.950 541.050 302.400 ;
        RECT 562.950 301.950 565.050 302.400 ;
        RECT 586.950 303.600 589.050 304.050 ;
        RECT 640.950 303.600 643.050 304.050 ;
        RECT 658.950 303.600 661.050 304.050 ;
        RECT 586.950 302.400 661.050 303.600 ;
        RECT 586.950 301.950 589.050 302.400 ;
        RECT 640.950 301.950 643.050 302.400 ;
        RECT 658.950 301.950 661.050 302.400 ;
        RECT 139.950 300.600 142.050 301.050 ;
        RECT 148.950 300.600 151.050 301.050 ;
        RECT 139.950 299.400 151.050 300.600 ;
        RECT 139.950 298.950 142.050 299.400 ;
        RECT 148.950 298.950 151.050 299.400 ;
        RECT 235.950 300.600 238.050 301.050 ;
        RECT 244.950 300.600 247.050 301.050 ;
        RECT 250.950 300.600 253.050 301.050 ;
        RECT 235.950 299.400 253.050 300.600 ;
        RECT 235.950 298.950 238.050 299.400 ;
        RECT 244.950 298.950 247.050 299.400 ;
        RECT 250.950 298.950 253.050 299.400 ;
        RECT 400.950 300.600 403.050 301.050 ;
        RECT 478.950 300.600 481.050 301.050 ;
        RECT 400.950 299.400 481.050 300.600 ;
        RECT 400.950 298.950 403.050 299.400 ;
        RECT 478.950 298.950 481.050 299.400 ;
        RECT 562.950 300.600 565.050 301.050 ;
        RECT 595.950 300.600 598.050 301.050 ;
        RECT 610.950 300.600 613.050 301.050 ;
        RECT 562.950 299.400 613.050 300.600 ;
        RECT 562.950 298.950 565.050 299.400 ;
        RECT 595.950 298.950 598.050 299.400 ;
        RECT 610.950 298.950 613.050 299.400 ;
        RECT 10.950 297.600 13.050 298.050 ;
        RECT 43.950 297.600 46.050 298.050 ;
        RECT 10.950 296.400 46.050 297.600 ;
        RECT 10.950 295.950 13.050 296.400 ;
        RECT 43.950 295.950 46.050 296.400 ;
        RECT 235.950 297.600 238.050 298.050 ;
        RECT 241.950 297.600 244.050 298.050 ;
        RECT 235.950 296.400 244.050 297.600 ;
        RECT 235.950 295.950 238.050 296.400 ;
        RECT 241.950 295.950 244.050 296.400 ;
        RECT 799.950 297.600 802.050 298.050 ;
        RECT 826.950 297.600 829.050 298.050 ;
        RECT 799.950 296.400 829.050 297.600 ;
        RECT 799.950 295.950 802.050 296.400 ;
        RECT 826.950 295.950 829.050 296.400 ;
        RECT 175.950 291.600 178.050 292.050 ;
        RECT 256.950 291.600 259.050 292.050 ;
        RECT 175.950 290.400 259.050 291.600 ;
        RECT 175.950 289.950 178.050 290.400 ;
        RECT 256.950 289.950 259.050 290.400 ;
        RECT 307.950 291.600 310.050 292.050 ;
        RECT 385.950 291.600 388.050 292.050 ;
        RECT 400.950 291.600 403.050 292.050 ;
        RECT 307.950 290.400 403.050 291.600 ;
        RECT 307.950 289.950 310.050 290.400 ;
        RECT 385.950 289.950 388.050 290.400 ;
        RECT 400.950 289.950 403.050 290.400 ;
        RECT 496.950 288.600 499.050 289.050 ;
        RECT 526.950 288.600 529.050 289.050 ;
        RECT 535.950 288.600 538.050 289.050 ;
        RECT 496.950 287.400 538.050 288.600 ;
        RECT 496.950 286.950 499.050 287.400 ;
        RECT 526.950 286.950 529.050 287.400 ;
        RECT 535.950 286.950 538.050 287.400 ;
        RECT 601.950 285.600 604.050 286.050 ;
        RECT 607.950 285.600 610.050 286.050 ;
        RECT 601.950 284.400 610.050 285.600 ;
        RECT 601.950 283.950 604.050 284.400 ;
        RECT 607.950 283.950 610.050 284.400 ;
        RECT 379.950 282.600 382.050 283.050 ;
        RECT 409.950 282.600 412.050 283.050 ;
        RECT 379.950 281.400 412.050 282.600 ;
        RECT 379.950 280.950 382.050 281.400 ;
        RECT 409.950 280.950 412.050 281.400 ;
        RECT 589.950 282.600 592.050 283.050 ;
        RECT 652.950 282.600 655.050 283.050 ;
        RECT 670.950 282.600 673.050 283.050 ;
        RECT 589.950 281.400 673.050 282.600 ;
        RECT 589.950 280.950 592.050 281.400 ;
        RECT 652.950 280.950 655.050 281.400 ;
        RECT 670.950 280.950 673.050 281.400 ;
        RECT 856.950 282.600 859.050 283.050 ;
        RECT 868.950 282.600 871.050 283.050 ;
        RECT 856.950 281.400 871.050 282.600 ;
        RECT 856.950 280.950 859.050 281.400 ;
        RECT 868.950 280.950 871.050 281.400 ;
        RECT 67.950 279.600 70.050 280.050 ;
        RECT 82.950 279.600 85.050 280.050 ;
        RECT 67.950 278.400 85.050 279.600 ;
        RECT 67.950 277.950 70.050 278.400 ;
        RECT 82.950 277.950 85.050 278.400 ;
        RECT 316.950 279.600 319.050 280.050 ;
        RECT 505.950 279.600 508.050 280.050 ;
        RECT 316.950 278.400 508.050 279.600 ;
        RECT 316.950 277.950 319.050 278.400 ;
        RECT 505.950 277.950 508.050 278.400 ;
        RECT 664.950 279.600 667.050 280.050 ;
        RECT 847.950 279.600 850.050 280.050 ;
        RECT 856.950 279.600 859.050 280.050 ;
        RECT 664.950 278.400 859.050 279.600 ;
        RECT 664.950 277.950 667.050 278.400 ;
        RECT 847.950 277.950 850.050 278.400 ;
        RECT 856.950 277.950 859.050 278.400 ;
        RECT 70.950 276.600 73.050 277.050 ;
        RECT 91.950 276.600 94.050 277.050 ;
        RECT 70.950 275.400 94.050 276.600 ;
        RECT 70.950 274.950 73.050 275.400 ;
        RECT 91.950 274.950 94.050 275.400 ;
        RECT 133.950 276.600 136.050 277.050 ;
        RECT 139.950 276.600 142.050 277.050 ;
        RECT 133.950 275.400 142.050 276.600 ;
        RECT 133.950 274.950 136.050 275.400 ;
        RECT 139.950 274.950 142.050 275.400 ;
        RECT 172.950 276.600 175.050 277.050 ;
        RECT 244.950 276.600 247.050 277.050 ;
        RECT 172.950 275.400 247.050 276.600 ;
        RECT 172.950 274.950 175.050 275.400 ;
        RECT 244.950 274.950 247.050 275.400 ;
        RECT 265.950 276.600 268.050 277.050 ;
        RECT 304.950 276.600 307.050 277.050 ;
        RECT 265.950 275.400 307.050 276.600 ;
        RECT 265.950 274.950 268.050 275.400 ;
        RECT 304.950 274.950 307.050 275.400 ;
        RECT 310.950 276.600 313.050 277.050 ;
        RECT 316.950 276.600 319.050 277.050 ;
        RECT 310.950 275.400 319.050 276.600 ;
        RECT 310.950 274.950 313.050 275.400 ;
        RECT 316.950 274.950 319.050 275.400 ;
        RECT 370.950 276.600 373.050 277.050 ;
        RECT 439.950 276.600 442.050 277.050 ;
        RECT 370.950 275.400 442.050 276.600 ;
        RECT 370.950 274.950 373.050 275.400 ;
        RECT 439.950 274.950 442.050 275.400 ;
        RECT 526.950 276.600 529.050 277.050 ;
        RECT 730.950 276.600 733.050 277.050 ;
        RECT 526.950 275.400 733.050 276.600 ;
        RECT 526.950 274.950 529.050 275.400 ;
        RECT 730.950 274.950 733.050 275.400 ;
        RECT 835.950 276.600 838.050 277.050 ;
        RECT 847.950 276.600 850.050 277.050 ;
        RECT 835.950 275.400 850.050 276.600 ;
        RECT 835.950 274.950 838.050 275.400 ;
        RECT 847.950 274.950 850.050 275.400 ;
        RECT 73.950 273.600 76.050 274.050 ;
        RECT 79.950 273.600 82.050 274.050 ;
        RECT 73.950 272.400 82.050 273.600 ;
        RECT 73.950 271.950 76.050 272.400 ;
        RECT 79.950 271.950 82.050 272.400 ;
        RECT 103.950 273.600 106.050 274.050 ;
        RECT 118.950 273.600 121.050 274.050 ;
        RECT 127.950 273.600 130.050 274.050 ;
        RECT 148.950 273.600 151.050 274.050 ;
        RECT 193.950 273.600 196.050 274.050 ;
        RECT 103.950 272.400 196.050 273.600 ;
        RECT 103.950 271.950 106.050 272.400 ;
        RECT 118.950 271.950 121.050 272.400 ;
        RECT 127.950 271.950 130.050 272.400 ;
        RECT 148.950 271.950 151.050 272.400 ;
        RECT 193.950 271.950 196.050 272.400 ;
        RECT 196.950 273.600 199.050 274.050 ;
        RECT 220.950 273.600 223.050 274.050 ;
        RECT 196.950 272.400 223.050 273.600 ;
        RECT 196.950 271.950 199.050 272.400 ;
        RECT 220.950 271.950 223.050 272.400 ;
        RECT 277.950 273.600 280.050 274.050 ;
        RECT 316.950 273.600 319.050 274.050 ;
        RECT 331.950 273.600 334.050 274.050 ;
        RECT 277.950 272.400 285.600 273.600 ;
        RECT 277.950 271.950 280.050 272.400 ;
        RECT 70.950 270.600 73.050 271.050 ;
        RECT 85.950 270.600 88.050 271.050 ;
        RECT 70.950 269.400 88.050 270.600 ;
        RECT 70.950 268.950 73.050 269.400 ;
        RECT 85.950 268.950 88.050 269.400 ;
        RECT 121.950 270.600 124.050 271.050 ;
        RECT 133.950 270.600 136.050 271.050 ;
        RECT 154.950 270.600 157.050 271.050 ;
        RECT 121.950 269.400 157.050 270.600 ;
        RECT 121.950 268.950 124.050 269.400 ;
        RECT 133.950 268.950 136.050 269.400 ;
        RECT 154.950 268.950 157.050 269.400 ;
        RECT 187.950 268.950 190.050 271.050 ;
        RECT 223.950 270.600 226.050 271.050 ;
        RECT 238.950 270.600 241.050 271.050 ;
        RECT 223.950 269.400 241.050 270.600 ;
        RECT 223.950 268.950 226.050 269.400 ;
        RECT 238.950 268.950 241.050 269.400 ;
        RECT 280.950 268.950 283.050 271.050 ;
        RECT 284.400 270.600 285.600 272.400 ;
        RECT 316.950 272.400 334.050 273.600 ;
        RECT 316.950 271.950 319.050 272.400 ;
        RECT 331.950 271.950 334.050 272.400 ;
        RECT 391.950 273.600 394.050 274.050 ;
        RECT 397.950 273.600 400.050 274.050 ;
        RECT 391.950 272.400 400.050 273.600 ;
        RECT 391.950 271.950 394.050 272.400 ;
        RECT 397.950 271.950 400.050 272.400 ;
        RECT 403.950 273.600 406.050 274.050 ;
        RECT 415.950 273.600 418.050 274.050 ;
        RECT 403.950 272.400 418.050 273.600 ;
        RECT 403.950 271.950 406.050 272.400 ;
        RECT 415.950 271.950 418.050 272.400 ;
        RECT 487.950 273.600 490.050 274.050 ;
        RECT 526.950 273.600 529.050 274.050 ;
        RECT 487.950 272.400 529.050 273.600 ;
        RECT 487.950 271.950 490.050 272.400 ;
        RECT 526.950 271.950 529.050 272.400 ;
        RECT 568.950 273.600 571.050 274.050 ;
        RECT 577.950 273.600 580.050 274.050 ;
        RECT 592.950 273.600 595.050 274.050 ;
        RECT 568.950 272.400 595.050 273.600 ;
        RECT 568.950 271.950 571.050 272.400 ;
        RECT 577.950 271.950 580.050 272.400 ;
        RECT 592.950 271.950 595.050 272.400 ;
        RECT 685.950 273.600 688.050 274.050 ;
        RECT 700.950 273.600 703.050 274.050 ;
        RECT 685.950 272.400 703.050 273.600 ;
        RECT 685.950 271.950 688.050 272.400 ;
        RECT 700.950 271.950 703.050 272.400 ;
        RECT 733.950 273.600 736.050 274.050 ;
        RECT 748.950 273.600 751.050 274.050 ;
        RECT 784.950 273.600 787.050 274.050 ;
        RECT 733.950 272.400 738.600 273.600 ;
        RECT 733.950 271.950 736.050 272.400 ;
        RECT 737.400 271.050 738.600 272.400 ;
        RECT 748.950 272.400 787.050 273.600 ;
        RECT 748.950 271.950 751.050 272.400 ;
        RECT 784.950 271.950 787.050 272.400 ;
        RECT 295.950 270.600 298.050 271.050 ;
        RECT 284.400 269.400 298.050 270.600 ;
        RECT 295.950 268.950 298.050 269.400 ;
        RECT 322.950 270.600 325.050 271.050 ;
        RECT 394.950 270.600 397.050 271.050 ;
        RECT 406.950 270.600 409.050 271.050 ;
        RECT 412.950 270.600 415.050 271.050 ;
        RECT 322.950 269.400 402.600 270.600 ;
        RECT 322.950 268.950 325.050 269.400 ;
        RECT 394.950 268.950 397.050 269.400 ;
        RECT 31.950 265.950 34.050 268.050 ;
        RECT 79.950 267.600 82.050 268.050 ;
        RECT 94.950 267.600 97.050 268.050 ;
        RECT 79.950 266.400 97.050 267.600 ;
        RECT 79.950 265.950 82.050 266.400 ;
        RECT 94.950 265.950 97.050 266.400 ;
        RECT 166.950 267.600 169.050 268.050 ;
        RECT 175.950 267.600 178.050 268.050 ;
        RECT 166.950 266.400 178.050 267.600 ;
        RECT 188.400 267.600 189.600 268.950 ;
        RECT 202.950 267.600 205.050 268.050 ;
        RECT 188.400 266.400 205.050 267.600 ;
        RECT 166.950 265.950 169.050 266.400 ;
        RECT 175.950 265.950 178.050 266.400 ;
        RECT 202.950 265.950 205.050 266.400 ;
        RECT 226.950 267.600 229.050 268.050 ;
        RECT 235.950 267.600 238.050 268.050 ;
        RECT 265.950 267.600 268.050 268.050 ;
        RECT 281.400 267.600 282.600 268.950 ;
        RECT 373.950 267.600 376.050 268.050 ;
        RECT 226.950 266.400 376.050 267.600 ;
        RECT 226.950 265.950 229.050 266.400 ;
        RECT 235.950 265.950 238.050 266.400 ;
        RECT 265.950 265.950 268.050 266.400 ;
        RECT 373.950 265.950 376.050 266.400 ;
        RECT 391.950 267.600 394.050 268.050 ;
        RECT 397.950 267.600 400.050 268.050 ;
        RECT 391.950 266.400 400.050 267.600 ;
        RECT 401.400 267.600 402.600 269.400 ;
        RECT 406.950 269.400 415.050 270.600 ;
        RECT 406.950 268.950 409.050 269.400 ;
        RECT 412.950 268.950 415.050 269.400 ;
        RECT 418.950 270.600 421.050 271.050 ;
        RECT 427.950 270.600 430.050 271.050 ;
        RECT 448.950 270.600 451.050 271.050 ;
        RECT 418.950 269.400 451.050 270.600 ;
        RECT 418.950 268.950 421.050 269.400 ;
        RECT 427.950 268.950 430.050 269.400 ;
        RECT 448.950 268.950 451.050 269.400 ;
        RECT 484.950 270.600 487.050 271.050 ;
        RECT 499.950 270.600 502.050 271.050 ;
        RECT 484.950 269.400 502.050 270.600 ;
        RECT 484.950 268.950 487.050 269.400 ;
        RECT 499.950 268.950 502.050 269.400 ;
        RECT 547.950 270.600 550.050 271.050 ;
        RECT 598.950 270.600 601.050 271.050 ;
        RECT 547.950 269.400 601.050 270.600 ;
        RECT 547.950 268.950 550.050 269.400 ;
        RECT 598.950 268.950 601.050 269.400 ;
        RECT 619.950 270.600 622.050 271.050 ;
        RECT 640.950 270.600 643.050 271.050 ;
        RECT 619.950 269.400 643.050 270.600 ;
        RECT 619.950 268.950 622.050 269.400 ;
        RECT 640.950 268.950 643.050 269.400 ;
        RECT 655.950 270.600 658.050 271.050 ;
        RECT 670.950 270.600 673.050 271.050 ;
        RECT 655.950 269.400 673.050 270.600 ;
        RECT 655.950 268.950 658.050 269.400 ;
        RECT 670.950 268.950 673.050 269.400 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 754.950 270.600 757.050 271.050 ;
        RECT 769.950 270.600 772.050 271.050 ;
        RECT 793.950 270.600 796.050 271.050 ;
        RECT 754.950 269.400 772.050 270.600 ;
        RECT 754.950 268.950 757.050 269.400 ;
        RECT 769.950 268.950 772.050 269.400 ;
        RECT 782.400 269.400 796.050 270.600 ;
        RECT 430.950 267.600 433.050 268.050 ;
        RECT 401.400 266.400 433.050 267.600 ;
        RECT 391.950 265.950 394.050 266.400 ;
        RECT 397.950 265.950 400.050 266.400 ;
        RECT 430.950 265.950 433.050 266.400 ;
        RECT 511.950 267.600 514.050 268.050 ;
        RECT 529.950 267.600 532.050 268.050 ;
        RECT 511.950 266.400 532.050 267.600 ;
        RECT 511.950 265.950 514.050 266.400 ;
        RECT 529.950 265.950 532.050 266.400 ;
        RECT 538.950 267.600 541.050 268.050 ;
        RECT 544.950 267.600 547.050 268.050 ;
        RECT 538.950 266.400 547.050 267.600 ;
        RECT 538.950 265.950 541.050 266.400 ;
        RECT 544.950 265.950 547.050 266.400 ;
        RECT 550.950 267.600 553.050 268.050 ;
        RECT 559.950 267.600 562.050 268.050 ;
        RECT 550.950 266.400 562.050 267.600 ;
        RECT 550.950 265.950 553.050 266.400 ;
        RECT 559.950 265.950 562.050 266.400 ;
        RECT 565.950 267.600 568.050 268.050 ;
        RECT 571.950 267.600 574.050 268.050 ;
        RECT 565.950 266.400 574.050 267.600 ;
        RECT 565.950 265.950 568.050 266.400 ;
        RECT 571.950 265.950 574.050 266.400 ;
        RECT 595.950 267.600 598.050 268.050 ;
        RECT 637.950 267.600 640.050 268.050 ;
        RECT 595.950 266.400 640.050 267.600 ;
        RECT 595.950 265.950 598.050 266.400 ;
        RECT 637.950 265.950 640.050 266.400 ;
        RECT 643.950 267.600 646.050 268.050 ;
        RECT 664.950 267.600 667.050 268.050 ;
        RECT 643.950 266.400 667.050 267.600 ;
        RECT 643.950 265.950 646.050 266.400 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 673.950 267.600 676.050 268.050 ;
        RECT 694.950 267.600 697.050 268.050 ;
        RECT 712.950 267.600 715.050 268.050 ;
        RECT 727.950 267.600 730.050 268.050 ;
        RECT 673.950 266.400 697.050 267.600 ;
        RECT 673.950 265.950 676.050 266.400 ;
        RECT 694.950 265.950 697.050 266.400 ;
        RECT 698.400 266.400 730.050 267.600 ;
        RECT 32.400 264.600 33.600 265.950 ;
        RECT 46.950 264.600 49.050 265.050 ;
        RECT 64.950 264.600 67.050 265.050 ;
        RECT 32.400 263.400 67.050 264.600 ;
        RECT 46.950 262.950 49.050 263.400 ;
        RECT 64.950 262.950 67.050 263.400 ;
        RECT 73.950 264.600 76.050 265.050 ;
        RECT 100.950 264.600 103.050 265.050 ;
        RECT 73.950 263.400 103.050 264.600 ;
        RECT 73.950 262.950 76.050 263.400 ;
        RECT 100.950 262.950 103.050 263.400 ;
        RECT 112.950 264.600 115.050 265.050 ;
        RECT 121.950 264.600 124.050 265.050 ;
        RECT 112.950 263.400 124.050 264.600 ;
        RECT 112.950 262.950 115.050 263.400 ;
        RECT 121.950 262.950 124.050 263.400 ;
        RECT 124.950 264.600 127.050 265.050 ;
        RECT 151.950 264.600 154.050 265.050 ;
        RECT 172.950 264.600 175.050 265.050 ;
        RECT 124.950 263.400 175.050 264.600 ;
        RECT 124.950 262.950 127.050 263.400 ;
        RECT 151.950 262.950 154.050 263.400 ;
        RECT 172.950 262.950 175.050 263.400 ;
        RECT 184.950 264.600 187.050 265.050 ;
        RECT 217.950 264.600 220.050 265.050 ;
        RECT 184.950 263.400 220.050 264.600 ;
        RECT 184.950 262.950 187.050 263.400 ;
        RECT 217.950 262.950 220.050 263.400 ;
        RECT 253.950 264.600 256.050 265.050 ;
        RECT 265.950 264.600 268.050 265.050 ;
        RECT 253.950 263.400 268.050 264.600 ;
        RECT 253.950 262.950 256.050 263.400 ;
        RECT 265.950 262.950 268.050 263.400 ;
        RECT 523.950 264.600 526.050 265.050 ;
        RECT 586.950 264.600 589.050 265.050 ;
        RECT 523.950 263.400 589.050 264.600 ;
        RECT 523.950 262.950 526.050 263.400 ;
        RECT 586.950 262.950 589.050 263.400 ;
        RECT 592.950 264.600 595.050 265.050 ;
        RECT 616.950 264.600 619.050 265.050 ;
        RECT 592.950 263.400 619.050 264.600 ;
        RECT 592.950 262.950 595.050 263.400 ;
        RECT 616.950 262.950 619.050 263.400 ;
        RECT 658.950 264.600 661.050 265.050 ;
        RECT 698.400 264.600 699.600 266.400 ;
        RECT 712.950 265.950 715.050 266.400 ;
        RECT 727.950 265.950 730.050 266.400 ;
        RECT 757.950 267.600 760.050 268.050 ;
        RECT 782.400 267.600 783.600 269.400 ;
        RECT 793.950 268.950 796.050 269.400 ;
        RECT 826.950 270.600 829.050 271.050 ;
        RECT 853.950 270.600 856.050 271.050 ;
        RECT 826.950 269.400 856.050 270.600 ;
        RECT 826.950 268.950 829.050 269.400 ;
        RECT 853.950 268.950 856.050 269.400 ;
        RECT 757.950 266.400 783.600 267.600 ;
        RECT 784.950 267.600 787.050 268.050 ;
        RECT 790.950 267.600 793.050 268.050 ;
        RECT 784.950 266.400 793.050 267.600 ;
        RECT 757.950 265.950 760.050 266.400 ;
        RECT 784.950 265.950 787.050 266.400 ;
        RECT 790.950 265.950 793.050 266.400 ;
        RECT 796.950 267.600 799.050 268.050 ;
        RECT 817.950 267.600 820.050 268.050 ;
        RECT 796.950 266.400 820.050 267.600 ;
        RECT 796.950 265.950 799.050 266.400 ;
        RECT 817.950 265.950 820.050 266.400 ;
        RECT 658.950 263.400 699.600 264.600 ;
        RECT 733.950 264.600 736.050 265.050 ;
        RECT 751.950 264.600 754.050 265.050 ;
        RECT 733.950 263.400 754.050 264.600 ;
        RECT 658.950 262.950 661.050 263.400 ;
        RECT 733.950 262.950 736.050 263.400 ;
        RECT 751.950 262.950 754.050 263.400 ;
        RECT 826.950 264.600 829.050 265.050 ;
        RECT 844.950 264.600 847.050 265.050 ;
        RECT 826.950 263.400 847.050 264.600 ;
        RECT 826.950 262.950 829.050 263.400 ;
        RECT 844.950 262.950 847.050 263.400 ;
        RECT 874.950 264.600 877.050 265.050 ;
        RECT 880.950 264.600 883.050 265.050 ;
        RECT 874.950 263.400 883.050 264.600 ;
        RECT 874.950 262.950 877.050 263.400 ;
        RECT 880.950 262.950 883.050 263.400 ;
        RECT 88.950 261.600 91.050 262.050 ;
        RECT 130.950 261.600 133.050 262.050 ;
        RECT 88.950 260.400 133.050 261.600 ;
        RECT 88.950 259.950 91.050 260.400 ;
        RECT 130.950 259.950 133.050 260.400 ;
        RECT 265.950 261.600 268.050 262.050 ;
        RECT 382.950 261.600 385.050 262.050 ;
        RECT 265.950 260.400 385.050 261.600 ;
        RECT 265.950 259.950 268.050 260.400 ;
        RECT 382.950 259.950 385.050 260.400 ;
        RECT 541.950 261.600 544.050 262.050 ;
        RECT 547.950 261.600 550.050 262.050 ;
        RECT 541.950 260.400 550.050 261.600 ;
        RECT 541.950 259.950 544.050 260.400 ;
        RECT 547.950 259.950 550.050 260.400 ;
        RECT 700.950 261.600 703.050 262.050 ;
        RECT 823.950 261.600 826.050 262.050 ;
        RECT 700.950 260.400 826.050 261.600 ;
        RECT 700.950 259.950 703.050 260.400 ;
        RECT 823.950 259.950 826.050 260.400 ;
        RECT 214.950 258.600 217.050 259.050 ;
        RECT 262.950 258.600 265.050 259.050 ;
        RECT 274.950 258.600 277.050 259.050 ;
        RECT 214.950 257.400 277.050 258.600 ;
        RECT 214.950 256.950 217.050 257.400 ;
        RECT 262.950 256.950 265.050 257.400 ;
        RECT 274.950 256.950 277.050 257.400 ;
        RECT 301.950 258.600 304.050 259.050 ;
        RECT 334.950 258.600 337.050 259.050 ;
        RECT 301.950 257.400 337.050 258.600 ;
        RECT 301.950 256.950 304.050 257.400 ;
        RECT 334.950 256.950 337.050 257.400 ;
        RECT 343.950 258.600 346.050 259.050 ;
        RECT 415.950 258.600 418.050 259.050 ;
        RECT 343.950 257.400 418.050 258.600 ;
        RECT 343.950 256.950 346.050 257.400 ;
        RECT 415.950 256.950 418.050 257.400 ;
        RECT 202.950 255.600 205.050 256.050 ;
        RECT 319.950 255.600 322.050 256.050 ;
        RECT 202.950 254.400 322.050 255.600 ;
        RECT 202.950 253.950 205.050 254.400 ;
        RECT 319.950 253.950 322.050 254.400 ;
        RECT 334.950 255.600 337.050 256.050 ;
        RECT 343.950 255.600 346.050 256.050 ;
        RECT 334.950 254.400 346.050 255.600 ;
        RECT 334.950 253.950 337.050 254.400 ;
        RECT 343.950 253.950 346.050 254.400 ;
        RECT 703.950 255.600 706.050 256.050 ;
        RECT 778.950 255.600 781.050 256.050 ;
        RECT 781.950 255.600 784.050 256.050 ;
        RECT 703.950 254.400 784.050 255.600 ;
        RECT 703.950 253.950 706.050 254.400 ;
        RECT 778.950 253.950 781.050 254.400 ;
        RECT 781.950 253.950 784.050 254.400 ;
        RECT 181.950 252.600 184.050 253.050 ;
        RECT 202.950 252.600 205.050 253.050 ;
        RECT 181.950 251.400 205.050 252.600 ;
        RECT 181.950 250.950 184.050 251.400 ;
        RECT 202.950 250.950 205.050 251.400 ;
        RECT 283.950 252.600 286.050 253.050 ;
        RECT 394.950 252.600 397.050 253.050 ;
        RECT 283.950 251.400 397.050 252.600 ;
        RECT 283.950 250.950 286.050 251.400 ;
        RECT 394.950 250.950 397.050 251.400 ;
        RECT 778.950 252.600 781.050 253.050 ;
        RECT 802.950 252.600 805.050 253.050 ;
        RECT 778.950 251.400 805.050 252.600 ;
        RECT 778.950 250.950 781.050 251.400 ;
        RECT 802.950 250.950 805.050 251.400 ;
        RECT 823.950 252.600 826.050 253.050 ;
        RECT 850.950 252.600 853.050 253.050 ;
        RECT 823.950 251.400 853.050 252.600 ;
        RECT 823.950 250.950 826.050 251.400 ;
        RECT 850.950 250.950 853.050 251.400 ;
        RECT 58.950 249.600 61.050 250.050 ;
        RECT 97.950 249.600 100.050 250.050 ;
        RECT 190.950 249.600 193.050 250.050 ;
        RECT 58.950 248.400 193.050 249.600 ;
        RECT 58.950 247.950 61.050 248.400 ;
        RECT 97.950 247.950 100.050 248.400 ;
        RECT 190.950 247.950 193.050 248.400 ;
        RECT 502.950 249.600 505.050 250.050 ;
        RECT 559.950 249.600 562.050 250.050 ;
        RECT 502.950 248.400 562.050 249.600 ;
        RECT 502.950 247.950 505.050 248.400 ;
        RECT 559.950 247.950 562.050 248.400 ;
        RECT 586.950 249.600 589.050 250.050 ;
        RECT 712.950 249.600 715.050 250.050 ;
        RECT 754.950 249.600 757.050 250.050 ;
        RECT 772.950 249.600 775.050 250.050 ;
        RECT 586.950 248.400 775.050 249.600 ;
        RECT 586.950 247.950 589.050 248.400 ;
        RECT 712.950 247.950 715.050 248.400 ;
        RECT 754.950 247.950 757.050 248.400 ;
        RECT 772.950 247.950 775.050 248.400 ;
        RECT 52.950 246.600 55.050 247.050 ;
        RECT 91.950 246.600 94.050 247.050 ;
        RECT 109.950 246.600 112.050 247.050 ;
        RECT 52.950 245.400 112.050 246.600 ;
        RECT 52.950 244.950 55.050 245.400 ;
        RECT 91.950 244.950 94.050 245.400 ;
        RECT 109.950 244.950 112.050 245.400 ;
        RECT 112.950 246.600 115.050 247.050 ;
        RECT 136.950 246.600 139.050 247.050 ;
        RECT 217.950 246.600 220.050 247.050 ;
        RECT 112.950 245.400 220.050 246.600 ;
        RECT 112.950 244.950 115.050 245.400 ;
        RECT 136.950 244.950 139.050 245.400 ;
        RECT 217.950 244.950 220.050 245.400 ;
        RECT 244.950 246.600 247.050 247.050 ;
        RECT 259.950 246.600 262.050 247.050 ;
        RECT 244.950 245.400 262.050 246.600 ;
        RECT 244.950 244.950 247.050 245.400 ;
        RECT 259.950 244.950 262.050 245.400 ;
        RECT 271.950 246.600 274.050 247.050 ;
        RECT 286.950 246.600 289.050 247.050 ;
        RECT 295.950 246.600 298.050 247.050 ;
        RECT 271.950 245.400 298.050 246.600 ;
        RECT 271.950 244.950 274.050 245.400 ;
        RECT 286.950 244.950 289.050 245.400 ;
        RECT 295.950 244.950 298.050 245.400 ;
        RECT 337.950 246.600 340.050 247.050 ;
        RECT 361.950 246.600 364.050 247.050 ;
        RECT 337.950 245.400 364.050 246.600 ;
        RECT 337.950 244.950 340.050 245.400 ;
        RECT 361.950 244.950 364.050 245.400 ;
        RECT 367.950 246.600 370.050 247.050 ;
        RECT 376.950 246.600 379.050 247.050 ;
        RECT 367.950 245.400 379.050 246.600 ;
        RECT 367.950 244.950 370.050 245.400 ;
        RECT 376.950 244.950 379.050 245.400 ;
        RECT 388.950 246.600 391.050 247.050 ;
        RECT 433.950 246.600 436.050 247.050 ;
        RECT 451.950 246.600 454.050 247.050 ;
        RECT 520.950 246.600 523.050 247.050 ;
        RECT 388.950 245.400 523.050 246.600 ;
        RECT 388.950 244.950 391.050 245.400 ;
        RECT 433.950 244.950 436.050 245.400 ;
        RECT 451.950 244.950 454.050 245.400 ;
        RECT 520.950 244.950 523.050 245.400 ;
        RECT 565.950 246.600 568.050 247.050 ;
        RECT 604.950 246.600 607.050 247.050 ;
        RECT 565.950 245.400 607.050 246.600 ;
        RECT 565.950 244.950 568.050 245.400 ;
        RECT 604.950 244.950 607.050 245.400 ;
        RECT 775.950 246.600 778.050 247.050 ;
        RECT 787.950 246.600 790.050 247.050 ;
        RECT 775.950 245.400 790.050 246.600 ;
        RECT 775.950 244.950 778.050 245.400 ;
        RECT 787.950 244.950 790.050 245.400 ;
        RECT 865.950 246.600 868.050 247.050 ;
        RECT 865.950 245.400 873.600 246.600 ;
        RECT 865.950 244.950 868.050 245.400 ;
        RECT 55.950 243.600 58.050 244.050 ;
        RECT 64.950 243.600 67.050 244.050 ;
        RECT 55.950 242.400 67.050 243.600 ;
        RECT 55.950 241.950 58.050 242.400 ;
        RECT 64.950 241.950 67.050 242.400 ;
        RECT 94.950 243.600 97.050 244.050 ;
        RECT 106.950 243.600 109.050 244.050 ;
        RECT 94.950 242.400 109.050 243.600 ;
        RECT 94.950 241.950 97.050 242.400 ;
        RECT 106.950 241.950 109.050 242.400 ;
        RECT 121.950 243.600 124.050 244.050 ;
        RECT 139.950 243.600 142.050 244.050 ;
        RECT 121.950 242.400 142.050 243.600 ;
        RECT 121.950 241.950 124.050 242.400 ;
        RECT 139.950 241.950 142.050 242.400 ;
        RECT 148.950 243.600 151.050 244.050 ;
        RECT 166.950 243.600 169.050 244.050 ;
        RECT 148.950 242.400 169.050 243.600 ;
        RECT 148.950 241.950 151.050 242.400 ;
        RECT 166.950 241.950 169.050 242.400 ;
        RECT 190.950 243.600 193.050 244.050 ;
        RECT 220.950 243.600 223.050 244.050 ;
        RECT 190.950 242.400 223.050 243.600 ;
        RECT 190.950 241.950 193.050 242.400 ;
        RECT 220.950 241.950 223.050 242.400 ;
        RECT 235.950 243.600 238.050 244.050 ;
        RECT 277.950 243.600 280.050 244.050 ;
        RECT 280.950 243.600 283.050 244.050 ;
        RECT 286.950 243.600 289.050 244.050 ;
        RECT 235.950 242.400 289.050 243.600 ;
        RECT 235.950 241.950 238.050 242.400 ;
        RECT 277.950 241.950 280.050 242.400 ;
        RECT 280.950 241.950 283.050 242.400 ;
        RECT 286.950 241.950 289.050 242.400 ;
        RECT 313.950 243.600 316.050 244.050 ;
        RECT 439.950 243.600 442.050 244.050 ;
        RECT 475.950 243.600 478.050 244.050 ;
        RECT 481.950 243.600 484.050 244.050 ;
        RECT 313.950 242.400 484.050 243.600 ;
        RECT 313.950 241.950 316.050 242.400 ;
        RECT 439.950 241.950 442.050 242.400 ;
        RECT 475.950 241.950 478.050 242.400 ;
        RECT 481.950 241.950 484.050 242.400 ;
        RECT 499.950 243.600 502.050 244.050 ;
        RECT 532.950 243.600 535.050 244.050 ;
        RECT 544.950 243.600 547.050 244.050 ;
        RECT 550.950 243.600 553.050 244.050 ;
        RECT 499.950 242.400 553.050 243.600 ;
        RECT 499.950 241.950 502.050 242.400 ;
        RECT 532.950 241.950 535.050 242.400 ;
        RECT 544.950 241.950 547.050 242.400 ;
        RECT 550.950 241.950 553.050 242.400 ;
        RECT 562.950 243.600 565.050 244.050 ;
        RECT 580.950 243.600 583.050 244.050 ;
        RECT 562.950 242.400 583.050 243.600 ;
        RECT 562.950 241.950 565.050 242.400 ;
        RECT 580.950 241.950 583.050 242.400 ;
        RECT 598.950 243.600 601.050 244.050 ;
        RECT 652.950 243.600 655.050 244.050 ;
        RECT 598.950 242.400 655.050 243.600 ;
        RECT 598.950 241.950 601.050 242.400 ;
        RECT 652.950 241.950 655.050 242.400 ;
        RECT 667.950 243.600 670.050 244.050 ;
        RECT 679.950 243.600 682.050 244.050 ;
        RECT 667.950 242.400 682.050 243.600 ;
        RECT 667.950 241.950 670.050 242.400 ;
        RECT 679.950 241.950 682.050 242.400 ;
        RECT 688.950 243.600 691.050 244.050 ;
        RECT 796.950 243.600 799.050 244.050 ;
        RECT 688.950 242.400 799.050 243.600 ;
        RECT 688.950 241.950 691.050 242.400 ;
        RECT 796.950 241.950 799.050 242.400 ;
        RECT 805.950 243.600 808.050 244.050 ;
        RECT 820.950 243.600 823.050 244.050 ;
        RECT 805.950 242.400 823.050 243.600 ;
        RECT 805.950 241.950 808.050 242.400 ;
        RECT 820.950 241.950 823.050 242.400 ;
        RECT 829.950 243.600 832.050 244.050 ;
        RECT 868.950 243.600 871.050 244.050 ;
        RECT 829.950 242.400 871.050 243.600 ;
        RECT 829.950 241.950 832.050 242.400 ;
        RECT 868.950 241.950 871.050 242.400 ;
        RECT 19.950 240.600 22.050 241.050 ;
        RECT 28.950 240.600 31.050 241.050 ;
        RECT 52.950 240.600 55.050 241.050 ;
        RECT 19.950 239.400 55.050 240.600 ;
        RECT 19.950 238.950 22.050 239.400 ;
        RECT 28.950 238.950 31.050 239.400 ;
        RECT 52.950 238.950 55.050 239.400 ;
        RECT 61.950 240.600 64.050 241.050 ;
        RECT 79.950 240.600 82.050 241.050 ;
        RECT 124.950 240.600 127.050 241.050 ;
        RECT 61.950 239.400 127.050 240.600 ;
        RECT 61.950 238.950 64.050 239.400 ;
        RECT 79.950 238.950 82.050 239.400 ;
        RECT 124.950 238.950 127.050 239.400 ;
        RECT 133.950 240.600 136.050 241.050 ;
        RECT 148.950 240.600 151.050 241.050 ;
        RECT 133.950 239.400 151.050 240.600 ;
        RECT 133.950 238.950 136.050 239.400 ;
        RECT 148.950 238.950 151.050 239.400 ;
        RECT 154.950 240.600 157.050 241.050 ;
        RECT 223.950 240.600 226.050 241.050 ;
        RECT 229.950 240.600 232.050 241.050 ;
        RECT 154.950 239.400 222.600 240.600 ;
        RECT 154.950 238.950 157.050 239.400 ;
        RECT 4.950 237.600 7.050 238.050 ;
        RECT 10.950 237.600 13.050 238.050 ;
        RECT 4.950 236.400 13.050 237.600 ;
        RECT 4.950 235.950 7.050 236.400 ;
        RECT 10.950 235.950 13.050 236.400 ;
        RECT 16.950 237.600 19.050 238.050 ;
        RECT 40.950 237.600 43.050 238.050 ;
        RECT 16.950 236.400 43.050 237.600 ;
        RECT 16.950 235.950 19.050 236.400 ;
        RECT 40.950 235.950 43.050 236.400 ;
        RECT 55.950 237.600 58.050 238.050 ;
        RECT 70.950 237.600 73.050 238.050 ;
        RECT 55.950 236.400 73.050 237.600 ;
        RECT 55.950 235.950 58.050 236.400 ;
        RECT 70.950 235.950 73.050 236.400 ;
        RECT 115.950 237.600 118.050 238.050 ;
        RECT 130.950 237.600 133.050 238.050 ;
        RECT 115.950 236.400 133.050 237.600 ;
        RECT 115.950 235.950 118.050 236.400 ;
        RECT 130.950 235.950 133.050 236.400 ;
        RECT 136.950 237.600 139.050 238.050 ;
        RECT 175.950 237.600 178.050 238.050 ;
        RECT 136.950 236.400 178.050 237.600 ;
        RECT 136.950 235.950 139.050 236.400 ;
        RECT 175.950 235.950 178.050 236.400 ;
        RECT 208.950 237.600 211.050 238.050 ;
        RECT 214.950 237.600 217.050 238.050 ;
        RECT 208.950 236.400 217.050 237.600 ;
        RECT 221.400 237.600 222.600 239.400 ;
        RECT 223.950 239.400 232.050 240.600 ;
        RECT 223.950 238.950 226.050 239.400 ;
        RECT 229.950 238.950 232.050 239.400 ;
        RECT 250.950 240.600 253.050 241.050 ;
        RECT 277.950 240.600 280.050 241.050 ;
        RECT 250.950 239.400 280.050 240.600 ;
        RECT 250.950 238.950 253.050 239.400 ;
        RECT 277.950 238.950 280.050 239.400 ;
        RECT 292.950 240.600 295.050 241.050 ;
        RECT 319.950 240.600 322.050 241.050 ;
        RECT 328.950 240.600 331.050 241.050 ;
        RECT 292.950 239.400 331.050 240.600 ;
        RECT 292.950 238.950 295.050 239.400 ;
        RECT 319.950 238.950 322.050 239.400 ;
        RECT 328.950 238.950 331.050 239.400 ;
        RECT 331.950 240.600 334.050 241.050 ;
        RECT 346.950 240.600 349.050 241.050 ;
        RECT 331.950 239.400 349.050 240.600 ;
        RECT 331.950 238.950 334.050 239.400 ;
        RECT 346.950 238.950 349.050 239.400 ;
        RECT 355.950 240.600 358.050 241.050 ;
        RECT 364.950 240.600 367.050 241.050 ;
        RECT 355.950 239.400 367.050 240.600 ;
        RECT 355.950 238.950 358.050 239.400 ;
        RECT 364.950 238.950 367.050 239.400 ;
        RECT 382.950 240.600 385.050 241.050 ;
        RECT 457.950 240.600 460.050 241.050 ;
        RECT 463.950 240.600 466.050 241.050 ;
        RECT 382.950 239.400 466.050 240.600 ;
        RECT 382.950 238.950 385.050 239.400 ;
        RECT 457.950 238.950 460.050 239.400 ;
        RECT 463.950 238.950 466.050 239.400 ;
        RECT 469.950 240.600 472.050 241.050 ;
        RECT 478.950 240.600 481.050 241.050 ;
        RECT 469.950 239.400 481.050 240.600 ;
        RECT 469.950 238.950 472.050 239.400 ;
        RECT 478.950 238.950 481.050 239.400 ;
        RECT 484.950 240.600 487.050 241.050 ;
        RECT 562.950 240.600 565.050 241.050 ;
        RECT 484.950 239.400 565.050 240.600 ;
        RECT 484.950 238.950 487.050 239.400 ;
        RECT 562.950 238.950 565.050 239.400 ;
        RECT 589.950 240.600 592.050 241.050 ;
        RECT 622.950 240.600 625.050 241.050 ;
        RECT 589.950 239.400 625.050 240.600 ;
        RECT 589.950 238.950 592.050 239.400 ;
        RECT 622.950 238.950 625.050 239.400 ;
        RECT 628.950 240.600 631.050 241.050 ;
        RECT 658.950 240.600 661.050 241.050 ;
        RECT 628.950 239.400 661.050 240.600 ;
        RECT 628.950 238.950 631.050 239.400 ;
        RECT 658.950 238.950 661.050 239.400 ;
        RECT 718.950 238.950 721.050 241.050 ;
        RECT 724.950 240.600 727.050 241.050 ;
        RECT 745.950 240.600 748.050 241.050 ;
        RECT 724.950 239.400 748.050 240.600 ;
        RECT 724.950 238.950 727.050 239.400 ;
        RECT 745.950 238.950 748.050 239.400 ;
        RECT 799.950 238.950 802.050 241.050 ;
        RECT 802.950 240.600 805.050 241.050 ;
        RECT 817.950 240.600 820.050 241.050 ;
        RECT 802.950 239.400 820.050 240.600 ;
        RECT 802.950 238.950 805.050 239.400 ;
        RECT 817.950 238.950 820.050 239.400 ;
        RECT 838.950 240.600 841.050 241.050 ;
        RECT 838.950 239.400 861.600 240.600 ;
        RECT 838.950 238.950 841.050 239.400 ;
        RECT 226.950 237.600 229.050 238.050 ;
        RECT 221.400 236.400 229.050 237.600 ;
        RECT 208.950 235.950 211.050 236.400 ;
        RECT 214.950 235.950 217.050 236.400 ;
        RECT 226.950 235.950 229.050 236.400 ;
        RECT 232.950 237.600 235.050 238.050 ;
        RECT 238.950 237.600 241.050 238.050 ;
        RECT 232.950 236.400 241.050 237.600 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 238.950 235.950 241.050 236.400 ;
        RECT 241.950 237.600 244.050 238.050 ;
        RECT 247.950 237.600 250.050 238.050 ;
        RECT 241.950 236.400 250.050 237.600 ;
        RECT 241.950 235.950 244.050 236.400 ;
        RECT 247.950 235.950 250.050 236.400 ;
        RECT 253.950 237.600 256.050 238.050 ;
        RECT 268.950 237.600 271.050 238.050 ;
        RECT 253.950 236.400 271.050 237.600 ;
        RECT 253.950 235.950 256.050 236.400 ;
        RECT 268.950 235.950 271.050 236.400 ;
        RECT 289.950 237.600 292.050 238.050 ;
        RECT 295.950 237.600 298.050 238.050 ;
        RECT 289.950 236.400 298.050 237.600 ;
        RECT 289.950 235.950 292.050 236.400 ;
        RECT 295.950 235.950 298.050 236.400 ;
        RECT 334.950 237.600 337.050 238.050 ;
        RECT 349.950 237.600 352.050 238.050 ;
        RECT 334.950 236.400 352.050 237.600 ;
        RECT 365.400 237.600 366.600 238.950 ;
        RECT 388.950 237.600 391.050 238.050 ;
        RECT 400.950 237.600 403.050 238.050 ;
        RECT 365.400 236.400 403.050 237.600 ;
        RECT 334.950 235.950 337.050 236.400 ;
        RECT 349.950 235.950 352.050 236.400 ;
        RECT 388.950 235.950 391.050 236.400 ;
        RECT 400.950 235.950 403.050 236.400 ;
        RECT 409.950 237.600 412.050 238.050 ;
        RECT 445.950 237.600 448.050 238.050 ;
        RECT 409.950 236.400 448.050 237.600 ;
        RECT 409.950 235.950 412.050 236.400 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 448.950 237.600 451.050 238.050 ;
        RECT 457.950 237.600 460.050 238.050 ;
        RECT 448.950 236.400 460.050 237.600 ;
        RECT 448.950 235.950 451.050 236.400 ;
        RECT 457.950 235.950 460.050 236.400 ;
        RECT 463.950 237.600 466.050 238.050 ;
        RECT 472.950 237.600 475.050 238.050 ;
        RECT 463.950 236.400 475.050 237.600 ;
        RECT 463.950 235.950 466.050 236.400 ;
        RECT 472.950 235.950 475.050 236.400 ;
        RECT 508.950 237.600 511.050 238.050 ;
        RECT 517.950 237.600 520.050 238.050 ;
        RECT 508.950 236.400 520.050 237.600 ;
        RECT 508.950 235.950 511.050 236.400 ;
        RECT 517.950 235.950 520.050 236.400 ;
        RECT 535.950 235.950 538.050 238.050 ;
        RECT 559.950 237.600 562.050 238.050 ;
        RECT 565.950 237.600 568.050 238.050 ;
        RECT 583.950 237.600 586.050 238.050 ;
        RECT 610.950 237.600 613.050 238.050 ;
        RECT 559.950 236.400 564.600 237.600 ;
        RECT 559.950 235.950 562.050 236.400 ;
        RECT 37.950 234.600 40.050 235.050 ;
        RECT 52.950 234.600 55.050 235.050 ;
        RECT 73.950 234.600 76.050 235.050 ;
        RECT 37.950 233.400 76.050 234.600 ;
        RECT 37.950 232.950 40.050 233.400 ;
        RECT 52.950 232.950 55.050 233.400 ;
        RECT 73.950 232.950 76.050 233.400 ;
        RECT 88.950 234.600 91.050 235.050 ;
        RECT 112.950 234.600 115.050 235.050 ;
        RECT 88.950 233.400 115.050 234.600 ;
        RECT 88.950 232.950 91.050 233.400 ;
        RECT 112.950 232.950 115.050 233.400 ;
        RECT 196.950 234.600 199.050 235.050 ;
        RECT 283.950 234.600 286.050 235.050 ;
        RECT 196.950 233.400 286.050 234.600 ;
        RECT 196.950 232.950 199.050 233.400 ;
        RECT 283.950 232.950 286.050 233.400 ;
        RECT 313.950 234.600 316.050 235.050 ;
        RECT 319.950 234.600 322.050 235.050 ;
        RECT 313.950 233.400 322.050 234.600 ;
        RECT 313.950 232.950 316.050 233.400 ;
        RECT 319.950 232.950 322.050 233.400 ;
        RECT 373.950 234.600 376.050 235.050 ;
        RECT 385.950 234.600 388.050 235.050 ;
        RECT 373.950 233.400 388.050 234.600 ;
        RECT 373.950 232.950 376.050 233.400 ;
        RECT 385.950 232.950 388.050 233.400 ;
        RECT 391.950 234.600 394.050 235.050 ;
        RECT 406.950 234.600 409.050 235.050 ;
        RECT 391.950 233.400 409.050 234.600 ;
        RECT 391.950 232.950 394.050 233.400 ;
        RECT 406.950 232.950 409.050 233.400 ;
        RECT 436.950 234.600 439.050 235.050 ;
        RECT 460.950 234.600 463.050 235.050 ;
        RECT 487.950 234.600 490.050 235.050 ;
        RECT 436.950 233.400 490.050 234.600 ;
        RECT 536.400 234.600 537.600 235.950 ;
        RECT 538.950 234.600 541.050 235.050 ;
        RECT 536.400 233.400 541.050 234.600 ;
        RECT 563.400 234.600 564.600 236.400 ;
        RECT 565.950 236.400 613.050 237.600 ;
        RECT 565.950 235.950 568.050 236.400 ;
        RECT 583.950 235.950 586.050 236.400 ;
        RECT 610.950 235.950 613.050 236.400 ;
        RECT 661.950 237.600 664.050 238.050 ;
        RECT 697.950 237.600 700.050 238.050 ;
        RECT 661.950 236.400 700.050 237.600 ;
        RECT 661.950 235.950 664.050 236.400 ;
        RECT 697.950 235.950 700.050 236.400 ;
        RECT 703.950 237.600 706.050 238.050 ;
        RECT 715.950 237.600 718.050 238.050 ;
        RECT 703.950 236.400 718.050 237.600 ;
        RECT 703.950 235.950 706.050 236.400 ;
        RECT 715.950 235.950 718.050 236.400 ;
        RECT 719.400 235.050 720.600 238.950 ;
        RECT 736.950 237.600 739.050 238.050 ;
        RECT 748.950 237.600 751.050 238.050 ;
        RECT 775.950 237.600 778.050 238.050 ;
        RECT 736.950 236.400 778.050 237.600 ;
        RECT 800.400 237.600 801.600 238.950 ;
        RECT 860.400 238.050 861.600 239.400 ;
        RECT 838.950 237.600 841.050 238.050 ;
        RECT 859.950 237.600 862.050 238.050 ;
        RECT 800.400 236.400 841.050 237.600 ;
        RECT 736.950 235.950 739.050 236.400 ;
        RECT 748.950 235.950 751.050 236.400 ;
        RECT 775.950 235.950 778.050 236.400 ;
        RECT 838.950 235.950 841.050 236.400 ;
        RECT 842.400 236.400 862.050 237.600 ;
        RECT 577.950 234.600 580.050 235.050 ;
        RECT 563.400 233.400 580.050 234.600 ;
        RECT 436.950 232.950 439.050 233.400 ;
        RECT 460.950 232.950 463.050 233.400 ;
        RECT 487.950 232.950 490.050 233.400 ;
        RECT 538.950 232.950 541.050 233.400 ;
        RECT 577.950 232.950 580.050 233.400 ;
        RECT 649.950 234.600 652.050 235.050 ;
        RECT 664.950 234.600 667.050 235.050 ;
        RECT 676.950 234.600 679.050 235.050 ;
        RECT 649.950 233.400 679.050 234.600 ;
        RECT 649.950 232.950 652.050 233.400 ;
        RECT 664.950 232.950 667.050 233.400 ;
        RECT 676.950 232.950 679.050 233.400 ;
        RECT 718.950 232.950 721.050 235.050 ;
        RECT 739.950 234.600 742.050 235.050 ;
        RECT 799.950 234.600 802.050 235.050 ;
        RECT 811.950 234.600 814.050 235.050 ;
        RECT 739.950 233.400 814.050 234.600 ;
        RECT 739.950 232.950 742.050 233.400 ;
        RECT 799.950 232.950 802.050 233.400 ;
        RECT 811.950 232.950 814.050 233.400 ;
        RECT 835.950 234.600 838.050 235.050 ;
        RECT 842.400 234.600 843.600 236.400 ;
        RECT 859.950 235.950 862.050 236.400 ;
        RECT 835.950 233.400 843.600 234.600 ;
        RECT 859.950 234.600 862.050 235.050 ;
        RECT 865.950 234.600 868.050 235.050 ;
        RECT 859.950 233.400 868.050 234.600 ;
        RECT 835.950 232.950 838.050 233.400 ;
        RECT 859.950 232.950 862.050 233.400 ;
        RECT 865.950 232.950 868.050 233.400 ;
        RECT 106.950 231.600 109.050 232.050 ;
        RECT 187.950 231.600 190.050 232.050 ;
        RECT 196.950 231.600 199.050 232.050 ;
        RECT 106.950 230.400 199.050 231.600 ;
        RECT 106.950 229.950 109.050 230.400 ;
        RECT 187.950 229.950 190.050 230.400 ;
        RECT 196.950 229.950 199.050 230.400 ;
        RECT 277.950 231.600 280.050 232.050 ;
        RECT 373.950 231.600 376.050 232.050 ;
        RECT 277.950 230.400 376.050 231.600 ;
        RECT 277.950 229.950 280.050 230.400 ;
        RECT 373.950 229.950 376.050 230.400 ;
        RECT 400.950 231.600 403.050 232.050 ;
        RECT 430.950 231.600 433.050 232.050 ;
        RECT 400.950 230.400 433.050 231.600 ;
        RECT 400.950 229.950 403.050 230.400 ;
        RECT 430.950 229.950 433.050 230.400 ;
        RECT 457.950 231.600 460.050 232.050 ;
        RECT 463.950 231.600 466.050 232.050 ;
        RECT 457.950 230.400 466.050 231.600 ;
        RECT 457.950 229.950 460.050 230.400 ;
        RECT 463.950 229.950 466.050 230.400 ;
        RECT 556.950 231.600 559.050 232.050 ;
        RECT 724.950 231.600 727.050 232.050 ;
        RECT 730.950 231.600 733.050 232.050 ;
        RECT 556.950 230.400 733.050 231.600 ;
        RECT 556.950 229.950 559.050 230.400 ;
        RECT 724.950 229.950 727.050 230.400 ;
        RECT 730.950 229.950 733.050 230.400 ;
        RECT 862.950 231.600 865.050 232.050 ;
        RECT 872.400 231.600 873.600 245.400 ;
        RECT 862.950 230.400 873.600 231.600 ;
        RECT 862.950 229.950 865.050 230.400 ;
        RECT 25.950 228.600 28.050 229.050 ;
        RECT 76.950 228.600 79.050 229.050 ;
        RECT 118.950 228.600 121.050 229.050 ;
        RECT 25.950 227.400 121.050 228.600 ;
        RECT 25.950 226.950 28.050 227.400 ;
        RECT 76.950 226.950 79.050 227.400 ;
        RECT 118.950 226.950 121.050 227.400 ;
        RECT 211.950 228.600 214.050 229.050 ;
        RECT 235.950 228.600 238.050 229.050 ;
        RECT 259.950 228.600 262.050 229.050 ;
        RECT 211.950 227.400 262.050 228.600 ;
        RECT 211.950 226.950 214.050 227.400 ;
        RECT 235.950 226.950 238.050 227.400 ;
        RECT 259.950 226.950 262.050 227.400 ;
        RECT 346.950 228.600 349.050 229.050 ;
        RECT 412.950 228.600 415.050 229.050 ;
        RECT 346.950 227.400 415.050 228.600 ;
        RECT 346.950 226.950 349.050 227.400 ;
        RECT 412.950 226.950 415.050 227.400 ;
        RECT 448.950 228.600 451.050 229.050 ;
        RECT 469.950 228.600 472.050 229.050 ;
        RECT 448.950 227.400 472.050 228.600 ;
        RECT 448.950 226.950 451.050 227.400 ;
        RECT 469.950 226.950 472.050 227.400 ;
        RECT 547.950 228.600 550.050 229.050 ;
        RECT 610.950 228.600 613.050 229.050 ;
        RECT 547.950 227.400 613.050 228.600 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 610.950 226.950 613.050 227.400 ;
        RECT 655.950 228.600 658.050 229.050 ;
        RECT 700.950 228.600 703.050 229.050 ;
        RECT 829.950 228.600 832.050 229.050 ;
        RECT 655.950 227.400 832.050 228.600 ;
        RECT 655.950 226.950 658.050 227.400 ;
        RECT 700.950 226.950 703.050 227.400 ;
        RECT 829.950 226.950 832.050 227.400 ;
        RECT 211.950 225.600 214.050 226.050 ;
        RECT 256.950 225.600 259.050 226.050 ;
        RECT 211.950 224.400 259.050 225.600 ;
        RECT 211.950 223.950 214.050 224.400 ;
        RECT 256.950 223.950 259.050 224.400 ;
        RECT 541.950 216.600 544.050 217.050 ;
        RECT 661.950 216.600 664.050 217.050 ;
        RECT 541.950 215.400 664.050 216.600 ;
        RECT 541.950 214.950 544.050 215.400 ;
        RECT 661.950 214.950 664.050 215.400 ;
        RECT 355.950 213.600 358.050 214.050 ;
        RECT 361.950 213.600 364.050 214.050 ;
        RECT 355.950 212.400 364.050 213.600 ;
        RECT 355.950 211.950 358.050 212.400 ;
        RECT 361.950 211.950 364.050 212.400 ;
        RECT 163.950 210.600 166.050 211.050 ;
        RECT 241.950 210.600 244.050 211.050 ;
        RECT 163.950 209.400 244.050 210.600 ;
        RECT 163.950 208.950 166.050 209.400 ;
        RECT 241.950 208.950 244.050 209.400 ;
        RECT 493.950 210.600 496.050 211.050 ;
        RECT 532.950 210.600 535.050 211.050 ;
        RECT 619.950 210.600 622.050 211.050 ;
        RECT 493.950 209.400 622.050 210.600 ;
        RECT 493.950 208.950 496.050 209.400 ;
        RECT 532.950 208.950 535.050 209.400 ;
        RECT 619.950 208.950 622.050 209.400 ;
        RECT 769.950 210.600 772.050 211.050 ;
        RECT 799.950 210.600 802.050 211.050 ;
        RECT 769.950 209.400 802.050 210.600 ;
        RECT 769.950 208.950 772.050 209.400 ;
        RECT 799.950 208.950 802.050 209.400 ;
        RECT 223.950 207.600 226.050 208.050 ;
        RECT 292.950 207.600 295.050 208.050 ;
        RECT 223.950 206.400 295.050 207.600 ;
        RECT 223.950 205.950 226.050 206.400 ;
        RECT 292.950 205.950 295.050 206.400 ;
        RECT 301.950 207.600 304.050 208.050 ;
        RECT 307.950 207.600 310.050 208.050 ;
        RECT 301.950 206.400 310.050 207.600 ;
        RECT 301.950 205.950 304.050 206.400 ;
        RECT 307.950 205.950 310.050 206.400 ;
        RECT 445.950 207.600 448.050 208.050 ;
        RECT 652.950 207.600 655.050 208.050 ;
        RECT 445.950 206.400 655.050 207.600 ;
        RECT 445.950 205.950 448.050 206.400 ;
        RECT 652.950 205.950 655.050 206.400 ;
        RECT 736.950 207.600 739.050 208.050 ;
        RECT 742.950 207.600 745.050 208.050 ;
        RECT 814.950 207.600 817.050 208.050 ;
        RECT 736.950 206.400 817.050 207.600 ;
        RECT 736.950 205.950 739.050 206.400 ;
        RECT 742.950 205.950 745.050 206.400 ;
        RECT 814.950 205.950 817.050 206.400 ;
        RECT 505.950 204.600 508.050 205.050 ;
        RECT 514.950 204.600 517.050 205.050 ;
        RECT 580.950 204.600 583.050 205.050 ;
        RECT 607.950 204.600 610.050 205.050 ;
        RECT 505.950 203.400 610.050 204.600 ;
        RECT 505.950 202.950 508.050 203.400 ;
        RECT 514.950 202.950 517.050 203.400 ;
        RECT 580.950 202.950 583.050 203.400 ;
        RECT 607.950 202.950 610.050 203.400 ;
        RECT 676.950 204.600 679.050 205.050 ;
        RECT 700.950 204.600 703.050 205.050 ;
        RECT 676.950 203.400 703.050 204.600 ;
        RECT 676.950 202.950 679.050 203.400 ;
        RECT 700.950 202.950 703.050 203.400 ;
        RECT 778.950 204.600 781.050 205.050 ;
        RECT 817.950 204.600 820.050 205.050 ;
        RECT 778.950 203.400 820.050 204.600 ;
        RECT 778.950 202.950 781.050 203.400 ;
        RECT 817.950 202.950 820.050 203.400 ;
        RECT 112.950 201.600 115.050 202.050 ;
        RECT 142.950 201.600 145.050 202.050 ;
        RECT 112.950 200.400 145.050 201.600 ;
        RECT 112.950 199.950 115.050 200.400 ;
        RECT 142.950 199.950 145.050 200.400 ;
        RECT 145.950 199.950 148.050 202.050 ;
        RECT 181.950 201.600 184.050 202.050 ;
        RECT 187.950 201.600 190.050 202.050 ;
        RECT 181.950 200.400 190.050 201.600 ;
        RECT 181.950 199.950 184.050 200.400 ;
        RECT 187.950 199.950 190.050 200.400 ;
        RECT 214.950 201.600 217.050 202.050 ;
        RECT 304.950 201.600 307.050 202.050 ;
        RECT 328.950 201.600 331.050 202.050 ;
        RECT 424.950 201.600 427.050 202.050 ;
        RECT 448.950 201.600 451.050 202.050 ;
        RECT 214.950 200.400 225.600 201.600 ;
        RECT 214.950 199.950 217.050 200.400 ;
        RECT 4.950 198.600 7.050 199.050 ;
        RECT 13.950 198.600 16.050 199.050 ;
        RECT 4.950 197.400 16.050 198.600 ;
        RECT 4.950 196.950 7.050 197.400 ;
        RECT 13.950 196.950 16.050 197.400 ;
        RECT 22.950 198.600 25.050 199.050 ;
        RECT 28.950 198.600 31.050 199.050 ;
        RECT 52.950 198.600 55.050 199.050 ;
        RECT 64.950 198.600 67.050 199.050 ;
        RECT 22.950 197.400 51.600 198.600 ;
        RECT 22.950 196.950 25.050 197.400 ;
        RECT 28.950 196.950 31.050 197.400 ;
        RECT 50.400 195.600 51.600 197.400 ;
        RECT 52.950 197.400 67.050 198.600 ;
        RECT 52.950 196.950 55.050 197.400 ;
        RECT 64.950 196.950 67.050 197.400 ;
        RECT 121.950 198.600 124.050 199.050 ;
        RECT 136.950 198.600 139.050 199.050 ;
        RECT 121.950 197.400 139.050 198.600 ;
        RECT 121.950 196.950 124.050 197.400 ;
        RECT 136.950 196.950 139.050 197.400 ;
        RECT 85.950 195.600 88.050 196.050 ;
        RECT 50.400 194.400 88.050 195.600 ;
        RECT 85.950 193.950 88.050 194.400 ;
        RECT 139.950 195.600 142.050 196.050 ;
        RECT 146.400 195.600 147.600 199.950 ;
        RECT 224.400 199.050 225.600 200.400 ;
        RECT 304.950 200.400 451.050 201.600 ;
        RECT 304.950 199.950 307.050 200.400 ;
        RECT 328.950 199.950 331.050 200.400 ;
        RECT 424.950 199.950 427.050 200.400 ;
        RECT 448.950 199.950 451.050 200.400 ;
        RECT 463.950 201.600 466.050 202.050 ;
        RECT 472.950 201.600 475.050 202.050 ;
        RECT 463.950 200.400 475.050 201.600 ;
        RECT 463.950 199.950 466.050 200.400 ;
        RECT 472.950 199.950 475.050 200.400 ;
        RECT 475.950 201.600 478.050 202.050 ;
        RECT 487.950 201.600 490.050 202.050 ;
        RECT 475.950 200.400 490.050 201.600 ;
        RECT 475.950 199.950 478.050 200.400 ;
        RECT 487.950 199.950 490.050 200.400 ;
        RECT 508.950 201.600 511.050 202.050 ;
        RECT 526.950 201.600 529.050 202.050 ;
        RECT 535.950 201.600 538.050 202.050 ;
        RECT 508.950 200.400 513.600 201.600 ;
        RECT 508.950 199.950 511.050 200.400 ;
        RECT 512.400 199.050 513.600 200.400 ;
        RECT 526.950 200.400 538.050 201.600 ;
        RECT 526.950 199.950 529.050 200.400 ;
        RECT 535.950 199.950 538.050 200.400 ;
        RECT 763.950 201.600 766.050 202.050 ;
        RECT 781.950 201.600 784.050 202.050 ;
        RECT 763.950 200.400 784.050 201.600 ;
        RECT 763.950 199.950 766.050 200.400 ;
        RECT 781.950 199.950 784.050 200.400 ;
        RECT 784.950 201.600 787.050 202.050 ;
        RECT 790.950 201.600 793.050 202.050 ;
        RECT 784.950 200.400 793.050 201.600 ;
        RECT 784.950 199.950 787.050 200.400 ;
        RECT 790.950 199.950 793.050 200.400 ;
        RECT 796.950 201.600 799.050 202.050 ;
        RECT 802.950 201.600 805.050 202.050 ;
        RECT 796.950 200.400 805.050 201.600 ;
        RECT 796.950 199.950 799.050 200.400 ;
        RECT 802.950 199.950 805.050 200.400 ;
        RECT 811.950 201.600 814.050 202.050 ;
        RECT 832.950 201.600 835.050 202.050 ;
        RECT 811.950 200.400 835.050 201.600 ;
        RECT 811.950 199.950 814.050 200.400 ;
        RECT 832.950 199.950 835.050 200.400 ;
        RECT 169.950 198.600 172.050 199.050 ;
        RECT 178.950 198.600 181.050 199.050 ;
        RECT 169.950 197.400 181.050 198.600 ;
        RECT 169.950 196.950 172.050 197.400 ;
        RECT 178.950 196.950 181.050 197.400 ;
        RECT 184.950 198.600 187.050 199.050 ;
        RECT 202.950 198.600 205.050 199.050 ;
        RECT 184.950 197.400 205.050 198.600 ;
        RECT 184.950 196.950 187.050 197.400 ;
        RECT 202.950 196.950 205.050 197.400 ;
        RECT 223.950 196.950 226.050 199.050 ;
        RECT 247.950 198.600 250.050 199.050 ;
        RECT 262.950 198.600 265.050 199.050 ;
        RECT 247.950 197.400 265.050 198.600 ;
        RECT 247.950 196.950 250.050 197.400 ;
        RECT 262.950 196.950 265.050 197.400 ;
        RECT 307.950 198.600 310.050 199.050 ;
        RECT 322.950 198.600 325.050 199.050 ;
        RECT 307.950 197.400 325.050 198.600 ;
        RECT 307.950 196.950 310.050 197.400 ;
        RECT 322.950 196.950 325.050 197.400 ;
        RECT 385.950 198.600 388.050 199.050 ;
        RECT 400.950 198.600 403.050 199.050 ;
        RECT 385.950 197.400 403.050 198.600 ;
        RECT 385.950 196.950 388.050 197.400 ;
        RECT 400.950 196.950 403.050 197.400 ;
        RECT 406.950 198.600 409.050 199.050 ;
        RECT 415.950 198.600 418.050 199.050 ;
        RECT 406.950 197.400 418.050 198.600 ;
        RECT 406.950 196.950 409.050 197.400 ;
        RECT 415.950 196.950 418.050 197.400 ;
        RECT 430.950 198.600 433.050 199.050 ;
        RECT 445.950 198.600 448.050 199.050 ;
        RECT 430.950 197.400 448.050 198.600 ;
        RECT 430.950 196.950 433.050 197.400 ;
        RECT 445.950 196.950 448.050 197.400 ;
        RECT 469.950 198.600 472.050 199.050 ;
        RECT 490.950 198.600 493.050 199.050 ;
        RECT 469.950 197.400 493.050 198.600 ;
        RECT 469.950 196.950 472.050 197.400 ;
        RECT 490.950 196.950 493.050 197.400 ;
        RECT 511.950 196.950 514.050 199.050 ;
        RECT 529.950 198.600 532.050 199.050 ;
        RECT 538.950 198.600 541.050 199.050 ;
        RECT 529.950 197.400 541.050 198.600 ;
        RECT 529.950 196.950 532.050 197.400 ;
        RECT 538.950 196.950 541.050 197.400 ;
        RECT 544.950 198.600 547.050 199.050 ;
        RECT 571.950 198.600 574.050 199.050 ;
        RECT 574.950 198.600 577.050 199.050 ;
        RECT 544.950 197.400 577.050 198.600 ;
        RECT 544.950 196.950 547.050 197.400 ;
        RECT 571.950 196.950 574.050 197.400 ;
        RECT 574.950 196.950 577.050 197.400 ;
        RECT 586.950 198.600 589.050 199.050 ;
        RECT 604.950 198.600 607.050 199.050 ;
        RECT 586.950 197.400 607.050 198.600 ;
        RECT 586.950 196.950 589.050 197.400 ;
        RECT 604.950 196.950 607.050 197.400 ;
        RECT 610.950 198.600 613.050 199.050 ;
        RECT 622.950 198.600 625.050 199.050 ;
        RECT 610.950 197.400 625.050 198.600 ;
        RECT 610.950 196.950 613.050 197.400 ;
        RECT 622.950 196.950 625.050 197.400 ;
        RECT 637.950 198.600 640.050 199.050 ;
        RECT 646.950 198.600 649.050 199.050 ;
        RECT 637.950 197.400 649.050 198.600 ;
        RECT 637.950 196.950 640.050 197.400 ;
        RECT 646.950 196.950 649.050 197.400 ;
        RECT 661.950 198.600 664.050 199.050 ;
        RECT 670.950 198.600 673.050 199.050 ;
        RECT 661.950 197.400 673.050 198.600 ;
        RECT 661.950 196.950 664.050 197.400 ;
        RECT 670.950 196.950 673.050 197.400 ;
        RECT 682.950 198.600 685.050 199.050 ;
        RECT 697.950 198.600 700.050 199.050 ;
        RECT 682.950 197.400 700.050 198.600 ;
        RECT 682.950 196.950 685.050 197.400 ;
        RECT 697.950 196.950 700.050 197.400 ;
        RECT 703.950 198.600 706.050 199.050 ;
        RECT 715.950 198.600 718.050 199.050 ;
        RECT 703.950 197.400 718.050 198.600 ;
        RECT 703.950 196.950 706.050 197.400 ;
        RECT 715.950 196.950 718.050 197.400 ;
        RECT 733.950 198.600 736.050 199.050 ;
        RECT 748.950 198.600 751.050 199.050 ;
        RECT 733.950 197.400 751.050 198.600 ;
        RECT 733.950 196.950 736.050 197.400 ;
        RECT 748.950 196.950 751.050 197.400 ;
        RECT 754.950 198.600 757.050 199.050 ;
        RECT 760.950 198.600 763.050 199.050 ;
        RECT 754.950 197.400 763.050 198.600 ;
        RECT 754.950 196.950 757.050 197.400 ;
        RECT 760.950 196.950 763.050 197.400 ;
        RECT 763.950 198.600 766.050 199.050 ;
        RECT 769.950 198.600 772.050 199.050 ;
        RECT 763.950 197.400 772.050 198.600 ;
        RECT 763.950 196.950 766.050 197.400 ;
        RECT 769.950 196.950 772.050 197.400 ;
        RECT 775.950 198.600 778.050 199.050 ;
        RECT 793.950 198.600 796.050 199.050 ;
        RECT 775.950 197.400 796.050 198.600 ;
        RECT 775.950 196.950 778.050 197.400 ;
        RECT 793.950 196.950 796.050 197.400 ;
        RECT 823.950 198.600 826.050 199.050 ;
        RECT 838.950 198.600 841.050 199.050 ;
        RECT 823.950 197.400 841.050 198.600 ;
        RECT 823.950 196.950 826.050 197.400 ;
        RECT 838.950 196.950 841.050 197.400 ;
        RECT 856.950 198.600 859.050 199.050 ;
        RECT 865.950 198.600 868.050 199.050 ;
        RECT 856.950 197.400 868.050 198.600 ;
        RECT 856.950 196.950 859.050 197.400 ;
        RECT 865.950 196.950 868.050 197.400 ;
        RECT 139.950 194.400 147.600 195.600 ;
        RECT 157.950 195.600 160.050 196.050 ;
        RECT 184.950 195.600 187.050 196.050 ;
        RECT 157.950 194.400 187.050 195.600 ;
        RECT 139.950 193.950 142.050 194.400 ;
        RECT 157.950 193.950 160.050 194.400 ;
        RECT 184.950 193.950 187.050 194.400 ;
        RECT 325.950 195.600 328.050 196.050 ;
        RECT 346.950 195.600 349.050 196.050 ;
        RECT 325.950 194.400 349.050 195.600 ;
        RECT 325.950 193.950 328.050 194.400 ;
        RECT 346.950 193.950 349.050 194.400 ;
        RECT 364.950 195.600 367.050 196.050 ;
        RECT 379.950 195.600 382.050 196.050 ;
        RECT 364.950 194.400 382.050 195.600 ;
        RECT 364.950 193.950 367.050 194.400 ;
        RECT 379.950 193.950 382.050 194.400 ;
        RECT 397.950 195.600 400.050 196.050 ;
        RECT 403.950 195.600 406.050 196.050 ;
        RECT 397.950 194.400 406.050 195.600 ;
        RECT 397.950 193.950 400.050 194.400 ;
        RECT 403.950 193.950 406.050 194.400 ;
        RECT 412.950 195.600 415.050 196.050 ;
        RECT 466.950 195.600 469.050 196.050 ;
        RECT 412.950 194.400 469.050 195.600 ;
        RECT 412.950 193.950 415.050 194.400 ;
        RECT 466.950 193.950 469.050 194.400 ;
        RECT 508.950 195.600 511.050 196.050 ;
        RECT 556.950 195.600 559.050 196.050 ;
        RECT 508.950 194.400 559.050 195.600 ;
        RECT 508.950 193.950 511.050 194.400 ;
        RECT 556.950 193.950 559.050 194.400 ;
        RECT 742.950 195.600 745.050 196.050 ;
        RECT 757.950 195.600 760.050 196.050 ;
        RECT 742.950 194.400 760.050 195.600 ;
        RECT 742.950 193.950 745.050 194.400 ;
        RECT 757.950 193.950 760.050 194.400 ;
        RECT 766.950 195.600 769.050 196.050 ;
        RECT 802.950 195.600 805.050 196.050 ;
        RECT 766.950 194.400 805.050 195.600 ;
        RECT 766.950 193.950 769.050 194.400 ;
        RECT 802.950 193.950 805.050 194.400 ;
        RECT 820.950 195.600 823.050 196.050 ;
        RECT 826.950 195.600 829.050 196.050 ;
        RECT 820.950 194.400 829.050 195.600 ;
        RECT 820.950 193.950 823.050 194.400 ;
        RECT 826.950 193.950 829.050 194.400 ;
        RECT 841.950 195.600 844.050 196.050 ;
        RECT 847.950 195.600 850.050 196.050 ;
        RECT 841.950 194.400 850.050 195.600 ;
        RECT 841.950 193.950 844.050 194.400 ;
        RECT 847.950 193.950 850.050 194.400 ;
        RECT 127.950 192.600 130.050 193.050 ;
        RECT 145.950 192.600 148.050 193.050 ;
        RECT 127.950 191.400 148.050 192.600 ;
        RECT 127.950 190.950 130.050 191.400 ;
        RECT 145.950 190.950 148.050 191.400 ;
        RECT 214.950 192.600 217.050 193.050 ;
        RECT 235.950 192.600 238.050 193.050 ;
        RECT 214.950 191.400 238.050 192.600 ;
        RECT 214.950 190.950 217.050 191.400 ;
        RECT 235.950 190.950 238.050 191.400 ;
        RECT 352.950 192.600 355.050 193.050 ;
        RECT 418.950 192.600 421.050 193.050 ;
        RECT 352.950 191.400 421.050 192.600 ;
        RECT 352.950 190.950 355.050 191.400 ;
        RECT 418.950 190.950 421.050 191.400 ;
        RECT 421.950 192.600 424.050 193.050 ;
        RECT 439.950 192.600 442.050 193.050 ;
        RECT 421.950 191.400 442.050 192.600 ;
        RECT 421.950 190.950 424.050 191.400 ;
        RECT 439.950 190.950 442.050 191.400 ;
        RECT 493.950 192.600 496.050 193.050 ;
        RECT 550.950 192.600 553.050 193.050 ;
        RECT 589.950 192.600 592.050 193.050 ;
        RECT 493.950 191.400 592.050 192.600 ;
        RECT 493.950 190.950 496.050 191.400 ;
        RECT 550.950 190.950 553.050 191.400 ;
        RECT 589.950 190.950 592.050 191.400 ;
        RECT 628.950 192.600 631.050 193.050 ;
        RECT 658.950 192.600 661.050 193.050 ;
        RECT 628.950 191.400 661.050 192.600 ;
        RECT 628.950 190.950 631.050 191.400 ;
        RECT 658.950 190.950 661.050 191.400 ;
        RECT 694.950 192.600 697.050 193.050 ;
        RECT 712.950 192.600 715.050 193.050 ;
        RECT 727.950 192.600 730.050 193.050 ;
        RECT 694.950 191.400 730.050 192.600 ;
        RECT 694.950 190.950 697.050 191.400 ;
        RECT 712.950 190.950 715.050 191.400 ;
        RECT 727.950 190.950 730.050 191.400 ;
        RECT 772.950 192.600 775.050 193.050 ;
        RECT 835.950 192.600 838.050 193.050 ;
        RECT 772.950 191.400 838.050 192.600 ;
        RECT 772.950 190.950 775.050 191.400 ;
        RECT 835.950 190.950 838.050 191.400 ;
        RECT 55.950 189.600 58.050 190.050 ;
        RECT 91.950 189.600 94.050 190.050 ;
        RECT 55.950 188.400 94.050 189.600 ;
        RECT 55.950 187.950 58.050 188.400 ;
        RECT 91.950 187.950 94.050 188.400 ;
        RECT 103.950 189.600 106.050 190.050 ;
        RECT 154.950 189.600 157.050 190.050 ;
        RECT 166.950 189.600 169.050 190.050 ;
        RECT 175.950 189.600 178.050 190.050 ;
        RECT 280.950 189.600 283.050 190.050 ;
        RECT 103.950 188.400 283.050 189.600 ;
        RECT 103.950 187.950 106.050 188.400 ;
        RECT 154.950 187.950 157.050 188.400 ;
        RECT 166.950 187.950 169.050 188.400 ;
        RECT 175.950 187.950 178.050 188.400 ;
        RECT 280.950 187.950 283.050 188.400 ;
        RECT 301.950 186.600 304.050 187.050 ;
        RECT 454.950 186.600 457.050 187.050 ;
        RECT 487.950 186.600 490.050 187.050 ;
        RECT 301.950 185.400 490.050 186.600 ;
        RECT 301.950 184.950 304.050 185.400 ;
        RECT 454.950 184.950 457.050 185.400 ;
        RECT 487.950 184.950 490.050 185.400 ;
        RECT 517.950 186.600 520.050 187.050 ;
        RECT 574.950 186.600 577.050 187.050 ;
        RECT 577.950 186.600 580.050 187.050 ;
        RECT 517.950 185.400 580.050 186.600 ;
        RECT 517.950 184.950 520.050 185.400 ;
        RECT 574.950 184.950 577.050 185.400 ;
        RECT 577.950 184.950 580.050 185.400 ;
        RECT 589.950 186.600 592.050 187.050 ;
        RECT 703.950 186.600 706.050 187.050 ;
        RECT 589.950 185.400 706.050 186.600 ;
        RECT 589.950 184.950 592.050 185.400 ;
        RECT 703.950 184.950 706.050 185.400 ;
        RECT 751.950 186.600 754.050 187.050 ;
        RECT 814.950 186.600 817.050 187.050 ;
        RECT 751.950 185.400 817.050 186.600 ;
        RECT 751.950 184.950 754.050 185.400 ;
        RECT 814.950 184.950 817.050 185.400 ;
        RECT 376.950 183.600 379.050 184.050 ;
        RECT 430.950 183.600 433.050 184.050 ;
        RECT 376.950 182.400 433.050 183.600 ;
        RECT 376.950 181.950 379.050 182.400 ;
        RECT 430.950 181.950 433.050 182.400 ;
        RECT 292.950 180.600 295.050 181.050 ;
        RECT 451.950 180.600 454.050 181.050 ;
        RECT 292.950 179.400 454.050 180.600 ;
        RECT 292.950 178.950 295.050 179.400 ;
        RECT 451.950 178.950 454.050 179.400 ;
        RECT 472.950 180.600 475.050 181.050 ;
        RECT 502.950 180.600 505.050 181.050 ;
        RECT 520.950 180.600 523.050 181.050 ;
        RECT 472.950 179.400 523.050 180.600 ;
        RECT 472.950 178.950 475.050 179.400 ;
        RECT 502.950 178.950 505.050 179.400 ;
        RECT 520.950 178.950 523.050 179.400 ;
        RECT 526.950 180.600 529.050 181.050 ;
        RECT 535.950 180.600 538.050 181.050 ;
        RECT 553.950 180.600 556.050 181.050 ;
        RECT 526.950 179.400 556.050 180.600 ;
        RECT 526.950 178.950 529.050 179.400 ;
        RECT 535.950 178.950 538.050 179.400 ;
        RECT 553.950 178.950 556.050 179.400 ;
        RECT 604.950 180.600 607.050 181.050 ;
        RECT 679.950 180.600 682.050 181.050 ;
        RECT 604.950 179.400 682.050 180.600 ;
        RECT 604.950 178.950 607.050 179.400 ;
        RECT 679.950 178.950 682.050 179.400 ;
        RECT 772.950 180.600 775.050 181.050 ;
        RECT 817.950 180.600 820.050 181.050 ;
        RECT 772.950 179.400 820.050 180.600 ;
        RECT 772.950 178.950 775.050 179.400 ;
        RECT 817.950 178.950 820.050 179.400 ;
        RECT 94.950 177.600 97.050 178.050 ;
        RECT 157.950 177.600 160.050 178.050 ;
        RECT 94.950 176.400 160.050 177.600 ;
        RECT 94.950 175.950 97.050 176.400 ;
        RECT 157.950 175.950 160.050 176.400 ;
        RECT 391.950 177.600 394.050 178.050 ;
        RECT 409.950 177.600 412.050 178.050 ;
        RECT 391.950 176.400 412.050 177.600 ;
        RECT 391.950 175.950 394.050 176.400 ;
        RECT 409.950 175.950 412.050 176.400 ;
        RECT 610.950 177.600 613.050 178.050 ;
        RECT 670.950 177.600 673.050 178.050 ;
        RECT 739.950 177.600 742.050 178.050 ;
        RECT 610.950 176.400 742.050 177.600 ;
        RECT 610.950 175.950 613.050 176.400 ;
        RECT 670.950 175.950 673.050 176.400 ;
        RECT 739.950 175.950 742.050 176.400 ;
        RECT 781.950 177.600 784.050 178.050 ;
        RECT 796.950 177.600 799.050 178.050 ;
        RECT 781.950 176.400 799.050 177.600 ;
        RECT 781.950 175.950 784.050 176.400 ;
        RECT 796.950 175.950 799.050 176.400 ;
        RECT 802.950 177.600 805.050 178.050 ;
        RECT 880.950 177.600 883.050 178.050 ;
        RECT 802.950 176.400 883.050 177.600 ;
        RECT 802.950 175.950 805.050 176.400 ;
        RECT 880.950 175.950 883.050 176.400 ;
        RECT 85.950 174.600 88.050 175.050 ;
        RECT 88.950 174.600 91.050 175.050 ;
        RECT 139.950 174.600 142.050 175.050 ;
        RECT 85.950 173.400 142.050 174.600 ;
        RECT 85.950 172.950 88.050 173.400 ;
        RECT 88.950 172.950 91.050 173.400 ;
        RECT 139.950 172.950 142.050 173.400 ;
        RECT 244.950 174.600 247.050 175.050 ;
        RECT 295.950 174.600 298.050 175.050 ;
        RECT 322.950 174.600 325.050 175.050 ;
        RECT 244.950 173.400 325.050 174.600 ;
        RECT 244.950 172.950 247.050 173.400 ;
        RECT 295.950 172.950 298.050 173.400 ;
        RECT 322.950 172.950 325.050 173.400 ;
        RECT 409.950 174.600 412.050 175.050 ;
        RECT 460.950 174.600 463.050 175.050 ;
        RECT 409.950 173.400 463.050 174.600 ;
        RECT 409.950 172.950 412.050 173.400 ;
        RECT 460.950 172.950 463.050 173.400 ;
        RECT 499.950 174.600 502.050 175.050 ;
        RECT 583.950 174.600 586.050 175.050 ;
        RECT 499.950 173.400 586.050 174.600 ;
        RECT 499.950 172.950 502.050 173.400 ;
        RECT 583.950 172.950 586.050 173.400 ;
        RECT 616.950 174.600 619.050 175.050 ;
        RECT 772.950 174.600 775.050 175.050 ;
        RECT 616.950 173.400 775.050 174.600 ;
        RECT 616.950 172.950 619.050 173.400 ;
        RECT 772.950 172.950 775.050 173.400 ;
        RECT 808.950 174.600 811.050 175.050 ;
        RECT 835.950 174.600 838.050 175.050 ;
        RECT 808.950 173.400 838.050 174.600 ;
        RECT 808.950 172.950 811.050 173.400 ;
        RECT 835.950 172.950 838.050 173.400 ;
        RECT 10.950 171.600 13.050 172.050 ;
        RECT 25.950 171.600 28.050 172.050 ;
        RECT 10.950 170.400 28.050 171.600 ;
        RECT 10.950 169.950 13.050 170.400 ;
        RECT 25.950 169.950 28.050 170.400 ;
        RECT 106.950 171.600 109.050 172.050 ;
        RECT 112.950 171.600 115.050 172.050 ;
        RECT 106.950 170.400 115.050 171.600 ;
        RECT 106.950 169.950 109.050 170.400 ;
        RECT 112.950 169.950 115.050 170.400 ;
        RECT 331.950 171.600 334.050 172.050 ;
        RECT 394.950 171.600 397.050 172.050 ;
        RECT 331.950 170.400 397.050 171.600 ;
        RECT 331.950 169.950 334.050 170.400 ;
        RECT 394.950 169.950 397.050 170.400 ;
        RECT 400.950 171.600 403.050 172.050 ;
        RECT 448.950 171.600 451.050 172.050 ;
        RECT 457.950 171.600 460.050 172.050 ;
        RECT 466.950 171.600 469.050 172.050 ;
        RECT 535.950 171.600 538.050 172.050 ;
        RECT 400.950 170.400 538.050 171.600 ;
        RECT 400.950 169.950 403.050 170.400 ;
        RECT 448.950 169.950 451.050 170.400 ;
        RECT 457.950 169.950 460.050 170.400 ;
        RECT 466.950 169.950 469.050 170.400 ;
        RECT 535.950 169.950 538.050 170.400 ;
        RECT 541.950 171.600 544.050 172.050 ;
        RECT 556.950 171.600 559.050 172.050 ;
        RECT 541.950 170.400 559.050 171.600 ;
        RECT 541.950 169.950 544.050 170.400 ;
        RECT 556.950 169.950 559.050 170.400 ;
        RECT 583.950 171.600 586.050 172.050 ;
        RECT 664.950 171.600 667.050 172.050 ;
        RECT 583.950 170.400 667.050 171.600 ;
        RECT 583.950 169.950 586.050 170.400 ;
        RECT 664.950 169.950 667.050 170.400 ;
        RECT 706.950 171.600 709.050 172.050 ;
        RECT 751.950 171.600 754.050 172.050 ;
        RECT 706.950 170.400 754.050 171.600 ;
        RECT 706.950 169.950 709.050 170.400 ;
        RECT 751.950 169.950 754.050 170.400 ;
        RECT 769.950 171.600 772.050 172.050 ;
        RECT 787.950 171.600 790.050 172.050 ;
        RECT 769.950 170.400 790.050 171.600 ;
        RECT 769.950 169.950 772.050 170.400 ;
        RECT 787.950 169.950 790.050 170.400 ;
        RECT 799.950 171.600 802.050 172.050 ;
        RECT 811.950 171.600 814.050 172.050 ;
        RECT 799.950 170.400 814.050 171.600 ;
        RECT 799.950 169.950 802.050 170.400 ;
        RECT 811.950 169.950 814.050 170.400 ;
        RECT 16.950 168.600 19.050 169.050 ;
        RECT 22.950 168.600 25.050 169.050 ;
        RECT 16.950 167.400 25.050 168.600 ;
        RECT 16.950 166.950 19.050 167.400 ;
        RECT 22.950 166.950 25.050 167.400 ;
        RECT 61.950 168.600 64.050 169.050 ;
        RECT 97.950 168.600 100.050 169.050 ;
        RECT 61.950 167.400 100.050 168.600 ;
        RECT 61.950 166.950 64.050 167.400 ;
        RECT 97.950 166.950 100.050 167.400 ;
        RECT 133.950 168.600 136.050 169.050 ;
        RECT 169.950 168.600 172.050 169.050 ;
        RECT 133.950 167.400 172.050 168.600 ;
        RECT 133.950 166.950 136.050 167.400 ;
        RECT 169.950 166.950 172.050 167.400 ;
        RECT 199.950 168.600 202.050 169.050 ;
        RECT 217.950 168.600 220.050 169.050 ;
        RECT 238.950 168.600 241.050 169.050 ;
        RECT 250.950 168.600 253.050 169.050 ;
        RECT 280.950 168.600 283.050 169.050 ;
        RECT 337.950 168.600 340.050 169.050 ;
        RECT 358.950 168.600 361.050 169.050 ;
        RECT 391.950 168.600 394.050 169.050 ;
        RECT 199.950 167.400 394.050 168.600 ;
        RECT 199.950 166.950 202.050 167.400 ;
        RECT 217.950 166.950 220.050 167.400 ;
        RECT 238.950 166.950 241.050 167.400 ;
        RECT 250.950 166.950 253.050 167.400 ;
        RECT 280.950 166.950 283.050 167.400 ;
        RECT 337.950 166.950 340.050 167.400 ;
        RECT 358.950 166.950 361.050 167.400 ;
        RECT 391.950 166.950 394.050 167.400 ;
        RECT 421.950 168.600 424.050 169.050 ;
        RECT 493.950 168.600 496.050 169.050 ;
        RECT 421.950 167.400 496.050 168.600 ;
        RECT 421.950 166.950 424.050 167.400 ;
        RECT 493.950 166.950 496.050 167.400 ;
        RECT 532.950 168.600 535.050 169.050 ;
        RECT 577.950 168.600 580.050 169.050 ;
        RECT 532.950 167.400 580.050 168.600 ;
        RECT 532.950 166.950 535.050 167.400 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 622.950 168.600 625.050 169.050 ;
        RECT 628.950 168.600 631.050 169.050 ;
        RECT 622.950 167.400 631.050 168.600 ;
        RECT 622.950 166.950 625.050 167.400 ;
        RECT 628.950 166.950 631.050 167.400 ;
        RECT 637.950 168.600 640.050 169.050 ;
        RECT 643.950 168.600 646.050 169.050 ;
        RECT 637.950 167.400 646.050 168.600 ;
        RECT 637.950 166.950 640.050 167.400 ;
        RECT 643.950 166.950 646.050 167.400 ;
        RECT 649.950 168.600 652.050 169.050 ;
        RECT 655.950 168.600 658.050 169.050 ;
        RECT 649.950 167.400 658.050 168.600 ;
        RECT 649.950 166.950 652.050 167.400 ;
        RECT 655.950 166.950 658.050 167.400 ;
        RECT 682.950 168.600 685.050 169.050 ;
        RECT 694.950 168.600 697.050 169.050 ;
        RECT 682.950 167.400 697.050 168.600 ;
        RECT 682.950 166.950 685.050 167.400 ;
        RECT 694.950 166.950 697.050 167.400 ;
        RECT 700.950 166.950 703.050 169.050 ;
        RECT 712.950 168.600 715.050 169.050 ;
        RECT 721.950 168.600 724.050 169.050 ;
        RECT 712.950 167.400 724.050 168.600 ;
        RECT 712.950 166.950 715.050 167.400 ;
        RECT 721.950 166.950 724.050 167.400 ;
        RECT 739.950 168.600 742.050 169.050 ;
        RECT 745.950 168.600 748.050 169.050 ;
        RECT 766.950 168.600 769.050 169.050 ;
        RECT 739.950 167.400 769.050 168.600 ;
        RECT 739.950 166.950 742.050 167.400 ;
        RECT 745.950 166.950 748.050 167.400 ;
        RECT 766.950 166.950 769.050 167.400 ;
        RECT 784.950 168.600 787.050 169.050 ;
        RECT 790.950 168.600 793.050 169.050 ;
        RECT 784.950 167.400 793.050 168.600 ;
        RECT 784.950 166.950 787.050 167.400 ;
        RECT 790.950 166.950 793.050 167.400 ;
        RECT 808.950 168.600 811.050 169.050 ;
        RECT 829.950 168.600 832.050 169.050 ;
        RECT 865.950 168.600 868.050 169.050 ;
        RECT 808.950 167.400 846.600 168.600 ;
        RECT 808.950 166.950 811.050 167.400 ;
        RECT 829.950 166.950 832.050 167.400 ;
        RECT 7.950 165.600 10.050 166.050 ;
        RECT 13.950 165.600 16.050 166.050 ;
        RECT 7.950 164.400 16.050 165.600 ;
        RECT 7.950 163.950 10.050 164.400 ;
        RECT 13.950 163.950 16.050 164.400 ;
        RECT 19.950 165.600 22.050 166.050 ;
        RECT 37.950 165.600 40.050 166.050 ;
        RECT 19.950 164.400 40.050 165.600 ;
        RECT 19.950 163.950 22.050 164.400 ;
        RECT 37.950 163.950 40.050 164.400 ;
        RECT 58.950 165.600 61.050 166.050 ;
        RECT 76.950 165.600 79.050 166.050 ;
        RECT 58.950 164.400 79.050 165.600 ;
        RECT 58.950 163.950 61.050 164.400 ;
        RECT 76.950 163.950 79.050 164.400 ;
        RECT 100.950 165.600 103.050 166.050 ;
        RECT 109.950 165.600 112.050 166.050 ;
        RECT 100.950 164.400 112.050 165.600 ;
        RECT 100.950 163.950 103.050 164.400 ;
        RECT 109.950 163.950 112.050 164.400 ;
        RECT 160.950 165.600 163.050 166.050 ;
        RECT 166.950 165.600 169.050 166.050 ;
        RECT 160.950 164.400 169.050 165.600 ;
        RECT 160.950 163.950 163.050 164.400 ;
        RECT 166.950 163.950 169.050 164.400 ;
        RECT 193.950 165.600 196.050 166.050 ;
        RECT 208.950 165.600 211.050 166.050 ;
        RECT 193.950 164.400 211.050 165.600 ;
        RECT 193.950 163.950 196.050 164.400 ;
        RECT 208.950 163.950 211.050 164.400 ;
        RECT 232.950 165.600 235.050 166.050 ;
        RECT 271.950 165.600 274.050 166.050 ;
        RECT 232.950 164.400 274.050 165.600 ;
        RECT 232.950 163.950 235.050 164.400 ;
        RECT 271.950 163.950 274.050 164.400 ;
        RECT 346.950 165.600 349.050 166.050 ;
        RECT 364.950 165.600 367.050 166.050 ;
        RECT 346.950 164.400 367.050 165.600 ;
        RECT 346.950 163.950 349.050 164.400 ;
        RECT 364.950 163.950 367.050 164.400 ;
        RECT 415.950 165.600 418.050 166.050 ;
        RECT 472.950 165.600 475.050 166.050 ;
        RECT 517.950 165.600 520.050 166.050 ;
        RECT 415.950 164.400 520.050 165.600 ;
        RECT 415.950 163.950 418.050 164.400 ;
        RECT 472.950 163.950 475.050 164.400 ;
        RECT 517.950 163.950 520.050 164.400 ;
        RECT 559.950 165.600 562.050 166.050 ;
        RECT 580.950 165.600 583.050 166.050 ;
        RECT 640.950 165.600 643.050 166.050 ;
        RECT 559.950 164.400 643.050 165.600 ;
        RECT 559.950 163.950 562.050 164.400 ;
        RECT 580.950 163.950 583.050 164.400 ;
        RECT 640.950 163.950 643.050 164.400 ;
        RECT 682.950 165.600 685.050 166.050 ;
        RECT 701.400 165.600 702.600 166.950 ;
        RECT 845.400 166.050 846.600 167.400 ;
        RECT 854.400 167.400 868.050 168.600 ;
        RECT 854.400 166.050 855.600 167.400 ;
        RECT 865.950 166.950 868.050 167.400 ;
        RECT 871.950 168.600 874.050 169.050 ;
        RECT 880.950 168.600 883.050 169.050 ;
        RECT 871.950 167.400 883.050 168.600 ;
        RECT 871.950 166.950 874.050 167.400 ;
        RECT 880.950 166.950 883.050 167.400 ;
        RECT 682.950 164.400 702.600 165.600 ;
        RECT 748.950 165.600 751.050 166.050 ;
        RECT 781.950 165.600 784.050 166.050 ;
        RECT 748.950 164.400 784.050 165.600 ;
        RECT 682.950 163.950 685.050 164.400 ;
        RECT 748.950 163.950 751.050 164.400 ;
        RECT 781.950 163.950 784.050 164.400 ;
        RECT 793.950 165.600 796.050 166.050 ;
        RECT 799.950 165.600 802.050 166.050 ;
        RECT 793.950 164.400 802.050 165.600 ;
        RECT 793.950 163.950 796.050 164.400 ;
        RECT 799.950 163.950 802.050 164.400 ;
        RECT 844.950 163.950 847.050 166.050 ;
        RECT 853.950 163.950 856.050 166.050 ;
        RECT 13.950 162.600 16.050 163.050 ;
        RECT 34.950 162.600 37.050 163.050 ;
        RECT 52.950 162.600 55.050 163.050 ;
        RECT 73.950 162.600 76.050 163.050 ;
        RECT 13.950 161.400 76.050 162.600 ;
        RECT 13.950 160.950 16.050 161.400 ;
        RECT 34.950 160.950 37.050 161.400 ;
        RECT 52.950 160.950 55.050 161.400 ;
        RECT 73.950 160.950 76.050 161.400 ;
        RECT 115.950 162.600 118.050 163.050 ;
        RECT 190.950 162.600 193.050 163.050 ;
        RECT 115.950 161.400 193.050 162.600 ;
        RECT 115.950 160.950 118.050 161.400 ;
        RECT 190.950 160.950 193.050 161.400 ;
        RECT 214.950 162.600 217.050 163.050 ;
        RECT 217.950 162.600 220.050 163.050 ;
        RECT 229.950 162.600 232.050 163.050 ;
        RECT 214.950 161.400 232.050 162.600 ;
        RECT 214.950 160.950 217.050 161.400 ;
        RECT 217.950 160.950 220.050 161.400 ;
        RECT 229.950 160.950 232.050 161.400 ;
        RECT 367.950 162.600 370.050 163.050 ;
        RECT 409.950 162.600 412.050 163.050 ;
        RECT 424.950 162.600 427.050 163.050 ;
        RECT 367.950 161.400 427.050 162.600 ;
        RECT 367.950 160.950 370.050 161.400 ;
        RECT 409.950 160.950 412.050 161.400 ;
        RECT 424.950 160.950 427.050 161.400 ;
        RECT 451.950 162.600 454.050 163.050 ;
        RECT 493.950 162.600 496.050 163.050 ;
        RECT 451.950 161.400 496.050 162.600 ;
        RECT 451.950 160.950 454.050 161.400 ;
        RECT 493.950 160.950 496.050 161.400 ;
        RECT 496.950 162.600 499.050 163.050 ;
        RECT 523.950 162.600 526.050 163.050 ;
        RECT 538.950 162.600 541.050 163.050 ;
        RECT 496.950 161.400 541.050 162.600 ;
        RECT 496.950 160.950 499.050 161.400 ;
        RECT 523.950 160.950 526.050 161.400 ;
        RECT 538.950 160.950 541.050 161.400 ;
        RECT 643.950 162.600 646.050 163.050 ;
        RECT 655.950 162.600 658.050 163.050 ;
        RECT 643.950 161.400 658.050 162.600 ;
        RECT 643.950 160.950 646.050 161.400 ;
        RECT 655.950 160.950 658.050 161.400 ;
        RECT 724.950 162.600 727.050 163.050 ;
        RECT 775.950 162.600 778.050 163.050 ;
        RECT 724.950 161.400 778.050 162.600 ;
        RECT 724.950 160.950 727.050 161.400 ;
        RECT 775.950 160.950 778.050 161.400 ;
        RECT 781.950 162.600 784.050 163.050 ;
        RECT 826.950 162.600 829.050 163.050 ;
        RECT 781.950 161.400 829.050 162.600 ;
        RECT 781.950 160.950 784.050 161.400 ;
        RECT 826.950 160.950 829.050 161.400 ;
        RECT 151.950 159.600 154.050 160.050 ;
        RECT 214.950 159.600 217.050 160.050 ;
        RECT 151.950 158.400 217.050 159.600 ;
        RECT 151.950 157.950 154.050 158.400 ;
        RECT 214.950 157.950 217.050 158.400 ;
        RECT 277.950 159.600 280.050 160.050 ;
        RECT 439.950 159.600 442.050 160.050 ;
        RECT 277.950 158.400 442.050 159.600 ;
        RECT 277.950 157.950 280.050 158.400 ;
        RECT 439.950 157.950 442.050 158.400 ;
        RECT 763.950 159.600 766.050 160.050 ;
        RECT 772.950 159.600 775.050 160.050 ;
        RECT 763.950 158.400 775.050 159.600 ;
        RECT 763.950 157.950 766.050 158.400 ;
        RECT 772.950 157.950 775.050 158.400 ;
        RECT 334.950 156.600 337.050 157.050 ;
        RECT 340.950 156.600 343.050 157.050 ;
        RECT 382.950 156.600 385.050 157.050 ;
        RECT 334.950 155.400 385.050 156.600 ;
        RECT 334.950 154.950 337.050 155.400 ;
        RECT 340.950 154.950 343.050 155.400 ;
        RECT 382.950 154.950 385.050 155.400 ;
        RECT 637.950 156.600 640.050 157.050 ;
        RECT 793.950 156.600 796.050 157.050 ;
        RECT 637.950 155.400 796.050 156.600 ;
        RECT 637.950 154.950 640.050 155.400 ;
        RECT 793.950 154.950 796.050 155.400 ;
        RECT 43.950 153.600 46.050 154.050 ;
        RECT 124.950 153.600 127.050 154.050 ;
        RECT 43.950 152.400 127.050 153.600 ;
        RECT 43.950 151.950 46.050 152.400 ;
        RECT 124.950 151.950 127.050 152.400 ;
        RECT 169.950 153.600 172.050 154.050 ;
        RECT 172.950 153.600 175.050 154.050 ;
        RECT 688.950 153.600 691.050 154.050 ;
        RECT 169.950 152.400 691.050 153.600 ;
        RECT 169.950 151.950 172.050 152.400 ;
        RECT 172.950 151.950 175.050 152.400 ;
        RECT 688.950 151.950 691.050 152.400 ;
        RECT 703.950 153.600 706.050 154.050 ;
        RECT 769.950 153.600 772.050 154.050 ;
        RECT 703.950 152.400 772.050 153.600 ;
        RECT 703.950 151.950 706.050 152.400 ;
        RECT 769.950 151.950 772.050 152.400 ;
        RECT 820.950 153.600 823.050 154.050 ;
        RECT 832.950 153.600 835.050 154.050 ;
        RECT 820.950 152.400 835.050 153.600 ;
        RECT 820.950 151.950 823.050 152.400 ;
        RECT 832.950 151.950 835.050 152.400 ;
        RECT 586.950 150.600 589.050 151.050 ;
        RECT 670.950 150.600 673.050 151.050 ;
        RECT 709.950 150.600 712.050 151.050 ;
        RECT 841.950 150.600 844.050 151.050 ;
        RECT 586.950 149.400 844.050 150.600 ;
        RECT 586.950 148.950 589.050 149.400 ;
        RECT 670.950 148.950 673.050 149.400 ;
        RECT 709.950 148.950 712.050 149.400 ;
        RECT 841.950 148.950 844.050 149.400 ;
        RECT 628.950 147.600 631.050 148.050 ;
        RECT 730.950 147.600 733.050 148.050 ;
        RECT 628.950 146.400 733.050 147.600 ;
        RECT 628.950 145.950 631.050 146.400 ;
        RECT 730.950 145.950 733.050 146.400 ;
        RECT 652.950 144.600 655.050 145.050 ;
        RECT 688.950 144.600 691.050 145.050 ;
        RECT 652.950 143.400 691.050 144.600 ;
        RECT 652.950 142.950 655.050 143.400 ;
        RECT 688.950 142.950 691.050 143.400 ;
        RECT 661.950 141.600 664.050 142.050 ;
        RECT 760.950 141.600 763.050 142.050 ;
        RECT 802.950 141.600 805.050 142.050 ;
        RECT 661.950 140.400 805.050 141.600 ;
        RECT 661.950 139.950 664.050 140.400 ;
        RECT 760.950 139.950 763.050 140.400 ;
        RECT 802.950 139.950 805.050 140.400 ;
        RECT 307.950 135.600 310.050 136.050 ;
        RECT 346.950 135.600 349.050 136.050 ;
        RECT 307.950 134.400 349.050 135.600 ;
        RECT 307.950 133.950 310.050 134.400 ;
        RECT 346.950 133.950 349.050 134.400 ;
        RECT 571.950 135.600 574.050 136.050 ;
        RECT 778.950 135.600 781.050 136.050 ;
        RECT 805.950 135.600 808.050 136.050 ;
        RECT 826.950 135.600 829.050 136.050 ;
        RECT 571.950 134.400 829.050 135.600 ;
        RECT 571.950 133.950 574.050 134.400 ;
        RECT 778.950 133.950 781.050 134.400 ;
        RECT 805.950 133.950 808.050 134.400 ;
        RECT 826.950 133.950 829.050 134.400 ;
        RECT 178.950 132.600 181.050 133.050 ;
        RECT 223.950 132.600 226.050 133.050 ;
        RECT 178.950 131.400 226.050 132.600 ;
        RECT 178.950 130.950 181.050 131.400 ;
        RECT 223.950 130.950 226.050 131.400 ;
        RECT 325.950 132.600 328.050 133.050 ;
        RECT 403.950 132.600 406.050 133.050 ;
        RECT 325.950 131.400 406.050 132.600 ;
        RECT 325.950 130.950 328.050 131.400 ;
        RECT 403.950 130.950 406.050 131.400 ;
        RECT 667.950 132.600 670.050 133.050 ;
        RECT 736.950 132.600 739.050 133.050 ;
        RECT 667.950 131.400 739.050 132.600 ;
        RECT 667.950 130.950 670.050 131.400 ;
        RECT 736.950 130.950 739.050 131.400 ;
        RECT 58.950 129.600 61.050 130.050 ;
        RECT 70.950 129.600 73.050 130.050 ;
        RECT 58.950 128.400 73.050 129.600 ;
        RECT 58.950 127.950 61.050 128.400 ;
        RECT 70.950 127.950 73.050 128.400 ;
        RECT 76.950 129.600 79.050 130.050 ;
        RECT 82.950 129.600 85.050 130.050 ;
        RECT 76.950 128.400 85.050 129.600 ;
        RECT 76.950 127.950 79.050 128.400 ;
        RECT 82.950 127.950 85.050 128.400 ;
        RECT 124.950 129.600 127.050 130.050 ;
        RECT 151.950 129.600 154.050 130.050 ;
        RECT 169.950 129.600 172.050 130.050 ;
        RECT 124.950 128.400 172.050 129.600 ;
        RECT 124.950 127.950 127.050 128.400 ;
        RECT 151.950 127.950 154.050 128.400 ;
        RECT 169.950 127.950 172.050 128.400 ;
        RECT 187.950 129.600 190.050 130.050 ;
        RECT 193.950 129.600 196.050 130.050 ;
        RECT 283.950 129.600 286.050 130.050 ;
        RECT 307.950 129.600 310.050 130.050 ;
        RECT 187.950 128.400 310.050 129.600 ;
        RECT 187.950 127.950 190.050 128.400 ;
        RECT 193.950 127.950 196.050 128.400 ;
        RECT 283.950 127.950 286.050 128.400 ;
        RECT 307.950 127.950 310.050 128.400 ;
        RECT 328.950 129.600 331.050 130.050 ;
        RECT 334.950 129.600 337.050 130.050 ;
        RECT 367.950 129.600 370.050 130.050 ;
        RECT 328.950 128.400 370.050 129.600 ;
        RECT 328.950 127.950 331.050 128.400 ;
        RECT 334.950 127.950 337.050 128.400 ;
        RECT 367.950 127.950 370.050 128.400 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 388.950 129.600 391.050 130.050 ;
        RECT 373.950 128.400 391.050 129.600 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 388.950 127.950 391.050 128.400 ;
        RECT 394.950 129.600 397.050 130.050 ;
        RECT 400.950 129.600 403.050 130.050 ;
        RECT 430.950 129.600 433.050 130.050 ;
        RECT 394.950 128.400 403.050 129.600 ;
        RECT 394.950 127.950 397.050 128.400 ;
        RECT 400.950 127.950 403.050 128.400 ;
        RECT 413.400 128.400 433.050 129.600 ;
        RECT 413.400 127.050 414.600 128.400 ;
        RECT 430.950 127.950 433.050 128.400 ;
        RECT 457.950 129.600 460.050 130.050 ;
        RECT 511.950 129.600 514.050 130.050 ;
        RECT 457.950 128.400 514.050 129.600 ;
        RECT 457.950 127.950 460.050 128.400 ;
        RECT 511.950 127.950 514.050 128.400 ;
        RECT 553.950 129.600 556.050 130.050 ;
        RECT 595.950 129.600 598.050 130.050 ;
        RECT 655.950 129.600 658.050 130.050 ;
        RECT 667.950 129.600 670.050 130.050 ;
        RECT 553.950 128.400 558.600 129.600 ;
        RECT 553.950 127.950 556.050 128.400 ;
        RECT 557.400 127.050 558.600 128.400 ;
        RECT 595.950 128.400 654.600 129.600 ;
        RECT 595.950 127.950 598.050 128.400 ;
        RECT 46.950 126.600 49.050 127.050 ;
        RECT 67.950 126.600 70.050 127.050 ;
        RECT 46.950 125.400 70.050 126.600 ;
        RECT 46.950 124.950 49.050 125.400 ;
        RECT 67.950 124.950 70.050 125.400 ;
        RECT 94.950 126.600 97.050 127.050 ;
        RECT 130.950 126.600 133.050 127.050 ;
        RECT 148.950 126.600 151.050 127.050 ;
        RECT 94.950 125.400 120.600 126.600 ;
        RECT 94.950 124.950 97.050 125.400 ;
        RECT 4.950 123.600 7.050 124.050 ;
        RECT 10.950 123.600 13.050 124.050 ;
        RECT 4.950 122.400 13.050 123.600 ;
        RECT 4.950 121.950 7.050 122.400 ;
        RECT 10.950 121.950 13.050 122.400 ;
        RECT 13.950 123.600 16.050 124.050 ;
        RECT 25.950 123.600 28.050 124.050 ;
        RECT 13.950 122.400 28.050 123.600 ;
        RECT 13.950 121.950 16.050 122.400 ;
        RECT 25.950 121.950 28.050 122.400 ;
        RECT 52.950 123.600 55.050 124.050 ;
        RECT 82.950 123.600 85.050 124.050 ;
        RECT 52.950 122.400 85.050 123.600 ;
        RECT 52.950 121.950 55.050 122.400 ;
        RECT 82.950 121.950 85.050 122.400 ;
        RECT 88.950 123.600 91.050 124.050 ;
        RECT 97.950 123.600 100.050 124.050 ;
        RECT 88.950 122.400 100.050 123.600 ;
        RECT 88.950 121.950 91.050 122.400 ;
        RECT 97.950 121.950 100.050 122.400 ;
        RECT 109.950 123.600 112.050 124.050 ;
        RECT 115.950 123.600 118.050 124.050 ;
        RECT 109.950 122.400 118.050 123.600 ;
        RECT 119.400 123.600 120.600 125.400 ;
        RECT 130.950 125.400 151.050 126.600 ;
        RECT 130.950 124.950 133.050 125.400 ;
        RECT 148.950 124.950 151.050 125.400 ;
        RECT 160.950 126.600 163.050 127.050 ;
        RECT 166.950 126.600 169.050 127.050 ;
        RECT 160.950 125.400 169.050 126.600 ;
        RECT 160.950 124.950 163.050 125.400 ;
        RECT 166.950 124.950 169.050 125.400 ;
        RECT 178.950 126.600 181.050 127.050 ;
        RECT 187.950 126.600 190.050 127.050 ;
        RECT 178.950 125.400 190.050 126.600 ;
        RECT 178.950 124.950 181.050 125.400 ;
        RECT 187.950 124.950 190.050 125.400 ;
        RECT 190.950 126.600 193.050 127.050 ;
        RECT 205.950 126.600 208.050 127.050 ;
        RECT 190.950 125.400 208.050 126.600 ;
        RECT 190.950 124.950 193.050 125.400 ;
        RECT 205.950 124.950 208.050 125.400 ;
        RECT 232.950 126.600 235.050 127.050 ;
        RECT 247.950 126.600 250.050 127.050 ;
        RECT 232.950 125.400 250.050 126.600 ;
        RECT 232.950 124.950 235.050 125.400 ;
        RECT 247.950 124.950 250.050 125.400 ;
        RECT 310.950 126.600 313.050 127.050 ;
        RECT 322.950 126.600 325.050 127.050 ;
        RECT 346.950 126.600 349.050 127.050 ;
        RECT 310.950 125.400 349.050 126.600 ;
        RECT 310.950 124.950 313.050 125.400 ;
        RECT 322.950 124.950 325.050 125.400 ;
        RECT 346.950 124.950 349.050 125.400 ;
        RECT 376.950 126.600 379.050 127.050 ;
        RECT 385.950 126.600 388.050 127.050 ;
        RECT 376.950 125.400 388.050 126.600 ;
        RECT 376.950 124.950 379.050 125.400 ;
        RECT 385.950 124.950 388.050 125.400 ;
        RECT 412.950 124.950 415.050 127.050 ;
        RECT 418.950 126.600 421.050 127.050 ;
        RECT 436.950 126.600 439.050 127.050 ;
        RECT 454.950 126.600 457.050 127.050 ;
        RECT 418.950 125.400 457.050 126.600 ;
        RECT 418.950 124.950 421.050 125.400 ;
        RECT 436.950 124.950 439.050 125.400 ;
        RECT 454.950 124.950 457.050 125.400 ;
        RECT 475.950 126.600 478.050 127.050 ;
        RECT 487.950 126.600 490.050 127.050 ;
        RECT 493.950 126.600 496.050 127.050 ;
        RECT 475.950 125.400 490.050 126.600 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 487.950 124.950 490.050 125.400 ;
        RECT 491.400 125.400 496.050 126.600 ;
        RECT 127.950 123.600 130.050 124.050 ;
        RECT 119.400 122.400 130.050 123.600 ;
        RECT 109.950 121.950 112.050 122.400 ;
        RECT 115.950 121.950 118.050 122.400 ;
        RECT 127.950 121.950 130.050 122.400 ;
        RECT 208.950 123.600 211.050 124.050 ;
        RECT 235.950 123.600 238.050 124.050 ;
        RECT 208.950 122.400 238.050 123.600 ;
        RECT 208.950 121.950 211.050 122.400 ;
        RECT 235.950 121.950 238.050 122.400 ;
        RECT 274.950 123.600 277.050 124.050 ;
        RECT 286.950 123.600 289.050 124.050 ;
        RECT 289.950 123.600 292.050 124.050 ;
        RECT 274.950 122.400 292.050 123.600 ;
        RECT 274.950 121.950 277.050 122.400 ;
        RECT 286.950 121.950 289.050 122.400 ;
        RECT 289.950 121.950 292.050 122.400 ;
        RECT 295.950 123.600 298.050 124.050 ;
        RECT 331.950 123.600 334.050 124.050 ;
        RECT 295.950 122.400 334.050 123.600 ;
        RECT 295.950 121.950 298.050 122.400 ;
        RECT 331.950 121.950 334.050 122.400 ;
        RECT 349.950 123.600 352.050 124.050 ;
        RECT 391.950 123.600 394.050 124.050 ;
        RECT 349.950 122.400 394.050 123.600 ;
        RECT 349.950 121.950 352.050 122.400 ;
        RECT 391.950 121.950 394.050 122.400 ;
        RECT 403.950 123.600 406.050 124.050 ;
        RECT 415.950 123.600 418.050 124.050 ;
        RECT 448.950 123.600 451.050 124.050 ;
        RECT 403.950 122.400 451.050 123.600 ;
        RECT 403.950 121.950 406.050 122.400 ;
        RECT 415.950 121.950 418.050 122.400 ;
        RECT 448.950 121.950 451.050 122.400 ;
        RECT 460.950 123.600 463.050 124.050 ;
        RECT 478.950 123.600 481.050 124.050 ;
        RECT 491.400 123.600 492.600 125.400 ;
        RECT 493.950 124.950 496.050 125.400 ;
        RECT 502.950 126.600 505.050 127.050 ;
        RECT 508.950 126.600 511.050 127.050 ;
        RECT 502.950 125.400 511.050 126.600 ;
        RECT 502.950 124.950 505.050 125.400 ;
        RECT 508.950 124.950 511.050 125.400 ;
        RECT 535.950 126.600 538.050 127.050 ;
        RECT 550.950 126.600 553.050 127.050 ;
        RECT 535.950 125.400 553.050 126.600 ;
        RECT 535.950 124.950 538.050 125.400 ;
        RECT 550.950 124.950 553.050 125.400 ;
        RECT 556.950 124.950 559.050 127.050 ;
        RECT 571.950 126.600 574.050 127.050 ;
        RECT 577.950 126.600 580.050 127.050 ;
        RECT 583.950 126.600 586.050 127.050 ;
        RECT 571.950 125.400 586.050 126.600 ;
        RECT 571.950 124.950 574.050 125.400 ;
        RECT 577.950 124.950 580.050 125.400 ;
        RECT 583.950 124.950 586.050 125.400 ;
        RECT 610.950 124.950 613.050 127.050 ;
        RECT 616.950 126.600 619.050 127.050 ;
        RECT 631.950 126.600 634.050 127.050 ;
        RECT 616.950 125.400 634.050 126.600 ;
        RECT 616.950 124.950 619.050 125.400 ;
        RECT 631.950 124.950 634.050 125.400 ;
        RECT 640.950 126.600 643.050 127.050 ;
        RECT 649.950 126.600 652.050 127.050 ;
        RECT 640.950 125.400 652.050 126.600 ;
        RECT 653.400 126.600 654.600 128.400 ;
        RECT 655.950 128.400 670.050 129.600 ;
        RECT 655.950 127.950 658.050 128.400 ;
        RECT 667.950 127.950 670.050 128.400 ;
        RECT 673.950 127.950 676.050 130.050 ;
        RECT 700.950 129.600 703.050 130.050 ;
        RECT 718.950 129.600 721.050 130.050 ;
        RECT 724.950 129.600 727.050 130.050 ;
        RECT 700.950 128.400 717.600 129.600 ;
        RECT 700.950 127.950 703.050 128.400 ;
        RECT 674.400 126.600 675.600 127.950 ;
        RECT 653.400 125.400 675.600 126.600 ;
        RECT 697.950 126.600 700.050 127.050 ;
        RECT 709.950 126.600 712.050 127.050 ;
        RECT 697.950 125.400 712.050 126.600 ;
        RECT 716.400 126.600 717.600 128.400 ;
        RECT 718.950 128.400 727.050 129.600 ;
        RECT 718.950 127.950 721.050 128.400 ;
        RECT 724.950 127.950 727.050 128.400 ;
        RECT 742.950 126.600 745.050 127.050 ;
        RECT 716.400 125.400 745.050 126.600 ;
        RECT 640.950 124.950 643.050 125.400 ;
        RECT 649.950 124.950 652.050 125.400 ;
        RECT 697.950 124.950 700.050 125.400 ;
        RECT 709.950 124.950 712.050 125.400 ;
        RECT 742.950 124.950 745.050 125.400 ;
        RECT 757.950 124.950 760.050 127.050 ;
        RECT 763.950 126.600 766.050 127.050 ;
        RECT 769.950 126.600 772.050 127.050 ;
        RECT 763.950 125.400 772.050 126.600 ;
        RECT 763.950 124.950 766.050 125.400 ;
        RECT 769.950 124.950 772.050 125.400 ;
        RECT 832.950 126.600 835.050 127.050 ;
        RECT 880.950 126.600 883.050 127.050 ;
        RECT 832.950 125.400 883.050 126.600 ;
        RECT 832.950 124.950 835.050 125.400 ;
        RECT 880.950 124.950 883.050 125.400 ;
        RECT 460.950 122.400 492.600 123.600 ;
        RECT 496.950 123.600 499.050 124.050 ;
        RECT 547.950 123.600 550.050 124.050 ;
        RECT 496.950 122.400 550.050 123.600 ;
        RECT 460.950 121.950 463.050 122.400 ;
        RECT 478.950 121.950 481.050 122.400 ;
        RECT 496.950 121.950 499.050 122.400 ;
        RECT 547.950 121.950 550.050 122.400 ;
        RECT 592.950 123.600 595.050 124.050 ;
        RECT 611.400 123.600 612.600 124.950 ;
        RECT 592.950 122.400 612.600 123.600 ;
        RECT 646.950 123.600 649.050 124.050 ;
        RECT 652.950 123.600 655.050 124.050 ;
        RECT 646.950 122.400 655.050 123.600 ;
        RECT 592.950 121.950 595.050 122.400 ;
        RECT 646.950 121.950 649.050 122.400 ;
        RECT 652.950 121.950 655.050 122.400 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 694.950 123.600 697.050 124.050 ;
        RECT 706.950 123.600 709.050 124.050 ;
        RECT 676.950 122.400 709.050 123.600 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 694.950 121.950 697.050 122.400 ;
        RECT 706.950 121.950 709.050 122.400 ;
        RECT 721.950 123.600 724.050 124.050 ;
        RECT 739.950 123.600 742.050 124.050 ;
        RECT 758.400 123.600 759.600 124.950 ;
        RECT 721.950 122.400 738.600 123.600 ;
        RECT 721.950 121.950 724.050 122.400 ;
        RECT 16.950 120.600 19.050 121.050 ;
        RECT 88.950 120.600 91.050 121.050 ;
        RECT 16.950 119.400 91.050 120.600 ;
        RECT 16.950 118.950 19.050 119.400 ;
        RECT 88.950 118.950 91.050 119.400 ;
        RECT 214.950 120.600 217.050 121.050 ;
        RECT 244.950 120.600 247.050 121.050 ;
        RECT 262.950 120.600 265.050 121.050 ;
        RECT 214.950 119.400 265.050 120.600 ;
        RECT 214.950 118.950 217.050 119.400 ;
        RECT 244.950 118.950 247.050 119.400 ;
        RECT 262.950 118.950 265.050 119.400 ;
        RECT 289.950 120.600 292.050 121.050 ;
        RECT 364.950 120.600 367.050 121.050 ;
        RECT 373.950 120.600 376.050 121.050 ;
        RECT 289.950 119.400 376.050 120.600 ;
        RECT 289.950 118.950 292.050 119.400 ;
        RECT 364.950 118.950 367.050 119.400 ;
        RECT 373.950 118.950 376.050 119.400 ;
        RECT 469.950 120.600 472.050 121.050 ;
        RECT 490.950 120.600 493.050 121.050 ;
        RECT 469.950 119.400 493.050 120.600 ;
        RECT 469.950 118.950 472.050 119.400 ;
        RECT 490.950 118.950 493.050 119.400 ;
        RECT 511.950 120.600 514.050 121.050 ;
        RECT 538.950 120.600 541.050 121.050 ;
        RECT 511.950 119.400 541.050 120.600 ;
        RECT 511.950 118.950 514.050 119.400 ;
        RECT 538.950 118.950 541.050 119.400 ;
        RECT 553.950 120.600 556.050 121.050 ;
        RECT 619.950 120.600 622.050 121.050 ;
        RECT 634.950 120.600 637.050 121.050 ;
        RECT 553.950 119.400 637.050 120.600 ;
        RECT 553.950 118.950 556.050 119.400 ;
        RECT 619.950 118.950 622.050 119.400 ;
        RECT 634.950 118.950 637.050 119.400 ;
        RECT 658.950 120.600 661.050 121.050 ;
        RECT 685.950 120.600 688.050 121.050 ;
        RECT 733.950 120.600 736.050 121.050 ;
        RECT 658.950 119.400 736.050 120.600 ;
        RECT 737.400 120.600 738.600 122.400 ;
        RECT 739.950 122.400 759.600 123.600 ;
        RECT 760.950 123.600 763.050 124.050 ;
        RECT 820.950 123.600 823.050 124.050 ;
        RECT 760.950 122.400 823.050 123.600 ;
        RECT 739.950 121.950 742.050 122.400 ;
        RECT 760.950 121.950 763.050 122.400 ;
        RECT 820.950 121.950 823.050 122.400 ;
        RECT 823.950 123.600 826.050 124.050 ;
        RECT 844.950 123.600 847.050 124.050 ;
        RECT 823.950 122.400 847.050 123.600 ;
        RECT 823.950 121.950 826.050 122.400 ;
        RECT 844.950 121.950 847.050 122.400 ;
        RECT 862.950 123.600 865.050 124.050 ;
        RECT 862.950 122.400 879.600 123.600 ;
        RECT 862.950 121.950 865.050 122.400 ;
        RECT 878.400 121.050 879.600 122.400 ;
        RECT 754.950 120.600 757.050 121.050 ;
        RECT 737.400 119.400 757.050 120.600 ;
        RECT 658.950 118.950 661.050 119.400 ;
        RECT 685.950 118.950 688.050 119.400 ;
        RECT 733.950 118.950 736.050 119.400 ;
        RECT 754.950 118.950 757.050 119.400 ;
        RECT 877.950 118.950 880.050 121.050 ;
        RECT 184.950 117.600 187.050 118.050 ;
        RECT 217.950 117.600 220.050 118.050 ;
        RECT 184.950 116.400 220.050 117.600 ;
        RECT 184.950 115.950 187.050 116.400 ;
        RECT 217.950 115.950 220.050 116.400 ;
        RECT 268.950 117.600 271.050 118.050 ;
        RECT 316.950 117.600 319.050 118.050 ;
        RECT 268.950 116.400 319.050 117.600 ;
        RECT 268.950 115.950 271.050 116.400 ;
        RECT 316.950 115.950 319.050 116.400 ;
        RECT 343.950 117.600 346.050 118.050 ;
        RECT 355.950 117.600 358.050 118.050 ;
        RECT 343.950 116.400 358.050 117.600 ;
        RECT 343.950 115.950 346.050 116.400 ;
        RECT 355.950 115.950 358.050 116.400 ;
        RECT 361.950 117.600 364.050 118.050 ;
        RECT 370.950 117.600 373.050 118.050 ;
        RECT 406.950 117.600 409.050 118.050 ;
        RECT 361.950 116.400 409.050 117.600 ;
        RECT 361.950 115.950 364.050 116.400 ;
        RECT 370.950 115.950 373.050 116.400 ;
        RECT 406.950 115.950 409.050 116.400 ;
        RECT 433.950 117.600 436.050 118.050 ;
        RECT 514.950 117.600 517.050 118.050 ;
        RECT 433.950 116.400 517.050 117.600 ;
        RECT 433.950 115.950 436.050 116.400 ;
        RECT 514.950 115.950 517.050 116.400 ;
        RECT 634.950 117.600 637.050 118.050 ;
        RECT 691.950 117.600 694.050 118.050 ;
        RECT 715.950 117.600 718.050 118.050 ;
        RECT 634.950 116.400 718.050 117.600 ;
        RECT 634.950 115.950 637.050 116.400 ;
        RECT 691.950 115.950 694.050 116.400 ;
        RECT 715.950 115.950 718.050 116.400 ;
        RECT 154.950 114.600 157.050 115.050 ;
        RECT 196.950 114.600 199.050 115.050 ;
        RECT 268.950 114.600 271.050 115.050 ;
        RECT 154.950 113.400 271.050 114.600 ;
        RECT 154.950 112.950 157.050 113.400 ;
        RECT 196.950 112.950 199.050 113.400 ;
        RECT 268.950 112.950 271.050 113.400 ;
        RECT 502.950 114.600 505.050 115.050 ;
        RECT 568.950 114.600 571.050 115.050 ;
        RECT 502.950 113.400 571.050 114.600 ;
        RECT 502.950 112.950 505.050 113.400 ;
        RECT 568.950 112.950 571.050 113.400 ;
        RECT 697.950 114.600 700.050 115.050 ;
        RECT 799.950 114.600 802.050 115.050 ;
        RECT 697.950 113.400 802.050 114.600 ;
        RECT 697.950 112.950 700.050 113.400 ;
        RECT 799.950 112.950 802.050 113.400 ;
        RECT 127.950 111.600 130.050 112.050 ;
        RECT 202.950 111.600 205.050 112.050 ;
        RECT 127.950 110.400 205.050 111.600 ;
        RECT 127.950 109.950 130.050 110.400 ;
        RECT 202.950 109.950 205.050 110.400 ;
        RECT 265.950 111.600 268.050 112.050 ;
        RECT 325.950 111.600 328.050 112.050 ;
        RECT 352.950 111.600 355.050 112.050 ;
        RECT 265.950 110.400 355.050 111.600 ;
        RECT 265.950 109.950 268.050 110.400 ;
        RECT 325.950 109.950 328.050 110.400 ;
        RECT 352.950 109.950 355.050 110.400 ;
        RECT 355.950 111.600 358.050 112.050 ;
        RECT 427.950 111.600 430.050 112.050 ;
        RECT 355.950 110.400 430.050 111.600 ;
        RECT 355.950 109.950 358.050 110.400 ;
        RECT 427.950 109.950 430.050 110.400 ;
        RECT 121.950 108.600 124.050 109.050 ;
        RECT 142.950 108.600 145.050 109.050 ;
        RECT 121.950 107.400 145.050 108.600 ;
        RECT 121.950 106.950 124.050 107.400 ;
        RECT 142.950 106.950 145.050 107.400 ;
        RECT 190.950 108.600 193.050 109.050 ;
        RECT 271.950 108.600 274.050 109.050 ;
        RECT 190.950 107.400 274.050 108.600 ;
        RECT 190.950 106.950 193.050 107.400 ;
        RECT 271.950 106.950 274.050 107.400 ;
        RECT 352.950 108.600 355.050 109.050 ;
        RECT 364.950 108.600 367.050 109.050 ;
        RECT 391.950 108.600 394.050 109.050 ;
        RECT 352.950 107.400 394.050 108.600 ;
        RECT 352.950 106.950 355.050 107.400 ;
        RECT 364.950 106.950 367.050 107.400 ;
        RECT 391.950 106.950 394.050 107.400 ;
        RECT 451.950 108.600 454.050 109.050 ;
        RECT 502.950 108.600 505.050 109.050 ;
        RECT 451.950 107.400 505.050 108.600 ;
        RECT 451.950 106.950 454.050 107.400 ;
        RECT 502.950 106.950 505.050 107.400 ;
        RECT 565.950 108.600 568.050 109.050 ;
        RECT 586.950 108.600 589.050 109.050 ;
        RECT 565.950 107.400 589.050 108.600 ;
        RECT 565.950 106.950 568.050 107.400 ;
        RECT 586.950 106.950 589.050 107.400 ;
        RECT 634.950 108.600 637.050 109.050 ;
        RECT 667.950 108.600 670.050 109.050 ;
        RECT 634.950 107.400 670.050 108.600 ;
        RECT 634.950 106.950 637.050 107.400 ;
        RECT 667.950 106.950 670.050 107.400 ;
        RECT 835.950 108.600 838.050 109.050 ;
        RECT 853.950 108.600 856.050 109.050 ;
        RECT 835.950 107.400 856.050 108.600 ;
        RECT 835.950 106.950 838.050 107.400 ;
        RECT 853.950 106.950 856.050 107.400 ;
        RECT 97.950 105.600 100.050 106.050 ;
        RECT 295.950 105.600 298.050 106.050 ;
        RECT 97.950 104.400 298.050 105.600 ;
        RECT 97.950 103.950 100.050 104.400 ;
        RECT 295.950 103.950 298.050 104.400 ;
        RECT 349.950 105.600 352.050 106.050 ;
        RECT 415.950 105.600 418.050 106.050 ;
        RECT 349.950 104.400 418.050 105.600 ;
        RECT 349.950 103.950 352.050 104.400 ;
        RECT 415.950 103.950 418.050 104.400 ;
        RECT 496.950 105.600 499.050 106.050 ;
        RECT 595.950 105.600 598.050 106.050 ;
        RECT 496.950 104.400 598.050 105.600 ;
        RECT 496.950 103.950 499.050 104.400 ;
        RECT 595.950 103.950 598.050 104.400 ;
        RECT 655.950 105.600 658.050 106.050 ;
        RECT 676.950 105.600 679.050 106.050 ;
        RECT 655.950 104.400 679.050 105.600 ;
        RECT 655.950 103.950 658.050 104.400 ;
        RECT 676.950 103.950 679.050 104.400 ;
        RECT 682.950 105.600 685.050 106.050 ;
        RECT 766.950 105.600 769.050 106.050 ;
        RECT 682.950 104.400 769.050 105.600 ;
        RECT 682.950 103.950 685.050 104.400 ;
        RECT 766.950 103.950 769.050 104.400 ;
        RECT 826.950 105.600 829.050 106.050 ;
        RECT 841.950 105.600 844.050 106.050 ;
        RECT 826.950 104.400 844.050 105.600 ;
        RECT 826.950 103.950 829.050 104.400 ;
        RECT 841.950 103.950 844.050 104.400 ;
        RECT 34.950 102.600 37.050 103.050 ;
        RECT 55.950 102.600 58.050 103.050 ;
        RECT 91.950 102.600 94.050 103.050 ;
        RECT 34.950 101.400 94.050 102.600 ;
        RECT 34.950 100.950 37.050 101.400 ;
        RECT 55.950 100.950 58.050 101.400 ;
        RECT 91.950 100.950 94.050 101.400 ;
        RECT 118.950 102.600 121.050 103.050 ;
        RECT 130.950 102.600 133.050 103.050 ;
        RECT 118.950 101.400 133.050 102.600 ;
        RECT 118.950 100.950 121.050 101.400 ;
        RECT 130.950 100.950 133.050 101.400 ;
        RECT 148.950 102.600 151.050 103.050 ;
        RECT 172.950 102.600 175.050 103.050 ;
        RECT 244.950 102.600 247.050 103.050 ;
        RECT 148.950 101.400 247.050 102.600 ;
        RECT 148.950 100.950 151.050 101.400 ;
        RECT 172.950 100.950 175.050 101.400 ;
        RECT 244.950 100.950 247.050 101.400 ;
        RECT 247.950 102.600 250.050 103.050 ;
        RECT 268.950 102.600 271.050 103.050 ;
        RECT 247.950 101.400 271.050 102.600 ;
        RECT 247.950 100.950 250.050 101.400 ;
        RECT 268.950 100.950 271.050 101.400 ;
        RECT 304.950 102.600 307.050 103.050 ;
        RECT 334.950 102.600 337.050 103.050 ;
        RECT 352.950 102.600 355.050 103.050 ;
        RECT 304.950 101.400 355.050 102.600 ;
        RECT 304.950 100.950 307.050 101.400 ;
        RECT 334.950 100.950 337.050 101.400 ;
        RECT 352.950 100.950 355.050 101.400 ;
        RECT 454.950 102.600 457.050 103.050 ;
        RECT 463.950 102.600 466.050 103.050 ;
        RECT 472.950 102.600 475.050 103.050 ;
        RECT 454.950 101.400 475.050 102.600 ;
        RECT 454.950 100.950 457.050 101.400 ;
        RECT 463.950 100.950 466.050 101.400 ;
        RECT 472.950 100.950 475.050 101.400 ;
        RECT 562.950 102.600 565.050 103.050 ;
        RECT 574.950 102.600 577.050 103.050 ;
        RECT 562.950 101.400 577.050 102.600 ;
        RECT 562.950 100.950 565.050 101.400 ;
        RECT 574.950 100.950 577.050 101.400 ;
        RECT 763.950 102.600 766.050 103.050 ;
        RECT 766.950 102.600 769.050 103.050 ;
        RECT 805.950 102.600 808.050 103.050 ;
        RECT 850.950 102.600 853.050 103.050 ;
        RECT 763.950 101.400 853.050 102.600 ;
        RECT 763.950 100.950 766.050 101.400 ;
        RECT 766.950 100.950 769.050 101.400 ;
        RECT 805.950 100.950 808.050 101.400 ;
        RECT 850.950 100.950 853.050 101.400 ;
        RECT 121.950 99.600 124.050 100.050 ;
        RECT 151.950 99.600 154.050 100.050 ;
        RECT 121.950 98.400 154.050 99.600 ;
        RECT 121.950 97.950 124.050 98.400 ;
        RECT 151.950 97.950 154.050 98.400 ;
        RECT 172.950 99.600 175.050 100.050 ;
        RECT 181.950 99.600 184.050 100.050 ;
        RECT 172.950 98.400 184.050 99.600 ;
        RECT 172.950 97.950 175.050 98.400 ;
        RECT 181.950 97.950 184.050 98.400 ;
        RECT 220.950 99.600 223.050 100.050 ;
        RECT 265.950 99.600 268.050 100.050 ;
        RECT 220.950 98.400 268.050 99.600 ;
        RECT 220.950 97.950 223.050 98.400 ;
        RECT 265.950 97.950 268.050 98.400 ;
        RECT 271.950 99.600 274.050 100.050 ;
        RECT 361.950 99.600 364.050 100.050 ;
        RECT 271.950 98.400 364.050 99.600 ;
        RECT 271.950 97.950 274.050 98.400 ;
        RECT 361.950 97.950 364.050 98.400 ;
        RECT 421.950 99.600 424.050 100.050 ;
        RECT 424.950 99.600 427.050 100.050 ;
        RECT 430.950 99.600 433.050 100.050 ;
        RECT 421.950 98.400 433.050 99.600 ;
        RECT 421.950 97.950 424.050 98.400 ;
        RECT 424.950 97.950 427.050 98.400 ;
        RECT 430.950 97.950 433.050 98.400 ;
        RECT 472.950 99.600 475.050 100.050 ;
        RECT 517.950 99.600 520.050 100.050 ;
        RECT 529.950 99.600 532.050 100.050 ;
        RECT 664.950 99.600 667.050 100.050 ;
        RECT 472.950 98.400 528.600 99.600 ;
        RECT 472.950 97.950 475.050 98.400 ;
        RECT 517.950 97.950 520.050 98.400 ;
        RECT 46.950 96.600 49.050 97.050 ;
        RECT 61.950 96.600 64.050 97.050 ;
        RECT 32.400 95.400 64.050 96.600 ;
        RECT 32.400 94.050 33.600 95.400 ;
        RECT 46.950 94.950 49.050 95.400 ;
        RECT 61.950 94.950 64.050 95.400 ;
        RECT 73.950 96.600 76.050 97.050 ;
        RECT 91.950 96.600 94.050 97.050 ;
        RECT 124.950 96.600 127.050 97.050 ;
        RECT 127.950 96.600 130.050 97.050 ;
        RECT 73.950 95.400 78.600 96.600 ;
        RECT 73.950 94.950 76.050 95.400 ;
        RECT 31.950 93.600 34.050 94.050 ;
        RECT 34.950 93.600 37.050 94.050 ;
        RECT 31.950 92.400 37.050 93.600 ;
        RECT 31.950 91.950 34.050 92.400 ;
        RECT 34.950 91.950 37.050 92.400 ;
        RECT 73.950 91.950 76.050 94.050 ;
        RECT 74.400 87.600 75.600 91.950 ;
        RECT 77.400 91.050 78.600 95.400 ;
        RECT 91.950 95.400 130.050 96.600 ;
        RECT 91.950 94.950 94.050 95.400 ;
        RECT 124.950 94.950 127.050 95.400 ;
        RECT 127.950 94.950 130.050 95.400 ;
        RECT 136.950 96.600 139.050 97.050 ;
        RECT 148.950 96.600 151.050 97.050 ;
        RECT 154.950 96.600 157.050 97.050 ;
        RECT 136.950 95.400 151.050 96.600 ;
        RECT 136.950 94.950 139.050 95.400 ;
        RECT 148.950 94.950 151.050 95.400 ;
        RECT 152.400 95.400 157.050 96.600 ;
        RECT 79.950 93.600 82.050 94.050 ;
        RECT 109.950 93.600 112.050 94.050 ;
        RECT 79.950 92.400 112.050 93.600 ;
        RECT 79.950 91.950 82.050 92.400 ;
        RECT 109.950 91.950 112.050 92.400 ;
        RECT 133.950 93.600 136.050 94.050 ;
        RECT 152.400 93.600 153.600 95.400 ;
        RECT 154.950 94.950 157.050 95.400 ;
        RECT 187.950 96.600 190.050 97.050 ;
        RECT 247.950 96.600 250.050 97.050 ;
        RECT 187.950 95.400 250.050 96.600 ;
        RECT 187.950 94.950 190.050 95.400 ;
        RECT 247.950 94.950 250.050 95.400 ;
        RECT 256.950 96.600 259.050 97.050 ;
        RECT 289.950 96.600 292.050 97.050 ;
        RECT 256.950 95.400 292.050 96.600 ;
        RECT 256.950 94.950 259.050 95.400 ;
        RECT 289.950 94.950 292.050 95.400 ;
        RECT 295.950 96.600 298.050 97.050 ;
        RECT 322.950 96.600 325.050 97.050 ;
        RECT 370.950 96.600 373.050 97.050 ;
        RECT 379.950 96.600 382.050 97.050 ;
        RECT 295.950 95.400 309.600 96.600 ;
        RECT 295.950 94.950 298.050 95.400 ;
        RECT 308.400 94.050 309.600 95.400 ;
        RECT 322.950 95.400 348.600 96.600 ;
        RECT 322.950 94.950 325.050 95.400 ;
        RECT 347.400 94.050 348.600 95.400 ;
        RECT 370.950 95.400 382.050 96.600 ;
        RECT 370.950 94.950 373.050 95.400 ;
        RECT 379.950 94.950 382.050 95.400 ;
        RECT 382.950 96.600 385.050 97.050 ;
        RECT 409.950 96.600 412.050 97.050 ;
        RECT 382.950 95.400 412.050 96.600 ;
        RECT 382.950 94.950 385.050 95.400 ;
        RECT 409.950 94.950 412.050 95.400 ;
        RECT 448.950 96.600 451.050 97.050 ;
        RECT 466.950 96.600 469.050 97.050 ;
        RECT 448.950 95.400 469.050 96.600 ;
        RECT 527.400 96.600 528.600 98.400 ;
        RECT 529.950 98.400 667.050 99.600 ;
        RECT 529.950 97.950 532.050 98.400 ;
        RECT 664.950 97.950 667.050 98.400 ;
        RECT 820.950 99.600 823.050 100.050 ;
        RECT 856.950 99.600 859.050 100.050 ;
        RECT 859.950 99.600 862.050 100.050 ;
        RECT 820.950 98.400 862.050 99.600 ;
        RECT 820.950 97.950 823.050 98.400 ;
        RECT 856.950 97.950 859.050 98.400 ;
        RECT 859.950 97.950 862.050 98.400 ;
        RECT 565.950 96.600 568.050 97.050 ;
        RECT 527.400 95.400 568.050 96.600 ;
        RECT 448.950 94.950 451.050 95.400 ;
        RECT 466.950 94.950 469.050 95.400 ;
        RECT 565.950 94.950 568.050 95.400 ;
        RECT 574.950 96.600 577.050 97.050 ;
        RECT 592.950 96.600 595.050 97.050 ;
        RECT 613.950 96.600 616.050 97.050 ;
        RECT 631.950 96.600 634.050 97.050 ;
        RECT 667.950 96.600 670.050 97.050 ;
        RECT 574.950 95.400 630.600 96.600 ;
        RECT 574.950 94.950 577.050 95.400 ;
        RECT 592.950 94.950 595.050 95.400 ;
        RECT 613.950 94.950 616.050 95.400 ;
        RECT 133.950 92.400 153.600 93.600 ;
        RECT 211.950 93.600 214.050 94.050 ;
        RECT 250.950 93.600 253.050 94.050 ;
        RECT 211.950 92.400 253.050 93.600 ;
        RECT 133.950 91.950 136.050 92.400 ;
        RECT 211.950 91.950 214.050 92.400 ;
        RECT 250.950 91.950 253.050 92.400 ;
        RECT 286.950 93.600 289.050 94.050 ;
        RECT 304.950 93.600 307.050 94.050 ;
        RECT 286.950 92.400 307.050 93.600 ;
        RECT 286.950 91.950 289.050 92.400 ;
        RECT 304.950 91.950 307.050 92.400 ;
        RECT 307.950 91.950 310.050 94.050 ;
        RECT 328.950 93.600 331.050 94.050 ;
        RECT 311.400 92.400 331.050 93.600 ;
        RECT 76.950 88.950 79.050 91.050 ;
        RECT 112.950 90.600 115.050 91.050 ;
        RECT 121.950 90.600 124.050 91.050 ;
        RECT 130.950 90.600 133.050 91.050 ;
        RECT 112.950 89.400 133.050 90.600 ;
        RECT 112.950 88.950 115.050 89.400 ;
        RECT 121.950 88.950 124.050 89.400 ;
        RECT 130.950 88.950 133.050 89.400 ;
        RECT 169.950 90.600 172.050 91.050 ;
        RECT 190.950 90.600 193.050 91.050 ;
        RECT 169.950 89.400 193.050 90.600 ;
        RECT 169.950 88.950 172.050 89.400 ;
        RECT 190.950 88.950 193.050 89.400 ;
        RECT 208.950 90.600 211.050 91.050 ;
        RECT 232.950 90.600 235.050 91.050 ;
        RECT 208.950 89.400 235.050 90.600 ;
        RECT 208.950 88.950 211.050 89.400 ;
        RECT 232.950 88.950 235.050 89.400 ;
        RECT 292.950 90.600 295.050 91.050 ;
        RECT 295.950 90.600 298.050 91.050 ;
        RECT 311.400 90.600 312.600 92.400 ;
        RECT 328.950 91.950 331.050 92.400 ;
        RECT 346.950 91.950 349.050 94.050 ;
        RECT 361.950 93.600 364.050 94.050 ;
        RECT 367.950 93.600 370.050 94.050 ;
        RECT 361.950 92.400 370.050 93.600 ;
        RECT 361.950 91.950 364.050 92.400 ;
        RECT 367.950 91.950 370.050 92.400 ;
        RECT 373.950 93.600 376.050 94.050 ;
        RECT 388.950 93.600 391.050 94.050 ;
        RECT 373.950 92.400 391.050 93.600 ;
        RECT 373.950 91.950 376.050 92.400 ;
        RECT 388.950 91.950 391.050 92.400 ;
        RECT 394.950 93.600 397.050 94.050 ;
        RECT 406.950 93.600 409.050 94.050 ;
        RECT 394.950 92.400 409.050 93.600 ;
        RECT 394.950 91.950 397.050 92.400 ;
        RECT 406.950 91.950 409.050 92.400 ;
        RECT 433.950 93.600 436.050 94.050 ;
        RECT 439.950 93.600 442.050 94.050 ;
        RECT 433.950 92.400 442.050 93.600 ;
        RECT 433.950 91.950 436.050 92.400 ;
        RECT 439.950 91.950 442.050 92.400 ;
        RECT 481.950 93.600 484.050 94.050 ;
        RECT 493.950 93.600 496.050 94.050 ;
        RECT 481.950 92.400 496.050 93.600 ;
        RECT 481.950 91.950 484.050 92.400 ;
        RECT 493.950 91.950 496.050 92.400 ;
        RECT 499.950 93.600 502.050 94.050 ;
        RECT 514.950 93.600 517.050 94.050 ;
        RECT 499.950 92.400 517.050 93.600 ;
        RECT 499.950 91.950 502.050 92.400 ;
        RECT 514.950 91.950 517.050 92.400 ;
        RECT 568.950 93.600 571.050 94.050 ;
        RECT 577.950 93.600 580.050 94.050 ;
        RECT 589.950 93.600 592.050 94.050 ;
        RECT 568.950 92.400 580.050 93.600 ;
        RECT 568.950 91.950 571.050 92.400 ;
        RECT 577.950 91.950 580.050 92.400 ;
        RECT 581.400 92.400 592.050 93.600 ;
        RECT 292.950 89.400 312.600 90.600 ;
        RECT 397.950 90.600 400.050 91.050 ;
        RECT 412.950 90.600 415.050 91.050 ;
        RECT 397.950 89.400 415.050 90.600 ;
        RECT 292.950 88.950 295.050 89.400 ;
        RECT 295.950 88.950 298.050 89.400 ;
        RECT 397.950 88.950 400.050 89.400 ;
        RECT 412.950 88.950 415.050 89.400 ;
        RECT 463.950 90.600 466.050 91.050 ;
        RECT 475.950 90.600 478.050 91.050 ;
        RECT 463.950 89.400 478.050 90.600 ;
        RECT 463.950 88.950 466.050 89.400 ;
        RECT 475.950 88.950 478.050 89.400 ;
        RECT 541.950 90.600 544.050 91.050 ;
        RECT 581.400 90.600 582.600 92.400 ;
        RECT 589.950 91.950 592.050 92.400 ;
        RECT 595.950 93.600 598.050 94.050 ;
        RECT 607.950 93.600 610.050 94.050 ;
        RECT 595.950 92.400 610.050 93.600 ;
        RECT 595.950 91.950 598.050 92.400 ;
        RECT 607.950 91.950 610.050 92.400 ;
        RECT 613.950 93.600 616.050 94.050 ;
        RECT 622.950 93.600 625.050 94.050 ;
        RECT 613.950 92.400 625.050 93.600 ;
        RECT 629.400 93.600 630.600 95.400 ;
        RECT 631.950 95.400 670.050 96.600 ;
        RECT 631.950 94.950 634.050 95.400 ;
        RECT 667.950 94.950 670.050 95.400 ;
        RECT 718.950 96.600 721.050 97.050 ;
        RECT 727.950 96.600 730.050 97.050 ;
        RECT 718.950 95.400 730.050 96.600 ;
        RECT 718.950 94.950 721.050 95.400 ;
        RECT 727.950 94.950 730.050 95.400 ;
        RECT 772.950 96.600 775.050 97.050 ;
        RECT 781.950 96.600 784.050 97.050 ;
        RECT 772.950 95.400 784.050 96.600 ;
        RECT 772.950 94.950 775.050 95.400 ;
        RECT 781.950 94.950 784.050 95.400 ;
        RECT 799.950 96.600 802.050 97.050 ;
        RECT 838.950 96.600 841.050 97.050 ;
        RECT 799.950 95.400 841.050 96.600 ;
        RECT 799.950 94.950 802.050 95.400 ;
        RECT 838.950 94.950 841.050 95.400 ;
        RECT 634.950 93.600 637.050 94.050 ;
        RECT 629.400 92.400 637.050 93.600 ;
        RECT 613.950 91.950 616.050 92.400 ;
        RECT 622.950 91.950 625.050 92.400 ;
        RECT 634.950 91.950 637.050 92.400 ;
        RECT 658.950 93.600 661.050 94.050 ;
        RECT 673.950 93.600 676.050 94.050 ;
        RECT 658.950 92.400 676.050 93.600 ;
        RECT 658.950 91.950 661.050 92.400 ;
        RECT 673.950 91.950 676.050 92.400 ;
        RECT 688.950 93.600 691.050 94.050 ;
        RECT 730.950 93.600 733.050 94.050 ;
        RECT 688.950 92.400 733.050 93.600 ;
        RECT 688.950 91.950 691.050 92.400 ;
        RECT 730.950 91.950 733.050 92.400 ;
        RECT 745.950 93.600 748.050 94.050 ;
        RECT 775.950 93.600 778.050 94.050 ;
        RECT 745.950 92.400 778.050 93.600 ;
        RECT 745.950 91.950 748.050 92.400 ;
        RECT 775.950 91.950 778.050 92.400 ;
        RECT 790.950 93.600 793.050 94.050 ;
        RECT 817.950 93.600 820.050 94.050 ;
        RECT 790.950 92.400 820.050 93.600 ;
        RECT 790.950 91.950 793.050 92.400 ;
        RECT 817.950 91.950 820.050 92.400 ;
        RECT 826.950 93.600 829.050 94.050 ;
        RECT 841.950 93.600 844.050 94.050 ;
        RECT 826.950 92.400 844.050 93.600 ;
        RECT 826.950 91.950 829.050 92.400 ;
        RECT 841.950 91.950 844.050 92.400 ;
        RECT 847.950 93.600 850.050 94.050 ;
        RECT 856.950 93.600 859.050 94.050 ;
        RECT 847.950 92.400 859.050 93.600 ;
        RECT 847.950 91.950 850.050 92.400 ;
        RECT 856.950 91.950 859.050 92.400 ;
        RECT 871.950 93.600 874.050 94.050 ;
        RECT 877.950 93.600 880.050 94.050 ;
        RECT 871.950 92.400 880.050 93.600 ;
        RECT 871.950 91.950 874.050 92.400 ;
        RECT 877.950 91.950 880.050 92.400 ;
        RECT 541.950 89.400 582.600 90.600 ;
        RECT 625.950 90.600 628.050 91.050 ;
        RECT 652.950 90.600 655.050 91.050 ;
        RECT 769.950 90.600 772.050 91.050 ;
        RECT 835.950 90.600 838.050 91.050 ;
        RECT 625.950 89.400 838.050 90.600 ;
        RECT 541.950 88.950 544.050 89.400 ;
        RECT 625.950 88.950 628.050 89.400 ;
        RECT 652.950 88.950 655.050 89.400 ;
        RECT 769.950 88.950 772.050 89.400 ;
        RECT 835.950 88.950 838.050 89.400 ;
        RECT 865.950 90.600 868.050 91.050 ;
        RECT 874.950 90.600 877.050 91.050 ;
        RECT 865.950 89.400 877.050 90.600 ;
        RECT 865.950 88.950 868.050 89.400 ;
        RECT 874.950 88.950 877.050 89.400 ;
        RECT 253.950 87.600 256.050 88.050 ;
        RECT 74.400 86.400 256.050 87.600 ;
        RECT 253.950 85.950 256.050 86.400 ;
        RECT 520.950 87.600 523.050 88.050 ;
        RECT 547.950 87.600 550.050 88.050 ;
        RECT 646.950 87.600 649.050 88.050 ;
        RECT 520.950 86.400 649.050 87.600 ;
        RECT 520.950 85.950 523.050 86.400 ;
        RECT 547.950 85.950 550.050 86.400 ;
        RECT 646.950 85.950 649.050 86.400 ;
        RECT 829.950 87.600 832.050 88.050 ;
        RECT 838.950 87.600 841.050 88.050 ;
        RECT 829.950 86.400 841.050 87.600 ;
        RECT 829.950 85.950 832.050 86.400 ;
        RECT 838.950 85.950 841.050 86.400 ;
        RECT 853.950 87.600 856.050 88.050 ;
        RECT 868.950 87.600 871.050 88.050 ;
        RECT 853.950 86.400 871.050 87.600 ;
        RECT 853.950 85.950 856.050 86.400 ;
        RECT 868.950 85.950 871.050 86.400 ;
        RECT 37.950 84.600 40.050 85.050 ;
        RECT 49.950 84.600 52.050 85.050 ;
        RECT 79.950 84.600 82.050 85.050 ;
        RECT 37.950 83.400 82.050 84.600 ;
        RECT 37.950 82.950 40.050 83.400 ;
        RECT 49.950 82.950 52.050 83.400 ;
        RECT 79.950 82.950 82.050 83.400 ;
        RECT 493.950 84.600 496.050 85.050 ;
        RECT 532.950 84.600 535.050 85.050 ;
        RECT 493.950 83.400 535.050 84.600 ;
        RECT 493.950 82.950 496.050 83.400 ;
        RECT 532.950 82.950 535.050 83.400 ;
        RECT 628.950 84.600 631.050 85.050 ;
        RECT 703.950 84.600 706.050 85.050 ;
        RECT 628.950 83.400 706.050 84.600 ;
        RECT 628.950 82.950 631.050 83.400 ;
        RECT 703.950 82.950 706.050 83.400 ;
        RECT 292.950 81.600 295.050 82.050 ;
        RECT 637.950 81.600 640.050 82.050 ;
        RECT 292.950 80.400 640.050 81.600 ;
        RECT 292.950 79.950 295.050 80.400 ;
        RECT 637.950 79.950 640.050 80.400 ;
        RECT 157.950 75.600 160.050 76.050 ;
        RECT 340.950 75.600 343.050 76.050 ;
        RECT 157.950 74.400 343.050 75.600 ;
        RECT 157.950 73.950 160.050 74.400 ;
        RECT 340.950 73.950 343.050 74.400 ;
        RECT 361.950 72.600 364.050 73.050 ;
        RECT 526.950 72.600 529.050 73.050 ;
        RECT 361.950 71.400 529.050 72.600 ;
        RECT 361.950 70.950 364.050 71.400 ;
        RECT 526.950 70.950 529.050 71.400 ;
        RECT 604.950 69.600 607.050 70.050 ;
        RECT 622.950 69.600 625.050 70.050 ;
        RECT 604.950 68.400 625.050 69.600 ;
        RECT 604.950 67.950 607.050 68.400 ;
        RECT 622.950 67.950 625.050 68.400 ;
        RECT 307.950 66.600 310.050 67.050 ;
        RECT 352.950 66.600 355.050 67.050 ;
        RECT 307.950 65.400 355.050 66.600 ;
        RECT 307.950 64.950 310.050 65.400 ;
        RECT 352.950 64.950 355.050 65.400 ;
        RECT 418.950 66.600 421.050 67.050 ;
        RECT 478.950 66.600 481.050 67.050 ;
        RECT 418.950 65.400 481.050 66.600 ;
        RECT 418.950 64.950 421.050 65.400 ;
        RECT 478.950 64.950 481.050 65.400 ;
        RECT 586.950 66.600 589.050 67.050 ;
        RECT 637.950 66.600 640.050 67.050 ;
        RECT 586.950 65.400 640.050 66.600 ;
        RECT 586.950 64.950 589.050 65.400 ;
        RECT 637.950 64.950 640.050 65.400 ;
        RECT 730.950 66.600 733.050 67.050 ;
        RECT 757.950 66.600 760.050 67.050 ;
        RECT 778.950 66.600 781.050 67.050 ;
        RECT 730.950 65.400 781.050 66.600 ;
        RECT 730.950 64.950 733.050 65.400 ;
        RECT 757.950 64.950 760.050 65.400 ;
        RECT 778.950 64.950 781.050 65.400 ;
        RECT 109.950 63.600 112.050 64.050 ;
        RECT 118.950 63.600 121.050 64.050 ;
        RECT 109.950 62.400 121.050 63.600 ;
        RECT 109.950 61.950 112.050 62.400 ;
        RECT 118.950 61.950 121.050 62.400 ;
        RECT 304.950 63.600 307.050 64.050 ;
        RECT 325.950 63.600 328.050 64.050 ;
        RECT 304.950 62.400 328.050 63.600 ;
        RECT 304.950 61.950 307.050 62.400 ;
        RECT 325.950 61.950 328.050 62.400 ;
        RECT 397.950 63.600 400.050 64.050 ;
        RECT 475.950 63.600 478.050 64.050 ;
        RECT 397.950 62.400 478.050 63.600 ;
        RECT 397.950 61.950 400.050 62.400 ;
        RECT 475.950 61.950 478.050 62.400 ;
        RECT 478.950 63.600 481.050 64.050 ;
        RECT 610.950 63.600 613.050 64.050 ;
        RECT 613.950 63.600 616.050 64.050 ;
        RECT 478.950 62.400 616.050 63.600 ;
        RECT 478.950 61.950 481.050 62.400 ;
        RECT 610.950 61.950 613.050 62.400 ;
        RECT 613.950 61.950 616.050 62.400 ;
        RECT 619.950 63.600 622.050 64.050 ;
        RECT 652.950 63.600 655.050 64.050 ;
        RECT 619.950 62.400 655.050 63.600 ;
        RECT 619.950 61.950 622.050 62.400 ;
        RECT 652.950 61.950 655.050 62.400 ;
        RECT 658.950 63.600 661.050 64.050 ;
        RECT 664.950 63.600 667.050 64.050 ;
        RECT 670.950 63.600 673.050 64.050 ;
        RECT 811.950 63.600 814.050 64.050 ;
        RECT 658.950 62.400 814.050 63.600 ;
        RECT 658.950 61.950 661.050 62.400 ;
        RECT 664.950 61.950 667.050 62.400 ;
        RECT 670.950 61.950 673.050 62.400 ;
        RECT 811.950 61.950 814.050 62.400 ;
        RECT 10.950 60.600 13.050 61.050 ;
        RECT 61.950 60.600 64.050 61.050 ;
        RECT 10.950 59.400 64.050 60.600 ;
        RECT 10.950 58.950 13.050 59.400 ;
        RECT 61.950 58.950 64.050 59.400 ;
        RECT 118.950 60.600 121.050 61.050 ;
        RECT 124.950 60.600 127.050 61.050 ;
        RECT 118.950 59.400 127.050 60.600 ;
        RECT 118.950 58.950 121.050 59.400 ;
        RECT 124.950 58.950 127.050 59.400 ;
        RECT 229.950 60.600 232.050 61.050 ;
        RECT 262.950 60.600 265.050 61.050 ;
        RECT 373.950 60.600 376.050 61.050 ;
        RECT 229.950 59.400 265.050 60.600 ;
        RECT 229.950 58.950 232.050 59.400 ;
        RECT 262.950 58.950 265.050 59.400 ;
        RECT 329.400 59.400 376.050 60.600 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 139.950 57.600 142.050 58.050 ;
        RECT 145.950 57.600 148.050 58.050 ;
        RECT 139.950 56.400 148.050 57.600 ;
        RECT 139.950 55.950 142.050 56.400 ;
        RECT 145.950 55.950 148.050 56.400 ;
        RECT 151.950 57.600 154.050 58.050 ;
        RECT 163.950 57.600 166.050 58.050 ;
        RECT 151.950 56.400 166.050 57.600 ;
        RECT 151.950 55.950 154.050 56.400 ;
        RECT 163.950 55.950 166.050 56.400 ;
        RECT 232.950 57.600 235.050 58.050 ;
        RECT 238.950 57.600 241.050 58.050 ;
        RECT 232.950 56.400 241.050 57.600 ;
        RECT 232.950 55.950 235.050 56.400 ;
        RECT 238.950 55.950 241.050 56.400 ;
        RECT 283.950 57.600 286.050 58.050 ;
        RECT 310.950 57.600 313.050 58.050 ;
        RECT 329.400 57.600 330.600 59.400 ;
        RECT 373.950 58.950 376.050 59.400 ;
        RECT 400.950 60.600 403.050 61.050 ;
        RECT 487.950 60.600 490.050 61.050 ;
        RECT 517.950 60.600 520.050 61.050 ;
        RECT 400.950 59.400 520.050 60.600 ;
        RECT 400.950 58.950 403.050 59.400 ;
        RECT 487.950 58.950 490.050 59.400 ;
        RECT 517.950 58.950 520.050 59.400 ;
        RECT 526.950 60.600 529.050 61.050 ;
        RECT 625.950 60.600 628.050 61.050 ;
        RECT 526.950 59.400 628.050 60.600 ;
        RECT 526.950 58.950 529.050 59.400 ;
        RECT 625.950 58.950 628.050 59.400 ;
        RECT 736.950 60.600 739.050 61.050 ;
        RECT 751.950 60.600 754.050 61.050 ;
        RECT 766.950 60.600 769.050 61.050 ;
        RECT 736.950 59.400 769.050 60.600 ;
        RECT 736.950 58.950 739.050 59.400 ;
        RECT 751.950 58.950 754.050 59.400 ;
        RECT 766.950 58.950 769.050 59.400 ;
        RECT 811.950 60.600 814.050 61.050 ;
        RECT 829.950 60.600 832.050 61.050 ;
        RECT 811.950 59.400 832.050 60.600 ;
        RECT 811.950 58.950 814.050 59.400 ;
        RECT 829.950 58.950 832.050 59.400 ;
        RECT 283.950 56.400 330.600 57.600 ;
        RECT 331.950 57.600 334.050 58.050 ;
        RECT 352.950 57.600 355.050 58.050 ;
        RECT 331.950 56.400 355.050 57.600 ;
        RECT 283.950 55.950 286.050 56.400 ;
        RECT 310.950 55.950 313.050 56.400 ;
        RECT 331.950 55.950 334.050 56.400 ;
        RECT 352.950 55.950 355.050 56.400 ;
        RECT 358.950 57.600 361.050 58.050 ;
        RECT 379.950 57.600 382.050 58.050 ;
        RECT 358.950 56.400 382.050 57.600 ;
        RECT 358.950 55.950 361.050 56.400 ;
        RECT 379.950 55.950 382.050 56.400 ;
        RECT 412.950 57.600 415.050 58.050 ;
        RECT 436.950 57.600 439.050 58.050 ;
        RECT 469.950 57.600 472.050 58.050 ;
        RECT 499.950 57.600 502.050 58.050 ;
        RECT 412.950 56.400 468.600 57.600 ;
        RECT 412.950 55.950 415.050 56.400 ;
        RECT 436.950 55.950 439.050 56.400 ;
        RECT 4.950 54.600 7.050 55.050 ;
        RECT 10.950 54.600 13.050 55.050 ;
        RECT 4.950 53.400 13.050 54.600 ;
        RECT 4.950 52.950 7.050 53.400 ;
        RECT 10.950 52.950 13.050 53.400 ;
        RECT 16.950 52.950 19.050 55.050 ;
        RECT 31.950 54.600 34.050 55.050 ;
        RECT 52.950 54.600 55.050 55.050 ;
        RECT 67.950 54.600 70.050 55.050 ;
        RECT 31.950 53.400 51.600 54.600 ;
        RECT 31.950 52.950 34.050 53.400 ;
        RECT 17.400 49.050 18.600 52.950 ;
        RECT 19.950 51.600 22.050 52.050 ;
        RECT 25.950 51.600 28.050 52.050 ;
        RECT 19.950 50.400 28.050 51.600 ;
        RECT 50.400 51.600 51.600 53.400 ;
        RECT 52.950 53.400 70.050 54.600 ;
        RECT 52.950 52.950 55.050 53.400 ;
        RECT 67.950 52.950 70.050 53.400 ;
        RECT 88.950 54.600 91.050 55.050 ;
        RECT 107.400 54.600 108.600 55.950 ;
        RECT 467.400 55.050 468.600 56.400 ;
        RECT 469.950 56.400 502.050 57.600 ;
        RECT 469.950 55.950 472.050 56.400 ;
        RECT 499.950 55.950 502.050 56.400 ;
        RECT 517.950 57.600 520.050 58.050 ;
        RECT 601.950 57.600 604.050 58.050 ;
        RECT 604.950 57.600 607.050 58.050 ;
        RECT 517.950 56.400 607.050 57.600 ;
        RECT 517.950 55.950 520.050 56.400 ;
        RECT 601.950 55.950 604.050 56.400 ;
        RECT 604.950 55.950 607.050 56.400 ;
        RECT 631.950 57.600 634.050 58.050 ;
        RECT 664.950 57.600 667.050 58.050 ;
        RECT 694.950 57.600 697.050 58.050 ;
        RECT 721.950 57.600 724.050 58.050 ;
        RECT 631.950 56.400 724.050 57.600 ;
        RECT 631.950 55.950 634.050 56.400 ;
        RECT 664.950 55.950 667.050 56.400 ;
        RECT 694.950 55.950 697.050 56.400 ;
        RECT 721.950 55.950 724.050 56.400 ;
        RECT 793.950 57.600 796.050 58.050 ;
        RECT 811.950 57.600 814.050 58.050 ;
        RECT 793.950 56.400 814.050 57.600 ;
        RECT 793.950 55.950 796.050 56.400 ;
        RECT 811.950 55.950 814.050 56.400 ;
        RECT 124.950 54.600 127.050 55.050 ;
        RECT 88.950 53.400 127.050 54.600 ;
        RECT 88.950 52.950 91.050 53.400 ;
        RECT 101.400 52.050 102.600 53.400 ;
        RECT 124.950 52.950 127.050 53.400 ;
        RECT 187.950 54.600 190.050 55.050 ;
        RECT 214.950 54.600 217.050 55.050 ;
        RECT 220.950 54.600 223.050 55.050 ;
        RECT 187.950 53.400 223.050 54.600 ;
        RECT 187.950 52.950 190.050 53.400 ;
        RECT 214.950 52.950 217.050 53.400 ;
        RECT 220.950 52.950 223.050 53.400 ;
        RECT 226.950 54.600 229.050 55.050 ;
        RECT 238.950 54.600 241.050 55.050 ;
        RECT 256.950 54.600 259.050 55.050 ;
        RECT 226.950 53.400 259.050 54.600 ;
        RECT 226.950 52.950 229.050 53.400 ;
        RECT 238.950 52.950 241.050 53.400 ;
        RECT 256.950 52.950 259.050 53.400 ;
        RECT 295.950 54.600 298.050 55.050 ;
        RECT 313.950 54.600 316.050 55.050 ;
        RECT 334.950 54.600 337.050 55.050 ;
        RECT 295.950 53.400 337.050 54.600 ;
        RECT 295.950 52.950 298.050 53.400 ;
        RECT 313.950 52.950 316.050 53.400 ;
        RECT 334.950 52.950 337.050 53.400 ;
        RECT 355.950 54.600 358.050 55.050 ;
        RECT 400.950 54.600 403.050 55.050 ;
        RECT 415.950 54.600 418.050 55.050 ;
        RECT 355.950 53.400 418.050 54.600 ;
        RECT 355.950 52.950 358.050 53.400 ;
        RECT 400.950 52.950 403.050 53.400 ;
        RECT 415.950 52.950 418.050 53.400 ;
        RECT 433.950 54.600 436.050 55.050 ;
        RECT 442.950 54.600 445.050 55.050 ;
        RECT 460.950 54.600 463.050 55.050 ;
        RECT 433.950 53.400 463.050 54.600 ;
        RECT 433.950 52.950 436.050 53.400 ;
        RECT 442.950 52.950 445.050 53.400 ;
        RECT 460.950 52.950 463.050 53.400 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 475.950 54.600 478.050 55.050 ;
        RECT 505.950 54.600 508.050 55.050 ;
        RECT 529.950 54.600 532.050 55.050 ;
        RECT 475.950 53.400 532.050 54.600 ;
        RECT 475.950 52.950 478.050 53.400 ;
        RECT 505.950 52.950 508.050 53.400 ;
        RECT 529.950 52.950 532.050 53.400 ;
        RECT 535.950 54.600 538.050 55.050 ;
        RECT 541.950 54.600 544.050 55.050 ;
        RECT 535.950 53.400 544.050 54.600 ;
        RECT 535.950 52.950 538.050 53.400 ;
        RECT 541.950 52.950 544.050 53.400 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 559.950 54.600 562.050 55.050 ;
        RECT 574.950 54.600 577.050 55.050 ;
        RECT 559.950 53.400 577.050 54.600 ;
        RECT 559.950 52.950 562.050 53.400 ;
        RECT 574.950 52.950 577.050 53.400 ;
        RECT 667.950 54.600 670.050 55.050 ;
        RECT 676.950 54.600 679.050 55.050 ;
        RECT 712.950 54.600 715.050 55.050 ;
        RECT 667.950 53.400 679.050 54.600 ;
        RECT 667.950 52.950 670.050 53.400 ;
        RECT 676.950 52.950 679.050 53.400 ;
        RECT 701.400 53.400 715.050 54.600 ;
        RECT 70.950 51.600 73.050 52.050 ;
        RECT 50.400 50.400 73.050 51.600 ;
        RECT 19.950 49.950 22.050 50.400 ;
        RECT 25.950 49.950 28.050 50.400 ;
        RECT 70.950 49.950 73.050 50.400 ;
        RECT 100.950 49.950 103.050 52.050 ;
        RECT 133.950 51.600 136.050 52.050 ;
        RECT 157.950 51.600 160.050 52.050 ;
        RECT 133.950 50.400 160.050 51.600 ;
        RECT 133.950 49.950 136.050 50.400 ;
        RECT 157.950 49.950 160.050 50.400 ;
        RECT 169.950 51.600 172.050 52.050 ;
        RECT 217.950 51.600 220.050 52.050 ;
        RECT 229.950 51.600 232.050 52.050 ;
        RECT 169.950 50.400 216.600 51.600 ;
        RECT 169.950 49.950 172.050 50.400 ;
        RECT 16.950 46.950 19.050 49.050 ;
        RECT 76.950 48.600 79.050 49.050 ;
        RECT 139.950 48.600 142.050 49.050 ;
        RECT 160.950 48.600 163.050 49.050 ;
        RECT 76.950 47.400 163.050 48.600 ;
        RECT 76.950 46.950 79.050 47.400 ;
        RECT 139.950 46.950 142.050 47.400 ;
        RECT 160.950 46.950 163.050 47.400 ;
        RECT 199.950 48.600 202.050 49.050 ;
        RECT 208.950 48.600 211.050 49.050 ;
        RECT 199.950 47.400 211.050 48.600 ;
        RECT 215.400 48.600 216.600 50.400 ;
        RECT 217.950 50.400 232.050 51.600 ;
        RECT 217.950 49.950 220.050 50.400 ;
        RECT 229.950 49.950 232.050 50.400 ;
        RECT 241.950 51.600 244.050 52.050 ;
        RECT 280.950 51.600 283.050 52.050 ;
        RECT 241.950 50.400 283.050 51.600 ;
        RECT 241.950 49.950 244.050 50.400 ;
        RECT 280.950 49.950 283.050 50.400 ;
        RECT 319.950 51.600 322.050 52.050 ;
        RECT 403.950 51.600 406.050 52.050 ;
        RECT 490.950 51.600 493.050 52.050 ;
        RECT 508.950 51.600 511.050 52.050 ;
        RECT 319.950 50.400 420.600 51.600 ;
        RECT 319.950 49.950 322.050 50.400 ;
        RECT 403.950 49.950 406.050 50.400 ;
        RECT 419.400 49.050 420.600 50.400 ;
        RECT 490.950 50.400 511.050 51.600 ;
        RECT 490.950 49.950 493.050 50.400 ;
        RECT 508.950 49.950 511.050 50.400 ;
        RECT 532.950 51.600 535.050 52.050 ;
        RECT 554.400 51.600 555.600 52.950 ;
        RECT 532.950 50.400 555.600 51.600 ;
        RECT 589.950 51.600 592.050 52.050 ;
        RECT 607.950 51.600 610.050 52.050 ;
        RECT 589.950 50.400 610.050 51.600 ;
        RECT 532.950 49.950 535.050 50.400 ;
        RECT 589.950 49.950 592.050 50.400 ;
        RECT 607.950 49.950 610.050 50.400 ;
        RECT 640.950 51.600 643.050 52.050 ;
        RECT 646.950 51.600 649.050 52.050 ;
        RECT 640.950 50.400 649.050 51.600 ;
        RECT 640.950 49.950 643.050 50.400 ;
        RECT 646.950 49.950 649.050 50.400 ;
        RECT 673.950 51.600 676.050 52.050 ;
        RECT 688.950 51.600 691.050 52.050 ;
        RECT 673.950 50.400 691.050 51.600 ;
        RECT 673.950 49.950 676.050 50.400 ;
        RECT 688.950 49.950 691.050 50.400 ;
        RECT 697.950 51.600 700.050 52.050 ;
        RECT 701.400 51.600 702.600 53.400 ;
        RECT 712.950 52.950 715.050 53.400 ;
        RECT 718.950 54.600 721.050 55.050 ;
        RECT 727.950 54.600 730.050 55.050 ;
        RECT 718.950 53.400 730.050 54.600 ;
        RECT 718.950 52.950 721.050 53.400 ;
        RECT 727.950 52.950 730.050 53.400 ;
        RECT 754.950 54.600 757.050 55.050 ;
        RECT 802.950 54.600 805.050 55.050 ;
        RECT 754.950 53.400 805.050 54.600 ;
        RECT 754.950 52.950 757.050 53.400 ;
        RECT 802.950 52.950 805.050 53.400 ;
        RECT 808.950 54.600 811.050 55.050 ;
        RECT 823.950 54.600 826.050 55.050 ;
        RECT 850.950 54.600 853.050 55.050 ;
        RECT 808.950 53.400 853.050 54.600 ;
        RECT 808.950 52.950 811.050 53.400 ;
        RECT 823.950 52.950 826.050 53.400 ;
        RECT 850.950 52.950 853.050 53.400 ;
        RECT 868.950 54.600 871.050 55.050 ;
        RECT 874.950 54.600 877.050 55.050 ;
        RECT 868.950 53.400 877.050 54.600 ;
        RECT 868.950 52.950 871.050 53.400 ;
        RECT 874.950 52.950 877.050 53.400 ;
        RECT 697.950 50.400 702.600 51.600 ;
        RECT 703.950 51.600 706.050 52.050 ;
        RECT 709.950 51.600 712.050 52.050 ;
        RECT 703.950 50.400 712.050 51.600 ;
        RECT 697.950 49.950 700.050 50.400 ;
        RECT 703.950 49.950 706.050 50.400 ;
        RECT 709.950 49.950 712.050 50.400 ;
        RECT 721.950 51.600 724.050 52.050 ;
        RECT 739.950 51.600 742.050 52.050 ;
        RECT 721.950 50.400 742.050 51.600 ;
        RECT 721.950 49.950 724.050 50.400 ;
        RECT 739.950 49.950 742.050 50.400 ;
        RECT 832.950 51.600 835.050 52.050 ;
        RECT 856.950 51.600 859.050 52.050 ;
        RECT 832.950 50.400 859.050 51.600 ;
        RECT 832.950 49.950 835.050 50.400 ;
        RECT 856.950 49.950 859.050 50.400 ;
        RECT 223.950 48.600 226.050 49.050 ;
        RECT 235.950 48.600 238.050 49.050 ;
        RECT 215.400 47.400 238.050 48.600 ;
        RECT 199.950 46.950 202.050 47.400 ;
        RECT 208.950 46.950 211.050 47.400 ;
        RECT 223.950 46.950 226.050 47.400 ;
        RECT 235.950 46.950 238.050 47.400 ;
        RECT 253.950 48.600 256.050 49.050 ;
        RECT 259.950 48.600 262.050 49.050 ;
        RECT 253.950 47.400 262.050 48.600 ;
        RECT 253.950 46.950 256.050 47.400 ;
        RECT 259.950 46.950 262.050 47.400 ;
        RECT 271.950 48.600 274.050 49.050 ;
        RECT 289.950 48.600 292.050 49.050 ;
        RECT 271.950 47.400 292.050 48.600 ;
        RECT 271.950 46.950 274.050 47.400 ;
        RECT 289.950 46.950 292.050 47.400 ;
        RECT 376.950 48.600 379.050 49.050 ;
        RECT 412.950 48.600 415.050 49.050 ;
        RECT 376.950 47.400 415.050 48.600 ;
        RECT 376.950 46.950 379.050 47.400 ;
        RECT 412.950 46.950 415.050 47.400 ;
        RECT 418.950 46.950 421.050 49.050 ;
        RECT 439.950 48.600 442.050 49.050 ;
        RECT 463.950 48.600 466.050 49.050 ;
        RECT 439.950 47.400 466.050 48.600 ;
        RECT 439.950 46.950 442.050 47.400 ;
        RECT 463.950 46.950 466.050 47.400 ;
        RECT 517.950 48.600 520.050 49.050 ;
        RECT 538.950 48.600 541.050 49.050 ;
        RECT 517.950 47.400 541.050 48.600 ;
        RECT 517.950 46.950 520.050 47.400 ;
        RECT 538.950 46.950 541.050 47.400 ;
        RECT 556.950 48.600 559.050 49.050 ;
        RECT 616.950 48.600 619.050 49.050 ;
        RECT 556.950 47.400 619.050 48.600 ;
        RECT 556.950 46.950 559.050 47.400 ;
        RECT 616.950 46.950 619.050 47.400 ;
        RECT 649.950 48.600 652.050 49.050 ;
        RECT 667.950 48.600 670.050 49.050 ;
        RECT 697.950 48.600 700.050 49.050 ;
        RECT 649.950 47.400 700.050 48.600 ;
        RECT 649.950 46.950 652.050 47.400 ;
        RECT 667.950 46.950 670.050 47.400 ;
        RECT 697.950 46.950 700.050 47.400 ;
        RECT 715.950 48.600 718.050 49.050 ;
        RECT 733.950 48.600 736.050 49.050 ;
        RECT 754.950 48.600 757.050 49.050 ;
        RECT 715.950 47.400 757.050 48.600 ;
        RECT 715.950 46.950 718.050 47.400 ;
        RECT 733.950 46.950 736.050 47.400 ;
        RECT 754.950 46.950 757.050 47.400 ;
        RECT 772.950 48.600 775.050 49.050 ;
        RECT 790.950 48.600 793.050 49.050 ;
        RECT 772.950 47.400 793.050 48.600 ;
        RECT 772.950 46.950 775.050 47.400 ;
        RECT 790.950 46.950 793.050 47.400 ;
        RECT 838.950 48.600 841.050 49.050 ;
        RECT 853.950 48.600 856.050 49.050 ;
        RECT 838.950 47.400 856.050 48.600 ;
        RECT 838.950 46.950 841.050 47.400 ;
        RECT 853.950 46.950 856.050 47.400 ;
        RECT 13.950 45.600 16.050 46.050 ;
        RECT 163.950 45.600 166.050 46.050 ;
        RECT 190.950 45.600 193.050 46.050 ;
        RECT 13.950 44.400 193.050 45.600 ;
        RECT 13.950 43.950 16.050 44.400 ;
        RECT 163.950 43.950 166.050 44.400 ;
        RECT 190.950 43.950 193.050 44.400 ;
        RECT 214.950 45.600 217.050 46.050 ;
        RECT 316.950 45.600 319.050 46.050 ;
        RECT 214.950 44.400 319.050 45.600 ;
        RECT 214.950 43.950 217.050 44.400 ;
        RECT 316.950 43.950 319.050 44.400 ;
        RECT 340.950 45.600 343.050 46.050 ;
        RECT 439.950 45.600 442.050 46.050 ;
        RECT 340.950 44.400 442.050 45.600 ;
        RECT 340.950 43.950 343.050 44.400 ;
        RECT 439.950 43.950 442.050 44.400 ;
        RECT 445.950 45.600 448.050 46.050 ;
        RECT 580.950 45.600 583.050 46.050 ;
        RECT 589.950 45.600 592.050 46.050 ;
        RECT 445.950 44.400 592.050 45.600 ;
        RECT 445.950 43.950 448.050 44.400 ;
        RECT 580.950 43.950 583.050 44.400 ;
        RECT 589.950 43.950 592.050 44.400 ;
        RECT 643.950 45.600 646.050 46.050 ;
        RECT 664.950 45.600 667.050 46.050 ;
        RECT 643.950 44.400 667.050 45.600 ;
        RECT 643.950 43.950 646.050 44.400 ;
        RECT 664.950 43.950 667.050 44.400 ;
        RECT 685.950 45.600 688.050 46.050 ;
        RECT 691.950 45.600 694.050 46.050 ;
        RECT 685.950 44.400 694.050 45.600 ;
        RECT 685.950 43.950 688.050 44.400 ;
        RECT 691.950 43.950 694.050 44.400 ;
        RECT 730.950 45.600 733.050 46.050 ;
        RECT 826.950 45.600 829.050 46.050 ;
        RECT 847.950 45.600 850.050 46.050 ;
        RECT 730.950 44.400 850.050 45.600 ;
        RECT 730.950 43.950 733.050 44.400 ;
        RECT 826.950 43.950 829.050 44.400 ;
        RECT 847.950 43.950 850.050 44.400 ;
        RECT 244.950 42.600 247.050 43.050 ;
        RECT 268.950 42.600 271.050 43.050 ;
        RECT 439.950 42.600 442.050 43.050 ;
        RECT 457.950 42.600 460.050 43.050 ;
        RECT 244.950 41.400 460.050 42.600 ;
        RECT 244.950 40.950 247.050 41.400 ;
        RECT 268.950 40.950 271.050 41.400 ;
        RECT 439.950 40.950 442.050 41.400 ;
        RECT 457.950 40.950 460.050 41.400 ;
        RECT 523.950 42.600 526.050 43.050 ;
        RECT 784.950 42.600 787.050 43.050 ;
        RECT 523.950 41.400 787.050 42.600 ;
        RECT 523.950 40.950 526.050 41.400 ;
        RECT 784.950 40.950 787.050 41.400 ;
        RECT 817.950 42.600 820.050 43.050 ;
        RECT 826.950 42.600 829.050 43.050 ;
        RECT 868.950 42.600 871.050 43.050 ;
        RECT 817.950 41.400 871.050 42.600 ;
        RECT 817.950 40.950 820.050 41.400 ;
        RECT 826.950 40.950 829.050 41.400 ;
        RECT 868.950 40.950 871.050 41.400 ;
        RECT 277.950 39.600 280.050 40.050 ;
        RECT 286.950 39.600 289.050 40.050 ;
        RECT 325.950 39.600 328.050 40.050 ;
        RECT 277.950 38.400 328.050 39.600 ;
        RECT 277.950 37.950 280.050 38.400 ;
        RECT 286.950 37.950 289.050 38.400 ;
        RECT 325.950 37.950 328.050 38.400 ;
        RECT 424.950 39.600 427.050 40.050 ;
        RECT 541.950 39.600 544.050 40.050 ;
        RECT 583.950 39.600 586.050 40.050 ;
        RECT 586.950 39.600 589.050 40.050 ;
        RECT 424.950 38.400 589.050 39.600 ;
        RECT 424.950 37.950 427.050 38.400 ;
        RECT 541.950 37.950 544.050 38.400 ;
        RECT 583.950 37.950 586.050 38.400 ;
        RECT 586.950 37.950 589.050 38.400 ;
        RECT 616.950 39.600 619.050 40.050 ;
        RECT 628.950 39.600 631.050 40.050 ;
        RECT 616.950 38.400 631.050 39.600 ;
        RECT 616.950 37.950 619.050 38.400 ;
        RECT 628.950 37.950 631.050 38.400 ;
        RECT 13.950 36.600 16.050 37.050 ;
        RECT 43.950 36.600 46.050 37.050 ;
        RECT 52.950 36.600 55.050 37.050 ;
        RECT 13.950 35.400 55.050 36.600 ;
        RECT 13.950 34.950 16.050 35.400 ;
        RECT 43.950 34.950 46.050 35.400 ;
        RECT 52.950 34.950 55.050 35.400 ;
        RECT 58.950 36.600 61.050 37.050 ;
        RECT 85.950 36.600 88.050 37.050 ;
        RECT 121.950 36.600 124.050 37.050 ;
        RECT 154.950 36.600 157.050 37.050 ;
        RECT 58.950 35.400 157.050 36.600 ;
        RECT 58.950 34.950 61.050 35.400 ;
        RECT 85.950 34.950 88.050 35.400 ;
        RECT 121.950 34.950 124.050 35.400 ;
        RECT 154.950 34.950 157.050 35.400 ;
        RECT 259.950 36.600 262.050 37.050 ;
        RECT 286.950 36.600 289.050 37.050 ;
        RECT 259.950 35.400 289.050 36.600 ;
        RECT 259.950 34.950 262.050 35.400 ;
        RECT 286.950 34.950 289.050 35.400 ;
        RECT 289.950 36.600 292.050 37.050 ;
        RECT 550.950 36.600 553.050 37.050 ;
        RECT 289.950 35.400 553.050 36.600 ;
        RECT 289.950 34.950 292.050 35.400 ;
        RECT 550.950 34.950 553.050 35.400 ;
        RECT 607.950 36.600 610.050 37.050 ;
        RECT 685.950 36.600 688.050 37.050 ;
        RECT 703.950 36.600 706.050 37.050 ;
        RECT 607.950 35.400 706.050 36.600 ;
        RECT 607.950 34.950 610.050 35.400 ;
        RECT 685.950 34.950 688.050 35.400 ;
        RECT 703.950 34.950 706.050 35.400 ;
        RECT 49.950 33.600 52.050 34.050 ;
        RECT 73.950 33.600 76.050 34.050 ;
        RECT 118.950 33.600 121.050 34.050 ;
        RECT 49.950 32.400 121.050 33.600 ;
        RECT 49.950 31.950 52.050 32.400 ;
        RECT 73.950 31.950 76.050 32.400 ;
        RECT 118.950 31.950 121.050 32.400 ;
        RECT 127.950 33.600 130.050 34.050 ;
        RECT 145.950 33.600 148.050 34.050 ;
        RECT 160.950 33.600 163.050 34.050 ;
        RECT 127.950 32.400 163.050 33.600 ;
        RECT 127.950 31.950 130.050 32.400 ;
        RECT 145.950 31.950 148.050 32.400 ;
        RECT 160.950 31.950 163.050 32.400 ;
        RECT 205.950 33.600 208.050 34.050 ;
        RECT 412.950 33.600 415.050 34.050 ;
        RECT 205.950 32.400 415.050 33.600 ;
        RECT 205.950 31.950 208.050 32.400 ;
        RECT 412.950 31.950 415.050 32.400 ;
        RECT 415.950 33.600 418.050 34.050 ;
        RECT 472.950 33.600 475.050 34.050 ;
        RECT 415.950 32.400 475.050 33.600 ;
        RECT 415.950 31.950 418.050 32.400 ;
        RECT 472.950 31.950 475.050 32.400 ;
        RECT 502.950 33.600 505.050 34.050 ;
        RECT 571.950 33.600 574.050 34.050 ;
        RECT 502.950 32.400 574.050 33.600 ;
        RECT 502.950 31.950 505.050 32.400 ;
        RECT 571.950 31.950 574.050 32.400 ;
        RECT 613.950 33.600 616.050 34.050 ;
        RECT 622.950 33.600 625.050 34.050 ;
        RECT 613.950 32.400 625.050 33.600 ;
        RECT 613.950 31.950 616.050 32.400 ;
        RECT 622.950 31.950 625.050 32.400 ;
        RECT 796.950 33.600 799.050 34.050 ;
        RECT 868.950 33.600 871.050 34.050 ;
        RECT 796.950 32.400 871.050 33.600 ;
        RECT 796.950 31.950 799.050 32.400 ;
        RECT 868.950 31.950 871.050 32.400 ;
        RECT 67.950 30.600 70.050 31.050 ;
        RECT 124.950 30.600 127.050 31.050 ;
        RECT 184.950 30.600 187.050 31.050 ;
        RECT 217.950 30.600 220.050 31.050 ;
        RECT 67.950 29.400 187.050 30.600 ;
        RECT 67.950 28.950 70.050 29.400 ;
        RECT 124.950 28.950 127.050 29.400 ;
        RECT 184.950 28.950 187.050 29.400 ;
        RECT 188.400 29.400 220.050 30.600 ;
        RECT 136.950 27.600 139.050 28.050 ;
        RECT 166.950 27.600 169.050 28.050 ;
        RECT 136.950 26.400 169.050 27.600 ;
        RECT 136.950 25.950 139.050 26.400 ;
        RECT 166.950 25.950 169.050 26.400 ;
        RECT 175.950 27.600 178.050 28.050 ;
        RECT 188.400 27.600 189.600 29.400 ;
        RECT 217.950 28.950 220.050 29.400 ;
        RECT 232.950 30.600 235.050 31.050 ;
        RECT 379.950 30.600 382.050 31.050 ;
        RECT 394.950 30.600 397.050 31.050 ;
        RECT 430.950 30.600 433.050 31.050 ;
        RECT 232.950 29.400 433.050 30.600 ;
        RECT 232.950 28.950 235.050 29.400 ;
        RECT 379.950 28.950 382.050 29.400 ;
        RECT 394.950 28.950 397.050 29.400 ;
        RECT 430.950 28.950 433.050 29.400 ;
        RECT 436.950 30.600 439.050 31.050 ;
        RECT 454.950 30.600 457.050 31.050 ;
        RECT 436.950 29.400 457.050 30.600 ;
        RECT 436.950 28.950 439.050 29.400 ;
        RECT 454.950 28.950 457.050 29.400 ;
        RECT 457.950 30.600 460.050 31.050 ;
        RECT 505.950 30.600 508.050 31.050 ;
        RECT 520.950 30.600 523.050 31.050 ;
        RECT 676.950 30.600 679.050 31.050 ;
        RECT 457.950 29.400 523.050 30.600 ;
        RECT 457.950 28.950 460.050 29.400 ;
        RECT 505.950 28.950 508.050 29.400 ;
        RECT 520.950 28.950 523.050 29.400 ;
        RECT 545.400 29.400 679.050 30.600 ;
        RECT 175.950 26.400 189.600 27.600 ;
        RECT 175.950 25.950 178.050 26.400 ;
        RECT 193.950 25.950 196.050 28.050 ;
        RECT 208.950 27.600 211.050 28.050 ;
        RECT 283.950 27.600 286.050 28.050 ;
        RECT 289.950 27.600 292.050 28.050 ;
        RECT 376.950 27.600 379.050 28.050 ;
        RECT 475.950 27.600 478.050 28.050 ;
        RECT 496.950 27.600 499.050 28.050 ;
        RECT 208.950 26.400 282.600 27.600 ;
        RECT 208.950 25.950 211.050 26.400 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 79.950 24.600 82.050 25.050 ;
        RECT 94.950 24.600 97.050 25.050 ;
        RECT 79.950 23.400 97.050 24.600 ;
        RECT 79.950 22.950 82.050 23.400 ;
        RECT 94.950 22.950 97.050 23.400 ;
        RECT 100.950 24.600 103.050 25.050 ;
        RECT 142.950 24.600 145.050 25.050 ;
        RECT 172.950 24.600 175.050 25.050 ;
        RECT 100.950 23.400 141.600 24.600 ;
        RECT 100.950 22.950 103.050 23.400 ;
        RECT 20.400 21.600 21.600 22.950 ;
        RECT 31.950 21.600 34.050 22.050 ;
        RECT 46.950 21.600 49.050 22.050 ;
        RECT 20.400 20.400 49.050 21.600 ;
        RECT 31.950 19.950 34.050 20.400 ;
        RECT 46.950 19.950 49.050 20.400 ;
        RECT 55.950 21.600 58.050 22.050 ;
        RECT 67.950 21.600 70.050 22.050 ;
        RECT 55.950 20.400 70.050 21.600 ;
        RECT 55.950 19.950 58.050 20.400 ;
        RECT 67.950 19.950 70.050 20.400 ;
        RECT 76.950 21.600 79.050 22.050 ;
        RECT 85.950 21.600 88.050 22.050 ;
        RECT 76.950 20.400 88.050 21.600 ;
        RECT 76.950 19.950 79.050 20.400 ;
        RECT 85.950 19.950 88.050 20.400 ;
        RECT 103.950 21.600 106.050 22.050 ;
        RECT 115.950 21.600 118.050 22.050 ;
        RECT 103.950 20.400 118.050 21.600 ;
        RECT 140.400 21.600 141.600 23.400 ;
        RECT 142.950 23.400 171.600 24.600 ;
        RECT 142.950 22.950 145.050 23.400 ;
        RECT 170.400 22.050 171.600 23.400 ;
        RECT 172.950 23.400 192.600 24.600 ;
        RECT 172.950 22.950 175.050 23.400 ;
        RECT 191.400 22.050 192.600 23.400 ;
        RECT 166.950 21.600 169.050 22.050 ;
        RECT 140.400 20.400 169.050 21.600 ;
        RECT 103.950 19.950 106.050 20.400 ;
        RECT 115.950 19.950 118.050 20.400 ;
        RECT 166.950 19.950 169.050 20.400 ;
        RECT 169.950 19.950 172.050 22.050 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 97.950 18.600 100.050 19.050 ;
        RECT 106.950 18.600 109.050 19.050 ;
        RECT 97.950 17.400 109.050 18.600 ;
        RECT 97.950 16.950 100.050 17.400 ;
        RECT 106.950 16.950 109.050 17.400 ;
        RECT 127.950 18.600 130.050 19.050 ;
        RECT 136.950 18.600 139.050 19.050 ;
        RECT 142.950 18.600 145.050 19.050 ;
        RECT 127.950 17.400 145.050 18.600 ;
        RECT 127.950 16.950 130.050 17.400 ;
        RECT 136.950 16.950 139.050 17.400 ;
        RECT 142.950 16.950 145.050 17.400 ;
        RECT 148.950 18.600 151.050 19.050 ;
        RECT 194.400 18.600 195.600 25.950 ;
        RECT 217.950 24.600 220.050 25.050 ;
        RECT 281.400 24.600 282.600 26.400 ;
        RECT 283.950 26.400 292.050 27.600 ;
        RECT 283.950 25.950 286.050 26.400 ;
        RECT 289.950 25.950 292.050 26.400 ;
        RECT 344.400 26.400 499.050 27.600 ;
        RECT 344.400 24.600 345.600 26.400 ;
        RECT 376.950 25.950 379.050 26.400 ;
        RECT 475.950 25.950 478.050 26.400 ;
        RECT 496.950 25.950 499.050 26.400 ;
        RECT 514.950 27.600 517.050 28.050 ;
        RECT 541.950 27.600 544.050 28.050 ;
        RECT 514.950 26.400 544.050 27.600 ;
        RECT 514.950 25.950 517.050 26.400 ;
        RECT 541.950 25.950 544.050 26.400 ;
        RECT 217.950 23.400 234.600 24.600 ;
        RECT 281.400 23.400 345.600 24.600 ;
        RECT 217.950 22.950 220.050 23.400 ;
        RECT 196.950 21.600 199.050 22.050 ;
        RECT 205.950 21.600 208.050 22.050 ;
        RECT 196.950 20.400 208.050 21.600 ;
        RECT 196.950 19.950 199.050 20.400 ;
        RECT 205.950 19.950 208.050 20.400 ;
        RECT 229.950 19.950 232.050 22.050 ;
        RECT 211.950 18.600 214.050 19.050 ;
        RECT 230.400 18.600 231.600 19.950 ;
        RECT 233.400 19.050 234.600 23.400 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 352.950 24.600 355.050 25.050 ;
        RECT 388.950 24.600 391.050 25.050 ;
        RECT 352.950 23.400 391.050 24.600 ;
        RECT 352.950 22.950 355.050 23.400 ;
        RECT 388.950 22.950 391.050 23.400 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 400.950 24.600 403.050 25.050 ;
        RECT 418.950 24.600 421.050 25.050 ;
        RECT 448.950 24.600 451.050 25.050 ;
        RECT 400.950 23.400 451.050 24.600 ;
        RECT 400.950 22.950 403.050 23.400 ;
        RECT 418.950 22.950 421.050 23.400 ;
        RECT 448.950 22.950 451.050 23.400 ;
        RECT 472.950 24.600 475.050 25.050 ;
        RECT 502.950 24.600 505.050 25.050 ;
        RECT 517.950 24.600 520.050 25.050 ;
        RECT 472.950 23.400 501.600 24.600 ;
        RECT 472.950 22.950 475.050 23.400 ;
        RECT 253.950 21.600 256.050 22.050 ;
        RECT 271.950 21.600 274.050 22.050 ;
        RECT 253.950 20.400 274.050 21.600 ;
        RECT 253.950 19.950 256.050 20.400 ;
        RECT 271.950 19.950 274.050 20.400 ;
        RECT 286.950 21.600 289.050 22.050 ;
        RECT 301.950 21.600 304.050 22.050 ;
        RECT 322.950 21.600 325.050 22.050 ;
        RECT 286.950 20.400 291.600 21.600 ;
        RECT 286.950 19.950 289.050 20.400 ;
        RECT 148.950 17.400 231.600 18.600 ;
        RECT 148.950 16.950 151.050 17.400 ;
        RECT 211.950 16.950 214.050 17.400 ;
        RECT 232.950 16.950 235.050 19.050 ;
        RECT 238.950 18.600 241.050 19.050 ;
        RECT 247.950 18.600 250.050 19.050 ;
        RECT 238.950 17.400 250.050 18.600 ;
        RECT 238.950 16.950 241.050 17.400 ;
        RECT 247.950 16.950 250.050 17.400 ;
        RECT 262.950 18.600 265.050 19.050 ;
        RECT 286.950 18.600 289.050 19.050 ;
        RECT 262.950 17.400 289.050 18.600 ;
        RECT 290.400 18.600 291.600 20.400 ;
        RECT 301.950 20.400 325.050 21.600 ;
        RECT 301.950 19.950 304.050 20.400 ;
        RECT 322.950 19.950 325.050 20.400 ;
        RECT 331.950 21.600 334.050 22.050 ;
        RECT 347.400 21.600 348.600 22.950 ;
        RECT 331.950 20.400 348.600 21.600 ;
        RECT 355.950 21.600 358.050 22.050 ;
        RECT 361.950 21.600 364.050 22.050 ;
        RECT 355.950 20.400 364.050 21.600 ;
        RECT 331.950 19.950 334.050 20.400 ;
        RECT 355.950 19.950 358.050 20.400 ;
        RECT 361.950 19.950 364.050 20.400 ;
        RECT 373.950 21.600 376.050 22.050 ;
        RECT 392.400 21.600 393.600 22.950 ;
        RECT 500.400 22.050 501.600 23.400 ;
        RECT 502.950 23.400 520.050 24.600 ;
        RECT 502.950 22.950 505.050 23.400 ;
        RECT 517.950 22.950 520.050 23.400 ;
        RECT 545.400 22.050 546.600 29.400 ;
        RECT 676.950 28.950 679.050 29.400 ;
        RECT 763.950 30.600 766.050 31.050 ;
        RECT 769.950 30.600 772.050 31.050 ;
        RECT 847.950 30.600 850.050 31.050 ;
        RECT 763.950 29.400 850.050 30.600 ;
        RECT 763.950 28.950 766.050 29.400 ;
        RECT 769.950 28.950 772.050 29.400 ;
        RECT 847.950 28.950 850.050 29.400 ;
        RECT 586.950 27.600 589.050 28.050 ;
        RECT 652.950 27.600 655.050 28.050 ;
        RECT 661.950 27.600 664.050 28.050 ;
        RECT 586.950 26.400 664.050 27.600 ;
        RECT 586.950 25.950 589.050 26.400 ;
        RECT 652.950 25.950 655.050 26.400 ;
        RECT 661.950 25.950 664.050 26.400 ;
        RECT 745.950 27.600 748.050 28.050 ;
        RECT 763.950 27.600 766.050 28.050 ;
        RECT 814.950 27.600 817.050 28.050 ;
        RECT 871.950 27.600 874.050 28.050 ;
        RECT 745.950 26.400 766.050 27.600 ;
        RECT 745.950 25.950 748.050 26.400 ;
        RECT 763.950 25.950 766.050 26.400 ;
        RECT 770.400 26.400 817.050 27.600 ;
        RECT 547.950 24.600 550.050 25.050 ;
        RECT 553.950 24.600 556.050 25.050 ;
        RECT 565.950 24.600 568.050 25.050 ;
        RECT 547.950 23.400 556.050 24.600 ;
        RECT 547.950 22.950 550.050 23.400 ;
        RECT 553.950 22.950 556.050 23.400 ;
        RECT 557.400 23.400 568.050 24.600 ;
        RECT 433.950 21.600 436.050 22.050 ;
        RECT 373.950 20.400 436.050 21.600 ;
        RECT 373.950 19.950 376.050 20.400 ;
        RECT 433.950 19.950 436.050 20.400 ;
        RECT 460.950 21.600 463.050 22.050 ;
        RECT 493.950 21.600 496.050 22.050 ;
        RECT 460.950 20.400 496.050 21.600 ;
        RECT 460.950 19.950 463.050 20.400 ;
        RECT 493.950 19.950 496.050 20.400 ;
        RECT 499.950 19.950 502.050 22.050 ;
        RECT 544.950 19.950 547.050 22.050 ;
        RECT 550.950 21.600 553.050 22.050 ;
        RECT 557.400 21.600 558.600 23.400 ;
        RECT 565.950 22.950 568.050 23.400 ;
        RECT 628.950 24.600 631.050 25.050 ;
        RECT 640.950 24.600 643.050 25.050 ;
        RECT 667.950 24.600 670.050 25.050 ;
        RECT 628.950 23.400 670.050 24.600 ;
        RECT 628.950 22.950 631.050 23.400 ;
        RECT 640.950 22.950 643.050 23.400 ;
        RECT 667.950 22.950 670.050 23.400 ;
        RECT 709.950 24.600 712.050 25.050 ;
        RECT 770.400 24.600 771.600 26.400 ;
        RECT 814.950 25.950 817.050 26.400 ;
        RECT 869.400 26.400 874.050 27.600 ;
        RECT 709.950 23.400 771.600 24.600 ;
        RECT 820.950 24.600 823.050 25.050 ;
        RECT 841.950 24.600 844.050 25.050 ;
        RECT 820.950 23.400 844.050 24.600 ;
        RECT 709.950 22.950 712.050 23.400 ;
        RECT 820.950 22.950 823.050 23.400 ;
        RECT 841.950 22.950 844.050 23.400 ;
        RECT 859.950 24.600 862.050 25.050 ;
        RECT 869.400 24.600 870.600 26.400 ;
        RECT 871.950 25.950 874.050 26.400 ;
        RECT 859.950 23.400 870.600 24.600 ;
        RECT 871.950 24.600 874.050 25.050 ;
        RECT 877.950 24.600 880.050 25.050 ;
        RECT 871.950 23.400 880.050 24.600 ;
        RECT 859.950 22.950 862.050 23.400 ;
        RECT 871.950 22.950 874.050 23.400 ;
        RECT 877.950 22.950 880.050 23.400 ;
        RECT 550.950 20.400 558.600 21.600 ;
        RECT 568.950 21.600 571.050 22.050 ;
        RECT 580.950 21.600 583.050 22.050 ;
        RECT 568.950 20.400 583.050 21.600 ;
        RECT 550.950 19.950 553.050 20.400 ;
        RECT 568.950 19.950 571.050 20.400 ;
        RECT 580.950 19.950 583.050 20.400 ;
        RECT 607.950 21.600 610.050 22.050 ;
        RECT 625.950 21.600 628.050 22.050 ;
        RECT 607.950 20.400 628.050 21.600 ;
        RECT 607.950 19.950 610.050 20.400 ;
        RECT 625.950 19.950 628.050 20.400 ;
        RECT 676.950 21.600 679.050 22.050 ;
        RECT 682.950 21.600 685.050 22.050 ;
        RECT 706.950 21.600 709.050 22.050 ;
        RECT 676.950 20.400 709.050 21.600 ;
        RECT 676.950 19.950 679.050 20.400 ;
        RECT 682.950 19.950 685.050 20.400 ;
        RECT 706.950 19.950 709.050 20.400 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 751.950 21.600 754.050 22.050 ;
        RECT 796.950 21.600 799.050 22.050 ;
        RECT 751.950 20.400 799.050 21.600 ;
        RECT 751.950 19.950 754.050 20.400 ;
        RECT 796.950 19.950 799.050 20.400 ;
        RECT 817.950 21.600 820.050 22.050 ;
        RECT 832.950 21.600 835.050 22.050 ;
        RECT 817.950 20.400 835.050 21.600 ;
        RECT 817.950 19.950 820.050 20.400 ;
        RECT 832.950 19.950 835.050 20.400 ;
        RECT 862.950 21.600 865.050 22.050 ;
        RECT 877.950 21.600 880.050 22.050 ;
        RECT 862.950 20.400 880.050 21.600 ;
        RECT 862.950 19.950 865.050 20.400 ;
        RECT 877.950 19.950 880.050 20.400 ;
        RECT 370.950 18.600 373.050 19.050 ;
        RECT 290.400 17.400 373.050 18.600 ;
        RECT 262.950 16.950 265.050 17.400 ;
        RECT 286.950 16.950 289.050 17.400 ;
        RECT 370.950 16.950 373.050 17.400 ;
        RECT 433.950 18.600 436.050 19.050 ;
        RECT 553.950 18.600 556.050 19.050 ;
        RECT 433.950 17.400 556.050 18.600 ;
        RECT 433.950 16.950 436.050 17.400 ;
        RECT 553.950 16.950 556.050 17.400 ;
        RECT 574.950 18.600 577.050 19.050 ;
        RECT 607.950 18.600 610.050 19.050 ;
        RECT 574.950 17.400 610.050 18.600 ;
        RECT 574.950 16.950 577.050 17.400 ;
        RECT 607.950 16.950 610.050 17.400 ;
        RECT 658.950 18.600 661.050 19.050 ;
        RECT 688.950 18.600 691.050 19.050 ;
        RECT 658.950 17.400 691.050 18.600 ;
        RECT 658.950 16.950 661.050 17.400 ;
        RECT 688.950 16.950 691.050 17.400 ;
        RECT 694.950 18.600 697.050 19.050 ;
        RECT 713.400 18.600 714.600 19.950 ;
        RECT 694.950 17.400 714.600 18.600 ;
        RECT 781.950 18.600 784.050 19.050 ;
        RECT 787.950 18.600 790.050 19.050 ;
        RECT 793.950 18.600 796.050 19.050 ;
        RECT 781.950 17.400 796.050 18.600 ;
        RECT 694.950 16.950 697.050 17.400 ;
        RECT 781.950 16.950 784.050 17.400 ;
        RECT 787.950 16.950 790.050 17.400 ;
        RECT 793.950 16.950 796.050 17.400 ;
        RECT 799.950 18.600 802.050 19.050 ;
        RECT 823.950 18.600 826.050 19.050 ;
        RECT 838.950 18.600 841.050 19.050 ;
        RECT 799.950 17.400 841.050 18.600 ;
        RECT 799.950 16.950 802.050 17.400 ;
        RECT 823.950 16.950 826.050 17.400 ;
        RECT 838.950 16.950 841.050 17.400 ;
        RECT 871.950 18.600 874.050 19.050 ;
        RECT 880.950 18.600 883.050 19.050 ;
        RECT 871.950 17.400 883.050 18.600 ;
        RECT 871.950 16.950 874.050 17.400 ;
        RECT 880.950 16.950 883.050 17.400 ;
        RECT 184.950 15.600 187.050 16.050 ;
        RECT 262.950 15.600 265.050 16.050 ;
        RECT 184.950 14.400 265.050 15.600 ;
        RECT 184.950 13.950 187.050 14.400 ;
        RECT 262.950 13.950 265.050 14.400 ;
        RECT 265.950 15.600 268.050 16.050 ;
        RECT 349.950 15.600 352.050 16.050 ;
        RECT 265.950 14.400 352.050 15.600 ;
        RECT 265.950 13.950 268.050 14.400 ;
        RECT 349.950 13.950 352.050 14.400 ;
        RECT 484.950 15.600 487.050 16.050 ;
        RECT 520.950 15.600 523.050 16.050 ;
        RECT 484.950 14.400 523.050 15.600 ;
        RECT 484.950 13.950 487.050 14.400 ;
        RECT 520.950 13.950 523.050 14.400 ;
        RECT 868.950 15.600 871.050 16.050 ;
        RECT 874.950 15.600 877.050 16.050 ;
        RECT 868.950 14.400 877.050 15.600 ;
        RECT 868.950 13.950 871.050 14.400 ;
        RECT 874.950 13.950 877.050 14.400 ;
        RECT 151.950 12.600 154.050 13.050 ;
        RECT 280.950 12.600 283.050 13.050 ;
        RECT 151.950 11.400 283.050 12.600 ;
        RECT 151.950 10.950 154.050 11.400 ;
        RECT 280.950 10.950 283.050 11.400 ;
        RECT 388.950 12.600 391.050 13.050 ;
        RECT 742.950 12.600 745.050 13.050 ;
        RECT 388.950 11.400 745.050 12.600 ;
        RECT 388.950 10.950 391.050 11.400 ;
        RECT 742.950 10.950 745.050 11.400 ;
  END
END cordic_element
END LIBRARY

