* NGSPICE file created from output_terminal.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

.subckt output_terminal gnd vdd Dout[11] Dout[10] Dout[9] Dout[8] Dout[7] Dout[6]
+ Dout[5] Dout[4] Dout[3] Dout[2] Dout[1] Dout[0] ISin Rdy Vld Xin[1] Xin[0] Yin[1]
+ Yin[0] clk selSign selXY
XFILL_5__370_ vdd gnd FILL
XFILL_7__317_ vdd gnd FILL
XFILL_2__288_ vdd gnd FILL
XFILL_2__426_ vdd gnd FILL
XFILL_2__357_ vdd gnd FILL
X_501_ _625_/A _501_/B _501_/C _502_/C vdd gnd NAND3X1
XFILL_5__499_ vdd gnd FILL
X_432_ _432_/A _432_/B _433_/B vdd gnd NAND2X1
X_294_ _577_/Q _479_/A vdd gnd INVX1
X_363_ _590_/Q _591_/Q _367_/B vdd gnd NOR2X1
XFILL_9__615_ vdd gnd FILL
XFILL_6__404_ vdd gnd FILL
XFILL_0_CLKBUF1_insert6 vdd gnd FILL
XFILL_6__335_ vdd gnd FILL
XFILL_9__477_ vdd gnd FILL
XFILL_9__546_ vdd gnd FILL
XFILL_1__513_ vdd gnd FILL
XFILL_1__444_ vdd gnd FILL
XFILL_1__375_ vdd gnd FILL
XFILL_5__422_ vdd gnd FILL
XFILL_5__353_ vdd gnd FILL
XFILL_8__495_ vdd gnd FILL
XFILL_5__284_ vdd gnd FILL
XFILL_6_CLKBUF1_insert1 vdd gnd FILL
XFILL_0__462_ vdd gnd FILL
XFILL_7_BUFX2_insert7 vdd gnd FILL
XFILL_0__531_ vdd gnd FILL
XFILL_2__409_ vdd gnd FILL
XFILL_0__393_ vdd gnd FILL
XFILL_9__331_ vdd gnd FILL
X_415_ _415_/A _582_/Q _417_/B _419_/B vdd gnd NAND3X1
X_346_ _346_/A _346_/B _348_/B vdd gnd NAND2X1
X_277_ _286_/A _559_/Q _278_/C vdd gnd NAND2X1
XFILL_4__440_ vdd gnd FILL
XFILL_6__318_ vdd gnd FILL
XFILL_4__371_ vdd gnd FILL
XFILL_9__529_ vdd gnd FILL
XFILL_1__427_ vdd gnd FILL
XFILL_1__358_ vdd gnd FILL
XFILL_1__289_ vdd gnd FILL
XFILL_8__280_ vdd gnd FILL
XFILL_5__336_ vdd gnd FILL
XFILL_5__405_ vdd gnd FILL
XFILL_8__616_ vdd gnd FILL
XFILL_8__478_ vdd gnd FILL
XFILL_8__547_ vdd gnd FILL
XFILL_0__514_ vdd gnd FILL
XFILL_0__445_ vdd gnd FILL
XFILL_0__376_ vdd gnd FILL
X_329_ _554_/A _542_/B _329_/C _603_/D vdd gnd OAI21X1
XFILL_4__423_ vdd gnd FILL
XFILL_4__354_ vdd gnd FILL
XFILL_4__285_ vdd gnd FILL
XFILL_7__496_ vdd gnd FILL
XFILL74250x39750 vdd gnd FILL
XFILL_8__401_ vdd gnd FILL
XFILL_8__332_ vdd gnd FILL
XFILL_3__510_ vdd gnd FILL
XFILL_3__441_ vdd gnd FILL
XFILL_5__319_ vdd gnd FILL
XFILL_3__372_ vdd gnd FILL
XFILL_0__428_ vdd gnd FILL
XFILL_0__359_ vdd gnd FILL
XFILL_7__281_ vdd gnd FILL
XFILL_7__350_ vdd gnd FILL
XFILL_4__337_ vdd gnd FILL
XFILL_4__406_ vdd gnd FILL
XFILL_2__390_ vdd gnd FILL
XFILL_7__617_ vdd gnd FILL
XFILL_7__548_ vdd gnd FILL
XFILL_7__479_ vdd gnd FILL
XFILL_8__315_ vdd gnd FILL
X_594_ _594_/D _605_/CLK _594_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert16 vdd gnd FILL
XFILL_3__424_ vdd gnd FILL
XFILL_3__286_ vdd gnd FILL
XFILL_3__355_ vdd gnd FILL
XFILL_6__497_ vdd gnd FILL
XFILL75750x46950 vdd gnd FILL
XFILL_7__402_ vdd gnd FILL
XFILL_7__333_ vdd gnd FILL
XFILL_2__511_ vdd gnd FILL
XFILL_2__442_ vdd gnd FILL
XFILL_2__373_ vdd gnd FILL
XFILL_6__420_ vdd gnd FILL
XFILL_6__282_ vdd gnd FILL
XFILL_6__351_ vdd gnd FILL
XFILL_9__493_ vdd gnd FILL
X_577_ _577_/D _581_/CLK _577_/Q vdd gnd DFFPOSX1
XFILL_1__460_ vdd gnd FILL
XFILL_3__407_ vdd gnd FILL
XFILL_1__391_ vdd gnd FILL
XFILL_3__338_ vdd gnd FILL
XFILL_6__618_ vdd gnd FILL
XFILL_1_CLKBUF1_insert0 vdd gnd FILL
XFILL_6__549_ vdd gnd FILL
XFILL_2_BUFX2_insert25 vdd gnd FILL
XFILL_2_BUFX2_insert14 vdd gnd FILL
XFILL_7__316_ vdd gnd FILL
XFILL_2__425_ vdd gnd FILL
X_500_ _548_/A _510_/C _501_/C vdd gnd NAND2X1
XFILL_2__287_ vdd gnd FILL
XFILL_2__356_ vdd gnd FILL
XFILL_5__498_ vdd gnd FILL
X_362_ _410_/B _362_/B _362_/C _561_/D vdd gnd OAI21X1
X_431_ _431_/A _431_/B _431_/C _432_/B vdd gnd NAND3X1
X_293_ _308_/A _472_/A _293_/C _621_/A vdd gnd OAI21X1
XFILL_6__403_ vdd gnd FILL
XFILL_9_BUFX2_insert20 vdd gnd FILL
XFILL_6__334_ vdd gnd FILL
XFILL_1__512_ vdd gnd FILL
XFILL_9__545_ vdd gnd FILL
XFILL_1__443_ vdd gnd FILL
XFILL_1__374_ vdd gnd FILL
XFILL_5__283_ vdd gnd FILL
XFILL_5__421_ vdd gnd FILL
XFILL_5__352_ vdd gnd FILL
XFILL_8__494_ vdd gnd FILL
XFILL_6_CLKBUF1_insert2 vdd gnd FILL
XFILL_7_BUFX2_insert8 vdd gnd FILL
XFILL_0__461_ vdd gnd FILL
XFILL_2__408_ vdd gnd FILL
XFILL_0__530_ vdd gnd FILL
XFILL_0__392_ vdd gnd FILL
XFILL_5__619_ vdd gnd FILL
XFILL_2__339_ vdd gnd FILL
XFILL_9__330_ vdd gnd FILL
X_414_ _414_/A _414_/B _414_/C _417_/B vdd gnd NAND3X1
X_345_ _490_/A _544_/B _546_/B _346_/B vdd gnd OAI21X1
X_276_ _571_/Q _440_/A vdd gnd INVX1
XFILL_4__370_ vdd gnd FILL
XFILL_6__317_ vdd gnd FILL
XFILL_9__459_ vdd gnd FILL
XFILL_1__288_ vdd gnd FILL
XFILL_1__426_ vdd gnd FILL
XFILL_1__357_ vdd gnd FILL
XFILL_4__499_ vdd gnd FILL
XFILL_5__404_ vdd gnd FILL
XFILL_8__615_ vdd gnd FILL
XFILL_5__335_ vdd gnd FILL
XFILL_8__477_ vdd gnd FILL
XFILL_8__546_ vdd gnd FILL
XFILL_0__513_ vdd gnd FILL
XFILL_0__444_ vdd gnd FILL
XFILL_0__375_ vdd gnd FILL
XFILL_9__313_ vdd gnd FILL
X_328_ _607_/D _541_/B _603_/Q _329_/C vdd gnd OAI21X1
XFILL_4__422_ vdd gnd FILL
XFILL_4__353_ vdd gnd FILL
XFILL_7__495_ vdd gnd FILL
XFILL_4__284_ vdd gnd FILL
XFILL_1__409_ vdd gnd FILL
XFILL_8__400_ vdd gnd FILL
XFILL_8__331_ vdd gnd FILL
XFILL_3__440_ vdd gnd FILL
XFILL_3__371_ vdd gnd FILL
XFILL_5__318_ vdd gnd FILL
XFILL_8__529_ vdd gnd FILL
XFILL_0__427_ vdd gnd FILL
XFILL_0__358_ vdd gnd FILL
XFILL_0__289_ vdd gnd FILL
XFILL_7__280_ vdd gnd FILL
XFILL_4__336_ vdd gnd FILL
XFILL_4__405_ vdd gnd FILL
XFILL_7__616_ vdd gnd FILL
XFILL_7__478_ vdd gnd FILL
XFILL_7__547_ vdd gnd FILL
XFILL_8__314_ vdd gnd FILL
XFILL_3__423_ vdd gnd FILL
X_593_ _593_/D _595_/CLK _593_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert17 vdd gnd FILL
XFILL_3__354_ vdd gnd FILL
XFILL_3__285_ vdd gnd FILL
XFILL_6__496_ vdd gnd FILL
XFILL_7__401_ vdd gnd FILL
XFILL_7__332_ vdd gnd FILL
XFILL_2__510_ vdd gnd FILL
XFILL_2__441_ vdd gnd FILL
XFILL_4__319_ vdd gnd FILL
XFILL_2__372_ vdd gnd FILL
XFILL_6__281_ vdd gnd FILL
XFILL_6__350_ vdd gnd FILL
XFILL_9__492_ vdd gnd FILL
X_576_ _576_/D _601_/CLK _576_/Q vdd gnd DFFPOSX1
XFILL_3__337_ vdd gnd FILL
XFILL_3__406_ vdd gnd FILL
XFILL_1_CLKBUF1_insert1 vdd gnd FILL
XFILL_1__390_ vdd gnd FILL
XFILL_6__479_ vdd gnd FILL
XFILL_6__617_ vdd gnd FILL
XFILL_6__548_ vdd gnd FILL
XFILL_2_BUFX2_insert15 vdd gnd FILL
XFILL_7__315_ vdd gnd FILL
XFILL_2__424_ vdd gnd FILL
XFILL_2__286_ vdd gnd FILL
XFILL_2__355_ vdd gnd FILL
XFILL_5__497_ vdd gnd FILL
X_292_ _305_/A _564_/Q _293_/C vdd gnd NAND2X1
X_361_ _561_/Q _503_/B _362_/C vdd gnd NAND2X1
X_430_ _584_/Q _585_/Q _430_/C _431_/A vdd gnd OAI21X1
XFILL_6__402_ vdd gnd FILL
XFILL_6__333_ vdd gnd FILL
XFILL_9__613_ vdd gnd FILL
XFILL_9_BUFX2_insert21 vdd gnd FILL
XFILL_9__544_ vdd gnd FILL
XFILL_1__511_ vdd gnd FILL
XFILL_9__475_ vdd gnd FILL
XFILL_1__442_ vdd gnd FILL
XFILL_1__373_ vdd gnd FILL
X_559_ _559_/D _573_/CLK _559_/Q vdd gnd DFFPOSX1
XFILL_5__420_ vdd gnd FILL
XFILL_5__282_ vdd gnd FILL
XFILL_5__351_ vdd gnd FILL
XFILL_8__493_ vdd gnd FILL
XFILL_7_BUFX2_insert9 vdd gnd FILL
XFILL_6_CLKBUF1_insert3 vdd gnd FILL
XFILL_2__338_ vdd gnd FILL
XFILL_0__460_ vdd gnd FILL
XFILL_2__407_ vdd gnd FILL
XFILL_0__391_ vdd gnd FILL
XFILL_5__618_ vdd gnd FILL
XFILL_5__549_ vdd gnd FILL
X_413_ _584_/Q _585_/Q _414_/A vdd gnd NOR2X1
X_275_ _286_/A _436_/B _275_/C _613_/A vdd gnd OAI21X1
X_344_ _593_/Q _546_/B vdd gnd INVX1
XFILL_6__316_ vdd gnd FILL
XFILL_9__527_ vdd gnd FILL
XFILL_9__458_ vdd gnd FILL
XFILL_1__425_ vdd gnd FILL
XFILL_1__287_ vdd gnd FILL
XFILL_1__356_ vdd gnd FILL
XFILL_4__498_ vdd gnd FILL
XFILL_5__403_ vdd gnd FILL
XFILL_8__614_ vdd gnd FILL
XFILL_8__545_ vdd gnd FILL
XFILL_5__334_ vdd gnd FILL
XFILL_0__512_ vdd gnd FILL
XFILL_8__476_ vdd gnd FILL
XFILL_0__443_ vdd gnd FILL
XFILL_9__312_ vdd gnd FILL
XFILL_0__374_ vdd gnd FILL
X_327_ _556_/A _542_/B _327_/C _602_/D vdd gnd OAI21X1
XFILL_4__283_ vdd gnd FILL
XFILL_4__421_ vdd gnd FILL
XFILL_4__352_ vdd gnd FILL
XFILL_7__494_ vdd gnd FILL
XFILL_1__408_ vdd gnd FILL
XFILL_4__619_ vdd gnd FILL
XFILL_1__339_ vdd gnd FILL
XFILL_8__330_ vdd gnd FILL
XFILL_5__317_ vdd gnd FILL
XFILL_3__370_ vdd gnd FILL
XFILL_8__528_ vdd gnd FILL
XFILL_8__459_ vdd gnd FILL
XFILL_0__288_ vdd gnd FILL
XFILL_0__426_ vdd gnd FILL
XFILL_0__357_ vdd gnd FILL
XFILL_3__499_ vdd gnd FILL
XFILL_4__404_ vdd gnd FILL
XFILL_7__615_ vdd gnd FILL
XFILL_4__335_ vdd gnd FILL
XFILL_7__477_ vdd gnd FILL
XFILL_7__546_ vdd gnd FILL
XFILL_8__313_ vdd gnd FILL
XFILL_6_BUFX2_insert18 vdd gnd FILL
X_592_ _592_/D _595_/CLK _592_/Q vdd gnd DFFPOSX1
XFILL_3__284_ vdd gnd FILL
XFILL_3__422_ vdd gnd FILL
XFILL_3__353_ vdd gnd FILL
XFILL_6__495_ vdd gnd FILL
XFILL_0__409_ vdd gnd FILL
XFILL_7__400_ vdd gnd FILL
XFILL_7__331_ vdd gnd FILL
XFILL_2__440_ vdd gnd FILL
XFILL_2__371_ vdd gnd FILL
XFILL_4__318_ vdd gnd FILL
XFILL_7__529_ vdd gnd FILL
XFILL_6__280_ vdd gnd FILL
X_575_ _575_/D _581_/CLK _575_/Q vdd gnd DFFPOSX1
XFILL_6__616_ vdd gnd FILL
XFILL_3__336_ vdd gnd FILL
XFILL_3__405_ vdd gnd FILL
XFILL_1_CLKBUF1_insert2 vdd gnd FILL
XFILL75450x28950 vdd gnd FILL
XFILL_6__478_ vdd gnd FILL
XFILL_6__547_ vdd gnd FILL
XFILL_2_BUFX2_insert16 vdd gnd FILL
XFILL_7__314_ vdd gnd FILL
XFILL_2__423_ vdd gnd FILL
XFILL_2__354_ vdd gnd FILL
XFILL_5__496_ vdd gnd FILL
XFILL_2__285_ vdd gnd FILL
X_291_ _576_/Q _472_/A vdd gnd INVX1
X_360_ _360_/A _360_/B _362_/B vdd gnd NAND2X1
XFILL_9_BUFX2_insert11 vdd gnd FILL
XFILL_6__401_ vdd gnd FILL
XFILL_6__332_ vdd gnd FILL
XFILL_9__474_ vdd gnd FILL
XFILL_1__510_ vdd gnd FILL
XFILL_1__441_ vdd gnd FILL
X_558_ _558_/D _573_/CLK _558_/Q vdd gnd DFFPOSX1
X_489_ _597_/Q _492_/B vdd gnd INVX1
XFILL_3__319_ vdd gnd FILL
XFILL_1__372_ vdd gnd FILL
XFILL_5__350_ vdd gnd FILL
XFILL_5__281_ vdd gnd FILL
XFILL_8__492_ vdd gnd FILL
XFILL_6_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__337_ vdd gnd FILL
XFILL_2__406_ vdd gnd FILL
XFILL_0__390_ vdd gnd FILL
XFILL_5__479_ vdd gnd FILL
XFILL_5__617_ vdd gnd FILL
XFILL_5__548_ vdd gnd FILL
X_412_ _412_/A _412_/B _414_/C vdd gnd AND2X2
X_274_ _558_/Q _301_/A _275_/C vdd gnd NAND2X1
X_343_ _415_/A _592_/Q _593_/Q _346_/A vdd gnd NAND3X1
XFILL_6__315_ vdd gnd FILL
XFILL_9__526_ vdd gnd FILL
XFILL_5_BUFX2_insert20 vdd gnd FILL
XFILL_1__424_ vdd gnd FILL
XFILL_1__355_ vdd gnd FILL
XFILL_9__388_ vdd gnd FILL
XFILL_1__286_ vdd gnd FILL
XFILL_4__497_ vdd gnd FILL
XFILL_5__402_ vdd gnd FILL
XFILL_5__333_ vdd gnd FILL
XFILL_8__613_ vdd gnd FILL
XFILL_8__544_ vdd gnd FILL
XFILL_0__511_ vdd gnd FILL
XFILL_8__475_ vdd gnd FILL
XFILL_0__442_ vdd gnd FILL
XFILL_9__311_ vdd gnd FILL
XFILL_0__373_ vdd gnd FILL
X_326_ _607_/D _541_/B _602_/Q _327_/C vdd gnd OAI21X1
XFILL_4__420_ vdd gnd FILL
XFILL75150x25350 vdd gnd FILL
XFILL75750x72150 vdd gnd FILL
XFILL_4__282_ vdd gnd FILL
XFILL_4__351_ vdd gnd FILL
XFILL_7__493_ vdd gnd FILL
XFILL_1__338_ vdd gnd FILL
XFILL_1__407_ vdd gnd FILL
XFILL_4__618_ vdd gnd FILL
XFILL_4__549_ vdd gnd FILL
XFILL_5__316_ vdd gnd FILL
XFILL_8__458_ vdd gnd FILL
XFILL_8__527_ vdd gnd FILL
XFILL_0__425_ vdd gnd FILL
XFILL_8__389_ vdd gnd FILL
XFILL_0__287_ vdd gnd FILL
XFILL_0__356_ vdd gnd FILL
XFILL_3__498_ vdd gnd FILL
X_309_ Yin[1] _554_/A vdd gnd INVX1
XFILL_4__403_ vdd gnd FILL
XFILL_4__334_ vdd gnd FILL
XFILL_7__614_ vdd gnd FILL
XFILL_7__545_ vdd gnd FILL
XFILL_7__476_ vdd gnd FILL
XFILL_8__312_ vdd gnd FILL
XFILL_6_BUFX2_insert19 vdd gnd FILL
XFILL_3__421_ vdd gnd FILL
X_591_ _591_/D _606_/CLK _591_/Q vdd gnd DFFPOSX1
XFILL_3__283_ vdd gnd FILL
XFILL_3__352_ vdd gnd FILL
XFILL_6__494_ vdd gnd FILL
XFILL_0__408_ vdd gnd FILL
XFILL_0__339_ vdd gnd FILL
XFILL_3__619_ vdd gnd FILL
XFILL_7__330_ vdd gnd FILL
XFILL_4__317_ vdd gnd FILL
XFILL_2__370_ vdd gnd FILL
XFILL_7__528_ vdd gnd FILL
XFILL_7__459_ vdd gnd FILL
XFILL_9__490_ vdd gnd FILL
XFILL_2__499_ vdd gnd FILL
XFILL_3__404_ vdd gnd FILL
X_574_ _574_/D _581_/CLK _574_/Q vdd gnd DFFPOSX1
XFILL_6__615_ vdd gnd FILL
XFILL_1_CLKBUF1_insert3 vdd gnd FILL
XFILL_3__335_ vdd gnd FILL
XFILL_6__477_ vdd gnd FILL
XFILL_6__546_ vdd gnd FILL
XFILL_2_BUFX2_insert17 vdd gnd FILL
XFILL_7__313_ vdd gnd FILL
XFILL_2__284_ vdd gnd FILL
XFILL_2__422_ vdd gnd FILL
XFILL_2__353_ vdd gnd FILL
XFILL_5__495_ vdd gnd FILL
X_290_ _308_/A _464_/A _290_/C _620_/A vdd gnd OAI21X1
XFILL_6__400_ vdd gnd FILL
XFILL_9_BUFX2_insert12 vdd gnd FILL
XFILL_9_BUFX2_insert23 vdd gnd FILL
XFILL_6__331_ vdd gnd FILL
XFILL_9__473_ vdd gnd FILL
XFILL_9__542_ vdd gnd FILL
X_488_ _493_/B _488_/B _488_/C _578_/D vdd gnd OAI21X1
X_557_ _557_/D _601_/CLK _557_/Q vdd gnd DFFPOSX1
XFILL_4_BUFX2_insert7 vdd gnd FILL
XFILL_1__440_ vdd gnd FILL
XFILL_1__371_ vdd gnd FILL
XFILL_3__318_ vdd gnd FILL
XFILL_6__529_ vdd gnd FILL
XFILL_5__280_ vdd gnd FILL
XFILL_8__491_ vdd gnd FILL
XFILL_6_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__405_ vdd gnd FILL
XFILL_5__616_ vdd gnd FILL
XFILL_2__336_ vdd gnd FILL
XFILL_5__478_ vdd gnd FILL
XFILL_5__547_ vdd gnd FILL
X_411_ _568_/Q _420_/A vdd gnd INVX1
X_342_ _544_/B _378_/A _342_/C _558_/D vdd gnd OAI21X1
X_273_ _570_/Q _436_/B vdd gnd INVX1
XFILL_6__314_ vdd gnd FILL
XFILL_9__456_ vdd gnd FILL
XFILL_9__387_ vdd gnd FILL
X_609_ _609_/D _612_/CLK _610_/D vdd gnd DFFPOSX1
XFILL_9__525_ vdd gnd FILL
XFILL_5_BUFX2_insert10 vdd gnd FILL
XFILL_1__285_ vdd gnd FILL
XFILL_5_BUFX2_insert21 vdd gnd FILL
XFILL_1__423_ vdd gnd FILL
XFILL_1__354_ vdd gnd FILL
XFILL_4__496_ vdd gnd FILL
XFILL_5__401_ vdd gnd FILL
XFILL_5__332_ vdd gnd FILL
XFILL_8__474_ vdd gnd FILL
XFILL_8__543_ vdd gnd FILL
XFILL_0__510_ vdd gnd FILL
XFILL_0__441_ vdd gnd FILL
XFILL_0__372_ vdd gnd FILL
XFILL_2__319_ vdd gnd FILL
X_325_ _541_/B _607_/D _542_/B vdd gnd OR2X2
XFILL_4__350_ vdd gnd FILL
XFILL_9__508_ vdd gnd FILL
XFILL_4__281_ vdd gnd FILL
XFILL_7__492_ vdd gnd FILL
XFILL_9__439_ vdd gnd FILL
XFILL_1__337_ vdd gnd FILL
XFILL_1__406_ vdd gnd FILL
XFILL74550x28950 vdd gnd FILL
XFILL_4__479_ vdd gnd FILL
XFILL_4__617_ vdd gnd FILL
XFILL_4__548_ vdd gnd FILL
XFILL_5__315_ vdd gnd FILL
XFILL_8__457_ vdd gnd FILL
XFILL_8__526_ vdd gnd FILL
XFILL_8__388_ vdd gnd FILL
XFILL_0__424_ vdd gnd FILL
XFILL_0__355_ vdd gnd FILL
XFILL_0__286_ vdd gnd FILL
XFILL_3__497_ vdd gnd FILL
X_308_ _308_/A _308_/B _308_/C _616_/A vdd gnd OAI21X1
XFILL_4__402_ vdd gnd FILL
XFILL_4__333_ vdd gnd FILL
XFILL_7__475_ vdd gnd FILL
XFILL_7__613_ vdd gnd FILL
XFILL_7__544_ vdd gnd FILL
XFILL_8__311_ vdd gnd FILL
XFILL_3__420_ vdd gnd FILL
XFILL_3__351_ vdd gnd FILL
X_590_ _590_/D _606_/CLK _590_/Q vdd gnd DFFPOSX1
XFILL_3__282_ vdd gnd FILL
XFILL_6__493_ vdd gnd FILL
XFILL_8__509_ vdd gnd FILL
XFILL_0__338_ vdd gnd FILL
XFILL_0__407_ vdd gnd FILL
XFILL_3__618_ vdd gnd FILL
XFILL_3__549_ vdd gnd FILL
XFILL_4__316_ vdd gnd FILL
XFILL_7__458_ vdd gnd FILL
XFILL_7__527_ vdd gnd FILL
XFILL_7__389_ vdd gnd FILL
XFILL_2__498_ vdd gnd FILL
XFILL_3__403_ vdd gnd FILL
X_573_ _573_/D _573_/CLK _573_/Q vdd gnd DFFPOSX1
XFILL_3__334_ vdd gnd FILL
XFILL_6__614_ vdd gnd FILL
XFILL_6__545_ vdd gnd FILL
XFILL_1_CLKBUF1_insert4 vdd gnd FILL
XFILL_2_BUFX2_insert18 vdd gnd FILL
XFILL_6__476_ vdd gnd FILL
XFILL_7__312_ vdd gnd FILL
XFILL_2__421_ vdd gnd FILL
XFILL74250x25350 vdd gnd FILL
XFILL74850x72150 vdd gnd FILL
XFILL_2__283_ vdd gnd FILL
XFILL_2__352_ vdd gnd FILL
XFILL_5__494_ vdd gnd FILL
XFILL_2__619_ vdd gnd FILL
XFILL_9_BUFX2_insert24 vdd gnd FILL
XFILL_9_BUFX2_insert13 vdd gnd FILL
XFILL_9__541_ vdd gnd FILL
XFILL_6__330_ vdd gnd FILL
X_625_ _625_/A Vld vdd gnd BUFX2
X_487_ _578_/Q _493_/B _488_/C vdd gnd NAND2X1
XFILL_4_BUFX2_insert8 vdd gnd FILL
X_556_ _556_/A _556_/B _556_/C _598_/D vdd gnd OAI21X1
XFILL_3__317_ vdd gnd FILL
XFILL_1__370_ vdd gnd FILL
XFILL75750x57750 vdd gnd FILL
XFILL_6__459_ vdd gnd FILL
XFILL_6__528_ vdd gnd FILL
XFILL_8__490_ vdd gnd FILL
XFILL_1__499_ vdd gnd FILL
XFILL_6_CLKBUF1_insert6 vdd gnd FILL
XFILL_2__404_ vdd gnd FILL
XFILL_5__615_ vdd gnd FILL
XFILL_5__546_ vdd gnd FILL
XFILL_2__335_ vdd gnd FILL
XFILL_5__477_ vdd gnd FILL
X_410_ _410_/A _410_/B _410_/C _410_/D _567_/D vdd gnd AOI22X1
X_341_ _558_/Q _421_/B _342_/C vdd gnd NAND2X1
XFILL_6__313_ vdd gnd FILL
XFILL_9__455_ vdd gnd FILL
XFILL_9__386_ vdd gnd FILL
XFILL_1__422_ vdd gnd FILL
X_608_ _608_/D _612_/CLK _609_/D vdd gnd DFFPOSX1
XFILL_5_BUFX2_insert11 vdd gnd FILL
XFILL_1__284_ vdd gnd FILL
XFILL_5_BUFX2_insert22 vdd gnd FILL
XFILL_1__353_ vdd gnd FILL
X_539_ _607_/D _541_/B _590_/Q _540_/C vdd gnd OAI21X1
XFILL_4__495_ vdd gnd FILL
XFILL_5__400_ vdd gnd FILL
XFILL_5__331_ vdd gnd FILL
XFILL_8__473_ vdd gnd FILL
XFILL_8__542_ vdd gnd FILL
XFILL_2__318_ vdd gnd FILL
XFILL_0__440_ vdd gnd FILL
XFILL_0__371_ vdd gnd FILL
XFILL_5__529_ vdd gnd FILL
X_324_ _608_/D _541_/B vdd gnd INVX2
XFILL_4__280_ vdd gnd FILL
XFILL_7__491_ vdd gnd FILL
XFILL_9__507_ vdd gnd FILL
XFILL_1__405_ vdd gnd FILL
XFILL_9__369_ vdd gnd FILL
XFILL_4__616_ vdd gnd FILL
XFILL_1__336_ vdd gnd FILL
XFILL_4__478_ vdd gnd FILL
XFILL_1_BUFX2_insert20 vdd gnd FILL
XFILL_4__547_ vdd gnd FILL
XFILL_5__314_ vdd gnd FILL
XFILL_8__525_ vdd gnd FILL
XFILL_8__456_ vdd gnd FILL
XFILL_8__387_ vdd gnd FILL
XFILL_0__285_ vdd gnd FILL
XFILL_0__423_ vdd gnd FILL
XFILL_0__354_ vdd gnd FILL
XFILL_3__496_ vdd gnd FILL
X_307_ _308_/A _569_/Q _308_/C vdd gnd NAND2X1
XFILL75450x54150 vdd gnd FILL
XFILL_4__401_ vdd gnd FILL
XFILL_4__332_ vdd gnd FILL
XFILL_7__474_ vdd gnd FILL
XFILL_7__543_ vdd gnd FILL
XFILL_1__319_ vdd gnd FILL
XFILL_8__310_ vdd gnd FILL
XFILL_3__350_ vdd gnd FILL
XFILL_6__492_ vdd gnd FILL
XFILL_8__508_ vdd gnd FILL
XFILL_3__281_ vdd gnd FILL
XFILL_8__439_ vdd gnd FILL
XFILL_0__337_ vdd gnd FILL
XFILL_3__617_ vdd gnd FILL
XFILL_0__406_ vdd gnd FILL
XFILL_3__479_ vdd gnd FILL
XFILL_3__548_ vdd gnd FILL
XFILL_4__315_ vdd gnd FILL
XFILL_7__457_ vdd gnd FILL
XFILL_7__526_ vdd gnd FILL
XFILL_7__388_ vdd gnd FILL
XFILL_2__497_ vdd gnd FILL
X_572_ _572_/D _573_/CLK _572_/Q vdd gnd DFFPOSX1
XFILL_3__402_ vdd gnd FILL
XFILL_3__333_ vdd gnd FILL
XFILL_6__475_ vdd gnd FILL
XFILL_6__613_ vdd gnd FILL
XFILL_1_CLKBUF1_insert5 vdd gnd FILL
XFILL_6__544_ vdd gnd FILL
XFILL_2_BUFX2_insert19 vdd gnd FILL
XFILL_7__311_ vdd gnd FILL
XFILL_2__420_ vdd gnd FILL
XFILL_2__351_ vdd gnd FILL
XFILL_2__282_ vdd gnd FILL
XFILL_5__493_ vdd gnd FILL
XFILL_7__509_ vdd gnd FILL
XFILL_7_CLKBUF1_insert0 vdd gnd FILL
XFILL73650x28950 vdd gnd FILL
XFILL_9__471_ vdd gnd FILL
XFILL_2__618_ vdd gnd FILL
XFILL_9_BUFX2_insert25 vdd gnd FILL
XFILL_2__549_ vdd gnd FILL
XFILL_9__540_ vdd gnd FILL
X_624_ _624_/A Dout[9] vdd gnd BUFX2
X_555_ _598_/Q _556_/B _556_/C vdd gnd NAND2X1
X_486_ _486_/A _486_/B _488_/B vdd gnd NAND2X1
XFILL_4_BUFX2_insert9 vdd gnd FILL
XFILL_3__316_ vdd gnd FILL
XFILL_6__458_ vdd gnd FILL
XFILL_6__527_ vdd gnd FILL
XFILL_6__389_ vdd gnd FILL
XFILL_1__498_ vdd gnd FILL
XFILL_2__403_ vdd gnd FILL
XFILL_2__334_ vdd gnd FILL
XFILL_5__476_ vdd gnd FILL
XFILL_5__614_ vdd gnd FILL
XFILL_5__545_ vdd gnd FILL
X_340_ _452_/B _340_/Y vdd gnd INVX8
XFILL_6__312_ vdd gnd FILL
XFILL_9__454_ vdd gnd FILL
XFILL_9__523_ vdd gnd FILL
XFILL_5_BUFX2_insert12 vdd gnd FILL
XFILL_5_BUFX2_insert23 vdd gnd FILL
X_538_ _538_/A _538_/B _538_/C _589_/D vdd gnd OAI21X1
X_607_ _607_/D _612_/CLK _608_/D vdd gnd DFFPOSX1
XFILL_1__421_ vdd gnd FILL
X_469_ _511_/C _469_/B _477_/C vdd gnd NAND2X1
XFILL_1__283_ vdd gnd FILL
XFILL_1__352_ vdd gnd FILL
XFILL_4__494_ vdd gnd FILL
XFILL_5__330_ vdd gnd FILL
XFILL_1__619_ vdd gnd FILL
XFILL_8__541_ vdd gnd FILL
XFILL_8__472_ vdd gnd FILL
XFILL_2__317_ vdd gnd FILL
XFILL_0__370_ vdd gnd FILL
XFILL_5__459_ vdd gnd FILL
XFILL_5__528_ vdd gnd FILL
X_323_ Yin[0] _556_/A vdd gnd INVX1
XFILL_7__490_ vdd gnd FILL
XFILL_0__499_ vdd gnd FILL
XFILL_9__437_ vdd gnd FILL
XFILL_1__404_ vdd gnd FILL
XFILL_9__368_ vdd gnd FILL
XFILL_1__335_ vdd gnd FILL
XFILL_4__615_ vdd gnd FILL
XFILL_4__546_ vdd gnd FILL
XFILL_4__477_ vdd gnd FILL
XFILL_1_BUFX2_insert10 vdd gnd FILL
XFILL_1_BUFX2_insert21 vdd gnd FILL
XFILL_5__313_ vdd gnd FILL
XFILL_8__524_ vdd gnd FILL
XFILL_8__455_ vdd gnd FILL
XFILL_8__386_ vdd gnd FILL
XFILL_0__422_ vdd gnd FILL
XFILL73950x72150 vdd gnd FILL
XFILL_0__284_ vdd gnd FILL
XFILL_0__353_ vdd gnd FILL
X_306_ _581_/Q _308_/B vdd gnd INVX1
XFILL_3__495_ vdd gnd FILL
XFILL_4__400_ vdd gnd FILL
XFILL_7__542_ vdd gnd FILL
XFILL_4__331_ vdd gnd FILL
XFILL_7__473_ vdd gnd FILL
XFILL74850x57750 vdd gnd FILL
XFILL_1__318_ vdd gnd FILL
XFILL_4__529_ vdd gnd FILL
XFILL_3__280_ vdd gnd FILL
XFILL_6__491_ vdd gnd FILL
XFILL_8__507_ vdd gnd FILL
XFILL_8__438_ vdd gnd FILL
XFILL_0__405_ vdd gnd FILL
XFILL_8__369_ vdd gnd FILL
XFILL_3__616_ vdd gnd FILL
XFILL_0__336_ vdd gnd FILL
XFILL_3__547_ vdd gnd FILL
XFILL_3__478_ vdd gnd FILL
XFILL_4__314_ vdd gnd FILL
XFILL_7__525_ vdd gnd FILL
XFILL_7__456_ vdd gnd FILL
XFILL_7__387_ vdd gnd FILL
XFILL_2__496_ vdd gnd FILL
X_571_ _571_/D _605_/CLK _571_/Q vdd gnd DFFPOSX1
XFILL_3__401_ vdd gnd FILL
XFILL_1_CLKBUF1_insert6 vdd gnd FILL
XFILL_3__332_ vdd gnd FILL
XFILL_6__474_ vdd gnd FILL
XFILL_6__543_ vdd gnd FILL
XFILL_0__319_ vdd gnd FILL
XFILL_7__310_ vdd gnd FILL
XFILL_2__281_ vdd gnd FILL
XFILL_2__350_ vdd gnd FILL
XFILL_5__492_ vdd gnd FILL
XFILL_7__508_ vdd gnd FILL
XFILL_7__439_ vdd gnd FILL
XFILL_7_CLKBUF1_insert1 vdd gnd FILL
XFILL_2__617_ vdd gnd FILL
XFILL_9_BUFX2_insert15 vdd gnd FILL
XFILL_2__479_ vdd gnd FILL
XFILL_9__470_ vdd gnd FILL
XFILL_2__548_ vdd gnd FILL
X_485_ _490_/B _512_/C _486_/A vdd gnd NAND2X1
X_623_ _623_/A Dout[8] vdd gnd BUFX2
X_554_ _554_/A _554_/B _554_/C _597_/D vdd gnd OAI21X1
XFILL_3__315_ vdd gnd FILL
XFILL_6__457_ vdd gnd FILL
XFILL_6__526_ vdd gnd FILL
XFILL_6__388_ vdd gnd FILL
XFILL_1__497_ vdd gnd FILL
XFILL_5__613_ vdd gnd FILL
XFILL_2__402_ vdd gnd FILL
XFILL_2__333_ vdd gnd FILL
XFILL_5__475_ vdd gnd FILL
XFILL_5__544_ vdd gnd FILL
XFILL_6__311_ vdd gnd FILL
XFILL_9__522_ vdd gnd FILL
XFILL_9__384_ vdd gnd FILL
X_468_ _598_/Q _473_/A vdd gnd INVX1
XFILL_5_BUFX2_insert24 vdd gnd FILL
XFILL75450x39750 vdd gnd FILL
XFILL_1__420_ vdd gnd FILL
X_606_ Rdy _606_/CLK _607_/D vdd gnd DFFPOSX1
X_537_ Xin[1] _538_/B _538_/C vdd gnd NAND2X1
XFILL_5_BUFX2_insert13 vdd gnd FILL
XFILL_1__351_ vdd gnd FILL
XFILL_4__493_ vdd gnd FILL
XFILL_6__509_ vdd gnd FILL
XFILL_1__282_ vdd gnd FILL
X_399_ _399_/A _399_/B _442_/C _431_/C vdd gnd OAI21X1
XFILL_1__618_ vdd gnd FILL
XFILL_8__471_ vdd gnd FILL
XFILL_1__549_ vdd gnd FILL
XFILL_8__540_ vdd gnd FILL
XFILL_2__316_ vdd gnd FILL
XFILL_5__458_ vdd gnd FILL
X_322_ _463_/B _538_/B _322_/C _601_/D vdd gnd OAI21X1
XFILL_5__527_ vdd gnd FILL
XFILL_5__389_ vdd gnd FILL
XFILL_0__498_ vdd gnd FILL
XFILL_9__436_ vdd gnd FILL
XBUFX2_insert7 selXY _286_/A vdd gnd BUFX2
XFILL_9__505_ vdd gnd FILL
XFILL_9__298_ vdd gnd FILL
XFILL_1__403_ vdd gnd FILL
XFILL_1__334_ vdd gnd FILL
XFILL_4__476_ vdd gnd FILL
XFILL_4__614_ vdd gnd FILL
XFILL_4__545_ vdd gnd FILL
XFILL_1_BUFX2_insert11 vdd gnd FILL
XFILL_1_BUFX2_insert22 vdd gnd FILL
XFILL_5__312_ vdd gnd FILL
XFILL_8__454_ vdd gnd FILL
XFILL_8__523_ vdd gnd FILL
XFILL_8__385_ vdd gnd FILL
XFILL_0__421_ vdd gnd FILL
XFILL_0__352_ vdd gnd FILL
XFILL_0__283_ vdd gnd FILL
X_305_ _305_/A _502_/A _305_/C _615_/A vdd gnd OAI21X1
XFILL_3__494_ vdd gnd FILL
XFILL_4__330_ vdd gnd FILL
XFILL_0__619_ vdd gnd FILL
XFILL_7__541_ vdd gnd FILL
XFILL_7__472_ vdd gnd FILL
XFILL_1__317_ vdd gnd FILL
XFILL_4__459_ vdd gnd FILL
XFILL_4__528_ vdd gnd FILL
XFILL_6__490_ vdd gnd FILL
XFILL_8__437_ vdd gnd FILL
XFILL_8__506_ vdd gnd FILL
XFILL_8__299_ vdd gnd FILL
XFILL_0__404_ vdd gnd FILL
XFILL_8__368_ vdd gnd FILL
XFILL_0__335_ vdd gnd FILL
XFILL_3__615_ vdd gnd FILL
XFILL_2_CLKBUF1_insert0 vdd gnd FILL
XFILL_3__546_ vdd gnd FILL
XFILL_3__477_ vdd gnd FILL
XFILL75150x36150 vdd gnd FILL
XFILL_4__313_ vdd gnd FILL
XFILL_7__455_ vdd gnd FILL
XFILL_7__524_ vdd gnd FILL
XFILL_7__386_ vdd gnd FILL
XFILL_2__495_ vdd gnd FILL
XFILL75150x7350 vdd gnd FILL
X_570_ _570_/D _605_/CLK _570_/Q vdd gnd DFFPOSX1
XFILL_3__400_ vdd gnd FILL
XFILL_3__331_ vdd gnd FILL
XFILL_6__542_ vdd gnd FILL
XFILL_6__473_ vdd gnd FILL
XFILL_0__318_ vdd gnd FILL
XFILL_3__529_ vdd gnd FILL
XFILL_2__280_ vdd gnd FILL
XFILL_5__491_ vdd gnd FILL
XFILL_1_BUFX2_insert7 vdd gnd FILL
XFILL_7__507_ vdd gnd FILL
XFILL_7__438_ vdd gnd FILL
XFILL_7_CLKBUF1_insert2 vdd gnd FILL
XFILL_7__369_ vdd gnd FILL
XFILL_2__616_ vdd gnd FILL
XFILL_2__547_ vdd gnd FILL
XFILL_9_BUFX2_insert16 vdd gnd FILL
XFILL_2__478_ vdd gnd FILL
X_622_ _622_/A Dout[7] vdd gnd BUFX2
X_484_ _512_/C _490_/B _486_/B vdd gnd OR2X2
X_553_ _597_/Q _554_/B _554_/C vdd gnd NAND2X1
XFILL_3__314_ vdd gnd FILL
XFILL_6__525_ vdd gnd FILL
XFILL_6__456_ vdd gnd FILL
XFILL_6__387_ vdd gnd FILL
XFILL_1__496_ vdd gnd FILL
XFILL_2__401_ vdd gnd FILL
XFILL_2__332_ vdd gnd FILL
XFILL_5__474_ vdd gnd FILL
XFILL_5__543_ vdd gnd FILL
XFILL73950x57750 vdd gnd FILL
XFILL_6__310_ vdd gnd FILL
XFILL_9__452_ vdd gnd FILL
X_605_ _605_/D _605_/CLK _605_/Q vdd gnd DFFPOSX1
XFILL_9__383_ vdd gnd FILL
X_467_ _511_/C _598_/Q _469_/B _471_/B vdd gnd NAND3X1
XFILL_5_BUFX2_insert25 vdd gnd FILL
XFILL_1__281_ vdd gnd FILL
X_536_ _536_/A _538_/B _536_/C _588_/D vdd gnd OAI21X1
X_398_ _412_/A _412_/B _399_/B vdd gnd NAND2X1
XFILL_5_BUFX2_insert14 vdd gnd FILL
XFILL_1__350_ vdd gnd FILL
XFILL_4__492_ vdd gnd FILL
XFILL_6__508_ vdd gnd FILL
XFILL_6__439_ vdd gnd FILL
XFILL_1__617_ vdd gnd FILL
XFILL_1__479_ vdd gnd FILL
XFILL_8__470_ vdd gnd FILL
XFILL_1__548_ vdd gnd FILL
XFILL_2__315_ vdd gnd FILL
XFILL_5__526_ vdd gnd FILL
XFILL_5__457_ vdd gnd FILL
X_321_ Yin[1] _538_/B _322_/C vdd gnd NAND2X1
XFILL_5__388_ vdd gnd FILL
XFILL_0__497_ vdd gnd FILL
XFILL_9__504_ vdd gnd FILL
XFILL_9__297_ vdd gnd FILL
XBUFX2_insert8 selXY _308_/A vdd gnd BUFX2
XFILL_9__435_ vdd gnd FILL
XFILL_1__402_ vdd gnd FILL
XFILL_9__366_ vdd gnd FILL
XFILL_4__613_ vdd gnd FILL
X_519_ _611_/D _519_/B _550_/B vdd gnd NOR2X1
XFILL_1__333_ vdd gnd FILL
XFILL_4__475_ vdd gnd FILL
XFILL_4__544_ vdd gnd FILL
XFILL_1_BUFX2_insert12 vdd gnd FILL
XFILL_1_BUFX2_insert23 vdd gnd FILL
XFILL_5__311_ vdd gnd FILL
XFILL_8__453_ vdd gnd FILL
XFILL_8__522_ vdd gnd FILL
XFILL_8__384_ vdd gnd FILL
XFILL_0__420_ vdd gnd FILL
XFILL_0__351_ vdd gnd FILL
XFILL_3__493_ vdd gnd FILL
XFILL_5__509_ vdd gnd FILL
XFILL_0__282_ vdd gnd FILL
X_304_ _308_/A _568_/Q _305_/C vdd gnd NAND2X1
XFILL_0__618_ vdd gnd FILL
XFILL_7__471_ vdd gnd FILL
XFILL_0__549_ vdd gnd FILL
XFILL_7__540_ vdd gnd FILL
XFILL_9__418_ vdd gnd FILL
XFILL_9__349_ vdd gnd FILL
XFILL_1__316_ vdd gnd FILL
XFILL_4__458_ vdd gnd FILL
XFILL_4__527_ vdd gnd FILL
XFILL_4__389_ vdd gnd FILL
XFILL_8__505_ vdd gnd FILL
XFILL_8__436_ vdd gnd FILL
XFILL_8__367_ vdd gnd FILL
XFILL_8__298_ vdd gnd FILL
XFILL_0__403_ vdd gnd FILL
XFILL_0__334_ vdd gnd FILL
XFILL_3__476_ vdd gnd FILL
XFILL_3__614_ vdd gnd FILL
XFILL_3__545_ vdd gnd FILL
XFILL_2_CLKBUF1_insert1 vdd gnd FILL
XCLKBUF1_insert0 clk _581_/CLK vdd gnd CLKBUF1
XFILL_4__312_ vdd gnd FILL
XFILL_7__454_ vdd gnd FILL
XFILL_7__523_ vdd gnd FILL
XFILL74550x39750 vdd gnd FILL
XFILL_7__385_ vdd gnd FILL
XFILL_2__494_ vdd gnd FILL
XFILL_3__330_ vdd gnd FILL
XFILL_6__472_ vdd gnd FILL
XFILL_6__541_ vdd gnd FILL
XFILL_8__419_ vdd gnd FILL
XFILL_0__317_ vdd gnd FILL
XFILL_3__459_ vdd gnd FILL
XFILL_3__528_ vdd gnd FILL
XFILL_1_BUFX2_insert8 vdd gnd FILL
XFILL_5__490_ vdd gnd FILL
XFILL_7__437_ vdd gnd FILL
XFILL_7__506_ vdd gnd FILL
XFILL_7__368_ vdd gnd FILL
XFILL_7__299_ vdd gnd FILL
XFILL_7_CLKBUF1_insert3 vdd gnd FILL
XFILL_2__615_ vdd gnd FILL
XFILL_2__477_ vdd gnd FILL
XFILL_2__546_ vdd gnd FILL
XFILL_9_BUFX2_insert17 vdd gnd FILL
X_621_ _621_/A Dout[6] vdd gnd BUFX2
X_483_ _483_/A _483_/B _509_/A _512_/C vdd gnd OAI21X1
X_552_ _556_/A _554_/B _552_/C _596_/D vdd gnd OAI21X1
XFILL_3__313_ vdd gnd FILL
XFILL_6__455_ vdd gnd FILL
XFILL_6__524_ vdd gnd FILL
XFILL_6__386_ vdd gnd FILL
XFILL_1__495_ vdd gnd FILL
XFILL_2__400_ vdd gnd FILL
XFILL_2__331_ vdd gnd FILL
XFILL_5__542_ vdd gnd FILL
XFILL_5__473_ vdd gnd FILL
XFILL_9__451_ vdd gnd FILL
XFILL_9__520_ vdd gnd FILL
XFILL_2__529_ vdd gnd FILL
X_604_ _604_/D _605_/CLK _604_/Q vdd gnd DFFPOSX1
X_535_ Xin[0] _538_/B _536_/C vdd gnd NAND2X1
X_466_ _494_/A _496_/B _469_/B vdd gnd NAND2X1
X_397_ _586_/Q _587_/Q _412_/B vdd gnd NOR2X1
XFILL_5_BUFX2_insert15 vdd gnd FILL
XFILL_1__280_ vdd gnd FILL
XFILL_4__491_ vdd gnd FILL
XFILL_6__507_ vdd gnd FILL
XFILL_6__438_ vdd gnd FILL
XFILL_6__369_ vdd gnd FILL
XFILL_1__616_ vdd gnd FILL
XFILL_1__547_ vdd gnd FILL
XFILL_1__478_ vdd gnd FILL
XFILL_2__314_ vdd gnd FILL
XFILL_5__525_ vdd gnd FILL
XFILL_5__456_ vdd gnd FILL
X_320_ _601_/Q _463_/B vdd gnd INVX1
XFILL_5__387_ vdd gnd FILL
XFILL_9__503_ vdd gnd FILL
XFILL_0__496_ vdd gnd FILL
XFILL_9__296_ vdd gnd FILL
XBUFX2_insert9 selXY _305_/A vdd gnd BUFX2
X_518_ _612_/D _525_/B _519_/B vdd gnd NAND2X1
XFILL_9__365_ vdd gnd FILL
XFILL_1__401_ vdd gnd FILL
X_449_ _603_/Q _450_/A _451_/B vdd gnd NAND2X1
XFILL_4__543_ vdd gnd FILL
XFILL_1__332_ vdd gnd FILL
XFILL_4__474_ vdd gnd FILL
XFILL_1_BUFX2_insert24 vdd gnd FILL
XFILL_1_BUFX2_insert13 vdd gnd FILL
XFILL_5__310_ vdd gnd FILL
XFILL_8__521_ vdd gnd FILL
XFILL_8__452_ vdd gnd FILL
XFILL_8__383_ vdd gnd FILL
XFILL_0__281_ vdd gnd FILL
XFILL_0__350_ vdd gnd FILL
XFILL_3__492_ vdd gnd FILL
XFILL_5__508_ vdd gnd FILL
XFILL_5__439_ vdd gnd FILL
X_303_ _580_/Q _502_/A vdd gnd INVX1
XFILL_0__617_ vdd gnd FILL
XFILL_0__548_ vdd gnd FILL
XFILL_0__479_ vdd gnd FILL
XFILL_7__470_ vdd gnd FILL
XFILL_9__417_ vdd gnd FILL
XFILL_1__315_ vdd gnd FILL
XFILL_9__279_ vdd gnd FILL
XFILL_4__526_ vdd gnd FILL
XFILL_4__457_ vdd gnd FILL
XFILL_4__388_ vdd gnd FILL
XFILL_8__504_ vdd gnd FILL
XFILL_8__297_ vdd gnd FILL
XFILL_8__435_ vdd gnd FILL
XFILL_0__402_ vdd gnd FILL
XFILL_8__366_ vdd gnd FILL
XFILL_3__613_ vdd gnd FILL
XFILL_0__333_ vdd gnd FILL
XFILL_3__475_ vdd gnd FILL
XFILL_2_CLKBUF1_insert2 vdd gnd FILL
XFILL_3__544_ vdd gnd FILL
XCLKBUF1_insert1 clk _606_/CLK vdd gnd CLKBUF1
XFILL_4__311_ vdd gnd FILL
XFILL_7__522_ vdd gnd FILL
XFILL_7__453_ vdd gnd FILL
XFILL_7__384_ vdd gnd FILL
XFILL_2__493_ vdd gnd FILL
XFILL_4__509_ vdd gnd FILL
XFILL_6__471_ vdd gnd FILL
XFILL_8__418_ vdd gnd FILL
XFILL_6__540_ vdd gnd FILL
XFILL_8__349_ vdd gnd FILL
XFILL_0__316_ vdd gnd FILL
XFILL_3__458_ vdd gnd FILL
XFILL_3__527_ vdd gnd FILL
XFILL_3__389_ vdd gnd FILL
XFILL_1_BUFX2_insert9 vdd gnd FILL
XFILL_7__505_ vdd gnd FILL
XFILL_7__298_ vdd gnd FILL
XFILL_7__436_ vdd gnd FILL
XFILL_7_CLKBUF1_insert4 vdd gnd FILL
XFILL_7__367_ vdd gnd FILL
XFILL_2__614_ vdd gnd FILL
XFILL_2__476_ vdd gnd FILL
XFILL_2__545_ vdd gnd FILL
X_620_ _620_/A Dout[5] vdd gnd BUFX2
X_551_ _596_/Q _554_/B _552_/C vdd gnd NAND2X1
X_482_ _494_/A _494_/B _483_/B vdd gnd NAND2X1
XFILL_3__312_ vdd gnd FILL
XFILL_6__454_ vdd gnd FILL
XFILL_6__385_ vdd gnd FILL
XFILL_6__523_ vdd gnd FILL
XFILL_1__494_ vdd gnd FILL
XFILL_2__330_ vdd gnd FILL
XFILL_5__472_ vdd gnd FILL
XFILL_5__541_ vdd gnd FILL
XFILL_7__419_ vdd gnd FILL
XFILL_2__459_ vdd gnd FILL
XFILL_9__450_ vdd gnd FILL
XFILL_2__528_ vdd gnd FILL
X_465_ _600_/Q _601_/Q _494_/A vdd gnd NOR2X1
XFILL_5_BUFX2_insert16 vdd gnd FILL
X_603_ _603_/D _606_/CLK _603_/Q vdd gnd DFFPOSX1
X_534_ _542_/A _556_/B _534_/C _587_/D vdd gnd OAI21X1
XFILL_9__381_ vdd gnd FILL
X_396_ _584_/Q _407_/B vdd gnd INVX1
XFILL_4__490_ vdd gnd FILL
XFILL_6__437_ vdd gnd FILL
XFILL_6__506_ vdd gnd FILL
XFILL_6__368_ vdd gnd FILL
XFILL_6__299_ vdd gnd FILL
XFILL_1__615_ vdd gnd FILL
XFILL_1__477_ vdd gnd FILL
XFILL_1__546_ vdd gnd FILL
XFILL_2__313_ vdd gnd FILL
XFILL_5__455_ vdd gnd FILL
XFILL_5__524_ vdd gnd FILL
XFILL_5__386_ vdd gnd FILL
XFILL75750x7350 vdd gnd FILL
XFILL_0__495_ vdd gnd FILL
XFILL_9__433_ vdd gnd FILL
XFILL_9__364_ vdd gnd FILL
X_448_ _490_/A _448_/B _448_/C _450_/A vdd gnd OAI21X1
X_517_ _517_/A _517_/B _525_/B vdd gnd AND2X2
XFILL_1__400_ vdd gnd FILL
XFILL_1__331_ vdd gnd FILL
X_379_ _588_/Q _589_/Q _412_/A vdd gnd NOR2X1
XFILL_4__542_ vdd gnd FILL
XFILL_4__473_ vdd gnd FILL
XFILL_1_BUFX2_insert25 vdd gnd FILL
XFILL_1_BUFX2_insert14 vdd gnd FILL
XFILL_8__451_ vdd gnd FILL
XFILL_8__520_ vdd gnd FILL
XFILL_1__529_ vdd gnd FILL
XFILL_8__382_ vdd gnd FILL
XFILL73050x10950 vdd gnd FILL
XFILL_0__280_ vdd gnd FILL
X_302_ _305_/A _493_/A _302_/C _624_/A vdd gnd OAI21X1
XFILL_3__491_ vdd gnd FILL
XFILL_9_BUFX2_insert8 vdd gnd FILL
XFILL_5__507_ vdd gnd FILL
XFILL_5__369_ vdd gnd FILL
XFILL_5__438_ vdd gnd FILL
XFILL_0__616_ vdd gnd FILL
XFILL_8_BUFX2_insert20 vdd gnd FILL
XFILL_0__547_ vdd gnd FILL
XFILL_0__478_ vdd gnd FILL
XFILL_9__347_ vdd gnd FILL
XFILL_1__314_ vdd gnd FILL
XFILL_9__278_ vdd gnd FILL
XFILL_4__456_ vdd gnd FILL
XFILL_4__525_ vdd gnd FILL
XFILL_4__387_ vdd gnd FILL
XFILL_8__503_ vdd gnd FILL
XFILL_8__434_ vdd gnd FILL
XFILL_8__296_ vdd gnd FILL
XFILL_8__365_ vdd gnd FILL
XFILL_0__401_ vdd gnd FILL
XFILL_0__332_ vdd gnd FILL
XFILL_3__543_ vdd gnd FILL
XFILL_3__474_ vdd gnd FILL
XFILL_2_CLKBUF1_insert3 vdd gnd FILL
XCLKBUF1_insert2 clk _601_/CLK vdd gnd CLKBUF1
XFILL_4__310_ vdd gnd FILL
XFILL_7__521_ vdd gnd FILL
XFILL_7__452_ vdd gnd FILL
XFILL_7__383_ vdd gnd FILL
XFILL_2__492_ vdd gnd FILL
XFILL_4__508_ vdd gnd FILL
XFILL_4__439_ vdd gnd FILL
XFILL_6__470_ vdd gnd FILL
XFILL_8__417_ vdd gnd FILL
XFILL_0__315_ vdd gnd FILL
XFILL_8__279_ vdd gnd FILL
XFILL_8__348_ vdd gnd FILL
XFILL_3__526_ vdd gnd FILL
XFILL_3__457_ vdd gnd FILL
XFILL_3__388_ vdd gnd FILL
XFILL_7__435_ vdd gnd FILL
XFILL_7__504_ vdd gnd FILL
XFILL_7__297_ vdd gnd FILL
XFILL_7__366_ vdd gnd FILL
XFILL_7_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__613_ vdd gnd FILL
XFILL_9_BUFX2_insert19 vdd gnd FILL
XFILL_2__475_ vdd gnd FILL
XFILL_2__544_ vdd gnd FILL
X_481_ _598_/Q _599_/Q _494_/B vdd gnd NOR2X1
X_550_ _550_/A _550_/B _550_/C _595_/D vdd gnd OAI21X1
XFILL_3__311_ vdd gnd FILL
XFILL_6__522_ vdd gnd FILL
XFILL_6__453_ vdd gnd FILL
XFILL_6__384_ vdd gnd FILL
XFILL_1__493_ vdd gnd FILL
XFILL_3__509_ vdd gnd FILL
XFILL_5__471_ vdd gnd FILL
XFILL_7__418_ vdd gnd FILL
XFILL_5__540_ vdd gnd FILL
XFILL_7__349_ vdd gnd FILL
XFILL_2__527_ vdd gnd FILL
XFILL_2__458_ vdd gnd FILL
X_602_ _602_/D _606_/CLK _602_/Q vdd gnd DFFPOSX1
XFILL_9__380_ vdd gnd FILL
XFILL_2__389_ vdd gnd FILL
X_464_ _464_/A _503_/B _464_/C _464_/D _575_/D vdd gnd AOI22X1
X_533_ _587_/Q _556_/B _534_/C vdd gnd NAND2X1
XFILL_5_BUFX2_insert17 vdd gnd FILL
XFILL75750x28950 vdd gnd FILL
XFILL_6__505_ vdd gnd FILL
X_395_ _395_/A _439_/A _395_/C _565_/D vdd gnd OAI21X1
XFILL_6__298_ vdd gnd FILL
XFILL_6__436_ vdd gnd FILL
XFILL_6__367_ vdd gnd FILL
XFILL_1__614_ vdd gnd FILL
XFILL_1__476_ vdd gnd FILL
XFILL_1__545_ vdd gnd FILL
XFILL_2__312_ vdd gnd FILL
XFILL_5__454_ vdd gnd FILL
XFILL_5__385_ vdd gnd FILL
XFILL_5__523_ vdd gnd FILL
XFILL_9__501_ vdd gnd FILL
XFILL_0__494_ vdd gnd FILL
XFILL_9__432_ vdd gnd FILL
XFILL_9__294_ vdd gnd FILL
X_447_ _447_/A _452_/B _447_/C _572_/D vdd gnd OAI21X1
X_516_ _609_/D _610_/D _517_/B vdd gnd NOR2X1
XFILL_1__330_ vdd gnd FILL
X_378_ _378_/A _378_/B _378_/C _563_/D vdd gnd OAI21X1
XFILL_4__472_ vdd gnd FILL
XFILL_4__541_ vdd gnd FILL
XFILL_6__419_ vdd gnd FILL
XFILL_1_BUFX2_insert15 vdd gnd FILL
XFILL_1__459_ vdd gnd FILL
XFILL_8__450_ vdd gnd FILL
XFILL_1__528_ vdd gnd FILL
XFILL_8__381_ vdd gnd FILL
XFILL_5__506_ vdd gnd FILL
XFILL_3__490_ vdd gnd FILL
XFILL_9_BUFX2_insert9 vdd gnd FILL
X_301_ _301_/A _567_/Q _302_/C vdd gnd NAND2X1
XFILL_5__437_ vdd gnd FILL
XFILL_5__368_ vdd gnd FILL
XFILL_5__299_ vdd gnd FILL
XFILL_0__615_ vdd gnd FILL
XFILL_0__477_ vdd gnd FILL
XFILL_8_BUFX2_insert10 vdd gnd FILL
XFILL_8_BUFX2_insert21 vdd gnd FILL
XFILL_0__546_ vdd gnd FILL
XFILL_9__415_ vdd gnd FILL
XFILL_9__346_ vdd gnd FILL
XFILL_1__313_ vdd gnd FILL
XFILL_4__455_ vdd gnd FILL
XFILL_4__386_ vdd gnd FILL
XFILL_4__524_ vdd gnd FILL
XFILL_8__502_ vdd gnd FILL
XFILL_8__433_ vdd gnd FILL
XFILL_8__364_ vdd gnd FILL
XFILL_8__295_ vdd gnd FILL
XFILL_0__400_ vdd gnd FILL
XFILL_0__331_ vdd gnd FILL
XFILL_3__473_ vdd gnd FILL
XFILL_3__542_ vdd gnd FILL
XFILL_2_CLKBUF1_insert4 vdd gnd FILL
XCLKBUF1_insert3 clk _605_/CLK vdd gnd CLKBUF1
XFILL75450x25350 vdd gnd FILL
XFILL_7__451_ vdd gnd FILL
XFILL_7__520_ vdd gnd FILL
XFILL_0__529_ vdd gnd FILL
XFILL_7__382_ vdd gnd FILL
XFILL_2__491_ vdd gnd FILL
XFILL_4__507_ vdd gnd FILL
XFILL_4__369_ vdd gnd FILL
XFILL_4__438_ vdd gnd FILL
XFILL_8__416_ vdd gnd FILL
XFILL_8__347_ vdd gnd FILL
XFILL_0__314_ vdd gnd FILL
XFILL_8__278_ vdd gnd FILL
XFILL_3__456_ vdd gnd FILL
XFILL_3__525_ vdd gnd FILL
XFILL_3__387_ vdd gnd FILL
XFILL_7__503_ vdd gnd FILL
XFILL_7__434_ vdd gnd FILL
XFILL_7__296_ vdd gnd FILL
XFILL_7_CLKBUF1_insert6 vdd gnd FILL
XFILL_7__365_ vdd gnd FILL
XFILL_2__543_ vdd gnd FILL
XFILL_2__474_ vdd gnd FILL
X_480_ _596_/Q _490_/B vdd gnd INVX1
XFILL_3__310_ vdd gnd FILL
XFILL_6__452_ vdd gnd FILL
XFILL_6__521_ vdd gnd FILL
XFILL_6__383_ vdd gnd FILL
XFILL_1__492_ vdd gnd FILL
XFILL_3__508_ vdd gnd FILL
XFILL_3__439_ vdd gnd FILL
XFILL_5__470_ vdd gnd FILL
XFILL_7__417_ vdd gnd FILL
XFILL_7__348_ vdd gnd FILL
XFILL_7__279_ vdd gnd FILL
XFILL_2__457_ vdd gnd FILL
XFILL_2__526_ vdd gnd FILL
X_601_ _601_/D _601_/CLK _601_/Q vdd gnd DFFPOSX1
XFILL_2__388_ vdd gnd FILL
XFILL_5_BUFX2_insert18 vdd gnd FILL
X_463_ _463_/A _463_/B _503_/B _464_/D vdd gnd AOI21X1
X_532_ _540_/A _556_/B _532_/C _586_/D vdd gnd OAI21X1
X_394_ _439_/A _394_/B _394_/C _395_/C vdd gnd NAND3X1
XFILL_6__435_ vdd gnd FILL
XFILL_6__504_ vdd gnd FILL
XFILL_6__297_ vdd gnd FILL
XFILL_6__366_ vdd gnd FILL
XFILL_1__613_ vdd gnd FILL
XFILL_1__544_ vdd gnd FILL
XFILL_1__475_ vdd gnd FILL
XFILL_2__311_ vdd gnd FILL
XFILL_5__522_ vdd gnd FILL
XFILL_5__453_ vdd gnd FILL
XFILL_5__384_ vdd gnd FILL
XFILL_0__493_ vdd gnd FILL
XFILL_9__500_ vdd gnd FILL
XFILL_2__509_ vdd gnd FILL
XFILL_9__293_ vdd gnd FILL
X_515_ _515_/A _515_/B _581_/D vdd gnd NAND2X1
XFILL_9__362_ vdd gnd FILL
X_446_ _460_/B _446_/B _446_/C _447_/C vdd gnd NAND3X1
X_377_ _563_/Q _378_/A _378_/C vdd gnd NAND2X1
XFILL_4__471_ vdd gnd FILL
XFILL_6__418_ vdd gnd FILL
XFILL_4__540_ vdd gnd FILL
XFILL_1_BUFX2_insert16 vdd gnd FILL
XFILL_6__349_ vdd gnd FILL
XFILL_1__527_ vdd gnd FILL
XFILL_1__458_ vdd gnd FILL
XFILL_8__380_ vdd gnd FILL
XFILL_1__389_ vdd gnd FILL
XFILL_5__505_ vdd gnd FILL
X_300_ _579_/Q _493_/A vdd gnd INVX1
XFILL_5__298_ vdd gnd FILL
XFILL_5__436_ vdd gnd FILL
XFILL_5__367_ vdd gnd FILL
XFILL_0__614_ vdd gnd FILL
XFILL_8_BUFX2_insert11 vdd gnd FILL
XFILL_0__476_ vdd gnd FILL
XFILL_8_BUFX2_insert22 vdd gnd FILL
XFILL_0__545_ vdd gnd FILL
XFILL_9__414_ vdd gnd FILL
XFILL_9__345_ vdd gnd FILL
XFILL_9__276_ vdd gnd FILL
XFILL_4__523_ vdd gnd FILL
XFILL_1__312_ vdd gnd FILL
X_429_ _429_/A _431_/B _429_/C _433_/C vdd gnd NAND3X1
XFILL_4__454_ vdd gnd FILL
XFILL_4__385_ vdd gnd FILL
XFILL_8__501_ vdd gnd FILL
XFILL_8__294_ vdd gnd FILL
XFILL_8__432_ vdd gnd FILL
XFILL_8__363_ vdd gnd FILL
XFILL_0__330_ vdd gnd FILL
XFILL_3__472_ vdd gnd FILL
XFILL_2_CLKBUF1_insert5 vdd gnd FILL
XFILL_5__419_ vdd gnd FILL
XFILL_3__541_ vdd gnd FILL
XFILL_0__528_ vdd gnd FILL
XCLKBUF1_insert4 clk _595_/CLK vdd gnd CLKBUF1
XFILL_0__459_ vdd gnd FILL
XFILL_7__450_ vdd gnd FILL
XFILL_7__381_ vdd gnd FILL
XFILL_9__328_ vdd gnd FILL
XFILL_2__490_ vdd gnd FILL
XFILL_4_BUFX2_insert20 vdd gnd FILL
XFILL_4__506_ vdd gnd FILL
XFILL74850x28950 vdd gnd FILL
XFILL_4__299_ vdd gnd FILL
XFILL_4__437_ vdd gnd FILL
XFILL_4__368_ vdd gnd FILL
XFILL_8_CLKBUF1_insert0 vdd gnd FILL
XFILL_8__277_ vdd gnd FILL
XFILL_8__415_ vdd gnd FILL
XFILL_8__346_ vdd gnd FILL
XFILL_0__313_ vdd gnd FILL
XFILL_3__455_ vdd gnd FILL
XFILL_3__386_ vdd gnd FILL
XFILL_3__524_ vdd gnd FILL
XFILL_7__502_ vdd gnd FILL
XFILL_7__433_ vdd gnd FILL
XFILL_7__364_ vdd gnd FILL
XFILL_7__295_ vdd gnd FILL
XFILL_2__473_ vdd gnd FILL
XFILL_2__542_ vdd gnd FILL
XFILL_6__451_ vdd gnd FILL
XFILL_6__520_ vdd gnd FILL
XFILL_8__329_ vdd gnd FILL
XFILL_6__382_ vdd gnd FILL
XFILL_1__491_ vdd gnd FILL
XFILL_3__507_ vdd gnd FILL
XFILL_3__369_ vdd gnd FILL
XFILL_3__438_ vdd gnd FILL
XFILL_7__416_ vdd gnd FILL
XFILL_7__347_ vdd gnd FILL
XFILL_7__278_ vdd gnd FILL
XFILL_2__456_ vdd gnd FILL
XFILL_2__525_ vdd gnd FILL
X_600_ _600_/D _601_/CLK _600_/Q vdd gnd DFFPOSX1
XFILL_2__387_ vdd gnd FILL
X_531_ _586_/Q _556_/B _532_/C vdd gnd NAND2X1
XFILL_5_BUFX2_insert19 vdd gnd FILL
X_462_ _463_/A _463_/B _464_/C vdd gnd OR2X2
X_393_ _393_/A _393_/B _393_/C _394_/C vdd gnd NAND3X1
XFILL_6__503_ vdd gnd FILL
XFILL_6__365_ vdd gnd FILL
XFILL_6__434_ vdd gnd FILL
XFILL_6__296_ vdd gnd FILL
XFILL_1__474_ vdd gnd FILL
XFILL_1__543_ vdd gnd FILL
XFILL_2__310_ vdd gnd FILL
XFILL74550x25350 vdd gnd FILL
XFILL_5__452_ vdd gnd FILL
XFILL_5__521_ vdd gnd FILL
XFILL_5__383_ vdd gnd FILL
XFILL_0__492_ vdd gnd FILL
XFILL_2__508_ vdd gnd FILL
XFILL_2__439_ vdd gnd FILL
XFILL_9__430_ vdd gnd FILL
X_514_ _625_/A _514_/B _514_/C _515_/B vdd gnd NAND3X1
XFILL_9__361_ vdd gnd FILL
X_445_ _490_/A _457_/A _448_/B _446_/B vdd gnd OAI21X1
X_376_ _376_/A _376_/B _378_/B vdd gnd NAND2X1
XFILL_4__470_ vdd gnd FILL
XFILL_6__417_ vdd gnd FILL
XFILL_6__348_ vdd gnd FILL
XFILL_6_BUFX2_insert7 vdd gnd FILL
XFILL_6__279_ vdd gnd FILL
XFILL_1_BUFX2_insert17 vdd gnd FILL
XFILL_1__457_ vdd gnd FILL
XFILL_1__526_ vdd gnd FILL
XFILL_1__388_ vdd gnd FILL
XFILL_5__435_ vdd gnd FILL
XFILL_5__504_ vdd gnd FILL
XFILL_5__297_ vdd gnd FILL
XBUFX2_insert20 _612_/Q _460_/B vdd gnd BUFX2
XFILL_5__366_ vdd gnd FILL
XFILL_0__613_ vdd gnd FILL
XFILL_0__544_ vdd gnd FILL
XFILL_8_BUFX2_insert12 vdd gnd FILL
XFILL_0__475_ vdd gnd FILL
XFILL_8_BUFX2_insert23 vdd gnd FILL
XFILL_9__413_ vdd gnd FILL
XFILL_9__275_ vdd gnd FILL
XFILL_1__311_ vdd gnd FILL
X_428_ _442_/C _582_/Q _431_/B vdd gnd NAND2X1
XFILL_4__522_ vdd gnd FILL
X_359_ _359_/A _591_/Q _360_/B vdd gnd OR2X2
XFILL_4__453_ vdd gnd FILL
XFILL_4__384_ vdd gnd FILL
XFILL_8__500_ vdd gnd FILL
XFILL_1__509_ vdd gnd FILL
XFILL_8__431_ vdd gnd FILL
XFILL_8__293_ vdd gnd FILL
XFILL_8__362_ vdd gnd FILL
XFILL_3__540_ vdd gnd FILL
XFILL_3__471_ vdd gnd FILL
XFILL_2_CLKBUF1_insert6 vdd gnd FILL
XFILL_5__418_ vdd gnd FILL
XFILL_5__349_ vdd gnd FILL
XCLKBUF1_insert5 clk _612_/CLK vdd gnd CLKBUF1
XFILL_0__527_ vdd gnd FILL
XFILL_0__458_ vdd gnd FILL
XFILL_9__327_ vdd gnd FILL
XFILL_7__380_ vdd gnd FILL
XFILL_0__389_ vdd gnd FILL
XFILL_4_BUFX2_insert10 vdd gnd FILL
XFILL_4_BUFX2_insert21 vdd gnd FILL
XFILL_4__436_ vdd gnd FILL
XFILL_4__505_ vdd gnd FILL
XFILL_4__298_ vdd gnd FILL
XFILL_4__367_ vdd gnd FILL
XFILL_8_CLKBUF1_insert1 vdd gnd FILL
XFILL_8__414_ vdd gnd FILL
XFILL_0__312_ vdd gnd FILL
XFILL_8__345_ vdd gnd FILL
XFILL_8__276_ vdd gnd FILL
XFILL_3__523_ vdd gnd FILL
XFILL_3__454_ vdd gnd FILL
XFILL_3__385_ vdd gnd FILL
XFILL_7__501_ vdd gnd FILL
XFILL75750x54150 vdd gnd FILL
XFILL_7__294_ vdd gnd FILL
XFILL_7__432_ vdd gnd FILL
XFILL_7__363_ vdd gnd FILL
XFILL_2__472_ vdd gnd FILL
XFILL_4__419_ vdd gnd FILL
XFILL_2__541_ vdd gnd FILL
XFILL_6__450_ vdd gnd FILL
XFILL_6__381_ vdd gnd FILL
XFILL_8__328_ vdd gnd FILL
XFILL_1__490_ vdd gnd FILL
XFILL_3__506_ vdd gnd FILL
XFILL_3__299_ vdd gnd FILL
XFILL_3__437_ vdd gnd FILL
XFILL_3__368_ vdd gnd FILL
XFILL_7__415_ vdd gnd FILL
XFILL_7__277_ vdd gnd FILL
XFILL_7__346_ vdd gnd FILL
XFILL_2__455_ vdd gnd FILL
XFILL_2__386_ vdd gnd FILL
XFILL_2__524_ vdd gnd FILL
X_461_ _490_/A _461_/B _461_/C _463_/A vdd gnd OAI21X1
X_530_ _542_/A _554_/B _530_/C _585_/D vdd gnd OAI21X1
XFILL_6__502_ vdd gnd FILL
X_392_ _430_/C _586_/Q _393_/B vdd gnd NAND2X1
XFILL_6__433_ vdd gnd FILL
XFILL_6__364_ vdd gnd FILL
XFILL_6__295_ vdd gnd FILL
XFILL_1__473_ vdd gnd FILL
XFILL_1__542_ vdd gnd FILL
XFILL_5__451_ vdd gnd FILL
XFILL_5__520_ vdd gnd FILL
XFILL_5__382_ vdd gnd FILL
XFILL_7__329_ vdd gnd FILL
XFILL_0__491_ vdd gnd FILL
XFILL_2__507_ vdd gnd FILL
XFILL73950x28950 vdd gnd FILL
XFILL_2__369_ vdd gnd FILL
XFILL_9__360_ vdd gnd FILL
XFILL_2__438_ vdd gnd FILL
XFILL_9__291_ vdd gnd FILL
X_513_ _513_/A _513_/B _514_/B vdd gnd NAND2X1
X_444_ _604_/Q _605_/Q _457_/A vdd gnd NOR2X1
X_375_ _538_/A _375_/B _376_/A vdd gnd NAND2X1
XFILL_1_BUFX2_insert18 vdd gnd FILL
XFILL_6_BUFX2_insert8 vdd gnd FILL
XFILL_6__278_ vdd gnd FILL
XFILL_6__416_ vdd gnd FILL
XFILL_6__347_ vdd gnd FILL
XFILL_9__489_ vdd gnd FILL
XFILL_1__456_ vdd gnd FILL
XFILL_1__387_ vdd gnd FILL
XFILL_1__525_ vdd gnd FILL
XFILL_5__503_ vdd gnd FILL
XFILL_5__365_ vdd gnd FILL
XFILL_5__434_ vdd gnd FILL
XFILL_5__296_ vdd gnd FILL
XBUFX2_insert10 selXY _301_/A vdd gnd BUFX2
XBUFX2_insert21 _340_/Y _421_/B vdd gnd BUFX2
XFILL_0__474_ vdd gnd FILL
XFILL_8_BUFX2_insert24 vdd gnd FILL
XFILL_0__543_ vdd gnd FILL
XFILL_8_BUFX2_insert13 vdd gnd FILL
XFILL_3_CLKBUF1_insert0 vdd gnd FILL
XFILL_9__343_ vdd gnd FILL
XFILL_9__274_ vdd gnd FILL
X_427_ _432_/A _429_/A vdd gnd INVX1
XFILL_1__310_ vdd gnd FILL
X_358_ _591_/Q _359_/A _360_/A vdd gnd NAND2X1
X_289_ _301_/A _563_/Q _290_/C vdd gnd NAND2X1
XFILL_4__452_ vdd gnd FILL
XFILL_4__521_ vdd gnd FILL
XFILL_4__383_ vdd gnd FILL
XFILL_1__508_ vdd gnd FILL
XFILL_8__361_ vdd gnd FILL
XFILL_1__439_ vdd gnd FILL
XFILL_8__430_ vdd gnd FILL
XFILL_8__292_ vdd gnd FILL
XFILL_3__470_ vdd gnd FILL
XFILL_5__417_ vdd gnd FILL
XFILL_5__348_ vdd gnd FILL
XFILL_5__279_ vdd gnd FILL
XCLKBUF1_insert6 clk _573_/CLK vdd gnd CLKBUF1
XFILL_0__457_ vdd gnd FILL
XFILL_0__526_ vdd gnd FILL
XFILL_9__326_ vdd gnd FILL
XFILL_0__388_ vdd gnd FILL
XFILL_4_BUFX2_insert11 vdd gnd FILL
XFILL_4_BUFX2_insert22 vdd gnd FILL
XFILL_4__435_ vdd gnd FILL
XFILL_4__504_ vdd gnd FILL
XFILL_4__297_ vdd gnd FILL
XFILL_4__366_ vdd gnd FILL
XFILL_8_CLKBUF1_insert2 vdd gnd FILL
XFILL_8__413_ vdd gnd FILL
XFILL_8__344_ vdd gnd FILL
XFILL_8__275_ vdd gnd FILL
XFILL_0__311_ vdd gnd FILL
XFILL_3__453_ vdd gnd FILL
XFILL_3__522_ vdd gnd FILL
XFILL_3__384_ vdd gnd FILL
XFILL_7__500_ vdd gnd FILL
XFILL_0__509_ vdd gnd FILL
XFILL_7__431_ vdd gnd FILL
XFILL_7__293_ vdd gnd FILL
XFILL_7__362_ vdd gnd FILL
XFILL_9__309_ vdd gnd FILL
XFILL_2__540_ vdd gnd FILL
XFILL_2__471_ vdd gnd FILL
XFILL_4__418_ vdd gnd FILL
XFILL_4__349_ vdd gnd FILL
XFILL_0_BUFX2_insert20 vdd gnd FILL
XFILL_8__327_ vdd gnd FILL
XFILL_6__380_ vdd gnd FILL
XFILL_3__436_ vdd gnd FILL
XFILL_3__505_ vdd gnd FILL
XFILL_3__298_ vdd gnd FILL
XFILL_3__367_ vdd gnd FILL
XFILL_7__414_ vdd gnd FILL
XFILL_7__345_ vdd gnd FILL
XFILL_7__276_ vdd gnd FILL
XFILL_2__523_ vdd gnd FILL
XFILL_2__454_ vdd gnd FILL
XFILL_2__385_ vdd gnd FILL
X_460_ _460_/A _460_/B _460_/C _574_/D vdd gnd OAI21X1
X_391_ _587_/Q _393_/A vdd gnd INVX1
XFILL_6__501_ vdd gnd FILL
XFILL_6__432_ vdd gnd FILL
XFILL_6__294_ vdd gnd FILL
XFILL_6__363_ vdd gnd FILL
XFILL_1__472_ vdd gnd FILL
X_589_ _589_/D _595_/CLK _589_/Q vdd gnd DFFPOSX1
XFILL_3__419_ vdd gnd FILL
XFILL_1__541_ vdd gnd FILL
XFILL_5__450_ vdd gnd FILL
XFILL_7__328_ vdd gnd FILL
XFILL_5__381_ vdd gnd FILL
XFILL_0__490_ vdd gnd FILL
XFILL_2__437_ vdd gnd FILL
XFILL_2__506_ vdd gnd FILL
XFILL_2__299_ vdd gnd FILL
XFILL_9__290_ vdd gnd FILL
XFILL_2__368_ vdd gnd FILL
X_512_ _512_/A _512_/B _512_/C _513_/B vdd gnd NAND3X1
X_443_ _448_/C _448_/B _446_/C vdd gnd OR2X2
X_374_ _375_/B _538_/A _376_/B vdd gnd OR2X2
XFILL_6__415_ vdd gnd FILL
XFILL_6__277_ vdd gnd FILL
XFILL_1_BUFX2_insert19 vdd gnd FILL
XFILL_6_BUFX2_insert9 vdd gnd FILL
XFILL_6__346_ vdd gnd FILL
XFILL_9__488_ vdd gnd FILL
XFILL_1__524_ vdd gnd FILL
XFILL_1__455_ vdd gnd FILL
XFILL_1__386_ vdd gnd FILL
XFILL_5__502_ vdd gnd FILL
XFILL_5__295_ vdd gnd FILL
XFILL_5__433_ vdd gnd FILL
XFILL_5__364_ vdd gnd FILL
XBUFX2_insert11 _557_/Q _511_/C vdd gnd BUFX2
XBUFX2_insert22 _340_/Y _410_/B vdd gnd BUFX2
XFILL_0__473_ vdd gnd FILL
XFILL_8_BUFX2_insert25 vdd gnd FILL
XFILL_8_BUFX2_insert14 vdd gnd FILL
XFILL_0__542_ vdd gnd FILL
XFILL_9__411_ vdd gnd FILL
XFILL_3_CLKBUF1_insert1 vdd gnd FILL
XFILL_9__342_ vdd gnd FILL
XFILL75750x39750 vdd gnd FILL
X_426_ _426_/A _426_/B _432_/A vdd gnd NAND2X1
X_357_ _490_/A _357_/B _357_/C _359_/A vdd gnd OAI21X1
X_288_ _575_/Q _464_/A vdd gnd INVX1
XFILL_4__451_ vdd gnd FILL
XFILL_4__520_ vdd gnd FILL
XFILL_4__382_ vdd gnd FILL
XFILL_6__329_ vdd gnd FILL
XFILL_1__507_ vdd gnd FILL
XFILL_1__369_ vdd gnd FILL
XFILL_8__360_ vdd gnd FILL
XFILL_1__438_ vdd gnd FILL
XFILL_8__291_ vdd gnd FILL
XFILL_5__278_ vdd gnd FILL
XFILL_5__416_ vdd gnd FILL
XFILL_5__347_ vdd gnd FILL
XFILL_8__489_ vdd gnd FILL
XFILL_0__456_ vdd gnd FILL
XFILL_0__387_ vdd gnd FILL
XFILL_0__525_ vdd gnd FILL
XFILL75150x10950 vdd gnd FILL
XFILL75750x14550 vdd gnd FILL
XFILL_4_BUFX2_insert12 vdd gnd FILL
XFILL_4__503_ vdd gnd FILL
XFILL_4_BUFX2_insert23 vdd gnd FILL
X_409_ _409_/A _409_/B _410_/B _410_/D vdd gnd AOI21X1
XFILL_4__365_ vdd gnd FILL
XFILL_4__434_ vdd gnd FILL
XFILL_4__296_ vdd gnd FILL
XFILL_8_CLKBUF1_insert3 vdd gnd FILL
XFILL_8__274_ vdd gnd FILL
XFILL_8__412_ vdd gnd FILL
XFILL_8__343_ vdd gnd FILL
XFILL_0__310_ vdd gnd FILL
XFILL_3__452_ vdd gnd FILL
XFILL_3__521_ vdd gnd FILL
XFILL_3__383_ vdd gnd FILL
XFILL_0__508_ vdd gnd FILL
XFILL_7__361_ vdd gnd FILL
XFILL_0__439_ vdd gnd FILL
XFILL_7__430_ vdd gnd FILL
XFILL_7__292_ vdd gnd FILL
XFILL_9__308_ vdd gnd FILL
XFILL_2__470_ vdd gnd FILL
XFILL_4__279_ vdd gnd FILL
XFILL_4__417_ vdd gnd FILL
XFILL_4__348_ vdd gnd FILL
XFILL_0_BUFX2_insert10 vdd gnd FILL
XFILL_0_BUFX2_insert21 vdd gnd FILL
XFILL_8__326_ vdd gnd FILL
XFILL_3__435_ vdd gnd FILL
XFILL_3__366_ vdd gnd FILL
XFILL_3__504_ vdd gnd FILL
XFILL_3__297_ vdd gnd FILL
XFILL75450x36150 vdd gnd FILL
XFILL_7__413_ vdd gnd FILL
XFILL_7__344_ vdd gnd FILL
XFILL_7__275_ vdd gnd FILL
XFILL_2__453_ vdd gnd FILL
XFILL_2__522_ vdd gnd FILL
XFILL_2__384_ vdd gnd FILL
X_390_ _430_/C _587_/Q _390_/C _394_/B vdd gnd NAND3X1
XFILL_6__500_ vdd gnd FILL
XFILL_6__431_ vdd gnd FILL
XFILL_6__293_ vdd gnd FILL
XFILL_6__362_ vdd gnd FILL
XFILL_8__309_ vdd gnd FILL
XFILL_1__540_ vdd gnd FILL
XFILL_1__471_ vdd gnd FILL
X_588_ _588_/D _595_/CLK _588_/Q vdd gnd DFFPOSX1
XFILL_3__418_ vdd gnd FILL
XFILL_3__349_ vdd gnd FILL
XFILL_7__327_ vdd gnd FILL
XFILL_5__380_ vdd gnd FILL
XFILL_2__436_ vdd gnd FILL
XFILL_2__505_ vdd gnd FILL
XFILL_2__298_ vdd gnd FILL
X_511_ _596_/Q _597_/Q _511_/C _512_/A vdd gnd OAI21X1
XFILL_2__367_ vdd gnd FILL
X_442_ _604_/Q _605_/Q _442_/C _448_/C vdd gnd OAI21X1
X_373_ _588_/Q _399_/A _415_/A _375_/B vdd gnd OAI21X1
XFILL_6__414_ vdd gnd FILL
XFILL_6__345_ vdd gnd FILL
XFILL_9__625_ vdd gnd FILL
XFILL_9__556_ vdd gnd FILL
XFILL_6__276_ vdd gnd FILL
XFILL_1__523_ vdd gnd FILL
XFILL_1__454_ vdd gnd FILL
XFILL_1__385_ vdd gnd FILL
XFILL_5__501_ vdd gnd FILL
XFILL_5__432_ vdd gnd FILL
XFILL_5__294_ vdd gnd FILL
XFILL_5__363_ vdd gnd FILL
XBUFX2_insert12 _557_/Q _509_/A vdd gnd BUFX2
XBUFX2_insert23 _340_/Y _378_/A vdd gnd BUFX2
XFILL_0__541_ vdd gnd FILL
XFILL_0__472_ vdd gnd FILL
XFILL_9__410_ vdd gnd FILL
XFILL_2__419_ vdd gnd FILL
XFILL_8_BUFX2_insert15 vdd gnd FILL
XFILL_3_CLKBUF1_insert2 vdd gnd FILL
XFILL_9__341_ vdd gnd FILL
X_287_ _301_/A _460_/A _287_/C _619_/A vdd gnd OAI21X1
X_425_ _583_/Q _506_/B _426_/B vdd gnd NAND2X1
X_356_ _378_/A _356_/B _356_/C _560_/D vdd gnd OAI21X1
XFILL_4__450_ vdd gnd FILL
XFILL_6__328_ vdd gnd FILL
XFILL_4__381_ vdd gnd FILL
XFILL_1__437_ vdd gnd FILL
XFILL_1__506_ vdd gnd FILL
XFILL_1__299_ vdd gnd FILL
XFILL_8__290_ vdd gnd FILL
XFILL_1__368_ vdd gnd FILL
XFILL_5__415_ vdd gnd FILL
XFILL_5__277_ vdd gnd FILL
XFILL_5__346_ vdd gnd FILL
XFILL_8__488_ vdd gnd FILL
XFILL_0__524_ vdd gnd FILL
XFILL_0__455_ vdd gnd FILL
XFILL_0__386_ vdd gnd FILL
X_408_ _409_/A _409_/B _410_/C vdd gnd OR2X2
XFILL_9__324_ vdd gnd FILL
XFILL_4__502_ vdd gnd FILL
XFILL_4_BUFX2_insert24 vdd gnd FILL
XFILL_4_BUFX2_insert13 vdd gnd FILL
X_339_ _592_/Q _544_/B vdd gnd INVX1
XFILL_4__295_ vdd gnd FILL
XFILL_4__433_ vdd gnd FILL
XFILL_4__364_ vdd gnd FILL
XFILL_8_CLKBUF1_insert4 vdd gnd FILL
XFILL_8__411_ vdd gnd FILL
XFILL_8__273_ vdd gnd FILL
XFILL_8__342_ vdd gnd FILL
XFILL_3__520_ vdd gnd FILL
XFILL_3__451_ vdd gnd FILL
XFILL_3__382_ vdd gnd FILL
XFILL_5__329_ vdd gnd FILL
XFILL_0__507_ vdd gnd FILL
XFILL_7__291_ vdd gnd FILL
XFILL_0__369_ vdd gnd FILL
XFILL_7__360_ vdd gnd FILL
XFILL_0__438_ vdd gnd FILL
XFILL_4__416_ vdd gnd FILL
XFILL_0_BUFX2_insert11 vdd gnd FILL
XFILL_0_BUFX2_insert22 vdd gnd FILL
XFILL_4__278_ vdd gnd FILL
XFILL_4__347_ vdd gnd FILL
XFILL_7__489_ vdd gnd FILL
XFILL_8__325_ vdd gnd FILL
XFILL_3__503_ vdd gnd FILL
XFILL_3__296_ vdd gnd FILL
XFILL_3__365_ vdd gnd FILL
XFILL_3__434_ vdd gnd FILL
XFILL_7__274_ vdd gnd FILL
XFILL_7__412_ vdd gnd FILL
XFILL_7__343_ vdd gnd FILL
XFILL74850x39750 vdd gnd FILL
XFILL_2__452_ vdd gnd FILL
XFILL_2__521_ vdd gnd FILL
XFILL_2__383_ vdd gnd FILL
XFILL_6__361_ vdd gnd FILL
XFILL_6__430_ vdd gnd FILL
XFILL_6__292_ vdd gnd FILL
XFILL_8__308_ vdd gnd FILL
XFILL_1__470_ vdd gnd FILL
X_587_ _587_/D _612_/CLK _587_/Q vdd gnd DFFPOSX1
XFILL_3__279_ vdd gnd FILL
XFILL_3__417_ vdd gnd FILL
XFILL_3__348_ vdd gnd FILL
XFILL74250x10950 vdd gnd FILL
XFILL_7__326_ vdd gnd FILL
XFILL_3_BUFX2_insert7 vdd gnd FILL
XFILL_2__435_ vdd gnd FILL
XFILL_2__366_ vdd gnd FILL
XFILL_2__504_ vdd gnd FILL
XFILL_2__297_ vdd gnd FILL
X_510_ _510_/A _512_/B _510_/C _514_/C vdd gnd NAND3X1
X_441_ _602_/Q _448_/B vdd gnd INVX1
XFILL73050x72150 vdd gnd FILL
X_372_ _589_/Q _538_/A vdd gnd INVX1
XFILL_6__413_ vdd gnd FILL
XFILL_6__344_ vdd gnd FILL
XFILL_9__624_ vdd gnd FILL
XFILL_9__486_ vdd gnd FILL
XFILL_9__555_ vdd gnd FILL
XFILL_6__275_ vdd gnd FILL
XFILL_1__453_ vdd gnd FILL
XFILL_1__522_ vdd gnd FILL
XFILL_1__384_ vdd gnd FILL
XFILL_5__500_ vdd gnd FILL
XFILL_5__362_ vdd gnd FILL
XFILL_5__431_ vdd gnd FILL
XFILL_5__293_ vdd gnd FILL
XBUFX2_insert24 _340_/Y _503_/B vdd gnd BUFX2
XFILL_7__309_ vdd gnd FILL
XBUFX2_insert13 _557_/Q _442_/C vdd gnd BUFX2
XFILL_0__540_ vdd gnd FILL
XFILL_0__471_ vdd gnd FILL
XFILL_8_BUFX2_insert16 vdd gnd FILL
XFILL_2__418_ vdd gnd FILL
XFILL_2__349_ vdd gnd FILL
XFILL_3_CLKBUF1_insert3 vdd gnd FILL
X_424_ selSign _506_/B vdd gnd INVX1
X_286_ _286_/A _562_/Q _287_/C vdd gnd NAND2X1
X_355_ _560_/Q _378_/A _356_/C vdd gnd NAND2X1
XFILL_6__327_ vdd gnd FILL
XFILL_4__380_ vdd gnd FILL
XFILL_9__469_ vdd gnd FILL
XFILL_9__538_ vdd gnd FILL
XFILL_1__436_ vdd gnd FILL
XFILL_1__505_ vdd gnd FILL
XFILL_1__367_ vdd gnd FILL
XFILL_1__298_ vdd gnd FILL
XFILL74550x36150 vdd gnd FILL
XFILL_5__414_ vdd gnd FILL
XFILL_5__345_ vdd gnd FILL
XFILL_8__625_ vdd gnd FILL
XFILL_8__556_ vdd gnd FILL
XFILL_5__276_ vdd gnd FILL
XFILL_8__487_ vdd gnd FILL
XFILL_0__454_ vdd gnd FILL
XFILL_0__523_ vdd gnd FILL
XFILL_9__323_ vdd gnd FILL
XFILL_0__385_ vdd gnd FILL
X_338_ _478_/A _490_/A _338_/C _557_/D vdd gnd OAI21X1
X_407_ _490_/A _407_/B _431_/C _409_/A vdd gnd OAI21X1
XFILL_4_BUFX2_insert14 vdd gnd FILL
XFILL_4__501_ vdd gnd FILL
XFILL_4_BUFX2_insert25 vdd gnd FILL
XFILL_4__432_ vdd gnd FILL
XFILL_4__294_ vdd gnd FILL
XFILL_4__363_ vdd gnd FILL
XFILL_8_CLKBUF1_insert5 vdd gnd FILL
XFILL_8__410_ vdd gnd FILL
XFILL_1__419_ vdd gnd FILL
XFILL_8__341_ vdd gnd FILL
XFILL_3__450_ vdd gnd FILL
XFILL_5__328_ vdd gnd FILL
XFILL_3__381_ vdd gnd FILL
XFILL_8__539_ vdd gnd FILL
XFILL_0__437_ vdd gnd FILL
XFILL_0__506_ vdd gnd FILL
XFILL_0__299_ vdd gnd FILL
XFILL_7__290_ vdd gnd FILL
XFILL_9__306_ vdd gnd FILL
XFILL_0__368_ vdd gnd FILL
XFILL_4__415_ vdd gnd FILL
XFILL_4__277_ vdd gnd FILL
XFILL_0_BUFX2_insert12 vdd gnd FILL
XFILL_0_BUFX2_insert23 vdd gnd FILL
XFILL_4__346_ vdd gnd FILL
XFILL_7__488_ vdd gnd FILL
XFILL_8__324_ vdd gnd FILL
XFILL_3__502_ vdd gnd FILL
XFILL_3__433_ vdd gnd FILL
XFILL_3__295_ vdd gnd FILL
XFILL_3__364_ vdd gnd FILL
XFILL_7__411_ vdd gnd FILL
XFILL_7__273_ vdd gnd FILL
XFILL_7__342_ vdd gnd FILL
XFILL_2__520_ vdd gnd FILL
XFILL_2__451_ vdd gnd FILL
XFILL_4__329_ vdd gnd FILL
XFILL_2__382_ vdd gnd FILL
XFILL_6__291_ vdd gnd FILL
XFILL_8__307_ vdd gnd FILL
XFILL_6__360_ vdd gnd FILL
XFILL_3__416_ vdd gnd FILL
X_586_ _586_/D _606_/CLK _586_/Q vdd gnd DFFPOSX1
XFILL_3__278_ vdd gnd FILL
XFILL_3__347_ vdd gnd FILL
XFILL_6__489_ vdd gnd FILL
XFILL_7__325_ vdd gnd FILL
XFILL_3_BUFX2_insert8 vdd gnd FILL
XFILL_2__503_ vdd gnd FILL
XFILL_2__296_ vdd gnd FILL
XFILL_2__365_ vdd gnd FILL
XFILL_2__434_ vdd gnd FILL
X_440_ _440_/A _452_/B _440_/C _571_/D vdd gnd OAI21X1
X_371_ _421_/B _371_/B _371_/C _562_/D vdd gnd OAI21X1
XFILL_9__623_ vdd gnd FILL
XFILL_6__274_ vdd gnd FILL
XFILL_6__412_ vdd gnd FILL
XFILL_6__343_ vdd gnd FILL
XFILL_9__485_ vdd gnd FILL
XFILL_1__452_ vdd gnd FILL
XFILL_1__521_ vdd gnd FILL
X_569_ _569_/D _595_/CLK _569_/Q vdd gnd DFFPOSX1
XFILL_1__383_ vdd gnd FILL
XFILL_7__308_ vdd gnd FILL
XFILL_5__361_ vdd gnd FILL
XFILL_5__430_ vdd gnd FILL
XFILL_5__292_ vdd gnd FILL
XBUFX2_insert25 _340_/Y _493_/B vdd gnd BUFX2
XBUFX2_insert14 _557_/Q _415_/A vdd gnd BUFX2
XFILL_0__470_ vdd gnd FILL
XFILL_2__279_ vdd gnd FILL
XFILL_3_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__417_ vdd gnd FILL
XFILL_8_BUFX2_insert17 vdd gnd FILL
XFILL_2__348_ vdd gnd FILL
X_423_ selSign _523_/A _426_/A vdd gnd NAND2X1
X_354_ _354_/A _354_/B _356_/B vdd gnd NAND2X1
X_285_ _574_/Q _460_/A vdd gnd INVX1
XFILL_6__326_ vdd gnd FILL
XFILL_9__537_ vdd gnd FILL
XFILL_1__504_ vdd gnd FILL
XFILL_9__399_ vdd gnd FILL
XFILL_1__435_ vdd gnd FILL
XFILL_1__366_ vdd gnd FILL
XFILL_1__297_ vdd gnd FILL
XFILL_5__275_ vdd gnd FILL
XFILL_5__413_ vdd gnd FILL
XFILL_5__344_ vdd gnd FILL
XFILL_8__624_ vdd gnd FILL
XFILL_8__486_ vdd gnd FILL
XFILL_8__555_ vdd gnd FILL
XFILL_0__453_ vdd gnd FILL
XFILL_0__522_ vdd gnd FILL
XFILL_0__384_ vdd gnd FILL
X_337_ ISin _478_/A _338_/C vdd gnd NAND2X1
X_406_ _585_/Q _409_/B vdd gnd INVX1
XFILL_4_BUFX2_insert15 vdd gnd FILL
XFILL_4__500_ vdd gnd FILL
XFILL_4__362_ vdd gnd FILL
XFILL_4__431_ vdd gnd FILL
XFILL_4__293_ vdd gnd FILL
XFILL_6__309_ vdd gnd FILL
XFILL_8_CLKBUF1_insert6 vdd gnd FILL
XFILL_8__340_ vdd gnd FILL
XFILL_1__418_ vdd gnd FILL
XFILL_1__349_ vdd gnd FILL
XFILL73350x10950 vdd gnd FILL
XFILL_5__327_ vdd gnd FILL
XFILL_3__380_ vdd gnd FILL
XFILL_8__469_ vdd gnd FILL
XFILL_8__538_ vdd gnd FILL
XFILL_0__436_ vdd gnd FILL
XFILL_0__505_ vdd gnd FILL
XFILL_0__367_ vdd gnd FILL
XFILL_9__305_ vdd gnd FILL
XFILL_0__298_ vdd gnd FILL
XFILL_4__414_ vdd gnd FILL
XFILL_4__345_ vdd gnd FILL
XFILL_7__625_ vdd gnd FILL
XFILL_7__487_ vdd gnd FILL
XFILL_7__556_ vdd gnd FILL
XFILL_0_BUFX2_insert24 vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_4__276_ vdd gnd FILL
XFILL_8__323_ vdd gnd FILL
XFILL_3__501_ vdd gnd FILL
XFILL_3__432_ vdd gnd FILL
XFILL_3__294_ vdd gnd FILL
XFILL_3__363_ vdd gnd FILL
XFILL_7__410_ vdd gnd FILL
XFILL_0__419_ vdd gnd FILL
XFILL_7__341_ vdd gnd FILL
XFILL_2__450_ vdd gnd FILL
XFILL_4__328_ vdd gnd FILL
XFILL_2__381_ vdd gnd FILL
XFILL_7__539_ vdd gnd FILL
XFILL_6__290_ vdd gnd FILL
XFILL_8__306_ vdd gnd FILL
X_585_ _585_/D _612_/CLK _585_/Q vdd gnd DFFPOSX1
XFILL_3__415_ vdd gnd FILL
XFILL_3__346_ vdd gnd FILL
XFILL_3__277_ vdd gnd FILL
XFILL_6__488_ vdd gnd FILL
XFILL_7__324_ vdd gnd FILL
XFILL_2__502_ vdd gnd FILL
XFILL_3_BUFX2_insert9 vdd gnd FILL
XFILL_2__433_ vdd gnd FILL
XFILL_2__295_ vdd gnd FILL
XFILL_2__364_ vdd gnd FILL
X_370_ _562_/Q _421_/B _371_/C vdd gnd NAND2X1
XFILL_6__411_ vdd gnd FILL
XFILL_9__553_ vdd gnd FILL
XFILL_6__273_ vdd gnd FILL
XFILL_6__342_ vdd gnd FILL
XFILL_9__484_ vdd gnd FILL
XFILL_1__520_ vdd gnd FILL
X_499_ _509_/A _499_/B _510_/C vdd gnd NAND2X1
XFILL_1__451_ vdd gnd FILL
X_568_ _568_/D _605_/CLK _568_/Q vdd gnd DFFPOSX1
XFILL_3__329_ vdd gnd FILL
XFILL_1__382_ vdd gnd FILL
XFILL_5__291_ vdd gnd FILL
XFILL_7__307_ vdd gnd FILL
XFILL_5__360_ vdd gnd FILL
XBUFX2_insert15 _557_/Q _430_/C vdd gnd BUFX2
XFILL_8_BUFX2_insert18 vdd gnd FILL
XFILL_2__416_ vdd gnd FILL
XFILL_2__278_ vdd gnd FILL
XFILL_3_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__347_ vdd gnd FILL
XFILL_5__489_ vdd gnd FILL
X_284_ _301_/A _452_/A _284_/C _618_/A vdd gnd OAI21X1
X_422_ _583_/Q _523_/A vdd gnd INVX1
X_353_ _490_/A _367_/A _357_/B _354_/A vdd gnd OAI21X1
XFILL_6__325_ vdd gnd FILL
XFILL_9__467_ vdd gnd FILL
XFILL_1__503_ vdd gnd FILL
XFILL_9__398_ vdd gnd FILL
XFILL_1__296_ vdd gnd FILL
XFILL_1__365_ vdd gnd FILL
XFILL_1__434_ vdd gnd FILL
XFILL_9_CLKBUF1_insert0 vdd gnd FILL
XFILL_5__412_ vdd gnd FILL
XFILL_8__623_ vdd gnd FILL
XFILL_5__274_ vdd gnd FILL
XFILL_5__343_ vdd gnd FILL
XFILL_8__485_ vdd gnd FILL
XFILL_8__554_ vdd gnd FILL
XFILL_0__521_ vdd gnd FILL
XFILL_0__452_ vdd gnd FILL
XFILL_0__383_ vdd gnd FILL
XFILL_9__321_ vdd gnd FILL
X_336_ _511_/C _490_/A vdd gnd INVX4
X_405_ _567_/Q _410_/A vdd gnd INVX1
XFILL_4_BUFX2_insert16 vdd gnd FILL
XFILL_4__292_ vdd gnd FILL
XFILL_6__308_ vdd gnd FILL
XFILL_4__361_ vdd gnd FILL
XFILL_4__430_ vdd gnd FILL
XFILL_9__519_ vdd gnd FILL
XFILL_1__417_ vdd gnd FILL
XFILL_1__279_ vdd gnd FILL
XFILL_1__348_ vdd gnd FILL
XFILL_5__326_ vdd gnd FILL
XFILL_8__468_ vdd gnd FILL
XFILL_8__537_ vdd gnd FILL
XFILL_0__504_ vdd gnd FILL
XFILL_8__399_ vdd gnd FILL
XFILL_0__297_ vdd gnd FILL
XFILL_0__435_ vdd gnd FILL
XFILL_0__366_ vdd gnd FILL
XFILL_9__304_ vdd gnd FILL
X_319_ _461_/B _538_/B _319_/C _600_/D vdd gnd OAI21X1
XFILL75150x46950 vdd gnd FILL
XFILL_7__624_ vdd gnd FILL
XFILL_4__275_ vdd gnd FILL
XFILL_4__413_ vdd gnd FILL
XFILL_4__344_ vdd gnd FILL
XFILL_7__486_ vdd gnd FILL
XFILL_7__555_ vdd gnd FILL
XFILL_0_BUFX2_insert25 vdd gnd FILL
XFILL_0_BUFX2_insert14 vdd gnd FILL
XFILL_8__322_ vdd gnd FILL
XFILL_3__500_ vdd gnd FILL
XFILL_3__362_ vdd gnd FILL
XFILL_3__431_ vdd gnd FILL
XFILL_3__293_ vdd gnd FILL
XFILL_5__309_ vdd gnd FILL
XFILL75750x25350 vdd gnd FILL
XFILL_7__340_ vdd gnd FILL
XFILL_7_BUFX2_insert20 vdd gnd FILL
XFILL_0__418_ vdd gnd FILL
XFILL_0__349_ vdd gnd FILL
XFILL_4__327_ vdd gnd FILL
XFILL_2__380_ vdd gnd FILL
XFILL_7__469_ vdd gnd FILL
XFILL_7__538_ vdd gnd FILL
XFILL_8__305_ vdd gnd FILL
XFILL_3__414_ vdd gnd FILL
XFILL_3__345_ vdd gnd FILL
X_584_ _584_/D _606_/CLK _584_/Q vdd gnd DFFPOSX1
XFILL_6__625_ vdd gnd FILL
XFILL_6__487_ vdd gnd FILL
XFILL_6__556_ vdd gnd FILL
XFILL_3__276_ vdd gnd FILL
XFILL_7__323_ vdd gnd FILL
XFILL_2__501_ vdd gnd FILL
XFILL_2__432_ vdd gnd FILL
XFILL_2__363_ vdd gnd FILL
XFILL_2__294_ vdd gnd FILL
XFILL_6__410_ vdd gnd FILL
XFILL_6__341_ vdd gnd FILL
XFILL_9__621_ vdd gnd FILL
XFILL_9__552_ vdd gnd FILL
X_567_ _567_/D _605_/CLK _567_/Q vdd gnd DFFPOSX1
XFILL_1__450_ vdd gnd FILL
X_498_ _594_/Q _548_/A vdd gnd INVX1
XFILL_3__328_ vdd gnd FILL
XFILL_1__381_ vdd gnd FILL
XFILL_6__539_ vdd gnd FILL
XFILL_5__290_ vdd gnd FILL
XFILL_7__306_ vdd gnd FILL
XBUFX2_insert16 _612_/Q _452_/B vdd gnd BUFX2
XFILL_8_BUFX2_insert19 vdd gnd FILL
XFILL_2__415_ vdd gnd FILL
XFILL_2__346_ vdd gnd FILL
XFILL_2__277_ vdd gnd FILL
XFILL_3_CLKBUF1_insert6 vdd gnd FILL
X_421_ _569_/Q _421_/B _434_/A vdd gnd NAND2X1
XFILL_5__488_ vdd gnd FILL
X_283_ _301_/A _561_/Q _284_/C vdd gnd NAND2X1
X_352_ _592_/Q _593_/Q _367_/A vdd gnd NOR2X1
XFILL_6__324_ vdd gnd FILL
XFILL_9__466_ vdd gnd FILL
XFILL_9__535_ vdd gnd FILL
XFILL_1__502_ vdd gnd FILL
X_619_ _619_/A Dout[4] vdd gnd BUFX2
XFILL_1__433_ vdd gnd FILL
XFILL_1__295_ vdd gnd FILL
XFILL_1__364_ vdd gnd FILL
XFILL_5__411_ vdd gnd FILL
XFILL_9_CLKBUF1_insert1 vdd gnd FILL
XFILL_5__342_ vdd gnd FILL
XFILL_8__622_ vdd gnd FILL
XFILL_8__553_ vdd gnd FILL
XFILL_5__273_ vdd gnd FILL
XFILL_8__484_ vdd gnd FILL
XFILL_0__520_ vdd gnd FILL
XFILL_9__320_ vdd gnd FILL
XFILL_0__451_ vdd gnd FILL
XFILL_2__329_ vdd gnd FILL
XFILL_0__382_ vdd gnd FILL
X_404_ _493_/B _404_/B _404_/C _566_/D vdd gnd OAI21X1
XFILL_4_BUFX2_insert17 vdd gnd FILL
X_335_ _607_/D _438_/C _335_/C _605_/D vdd gnd OAI21X1
XFILL_4__291_ vdd gnd FILL
XFILL_6__307_ vdd gnd FILL
XFILL_4__360_ vdd gnd FILL
XFILL_9__518_ vdd gnd FILL
XFILL_1__416_ vdd gnd FILL
XFILL_1__347_ vdd gnd FILL
XFILL_1__278_ vdd gnd FILL
XFILL_4__489_ vdd gnd FILL
XFILL_5__325_ vdd gnd FILL
XFILL_8__536_ vdd gnd FILL
XFILL_8__467_ vdd gnd FILL
XFILL_0__503_ vdd gnd FILL
XFILL_8__398_ vdd gnd FILL
XFILL_0__434_ vdd gnd FILL
XFILL_0__296_ vdd gnd FILL
XFILL_0__365_ vdd gnd FILL
X_318_ Yin[0] _538_/B _319_/C vdd gnd NAND2X1
XFILL_4__412_ vdd gnd FILL
XFILL_7__623_ vdd gnd FILL
XFILL_4__274_ vdd gnd FILL
XFILL_4__343_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
XFILL_7__485_ vdd gnd FILL
XFILL_7__554_ vdd gnd FILL
XFILL_8__321_ vdd gnd FILL
XFILL_3__292_ vdd gnd FILL
XFILL_5__308_ vdd gnd FILL
XFILL_3__361_ vdd gnd FILL
XFILL_3__430_ vdd gnd FILL
XFILL_8__519_ vdd gnd FILL
XFILL_0__417_ vdd gnd FILL
XFILL_7_BUFX2_insert10 vdd gnd FILL
XFILL_0__279_ vdd gnd FILL
XFILL_7_BUFX2_insert21 vdd gnd FILL
XFILL_0__348_ vdd gnd FILL
XFILL_4__326_ vdd gnd FILL
XFILL_7__537_ vdd gnd FILL
XFILL_7__468_ vdd gnd FILL
XFILL_7__399_ vdd gnd FILL
XFILL_8__304_ vdd gnd FILL
XFILL_0_BUFX2_insert7 vdd gnd FILL
X_583_ _583_/D _595_/CLK _583_/Q vdd gnd DFFPOSX1
XFILL_3__413_ vdd gnd FILL
XFILL_6__624_ vdd gnd FILL
XFILL_3__275_ vdd gnd FILL
XFILL_3__344_ vdd gnd FILL
XFILL_6__486_ vdd gnd FILL
XFILL_6__555_ vdd gnd FILL
XFILL_7__322_ vdd gnd FILL
XFILL_2__500_ vdd gnd FILL
XFILL_2__362_ vdd gnd FILL
XFILL_4__309_ vdd gnd FILL
XFILL_2__431_ vdd gnd FILL
XFILL_2__293_ vdd gnd FILL
XFILL_6__340_ vdd gnd FILL
XFILL_9__482_ vdd gnd FILL
XFILL_9__620_ vdd gnd FILL
XFILL_4_CLKBUF1_insert0 vdd gnd FILL
X_566_ _566_/D _581_/CLK _566_/Q vdd gnd DFFPOSX1
XFILL_1__380_ vdd gnd FILL
X_497_ _509_/A _594_/Q _499_/B _501_/B vdd gnd NAND3X1
XFILL_3__327_ vdd gnd FILL
XFILL_6__469_ vdd gnd FILL
XFILL_6__538_ vdd gnd FILL
XFILL_7__305_ vdd gnd FILL
XBUFX2_insert17 _612_/Q _439_/A vdd gnd BUFX2
XFILL_2__414_ vdd gnd FILL
XFILL_2__345_ vdd gnd FILL
XFILL_2__276_ vdd gnd FILL
XFILL_5__625_ vdd gnd FILL
XFILL_5__487_ vdd gnd FILL
XFILL_5__556_ vdd gnd FILL
X_420_ _420_/A _452_/B _420_/C _568_/D vdd gnd OAI21X1
X_351_ _357_/C _357_/B _354_/B vdd gnd OR2X2
X_282_ _573_/Q _452_/A vdd gnd INVX1
XFILL_6__323_ vdd gnd FILL
XFILL_9__465_ vdd gnd FILL
XFILL_9__534_ vdd gnd FILL
XFILL_1__501_ vdd gnd FILL
X_618_ _618_/A Dout[3] vdd gnd BUFX2
X_549_ Yin[1] _550_/B _550_/C vdd gnd NAND2X1
XFILL_1__432_ vdd gnd FILL
XFILL_1__363_ vdd gnd FILL
XFILL_9__396_ vdd gnd FILL
XFILL_1__294_ vdd gnd FILL
XFILL_9_CLKBUF1_insert2 vdd gnd FILL
XFILL74850x25350 vdd gnd FILL
XFILL_5__410_ vdd gnd FILL
XFILL_5__341_ vdd gnd FILL
XFILL_8__621_ vdd gnd FILL
XFILL_8__483_ vdd gnd FILL
XFILL_8__552_ vdd gnd FILL
XFILL_0__450_ vdd gnd FILL
XFILL_2__328_ vdd gnd FILL
XFILL_0__381_ vdd gnd FILL
X_403_ _566_/Q _503_/B _404_/C vdd gnd NAND2X1
XFILL_5__539_ vdd gnd FILL
X_334_ _607_/D Yin[1] _335_/C vdd gnd NAND2X1
XFILL_4_BUFX2_insert18 vdd gnd FILL
XFILL_4__290_ vdd gnd FILL
XFILL_6__306_ vdd gnd FILL
XFILL_9__448_ vdd gnd FILL
XFILL_9__379_ vdd gnd FILL
XFILL_1__415_ vdd gnd FILL
XFILL_1__346_ vdd gnd FILL
XFILL_4__488_ vdd gnd FILL
XFILL_1__277_ vdd gnd FILL
XFILL_5__324_ vdd gnd FILL
XFILL_8__466_ vdd gnd FILL
XFILL_8__535_ vdd gnd FILL
XFILL_0__502_ vdd gnd FILL
XFILL_8__397_ vdd gnd FILL
XFILL_0__433_ vdd gnd FILL
XFILL_9__302_ vdd gnd FILL
XFILL_0__295_ vdd gnd FILL
XFILL_0__364_ vdd gnd FILL
X_317_ _317_/A _317_/B _538_/B vdd gnd NOR2X1
XFILL_4__411_ vdd gnd FILL
XFILL_4__342_ vdd gnd FILL
XFILL_7__622_ vdd gnd FILL
XFILL_7__553_ vdd gnd FILL
XFILL_4__273_ vdd gnd FILL
XFILL_0_BUFX2_insert16 vdd gnd FILL
XFILL_7__484_ vdd gnd FILL
XFILL_8__320_ vdd gnd FILL
XFILL_1__329_ vdd gnd FILL
XFILL_3__291_ vdd gnd FILL
XFILL_5__307_ vdd gnd FILL
XFILL_3__360_ vdd gnd FILL
XFILL_8__449_ vdd gnd FILL
XFILL_8__518_ vdd gnd FILL
XFILL_7_BUFX2_insert11 vdd gnd FILL
XFILL_7_BUFX2_insert22 vdd gnd FILL
XFILL_0__416_ vdd gnd FILL
XFILL_0__347_ vdd gnd FILL
XFILL_0__278_ vdd gnd FILL
XFILL_3__489_ vdd gnd FILL
XFILL_4__325_ vdd gnd FILL
XFILL_7__467_ vdd gnd FILL
XFILL_7__536_ vdd gnd FILL
XFILL_7__398_ vdd gnd FILL
XFILL_8__303_ vdd gnd FILL
XFILL_0_BUFX2_insert8 vdd gnd FILL
XFILL_3__412_ vdd gnd FILL
X_582_ _582_/D _595_/CLK _582_/Q vdd gnd DFFPOSX1
XFILL_6__623_ vdd gnd FILL
XFILL_6__554_ vdd gnd FILL
XFILL_3__274_ vdd gnd FILL
XFILL_3__343_ vdd gnd FILL
XFILL_6__485_ vdd gnd FILL
XFILL75450x50550 vdd gnd FILL
XFILL_7__321_ vdd gnd FILL
XFILL_3_BUFX2_insert20 vdd gnd FILL
XFILL_2__430_ vdd gnd FILL
XFILL_2__292_ vdd gnd FILL
XFILL_4__308_ vdd gnd FILL
XFILL_2__361_ vdd gnd FILL
XFILL_7__519_ vdd gnd FILL
XFILL_9__481_ vdd gnd FILL
XFILL_9__550_ vdd gnd FILL
XFILL_4_CLKBUF1_insert1 vdd gnd FILL
X_496_ _496_/A _496_/B _496_/C _499_/B vdd gnd NAND3X1
XFILL_3__326_ vdd gnd FILL
X_565_ _565_/D _573_/CLK _565_/Q vdd gnd DFFPOSX1
XFILL_6__537_ vdd gnd FILL
XFILL_6__468_ vdd gnd FILL
XFILL_6__399_ vdd gnd FILL
XFILL_7__304_ vdd gnd FILL
XBUFX2_insert18 _612_/Q _625_/A vdd gnd BUFX2
XFILL_2__413_ vdd gnd FILL
XFILL_5__624_ vdd gnd FILL
XFILL_2__275_ vdd gnd FILL
XFILL_2__344_ vdd gnd FILL
XFILL_5__486_ vdd gnd FILL
XFILL_5__555_ vdd gnd FILL
X_350_ _592_/Q _593_/Q _415_/A _357_/C vdd gnd OAI21X1
X_281_ _286_/A _447_/A _281_/C _617_/A vdd gnd OAI21X1
XFILL_6__322_ vdd gnd FILL
XFILL_9__533_ vdd gnd FILL
XFILL_1__500_ vdd gnd FILL
X_617_ _617_/A Dout[2] vdd gnd BUFX2
XFILL_9__395_ vdd gnd FILL
X_479_ _479_/A _625_/A _479_/C _577_/D vdd gnd OAI21X1
XFILL_1__293_ vdd gnd FILL
X_548_ _548_/A _550_/B _548_/C _594_/D vdd gnd OAI21X1
XFILL_1__362_ vdd gnd FILL
XFILL_3__309_ vdd gnd FILL
XFILL_1__431_ vdd gnd FILL
XFILL75150x72150 vdd gnd FILL
XFILL_8__620_ vdd gnd FILL
XFILL_5__340_ vdd gnd FILL
XFILL_8__482_ vdd gnd FILL
XFILL_8__551_ vdd gnd FILL
XFILL_0__380_ vdd gnd FILL
XFILL_2__327_ vdd gnd FILL
XFILL_5__538_ vdd gnd FILL
XFILL_4_BUFX2_insert19 vdd gnd FILL
XFILL_5__469_ vdd gnd FILL
X_402_ _402_/A _402_/B _404_/B vdd gnd NAND2X1
X_333_ _605_/Q _438_/C vdd gnd INVX1
XFILL_6__305_ vdd gnd FILL
XFILL_9__516_ vdd gnd FILL
XFILL_9__447_ vdd gnd FILL
XFILL_4__625_ vdd gnd FILL
XFILL_8_BUFX2_insert7 vdd gnd FILL
XFILL_1__414_ vdd gnd FILL
XFILL_1__345_ vdd gnd FILL
XFILL_1__276_ vdd gnd FILL
XFILL_4__487_ vdd gnd FILL
XFILL_4__556_ vdd gnd FILL
XFILL_5__323_ vdd gnd FILL
XFILL_0__501_ vdd gnd FILL
XFILL_8__465_ vdd gnd FILL
XFILL_8__534_ vdd gnd FILL
XFILL_8__396_ vdd gnd FILL
XFILL_0__432_ vdd gnd FILL
XFILL_0__363_ vdd gnd FILL
XFILL_0__294_ vdd gnd FILL
XFILL_9__301_ vdd gnd FILL
X_316_ _517_/A _317_/B vdd gnd INVX1
XFILL_4__410_ vdd gnd FILL
XFILL_4__341_ vdd gnd FILL
XFILL_7__621_ vdd gnd FILL
XFILL_7__483_ vdd gnd FILL
XFILL_7__552_ vdd gnd FILL
XFILL_0_BUFX2_insert17 vdd gnd FILL
XFILL_1__328_ vdd gnd FILL
XFILL_4__539_ vdd gnd FILL
XFILL_3__290_ vdd gnd FILL
XFILL_5__306_ vdd gnd FILL
XFILL_8__448_ vdd gnd FILL
XFILL_8__379_ vdd gnd FILL
XFILL_8__517_ vdd gnd FILL
XFILL_0__277_ vdd gnd FILL
XFILL_7_BUFX2_insert12 vdd gnd FILL
XFILL_7_BUFX2_insert23 vdd gnd FILL
XFILL_0__415_ vdd gnd FILL
XFILL_0__346_ vdd gnd FILL
XFILL_3__488_ vdd gnd FILL
XFILL_4__324_ vdd gnd FILL
XFILL_7__466_ vdd gnd FILL
XFILL_7__535_ vdd gnd FILL
XFILL_7__397_ vdd gnd FILL
XFILL_8__302_ vdd gnd FILL
XFILL_0_BUFX2_insert9 vdd gnd FILL
X_581_ _581_/D _581_/CLK _581_/Q vdd gnd DFFPOSX1
XFILL_3__411_ vdd gnd FILL
XFILL_3__342_ vdd gnd FILL
XFILL_6__622_ vdd gnd FILL
XFILL_6__553_ vdd gnd FILL
XFILL_3__273_ vdd gnd FILL
XFILL_6__484_ vdd gnd FILL
XFILL_7__320_ vdd gnd FILL
XFILL_0__329_ vdd gnd FILL
XFILL_3_BUFX2_insert10 vdd gnd FILL
XFILL_3_BUFX2_insert21 vdd gnd FILL
XFILL_2__291_ vdd gnd FILL
XFILL_4__307_ vdd gnd FILL
XFILL_2__360_ vdd gnd FILL
XFILL_7__449_ vdd gnd FILL
XFILL_7__518_ vdd gnd FILL
XFILL_2__489_ vdd gnd FILL
XFILL_9__480_ vdd gnd FILL
XFILL_4_CLKBUF1_insert2 vdd gnd FILL
X_495_ _596_/Q _597_/Q _496_/A vdd gnd NOR2X1
X_564_ _564_/D _606_/CLK _564_/Q vdd gnd DFFPOSX1
XFILL_3__325_ vdd gnd FILL
XFILL_6__467_ vdd gnd FILL
XFILL_6__536_ vdd gnd FILL
XFILL_6__398_ vdd gnd FILL
XFILL_7__303_ vdd gnd FILL
XBUFX2_insert19 _612_/Q _478_/A vdd gnd BUFX2
XFILL_2__412_ vdd gnd FILL
XFILL_2__343_ vdd gnd FILL
XFILL_5__623_ vdd gnd FILL
XFILL_5__554_ vdd gnd FILL
XFILL_2__274_ vdd gnd FILL
XFILL_5__485_ vdd gnd FILL
X_280_ _286_/A _560_/Q _281_/C vdd gnd NAND2X1
XFILL_6__321_ vdd gnd FILL
X_616_ _616_/A Dout[11] vdd gnd BUFX2
XFILL_9__463_ vdd gnd FILL
X_547_ Yin[0] _550_/B _548_/C vdd gnd NAND2X1
XFILL_1__430_ vdd gnd FILL
XFILL_9__394_ vdd gnd FILL
X_478_ _478_/A _478_/B _478_/C _479_/C vdd gnd NAND3X1
XFILL_1__292_ vdd gnd FILL
XFILL_3__308_ vdd gnd FILL
XFILL_1__361_ vdd gnd FILL
XFILL_6__519_ vdd gnd FILL
XFILL_9_CLKBUF1_insert4 vdd gnd FILL
XFILL_8__550_ vdd gnd FILL
XFILL_8__481_ vdd gnd FILL
XFILL_2__326_ vdd gnd FILL
XFILL_5__537_ vdd gnd FILL
X_401_ _407_/B _431_/C _402_/A vdd gnd NAND2X1
XFILL_5__468_ vdd gnd FILL
XFILL_5__399_ vdd gnd FILL
X_332_ _607_/D _438_/A _332_/C _604_/D vdd gnd OAI21X1
XFILL_6__304_ vdd gnd FILL
XFILL_9__515_ vdd gnd FILL
XFILL_9__377_ vdd gnd FILL
XFILL_1__413_ vdd gnd FILL
XFILL_4__624_ vdd gnd FILL
XFILL_8_BUFX2_insert8 vdd gnd FILL
XFILL_4__555_ vdd gnd FILL
XFILL_1__275_ vdd gnd FILL
XFILL_1__344_ vdd gnd FILL
XFILL_4__486_ vdd gnd FILL
XFILL_5__322_ vdd gnd FILL
XFILL_8__533_ vdd gnd FILL
XFILL_0__500_ vdd gnd FILL
XFILL_8__464_ vdd gnd FILL
XFILL_8__395_ vdd gnd FILL
XFILL_9__300_ vdd gnd FILL
XFILL_0__293_ vdd gnd FILL
XFILL_0__362_ vdd gnd FILL
XFILL_2__309_ vdd gnd FILL
XFILL_0__431_ vdd gnd FILL
X_315_ _600_/Q _461_/B vdd gnd INVX1
XFILL_7__620_ vdd gnd FILL
XFILL_4__340_ vdd gnd FILL
XFILL_0_BUFX2_insert18 vdd gnd FILL
XFILL_7__482_ vdd gnd FILL
XFILL_7__551_ vdd gnd FILL
XFILL_9__429_ vdd gnd FILL
XFILL_1__327_ vdd gnd FILL
XFILL_4__538_ vdd gnd FILL
XFILL_4__469_ vdd gnd FILL
XFILL_5__305_ vdd gnd FILL
XFILL_8__516_ vdd gnd FILL
XFILL_8__447_ vdd gnd FILL
XFILL_0__414_ vdd gnd FILL
XFILL_8__378_ vdd gnd FILL
XFILL_3__625_ vdd gnd FILL
XFILL_7_BUFX2_insert24 vdd gnd FILL
XFILL_0__345_ vdd gnd FILL
XFILL_7_BUFX2_insert13 vdd gnd FILL
XFILL_0__276_ vdd gnd FILL
XFILL_3__487_ vdd gnd FILL
XFILL_3__556_ vdd gnd FILL
XFILL75450x10950 vdd gnd FILL
XFILL_4__323_ vdd gnd FILL
XFILL_7__465_ vdd gnd FILL
XFILL_7__534_ vdd gnd FILL
XFILL_7__396_ vdd gnd FILL
XFILL74250x72150 vdd gnd FILL
XFILL_8__301_ vdd gnd FILL
X_580_ _580_/D _581_/CLK _580_/Q vdd gnd DFFPOSX1
XFILL_6__621_ vdd gnd FILL
XFILL_3__410_ vdd gnd FILL
XFILL_3__341_ vdd gnd FILL
XFILL_6__483_ vdd gnd FILL
XFILL_6__552_ vdd gnd FILL
XFILL_0__328_ vdd gnd FILL
XFILL75150x57750 vdd gnd FILL
XFILL_3__539_ vdd gnd FILL
XFILL_3_BUFX2_insert11 vdd gnd FILL
XFILL_3_BUFX2_insert22 vdd gnd FILL
XFILL_2__290_ vdd gnd FILL
XFILL_4__306_ vdd gnd FILL
XFILL_7__517_ vdd gnd FILL
XFILL_7__448_ vdd gnd FILL
XFILL_7__379_ vdd gnd FILL
XFILL_2__488_ vdd gnd FILL
XFILL_4_CLKBUF1_insert3 vdd gnd FILL
X_563_ _563_/D _573_/CLK _563_/Q vdd gnd DFFPOSX1
X_494_ _494_/A _494_/B _496_/C vdd gnd AND2X2
XFILL_3__324_ vdd gnd FILL
XFILL_6__466_ vdd gnd FILL
XFILL75750x36150 vdd gnd FILL
XFILL_6__397_ vdd gnd FILL
XFILL_6__535_ vdd gnd FILL
XFILL_7__302_ vdd gnd FILL
XFILL_2__411_ vdd gnd FILL
XFILL_2__342_ vdd gnd FILL
XFILL_5__484_ vdd gnd FILL
XFILL_5__622_ vdd gnd FILL
XFILL_5__553_ vdd gnd FILL
XFILL_2__273_ vdd gnd FILL
XFILL_6__320_ vdd gnd FILL
XFILL_9__462_ vdd gnd FILL
XFILL_9__531_ vdd gnd FILL
X_615_ _615_/A Dout[10] vdd gnd BUFX2
X_546_ _607_/D _546_/B _546_/C _593_/D vdd gnd OAI21X1
XFILL_1__360_ vdd gnd FILL
XFILL_1__291_ vdd gnd FILL
X_477_ _477_/A _477_/B _477_/C _478_/C vdd gnd NAND3X1
XFILL_3__307_ vdd gnd FILL
XFILL_6__449_ vdd gnd FILL
XFILL_6__518_ vdd gnd FILL
XFILL_9_CLKBUF1_insert5 vdd gnd FILL
XFILL_1__489_ vdd gnd FILL
XFILL_8__480_ vdd gnd FILL
XFILL_2__325_ vdd gnd FILL
XFILL_5__467_ vdd gnd FILL
XFILL_5__536_ vdd gnd FILL
X_400_ _431_/C _407_/B _402_/B vdd gnd OR2X2
X_331_ _607_/D Yin[0] _332_/C vdd gnd NAND2X1
XFILL_5__398_ vdd gnd FILL
XFILL_6__303_ vdd gnd FILL
XFILL_9__514_ vdd gnd FILL
XFILL_9__445_ vdd gnd FILL
XFILL_1__412_ vdd gnd FILL
X_529_ _585_/Q _554_/B _530_/C vdd gnd NAND2X1
XFILL_9__376_ vdd gnd FILL
XFILL_1__343_ vdd gnd FILL
XFILL_4__623_ vdd gnd FILL
XFILL_8_BUFX2_insert9 vdd gnd FILL
XFILL_4__554_ vdd gnd FILL
XFILL_1__274_ vdd gnd FILL
XFILL_4__485_ vdd gnd FILL
XFILL_5__321_ vdd gnd FILL
XFILL_8__463_ vdd gnd FILL
XFILL_8__532_ vdd gnd FILL
XFILL_0__430_ vdd gnd FILL
XFILL_8__394_ vdd gnd FILL
XFILL_0__292_ vdd gnd FILL
XFILL_2__308_ vdd gnd FILL
XFILL_0__361_ vdd gnd FILL
X_314_ _554_/A _556_/B _314_/C _599_/D vdd gnd OAI21X1
XFILL_5__519_ vdd gnd FILL
XFILL_7__550_ vdd gnd FILL
XFILL_0_BUFX2_insert19 vdd gnd FILL
XFILL_7__481_ vdd gnd FILL
XFILL_9__428_ vdd gnd FILL
XFILL_1__326_ vdd gnd FILL
XFILL_4__468_ vdd gnd FILL
XFILL_4__537_ vdd gnd FILL
XFILL_4__399_ vdd gnd FILL
XFILL_5__304_ vdd gnd FILL
XFILL_8__515_ vdd gnd FILL
XFILL_8__446_ vdd gnd FILL
XFILL_8__377_ vdd gnd FILL
XFILL_0__413_ vdd gnd FILL
XFILL_3__624_ vdd gnd FILL
XFILL_3__555_ vdd gnd FILL
XFILL_7_BUFX2_insert25 vdd gnd FILL
XFILL_0__275_ vdd gnd FILL
XFILL_0__344_ vdd gnd FILL
XFILL_7_BUFX2_insert14 vdd gnd FILL
XFILL_3__486_ vdd gnd FILL
XFILL_4__322_ vdd gnd FILL
XFILL_7__533_ vdd gnd FILL
XFILL_7__464_ vdd gnd FILL
XFILL_7__395_ vdd gnd FILL
XFILL_8__300_ vdd gnd FILL
XFILL_1__309_ vdd gnd FILL
XFILL_6__620_ vdd gnd FILL
XFILL_3__340_ vdd gnd FILL
XFILL73050x28950 vdd gnd FILL
XFILL_6__482_ vdd gnd FILL
XFILL_6__551_ vdd gnd FILL
XFILL_8__429_ vdd gnd FILL
XFILL_0__327_ vdd gnd FILL
XFILL_3__538_ vdd gnd FILL
XFILL_3_BUFX2_insert12 vdd gnd FILL
XFILL_3__469_ vdd gnd FILL
XFILL_4__305_ vdd gnd FILL
XFILL_3_BUFX2_insert23 vdd gnd FILL
XFILL_7__516_ vdd gnd FILL
XFILL_7__447_ vdd gnd FILL
XFILL_7__378_ vdd gnd FILL
XFILL_2__625_ vdd gnd FILL
XFILL_2__487_ vdd gnd FILL
XFILL_2__556_ vdd gnd FILL
XFILL_4_CLKBUF1_insert4 vdd gnd FILL
X_493_ _493_/A _493_/B _493_/C _493_/D _579_/D vdd gnd AOI22X1
X_562_ _562_/D _573_/CLK _562_/Q vdd gnd DFFPOSX1
XFILL_3__323_ vdd gnd FILL
XFILL_6__534_ vdd gnd FILL
XFILL_6__465_ vdd gnd FILL
XFILL_6__396_ vdd gnd FILL
XFILL_7__301_ vdd gnd FILL
XFILL_5__621_ vdd gnd FILL
XFILL_2__410_ vdd gnd FILL
XFILL_2__341_ vdd gnd FILL
XFILL_5__483_ vdd gnd FILL
XFILL_5__552_ vdd gnd FILL
XFILL_2__539_ vdd gnd FILL
XFILL_9__530_ vdd gnd FILL
XFILL_9__392_ vdd gnd FILL
X_476_ _511_/C _598_/Q _477_/B vdd gnd NAND2X1
XFILL_3__306_ vdd gnd FILL
X_614_ _614_/A Dout[1] vdd gnd BUFX2
X_545_ _607_/D Xin[1] _546_/C vdd gnd NAND2X1
XFILL_1__290_ vdd gnd FILL
XFILL_6__517_ vdd gnd FILL
XFILL_6__448_ vdd gnd FILL
XFILL_9_CLKBUF1_insert6 vdd gnd FILL
XFILL_6__379_ vdd gnd FILL
XFILL74550x10950 vdd gnd FILL
XFILL_1__488_ vdd gnd FILL
XFILL_2__324_ vdd gnd FILL
XFILL_5__466_ vdd gnd FILL
XFILL_5__397_ vdd gnd FILL
XFILL_5__535_ vdd gnd FILL
X_330_ _604_/Q _438_/A vdd gnd INVX1
XFILL73350x72150 vdd gnd FILL
XFILL_6__302_ vdd gnd FILL
XFILL_9__444_ vdd gnd FILL
XFILL_9__375_ vdd gnd FILL
X_459_ _460_/B _459_/B _459_/C _460_/C vdd gnd NAND3X1
XFILL_1__273_ vdd gnd FILL
XFILL_1__411_ vdd gnd FILL
X_528_ Xin[1] _542_/A vdd gnd INVX1
XFILL_1__342_ vdd gnd FILL
XFILL_4__484_ vdd gnd FILL
XFILL_4__622_ vdd gnd FILL
XFILL_4__553_ vdd gnd FILL
XFILL74250x57750 vdd gnd FILL
XFILL_5__320_ vdd gnd FILL
XFILL_8__462_ vdd gnd FILL
XFILL_8__531_ vdd gnd FILL
XFILL_8__393_ vdd gnd FILL
XFILL_0__360_ vdd gnd FILL
XFILL_0__291_ vdd gnd FILL
XFILL_2__307_ vdd gnd FILL
X_313_ _599_/Q _556_/B _314_/C vdd gnd NAND2X1
XFILL_5__449_ vdd gnd FILL
XFILL_5__518_ vdd gnd FILL
XFILL_0__489_ vdd gnd FILL
XFILL_7__480_ vdd gnd FILL
XFILL_9__289_ vdd gnd FILL
XFILL_9__358_ vdd gnd FILL
XFILL_1__325_ vdd gnd FILL
XFILL_4__467_ vdd gnd FILL
XFILL74850x36150 vdd gnd FILL
XFILL_4__536_ vdd gnd FILL
XFILL_4__398_ vdd gnd FILL
XFILL_5__303_ vdd gnd FILL
XFILL_8__514_ vdd gnd FILL
XFILL_8__445_ vdd gnd FILL
XFILL_8__376_ vdd gnd FILL
XFILL_0__412_ vdd gnd FILL
XFILL_0__343_ vdd gnd FILL
XFILL_3__485_ vdd gnd FILL
XFILL_3__623_ vdd gnd FILL
XFILL_3__554_ vdd gnd FILL
XFILL_0__274_ vdd gnd FILL
XFILL_7_BUFX2_insert15 vdd gnd FILL
XFILL_4__321_ vdd gnd FILL
XFILL_7__463_ vdd gnd FILL
XFILL_7__532_ vdd gnd FILL
XFILL_7__394_ vdd gnd FILL
XFILL_1__308_ vdd gnd FILL
XFILL_4__519_ vdd gnd FILL
XFILL_6__550_ vdd gnd FILL
XFILL_6__481_ vdd gnd FILL
XFILL_8__428_ vdd gnd FILL
XFILL_8__359_ vdd gnd FILL
XFILL_0__326_ vdd gnd FILL
XFILL_3__468_ vdd gnd FILL
XFILL_3__537_ vdd gnd FILL
XFILL_3_BUFX2_insert24 vdd gnd FILL
XFILL_3__399_ vdd gnd FILL
XFILL_3_BUFX2_insert13 vdd gnd FILL
XFILL_4__304_ vdd gnd FILL
XFILL_7__515_ vdd gnd FILL
XFILL_7__446_ vdd gnd FILL
XFILL_7__377_ vdd gnd FILL
XFILL_2__624_ vdd gnd FILL
XFILL_2__555_ vdd gnd FILL
XFILL_2__486_ vdd gnd FILL
XFILL_4_CLKBUF1_insert5 vdd gnd FILL
X_492_ _492_/A _492_/B _493_/B _493_/D vdd gnd AOI21X1
XFILL_3__322_ vdd gnd FILL
X_561_ _561_/D _605_/CLK _561_/Q vdd gnd DFFPOSX1
XFILL_6__533_ vdd gnd FILL
XFILL_6__464_ vdd gnd FILL
XFILL_6__395_ vdd gnd FILL
XFILL_7__300_ vdd gnd FILL
XFILL_0__309_ vdd gnd FILL
XFILL_5__620_ vdd gnd FILL
XFILL_5__551_ vdd gnd FILL
XFILL_2__340_ vdd gnd FILL
XFILL_5__482_ vdd gnd FILL
XFILL_7__429_ vdd gnd FILL
XFILL_2__538_ vdd gnd FILL
XFILL_2__469_ vdd gnd FILL
XFILL_9__460_ vdd gnd FILL
X_613_ _613_/A Dout[0] vdd gnd BUFX2
XFILL_9__391_ vdd gnd FILL
XFILL_3__305_ vdd gnd FILL
X_475_ _599_/Q _477_/A vdd gnd INVX1
X_544_ _607_/D _544_/B _544_/C _592_/D vdd gnd OAI21X1
XFILL_6__447_ vdd gnd FILL
XFILL_6__516_ vdd gnd FILL
XFILL75450x61350 vdd gnd FILL
XFILL_6__378_ vdd gnd FILL
XFILL_1__625_ vdd gnd FILL
XFILL_1__556_ vdd gnd FILL
XFILL_1__487_ vdd gnd FILL
XFILL_2__323_ vdd gnd FILL
XFILL_5_BUFX2_insert7 vdd gnd FILL
XFILL_5__534_ vdd gnd FILL
XFILL_5__465_ vdd gnd FILL
XFILL_5__396_ vdd gnd FILL
XFILL_6__301_ vdd gnd FILL
XFILL_9__512_ vdd gnd FILL
XFILL_9__443_ vdd gnd FILL
XFILL_1__410_ vdd gnd FILL
X_527_ _540_/A _554_/B _527_/C _584_/D vdd gnd OAI21X1
XFILL_4__621_ vdd gnd FILL
X_458_ _490_/A _496_/B _461_/B _459_/B vdd gnd OAI21X1
X_389_ _389_/A _412_/A _414_/B _390_/C vdd gnd NAND3X1
XFILL_1__341_ vdd gnd FILL
XFILL_4__483_ vdd gnd FILL
XFILL_4__552_ vdd gnd FILL
XFILL_1__539_ vdd gnd FILL
XFILL_8__461_ vdd gnd FILL
XFILL_8__530_ vdd gnd FILL
XFILL_8__392_ vdd gnd FILL
XFILL_0__290_ vdd gnd FILL
XFILL_2__306_ vdd gnd FILL
XFILL_5__517_ vdd gnd FILL
XFILL_5__448_ vdd gnd FILL
XFILL_5__379_ vdd gnd FILL
X_312_ _317_/A _610_/D _517_/A _556_/B vdd gnd NAND3X1
XFILL_0__488_ vdd gnd FILL
XFILL_9__426_ vdd gnd FILL
XFILL_9__357_ vdd gnd FILL
XFILL_1__324_ vdd gnd FILL
XFILL_4__466_ vdd gnd FILL
XFILL_4__397_ vdd gnd FILL
XFILL_4__535_ vdd gnd FILL
XFILL_5__302_ vdd gnd FILL
XFILL_8__513_ vdd gnd FILL
XFILL_8__444_ vdd gnd FILL
XFILL75450x7350 vdd gnd FILL
XFILL_8__375_ vdd gnd FILL
XFILL_3__622_ vdd gnd FILL
XFILL_0__273_ vdd gnd FILL
XFILL_7_BUFX2_insert16 vdd gnd FILL
XFILL_0__411_ vdd gnd FILL
XFILL_0__342_ vdd gnd FILL
XFILL_3__484_ vdd gnd FILL
XFILL_3__553_ vdd gnd FILL
XFILL_4__320_ vdd gnd FILL
XFILL_7__462_ vdd gnd FILL
XFILL_9__409_ vdd gnd FILL
XFILL_7__531_ vdd gnd FILL
XFILL_7__393_ vdd gnd FILL
XFILL_1__307_ vdd gnd FILL
XFILL_4__518_ vdd gnd FILL
XFILL_4__449_ vdd gnd FILL
XFILL73650x10950 vdd gnd FILL
XFILL_6__480_ vdd gnd FILL
XFILL_8__289_ vdd gnd FILL
XFILL_8__427_ vdd gnd FILL
XFILL_8__358_ vdd gnd FILL
XFILL_0__325_ vdd gnd FILL
XFILL_3__467_ vdd gnd FILL
XFILL_3__398_ vdd gnd FILL
XFILL_3__536_ vdd gnd FILL
XFILL_3_BUFX2_insert25 vdd gnd FILL
XFILL_3_BUFX2_insert14 vdd gnd FILL
XFILL_4__303_ vdd gnd FILL
XFILL_7__514_ vdd gnd FILL
XFILL_7__445_ vdd gnd FILL
XFILL_7__376_ vdd gnd FILL
XFILL_2__485_ vdd gnd FILL
XFILL_2__623_ vdd gnd FILL
XFILL_2__554_ vdd gnd FILL
XFILL_4_CLKBUF1_insert6 vdd gnd FILL
X_560_ _560_/D _573_/CLK _560_/Q vdd gnd DFFPOSX1
X_491_ _492_/A _492_/B _493_/C vdd gnd OR2X2
XFILL73350x57750 vdd gnd FILL
XFILL_3__321_ vdd gnd FILL
XFILL_6__463_ vdd gnd FILL
XFILL_6__532_ vdd gnd FILL
XFILL_6__394_ vdd gnd FILL
XFILL_0__308_ vdd gnd FILL
XFILL_3__519_ vdd gnd FILL
XFILL_5__550_ vdd gnd FILL
XFILL_5__481_ vdd gnd FILL
XFILL_7__428_ vdd gnd FILL
XFILL_7__359_ vdd gnd FILL
XFILL_2__468_ vdd gnd FILL
XFILL_2__537_ vdd gnd FILL
X_612_ _612_/D _612_/CLK _612_/Q vdd gnd DFFPOSX1
XFILL_2__399_ vdd gnd FILL
X_543_ _607_/D Xin[0] _544_/C vdd gnd NAND2X1
XFILL_9__390_ vdd gnd FILL
X_474_ _511_/C _599_/Q _474_/C _478_/B vdd gnd NAND3X1
XFILL_3__304_ vdd gnd FILL
XFILL_6__515_ vdd gnd FILL
XFILL_6__446_ vdd gnd FILL
XFILL_6__377_ vdd gnd FILL
XFILL_1__624_ vdd gnd FILL
XFILL_1__555_ vdd gnd FILL
XFILL_1__486_ vdd gnd FILL
XFILL_2__322_ vdd gnd FILL
XFILL_5_BUFX2_insert8 vdd gnd FILL
XFILL_5__464_ vdd gnd FILL
XFILL_5__533_ vdd gnd FILL
XFILL_5__395_ vdd gnd FILL
XFILL_6__300_ vdd gnd FILL
XFILL_9__511_ vdd gnd FILL
XFILL_1__340_ vdd gnd FILL
XFILL_9__373_ vdd gnd FILL
X_526_ _584_/Q _554_/B _527_/C vdd gnd NAND2X1
XFILL_4__620_ vdd gnd FILL
XFILL_4__551_ vdd gnd FILL
X_457_ _457_/A _457_/B _496_/B vdd gnd AND2X2
X_388_ _565_/Q _395_/A vdd gnd INVX1
XFILL_4__482_ vdd gnd FILL
XFILL_6__429_ vdd gnd FILL
XFILL_1__469_ vdd gnd FILL
XFILL_1__538_ vdd gnd FILL
XFILL_8__460_ vdd gnd FILL
XFILL_8__391_ vdd gnd FILL
XFILL_2__305_ vdd gnd FILL
XFILL_5__447_ vdd gnd FILL
XFILL_5__516_ vdd gnd FILL
X_311_ _607_/D _608_/D _517_/A vdd gnd NOR2X1
XFILL_5__378_ vdd gnd FILL
XFILL_0__625_ vdd gnd FILL
XFILL_0__556_ vdd gnd FILL
XFILL_0__487_ vdd gnd FILL
XFILL_9__425_ vdd gnd FILL
X_509_ _509_/A _594_/Q _512_/B vdd gnd NAND2X1
XFILL_9__287_ vdd gnd FILL
XFILL_1__323_ vdd gnd FILL
XFILL_9__356_ vdd gnd FILL
XFILL_4__534_ vdd gnd FILL
XFILL_4__465_ vdd gnd FILL
XFILL_4__396_ vdd gnd FILL
XFILL_5__301_ vdd gnd FILL
XFILL_8__512_ vdd gnd FILL
XFILL_8__443_ vdd gnd FILL
XFILL_0__410_ vdd gnd FILL
XFILL_8__374_ vdd gnd FILL
XFILL_3__621_ vdd gnd FILL
XFILL_7_BUFX2_insert17 vdd gnd FILL
XFILL_0__341_ vdd gnd FILL
XFILL_3__483_ vdd gnd FILL
XFILL_3__552_ vdd gnd FILL
XFILL_7__530_ vdd gnd FILL
XFILL_0__539_ vdd gnd FILL
XFILL_7__461_ vdd gnd FILL
XFILL_7__392_ vdd gnd FILL
XFILL_9__339_ vdd gnd FILL
XFILL_1__306_ vdd gnd FILL
XFILL_4__448_ vdd gnd FILL
XFILL_4__517_ vdd gnd FILL
XFILL_4__379_ vdd gnd FILL
XFILL_8__426_ vdd gnd FILL
XFILL_8__288_ vdd gnd FILL
XFILL_5_CLKBUF1_insert0 vdd gnd FILL
XFILL_8__357_ vdd gnd FILL
XFILL_3__535_ vdd gnd FILL
XFILL_0__324_ vdd gnd FILL
XFILL_3__466_ vdd gnd FILL
XFILL_3__397_ vdd gnd FILL
XFILL_4__302_ vdd gnd FILL
XFILL75450x46950 vdd gnd FILL
XFILL_3_BUFX2_insert15 vdd gnd FILL
XFILL_7__513_ vdd gnd FILL
XFILL_7__444_ vdd gnd FILL
XFILL_7__375_ vdd gnd FILL
XFILL_2__622_ vdd gnd FILL
XFILL_2__484_ vdd gnd FILL
XFILL_2__553_ vdd gnd FILL
X_490_ _490_/A _490_/B _512_/C _492_/A vdd gnd OAI21X1
XFILL_3__320_ vdd gnd FILL
XFILL_6__462_ vdd gnd FILL
XFILL_8__409_ vdd gnd FILL
XFILL_6__531_ vdd gnd FILL
XFILL_6__393_ vdd gnd FILL
XFILL_0__307_ vdd gnd FILL
XFILL_3__518_ vdd gnd FILL
XFILL_3__449_ vdd gnd FILL
XFILL_5__480_ vdd gnd FILL
XFILL_7__289_ vdd gnd FILL
XFILL_7__427_ vdd gnd FILL
XFILL_7__358_ vdd gnd FILL
XFILL_2__467_ vdd gnd FILL
XFILL_2__398_ vdd gnd FILL
XFILL_2__536_ vdd gnd FILL
X_473_ _473_/A _494_/A _496_/B _474_/C vdd gnd NAND3X1
X_611_ _611_/D _612_/CLK _612_/D vdd gnd DFFPOSX1
X_542_ _542_/A _542_/B _542_/C _591_/D vdd gnd OAI21X1
XFILL_3__303_ vdd gnd FILL
XFILL_6__514_ vdd gnd FILL
XFILL_6__445_ vdd gnd FILL
XFILL_6__376_ vdd gnd FILL
XFILL_1__485_ vdd gnd FILL
XFILL_1__623_ vdd gnd FILL
XFILL_1__554_ vdd gnd FILL
XFILL_2__321_ vdd gnd FILL
XFILL_5_BUFX2_insert9 vdd gnd FILL
XFILL_5__463_ vdd gnd FILL
XFILL_5__532_ vdd gnd FILL
XFILL_5__394_ vdd gnd FILL
XFILL_2__519_ vdd gnd FILL
XFILL_9__510_ vdd gnd FILL
XFILL_9__441_ vdd gnd FILL
XFILL_9__372_ vdd gnd FILL
X_456_ _461_/C _461_/B _459_/C vdd gnd OR2X2
X_525_ _611_/D _525_/B _554_/B vdd gnd NAND2X1
XFILL72750x10950 vdd gnd FILL
XFILL_4__481_ vdd gnd FILL
X_387_ _410_/B _387_/B _387_/C _564_/D vdd gnd OAI21X1
XFILL_4__550_ vdd gnd FILL
XFILL_6__428_ vdd gnd FILL
XFILL_6__359_ vdd gnd FILL
XFILL_1__468_ vdd gnd FILL
XFILL_1__537_ vdd gnd FILL
XFILL_1__399_ vdd gnd FILL
XFILL_8__390_ vdd gnd FILL
XFILL_2__304_ vdd gnd FILL
XFILL_5__515_ vdd gnd FILL
XFILL_5__446_ vdd gnd FILL
XFILL_5__377_ vdd gnd FILL
X_310_ _609_/D _317_/A vdd gnd INVX1
XFILL_0__624_ vdd gnd FILL
XFILL_0__486_ vdd gnd FILL
XFILL_0__555_ vdd gnd FILL
XFILL_9__424_ vdd gnd FILL
X_508_ _513_/A _510_/A vdd gnd INVX1
XFILL_1__322_ vdd gnd FILL
XFILL_9__286_ vdd gnd FILL
X_439_ _439_/A _439_/B _439_/C _440_/C vdd gnd NAND3X1
XFILL_4__464_ vdd gnd FILL
XFILL_4__533_ vdd gnd FILL
XFILL_4__395_ vdd gnd FILL
XFILL_5__300_ vdd gnd FILL
XFILL_8__511_ vdd gnd FILL
XFILL_8__442_ vdd gnd FILL
XFILL_0__340_ vdd gnd FILL
XFILL_8__373_ vdd gnd FILL
XFILL_7_BUFX2_insert18 vdd gnd FILL
XFILL_3__620_ vdd gnd FILL
XFILL_3__551_ vdd gnd FILL
XFILL_3__482_ vdd gnd FILL
XFILL_5__429_ vdd gnd FILL
XFILL_0__469_ vdd gnd FILL
XFILL_7__460_ vdd gnd FILL
XFILL_0__538_ vdd gnd FILL
XFILL_9__338_ vdd gnd FILL
XFILL_9__407_ vdd gnd FILL
XFILL_7__391_ vdd gnd FILL
XFILL_1__305_ vdd gnd FILL
XFILL_4__447_ vdd gnd FILL
XFILL_4__516_ vdd gnd FILL
XFILL_4__378_ vdd gnd FILL
XFILL_8__425_ vdd gnd FILL
XFILL_5_CLKBUF1_insert1 vdd gnd FILL
XFILL_8__356_ vdd gnd FILL
XFILL_8__287_ vdd gnd FILL
XFILL_0__323_ vdd gnd FILL
XFILL_3__465_ vdd gnd FILL
XFILL_3__534_ vdd gnd FILL
XFILL_3__396_ vdd gnd FILL
XFILL_4__301_ vdd gnd FILL
XFILL_3_BUFX2_insert16 vdd gnd FILL
XFILL_7__512_ vdd gnd FILL
XFILL_7__443_ vdd gnd FILL
XFILL_7__374_ vdd gnd FILL
XFILL_2__621_ vdd gnd FILL
XFILL_2__552_ vdd gnd FILL
XFILL_2__483_ vdd gnd FILL
XFILL_6__530_ vdd gnd FILL
XFILL_6__461_ vdd gnd FILL
XFILL_8__408_ vdd gnd FILL
XFILL_6__392_ vdd gnd FILL
XFILL_8__339_ vdd gnd FILL
XFILL_0__306_ vdd gnd FILL
XFILL_3__448_ vdd gnd FILL
XFILL_3__517_ vdd gnd FILL
XFILL_3__379_ vdd gnd FILL
XFILL_7__426_ vdd gnd FILL
XFILL_7__288_ vdd gnd FILL
XFILL_7__357_ vdd gnd FILL
XFILL_2__535_ vdd gnd FILL
XFILL_2__466_ vdd gnd FILL
XFILL_2__397_ vdd gnd FILL
X_610_ _610_/D _612_/CLK _611_/D vdd gnd DFFPOSX1
X_472_ _472_/A _478_/A _472_/C _576_/D vdd gnd OAI21X1
XFILL_3__302_ vdd gnd FILL
X_541_ _607_/D _541_/B _591_/Q _542_/C vdd gnd OAI21X1
XFILL_6__513_ vdd gnd FILL
XFILL_6__444_ vdd gnd FILL
XFILL_6__375_ vdd gnd FILL
XFILL_1__622_ vdd gnd FILL
XFILL_6_BUFX2_insert20 vdd gnd FILL
XFILL_1__484_ vdd gnd FILL
XFILL_1__553_ vdd gnd FILL
XFILL_2__320_ vdd gnd FILL
XFILL_5__531_ vdd gnd FILL
XFILL_5__462_ vdd gnd FILL
XFILL_7__409_ vdd gnd FILL
XFILL_5__393_ vdd gnd FILL
XFILL_2__518_ vdd gnd FILL
XFILL_2__449_ vdd gnd FILL
XFILL_9__440_ vdd gnd FILL
XFILL_9__371_ vdd gnd FILL
X_455_ _509_/A _483_/A _461_/C vdd gnd NAND2X1
X_386_ _564_/Q _410_/B _387_/C vdd gnd NAND2X1
X_524_ Xin[0] _540_/A vdd gnd INVX1
XFILL_4__480_ vdd gnd FILL
XFILL_6__427_ vdd gnd FILL
XFILL_6__289_ vdd gnd FILL
XFILL_6__358_ vdd gnd FILL
XFILL_1__536_ vdd gnd FILL
XFILL_1__467_ vdd gnd FILL
XFILL_1__398_ vdd gnd FILL
XFILL_2__303_ vdd gnd FILL
XFILL_5__514_ vdd gnd FILL
XFILL_5__445_ vdd gnd FILL
XFILL_5__376_ vdd gnd FILL
XFILL_0__623_ vdd gnd FILL
XFILL_0__485_ vdd gnd FILL
XFILL_0__554_ vdd gnd FILL
XFILL_9__285_ vdd gnd FILL
XFILL_9__354_ vdd gnd FILL
XFILL_1__321_ vdd gnd FILL
X_507_ _507_/A _507_/B _513_/A vdd gnd NAND2X1
X_369_ _369_/A _369_/B _371_/B vdd gnd NAND2X1
X_438_ _438_/A _490_/A _438_/C _439_/C vdd gnd OAI21X1
XFILL_4__463_ vdd gnd FILL
XFILL_0_CLKBUF1_insert0 vdd gnd FILL
XFILL_4__532_ vdd gnd FILL
XFILL_4__394_ vdd gnd FILL
XFILL_1__519_ vdd gnd FILL
XFILL_8__510_ vdd gnd FILL
XFILL_8__441_ vdd gnd FILL
XFILL_8__372_ vdd gnd FILL
XFILL_7_BUFX2_insert19 vdd gnd FILL
XFILL_3__481_ vdd gnd FILL
XFILL_3__550_ vdd gnd FILL
XFILL_5__428_ vdd gnd FILL
XFILL_5__359_ vdd gnd FILL
XFILL_0__468_ vdd gnd FILL
XFILL_9__406_ vdd gnd FILL
XFILL_0__537_ vdd gnd FILL
XFILL_0__399_ vdd gnd FILL
XFILL_7__390_ vdd gnd FILL
XFILL_1__304_ vdd gnd FILL
XFILL_4__515_ vdd gnd FILL
XFILL_4__446_ vdd gnd FILL
XFILL_4__377_ vdd gnd FILL
XFILL_5_CLKBUF1_insert2 vdd gnd FILL
XFILL_8__424_ vdd gnd FILL
XFILL_8__355_ vdd gnd FILL
XFILL_0__322_ vdd gnd FILL
XFILL_8__286_ vdd gnd FILL
XFILL_3__464_ vdd gnd FILL
XFILL_3__533_ vdd gnd FILL
XFILL_3_BUFX2_insert17 vdd gnd FILL
XFILL_3__395_ vdd gnd FILL
XFILL_4__300_ vdd gnd FILL
XFILL_7__511_ vdd gnd FILL
XFILL_7__442_ vdd gnd FILL
XFILL_7__373_ vdd gnd FILL
XFILL_2__620_ vdd gnd FILL
XFILL_2__551_ vdd gnd FILL
XFILL_2__482_ vdd gnd FILL
XFILL_4__429_ vdd gnd FILL
XFILL_6__460_ vdd gnd FILL
XFILL_8__338_ vdd gnd FILL
XFILL_8__407_ vdd gnd FILL
XFILL_6__391_ vdd gnd FILL
XFILL_0__305_ vdd gnd FILL
XFILL_3__447_ vdd gnd FILL
XFILL_3__516_ vdd gnd FILL
XFILL_3__378_ vdd gnd FILL
XFILL75150x28950 vdd gnd FILL
XFILL_7__425_ vdd gnd FILL
XFILL_7__356_ vdd gnd FILL
XFILL_7__287_ vdd gnd FILL
XFILL_2__465_ vdd gnd FILL
XFILL_2__534_ vdd gnd FILL
X_540_ _540_/A _542_/B _540_/C _590_/D vdd gnd OAI21X1
XFILL_2__396_ vdd gnd FILL
X_471_ _478_/A _471_/B _471_/C _472_/C vdd gnd NAND3X1
XFILL_3__301_ vdd gnd FILL
XFILL_6__512_ vdd gnd FILL
XFILL_6__443_ vdd gnd FILL
XFILL_2_BUFX2_insert7 vdd gnd FILL
XFILL_6__374_ vdd gnd FILL
XFILL_1__621_ vdd gnd FILL
XFILL_6_BUFX2_insert10 vdd gnd FILL
XFILL_1__552_ vdd gnd FILL
XFILL75750x50550 vdd gnd FILL
XFILL_6_BUFX2_insert21 vdd gnd FILL
XFILL_1__483_ vdd gnd FILL
XFILL_5__530_ vdd gnd FILL
XFILL_5__461_ vdd gnd FILL
XFILL_7__408_ vdd gnd FILL
XFILL_5__392_ vdd gnd FILL
XFILL_7__339_ vdd gnd FILL
XFILL_2__448_ vdd gnd FILL
XFILL_2__517_ vdd gnd FILL
X_523_ _523_/A _550_/B _523_/C _583_/D vdd gnd OAI21X1
XFILL_2__379_ vdd gnd FILL
X_454_ _457_/A _457_/B _483_/A vdd gnd NAND2X1
X_385_ _385_/A _385_/B _387_/B vdd gnd NAND2X1
XFILL_6__426_ vdd gnd FILL
XFILL_6__288_ vdd gnd FILL
XFILL_6__357_ vdd gnd FILL
XFILL_9__499_ vdd gnd FILL
XFILL_1__535_ vdd gnd FILL
XFILL_1__466_ vdd gnd FILL
XFILL_1__397_ vdd gnd FILL
XFILL_2__302_ vdd gnd FILL
XFILL_5__513_ vdd gnd FILL
XFILL_5__444_ vdd gnd FILL
XFILL_5__375_ vdd gnd FILL
XFILL_0__622_ vdd gnd FILL
XFILL_0__553_ vdd gnd FILL
XFILL_0__484_ vdd gnd FILL
XFILL_9__422_ vdd gnd FILL
X_506_ _595_/Q _506_/B _507_/B vdd gnd NAND2X1
XFILL_9__353_ vdd gnd FILL
X_299_ _305_/A _299_/B _299_/C _623_/A vdd gnd OAI21X1
XFILL_1__320_ vdd gnd FILL
X_437_ _604_/Q _605_/Q _442_/C _439_/B vdd gnd NAND3X1
X_368_ _490_/A _414_/B _536_/A _369_/B vdd gnd OAI21X1
XFILL_4__531_ vdd gnd FILL
XFILL75450x72150 vdd gnd FILL
XFILL_4__462_ vdd gnd FILL
XFILL_6__409_ vdd gnd FILL
XFILL_0_CLKBUF1_insert1 vdd gnd FILL
XFILL_4__393_ vdd gnd FILL
XFILL_1__449_ vdd gnd FILL
XFILL_1__518_ vdd gnd FILL
XFILL_8__440_ vdd gnd FILL
XFILL_8__371_ vdd gnd FILL
XFILL_3__480_ vdd gnd FILL
XFILL_5__427_ vdd gnd FILL
XFILL_5__289_ vdd gnd FILL
XFILL_5__358_ vdd gnd FILL
XFILL_0__536_ vdd gnd FILL
XFILL_0__467_ vdd gnd FILL
XFILL_9__405_ vdd gnd FILL
XFILL_0__398_ vdd gnd FILL
XFILL_9__336_ vdd gnd FILL
XFILL_1__303_ vdd gnd FILL
XFILL_4__514_ vdd gnd FILL
XFILL_4__445_ vdd gnd FILL
XFILL_4__376_ vdd gnd FILL
XFILL_8__285_ vdd gnd FILL
XFILL_5_CLKBUF1_insert3 vdd gnd FILL
XFILL_8__423_ vdd gnd FILL
XFILL_8__354_ vdd gnd FILL
XFILL_0__321_ vdd gnd FILL
XFILL_3__463_ vdd gnd FILL
XFILL_3__532_ vdd gnd FILL
XFILL_3__394_ vdd gnd FILL
XFILL_3_BUFX2_insert18 vdd gnd FILL
XFILL_7__510_ vdd gnd FILL
XFILL_0__519_ vdd gnd FILL
XFILL_9__319_ vdd gnd FILL
XFILL_7__441_ vdd gnd FILL
XFILL_7__372_ vdd gnd FILL
XFILL_2__481_ vdd gnd FILL
XFILL_2__550_ vdd gnd FILL
XFILL_4__428_ vdd gnd FILL
XFILL_4__359_ vdd gnd FILL
XFILL_8__406_ vdd gnd FILL
XFILL_6__390_ vdd gnd FILL
XFILL_8__337_ vdd gnd FILL
XFILL_3__515_ vdd gnd FILL
XFILL_0__304_ vdd gnd FILL
XFILL_3__446_ vdd gnd FILL
XFILL_3__377_ vdd gnd FILL
XFILL_7__286_ vdd gnd FILL
XFILL_7__424_ vdd gnd FILL
XFILL_7__355_ vdd gnd FILL
XFILL_2__464_ vdd gnd FILL
XFILL_2__533_ vdd gnd FILL
XFILL_2__395_ vdd gnd FILL
XFILL_3__300_ vdd gnd FILL
X_470_ _473_/A _477_/C _471_/C vdd gnd NAND2X1
XFILL_6__511_ vdd gnd FILL
XFILL_6__442_ vdd gnd FILL
XFILL_6__373_ vdd gnd FILL
XFILL_2_BUFX2_insert8 vdd gnd FILL
XFILL_6_BUFX2_insert11 vdd gnd FILL
XFILL_1__482_ vdd gnd FILL
XFILL_1__620_ vdd gnd FILL
XFILL_1__551_ vdd gnd FILL
X_599_ _599_/D _601_/CLK _599_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert22 vdd gnd FILL
XFILL_3__429_ vdd gnd FILL
XFILL_5__460_ vdd gnd FILL
XFILL_7__338_ vdd gnd FILL
XFILL_7__407_ vdd gnd FILL
XFILL_5__391_ vdd gnd FILL
XFILL_2__447_ vdd gnd FILL
XFILL_2__516_ vdd gnd FILL
XFILL_2__378_ vdd gnd FILL
X_453_ _602_/Q _603_/Q _457_/B vdd gnd NOR2X1
X_522_ Xin[1] _550_/B _523_/C vdd gnd NAND2X1
X_384_ _389_/A _393_/C _385_/B vdd gnd NAND2X1
XFILL_6__425_ vdd gnd FILL
XFILL_6__356_ vdd gnd FILL
XFILL_6__287_ vdd gnd FILL
XFILL_1__465_ vdd gnd FILL
XFILL_1__534_ vdd gnd FILL
XFILL_1__396_ vdd gnd FILL
XFILL_2__301_ vdd gnd FILL
XFILL_2_BUFX2_insert20 vdd gnd FILL
XFILL_5__512_ vdd gnd FILL
XFILL_5__443_ vdd gnd FILL
XFILL_5__374_ vdd gnd FILL
XFILL_0__621_ vdd gnd FILL
XFILL_0__552_ vdd gnd FILL
XFILL_0__483_ vdd gnd FILL
XFILL_9__421_ vdd gnd FILL
XFILL_9__283_ vdd gnd FILL
X_436_ _452_/B _436_/B _436_/C _570_/D vdd gnd OAI21X1
X_505_ selSign _550_/A _507_/A vdd gnd NAND2X1
X_298_ _305_/A _566_/Q _299_/C vdd gnd NAND2X1
XFILL_4__461_ vdd gnd FILL
XFILL_0_CLKBUF1_insert2 vdd gnd FILL
XFILL_4__530_ vdd gnd FILL
X_367_ _367_/A _367_/B _414_/B vdd gnd AND2X2
XFILL_6__408_ vdd gnd FILL
XFILL_4__392_ vdd gnd FILL
XFILL_6__339_ vdd gnd FILL
XFILL_9__619_ vdd gnd FILL
XFILL_1__448_ vdd gnd FILL
XFILL_1__517_ vdd gnd FILL
XFILL74250x28950 vdd gnd FILL
XFILL_1__379_ vdd gnd FILL
XFILL_8__370_ vdd gnd FILL
XFILL_5__426_ vdd gnd FILL
XFILL_5__357_ vdd gnd FILL
XFILL_5__288_ vdd gnd FILL
XFILL_8__499_ vdd gnd FILL
XFILL_0__466_ vdd gnd FILL
XFILL_0__535_ vdd gnd FILL
XFILL_0__397_ vdd gnd FILL
XFILL_9__335_ vdd gnd FILL
XFILL_1__302_ vdd gnd FILL
X_419_ _439_/A _419_/B _419_/C _420_/C vdd gnd NAND3X1
XFILL_4__513_ vdd gnd FILL
XFILL_4__444_ vdd gnd FILL
XFILL_4__375_ vdd gnd FILL
XFILL_8__422_ vdd gnd FILL
XFILL_0__320_ vdd gnd FILL
XFILL_8__284_ vdd gnd FILL
XFILL_5_CLKBUF1_insert4 vdd gnd FILL
XFILL_8__353_ vdd gnd FILL
XFILL_3__531_ vdd gnd FILL
XFILL_3__462_ vdd gnd FILL
XFILL_5__409_ vdd gnd FILL
XFILL_3__393_ vdd gnd FILL
XFILL_3_BUFX2_insert19 vdd gnd FILL
XFILL_0__449_ vdd gnd FILL
XFILL_0__518_ vdd gnd FILL
XFILL_7__440_ vdd gnd FILL
XFILL_7__371_ vdd gnd FILL
XFILL_2__480_ vdd gnd FILL
XFILL_4__427_ vdd gnd FILL
XFILL_4__289_ vdd gnd FILL
XFILL_4__358_ vdd gnd FILL
XFILL_8__336_ vdd gnd FILL
XFILL_8__405_ vdd gnd FILL
XFILL_0__303_ vdd gnd FILL
XFILL_3__514_ vdd gnd FILL
XFILL_3__445_ vdd gnd FILL
XFILL_3__376_ vdd gnd FILL
XFILL75750x10950 vdd gnd FILL
XFILL_7__423_ vdd gnd FILL
XFILL_7__285_ vdd gnd FILL
XFILL_7__354_ vdd gnd FILL
XFILL_2__532_ vdd gnd FILL
XFILL74550x72150 vdd gnd FILL
XFILL_2__463_ vdd gnd FILL
XFILL_2__394_ vdd gnd FILL
XFILL_6__510_ vdd gnd FILL
XFILL_2_BUFX2_insert9 vdd gnd FILL
XFILL_8__319_ vdd gnd FILL
XFILL_6__441_ vdd gnd FILL
XFILL_6__372_ vdd gnd FILL
XFILL_6_BUFX2_insert12 vdd gnd FILL
XFILL_1__481_ vdd gnd FILL
X_598_ _598_/D _601_/CLK _598_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert23 vdd gnd FILL
XFILL_1__550_ vdd gnd FILL
XFILL_3__428_ vdd gnd FILL
XFILL75450x57750 vdd gnd FILL
XFILL_3__359_ vdd gnd FILL
XFILL_7__406_ vdd gnd FILL
XFILL_5__390_ vdd gnd FILL
XFILL_7__337_ vdd gnd FILL
XFILL_2__515_ vdd gnd FILL
XFILL_2__446_ vdd gnd FILL
XFILL_2__377_ vdd gnd FILL
X_452_ _452_/A _452_/B _452_/C _573_/D vdd gnd OAI21X1
X_521_ _521_/A _550_/B _521_/C _582_/D vdd gnd OAI21X1
X_383_ _430_/C _383_/B _393_/C vdd gnd NAND2X1
XFILL_6__286_ vdd gnd FILL
XFILL_6__424_ vdd gnd FILL
XFILL_6__355_ vdd gnd FILL
XFILL_9__497_ vdd gnd FILL
XFILL_1__464_ vdd gnd FILL
XFILL_1__533_ vdd gnd FILL
XFILL_1__395_ vdd gnd FILL
XFILL_2_BUFX2_insert10 vdd gnd FILL
XFILL_2__300_ vdd gnd FILL
XFILL_2_BUFX2_insert21 vdd gnd FILL
XFILL_5__511_ vdd gnd FILL
XFILL_5__442_ vdd gnd FILL
XFILL_5__373_ vdd gnd FILL
XFILL_0__482_ vdd gnd FILL
XFILL_0__620_ vdd gnd FILL
XFILL_0__551_ vdd gnd FILL
XFILL_9__282_ vdd gnd FILL
XFILL_9__420_ vdd gnd FILL
XFILL_2__429_ vdd gnd FILL
XFILL_9__351_ vdd gnd FILL
X_435_ _604_/Q _460_/B _436_/C vdd gnd NAND2X1
X_366_ _588_/Q _536_/A vdd gnd INVX1
X_504_ _595_/Q _550_/A vdd gnd INVX1
X_297_ _578_/Q _299_/B vdd gnd INVX1
XFILL_4__460_ vdd gnd FILL
XFILL_0_CLKBUF1_insert3 vdd gnd FILL
XFILL_6__407_ vdd gnd FILL
XFILL_6__338_ vdd gnd FILL
XFILL_4__391_ vdd gnd FILL
XFILL_9__549_ vdd gnd FILL
XFILL_1__447_ vdd gnd FILL
XFILL_1__516_ vdd gnd FILL
XFILL_1__378_ vdd gnd FILL
XFILL_5__287_ vdd gnd FILL
XFILL_5__425_ vdd gnd FILL
XFILL_5__356_ vdd gnd FILL
XFILL_8__498_ vdd gnd FILL
XFILL_0__465_ vdd gnd FILL
XFILL_0__534_ vdd gnd FILL
XFILL_9__403_ vdd gnd FILL
XFILL_9__334_ vdd gnd FILL
XFILL_0__396_ vdd gnd FILL
XFILL_1__301_ vdd gnd FILL
X_418_ _521_/A _429_/C _419_/C vdd gnd NAND2X1
X_349_ _590_/Q _357_/B vdd gnd INVX1
XFILL_4__512_ vdd gnd FILL
XFILL_4__443_ vdd gnd FILL
XFILL_4__374_ vdd gnd FILL
XFILL_8__421_ vdd gnd FILL
XFILL_8__352_ vdd gnd FILL
XFILL_8__283_ vdd gnd FILL
XFILL_5_CLKBUF1_insert5 vdd gnd FILL
XFILL_3__461_ vdd gnd FILL
XFILL_3__530_ vdd gnd FILL
XFILL_5__408_ vdd gnd FILL
XFILL_3__392_ vdd gnd FILL
XFILL_5__339_ vdd gnd FILL
XFILL_8__619_ vdd gnd FILL
XFILL_0__448_ vdd gnd FILL
XFILL_0__379_ vdd gnd FILL
XFILL_0__517_ vdd gnd FILL
XFILL_9__317_ vdd gnd FILL
XFILL_7__370_ vdd gnd FILL
XFILL_4__426_ vdd gnd FILL
XFILL_4__357_ vdd gnd FILL
XFILL_4__288_ vdd gnd FILL
XFILL_7__499_ vdd gnd FILL
XFILL_8__404_ vdd gnd FILL
XFILL_8__335_ vdd gnd FILL
XFILL_0__302_ vdd gnd FILL
XFILL_3__513_ vdd gnd FILL
XFILL_3__444_ vdd gnd FILL
XFILL_3__375_ vdd gnd FILL
XFILL_7__422_ vdd gnd FILL
XFILL_7__353_ vdd gnd FILL
XFILL_7__284_ vdd gnd FILL
XFILL_2__531_ vdd gnd FILL
XFILL_2__462_ vdd gnd FILL
XFILL_4__409_ vdd gnd FILL
XFILL_2__393_ vdd gnd FILL
XFILL_6__440_ vdd gnd FILL
XFILL73350x28950 vdd gnd FILL
XFILL_8__318_ vdd gnd FILL
XFILL_6__371_ vdd gnd FILL
XFILL_1__480_ vdd gnd FILL
X_597_ _597_/D _601_/CLK _597_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert24 vdd gnd FILL
XFILL_3__427_ vdd gnd FILL
XFILL_6_BUFX2_insert13 vdd gnd FILL
XFILL_3__358_ vdd gnd FILL
XFILL_3__289_ vdd gnd FILL
XFILL_7__336_ vdd gnd FILL
XFILL_7__405_ vdd gnd FILL
XFILL_2__514_ vdd gnd FILL
XFILL_2__445_ vdd gnd FILL
X_520_ Xin[0] _550_/B _521_/C vdd gnd NAND2X1
XFILL_2__376_ vdd gnd FILL
X_451_ _460_/B _451_/B _451_/C _452_/C vdd gnd NAND3X1
X_382_ _586_/Q _389_/A vdd gnd INVX1
XFILL_6__423_ vdd gnd FILL
XFILL_6__285_ vdd gnd FILL
XFILL_6__354_ vdd gnd FILL
XFILL_9__496_ vdd gnd FILL
XFILL_1__532_ vdd gnd FILL
XFILL_1__463_ vdd gnd FILL
XFILL_1__394_ vdd gnd FILL
XFILL_2_BUFX2_insert11 vdd gnd FILL
XFILL_2_BUFX2_insert22 vdd gnd FILL
XFILL_5__510_ vdd gnd FILL
XFILL_7__319_ vdd gnd FILL
XFILL_5__441_ vdd gnd FILL
XFILL_5__372_ vdd gnd FILL
XFILL_0__481_ vdd gnd FILL
XFILL_0__550_ vdd gnd FILL
XFILL_2__428_ vdd gnd FILL
X_503_ _581_/Q _503_/B _515_/A vdd gnd NAND2X1
XFILL_9__281_ vdd gnd FILL
XFILL_9__350_ vdd gnd FILL
XFILL_2__359_ vdd gnd FILL
X_296_ _305_/A _479_/A _296_/C _622_/A vdd gnd OAI21X1
X_365_ _415_/A _588_/Q _399_/A _369_/A vdd gnd NAND3X1
X_434_ _434_/A _434_/B _569_/D vdd gnd NAND2X1
XFILL_6__406_ vdd gnd FILL
XFILL_0_CLKBUF1_insert4 vdd gnd FILL
XFILL_4__390_ vdd gnd FILL
XFILL_6__337_ vdd gnd FILL
XFILL_9__617_ vdd gnd FILL
XFILL_9__548_ vdd gnd FILL
XFILL_1__515_ vdd gnd FILL
XFILL74850x10950 vdd gnd FILL
XFILL_1__446_ vdd gnd FILL
XFILL_1__377_ vdd gnd FILL
XFILL_5__424_ vdd gnd FILL
XFILL_5__286_ vdd gnd FILL
XFILL_5__355_ vdd gnd FILL
XFILL_8__497_ vdd gnd FILL
XFILL73650x72150 vdd gnd FILL
XFILL_0__464_ vdd gnd FILL
XFILL_9__402_ vdd gnd FILL
XFILL_0__533_ vdd gnd FILL
XFILL_0__395_ vdd gnd FILL
XFILL_1__300_ vdd gnd FILL
XFILL_4__511_ vdd gnd FILL
X_279_ _572_/Q _447_/A vdd gnd INVX1
X_417_ _442_/C _417_/B _429_/C vdd gnd NAND2X1
X_348_ _421_/B _348_/B _348_/C _559_/D vdd gnd OAI21X1
XFILL_4__442_ vdd gnd FILL
XFILL_4__373_ vdd gnd FILL
XFILL74550x57750 vdd gnd FILL
XFILL_1__429_ vdd gnd FILL
XFILL_8__282_ vdd gnd FILL
XFILL_8__420_ vdd gnd FILL
XFILL_5_CLKBUF1_insert6 vdd gnd FILL
XFILL_8__351_ vdd gnd FILL
XFILL_3__460_ vdd gnd FILL
XFILL_5__407_ vdd gnd FILL
XFILL_3__391_ vdd gnd FILL
XFILL_5__338_ vdd gnd FILL
XFILL_8__618_ vdd gnd FILL
XFILL_8__549_ vdd gnd FILL
XFILL_0__516_ vdd gnd FILL
XFILL_0__447_ vdd gnd FILL
XFILL_0__378_ vdd gnd FILL
XFILL_9__316_ vdd gnd FILL
XFILL_4__287_ vdd gnd FILL
XFILL_4__425_ vdd gnd FILL
XFILL_4__356_ vdd gnd FILL
XFILL_7__498_ vdd gnd FILL
XFILL_8__403_ vdd gnd FILL
XFILL_8__334_ vdd gnd FILL
XFILL_0__301_ vdd gnd FILL
XFILL_3__512_ vdd gnd FILL
XFILL_3__443_ vdd gnd FILL
XFILL_3__374_ vdd gnd FILL
XFILL_7__421_ vdd gnd FILL
XFILL_7__352_ vdd gnd FILL
XFILL_7__283_ vdd gnd FILL
XFILL_2__461_ vdd gnd FILL
XFILL_2__530_ vdd gnd FILL
XFILL_7__619_ vdd gnd FILL
XFILL_4__408_ vdd gnd FILL
XFILL_2__392_ vdd gnd FILL
XFILL_4__339_ vdd gnd FILL
XFILL_6__370_ vdd gnd FILL
XFILL_8__317_ vdd gnd FILL
XFILL_6_BUFX2_insert25 vdd gnd FILL
XFILL_6_BUFX2_insert14 vdd gnd FILL
X_596_ _596_/D _601_/CLK _596_/Q vdd gnd DFFPOSX1
XFILL_3__426_ vdd gnd FILL
XFILL_3__357_ vdd gnd FILL
XFILL_6__499_ vdd gnd FILL
XFILL_3__288_ vdd gnd FILL
XFILL_7__404_ vdd gnd FILL
XFILL_7__335_ vdd gnd FILL
XFILL_2__513_ vdd gnd FILL
XFILL_2__444_ vdd gnd FILL
XFILL_2__375_ vdd gnd FILL
X_450_ _450_/A _603_/Q _451_/C vdd gnd OR2X2
X_381_ _430_/C _586_/Q _383_/B _385_/A vdd gnd NAND3X1
XFILL_6__422_ vdd gnd FILL
XFILL_6__353_ vdd gnd FILL
XFILL_6__284_ vdd gnd FILL
XFILL_1__462_ vdd gnd FILL
XFILL_9__495_ vdd gnd FILL
XFILL75150x39750 vdd gnd FILL
XFILL_1__531_ vdd gnd FILL
X_579_ _579_/D _581_/CLK _579_/Q vdd gnd DFFPOSX1
XFILL_3__409_ vdd gnd FILL
XFILL_1__393_ vdd gnd FILL
XFILL_2_BUFX2_insert12 vdd gnd FILL
XFILL_2_BUFX2_insert23 vdd gnd FILL
XFILL_5__440_ vdd gnd FILL
XFILL_7__318_ vdd gnd FILL
XFILL_5__371_ vdd gnd FILL
XFILL_0__480_ vdd gnd FILL
XFILL_2__427_ vdd gnd FILL
XFILL_2__358_ vdd gnd FILL
X_502_ _502_/A _625_/A _502_/C _580_/D vdd gnd OAI21X1
XFILL_2__289_ vdd gnd FILL
X_433_ _439_/A _433_/B _433_/C _434_/B vdd gnd NAND3X1
X_295_ _308_/A _565_/Q _296_/C vdd gnd NAND2X1
X_364_ _367_/A _367_/B _399_/A vdd gnd NAND2X1
XFILL_6__336_ vdd gnd FILL
XFILL_6__405_ vdd gnd FILL
XFILL_0_CLKBUF1_insert5 vdd gnd FILL
XFILL75750x18150 vdd gnd FILL
XFILL_9__616_ vdd gnd FILL
XFILL_9__478_ vdd gnd FILL
XFILL75750x61350 vdd gnd FILL
XFILL_1__514_ vdd gnd FILL
XFILL_1__445_ vdd gnd FILL
XFILL_1__376_ vdd gnd FILL
XFILL_5__423_ vdd gnd FILL
XFILL_6_CLKBUF1_insert0 vdd gnd FILL
XFILL_5__285_ vdd gnd FILL
XFILL_5__354_ vdd gnd FILL
XFILL_8__496_ vdd gnd FILL
XFILL_0__532_ vdd gnd FILL
XFILL_0__463_ vdd gnd FILL
XFILL_0__394_ vdd gnd FILL
XFILL_9__401_ vdd gnd FILL
XFILL_9__332_ vdd gnd FILL
X_416_ _582_/Q _521_/A vdd gnd INVX1
XFILL_4__510_ vdd gnd FILL
XFILL_4__441_ vdd gnd FILL
X_278_ _286_/A _440_/A _278_/C _614_/A vdd gnd OAI21X1
X_347_ _559_/Q _421_/B _348_/C vdd gnd NAND2X1
XFILL_6__319_ vdd gnd FILL
XFILL_4__372_ vdd gnd FILL
XFILL_1__428_ vdd gnd FILL
XFILL_8__281_ vdd gnd FILL
XFILL_8__350_ vdd gnd FILL
XFILL_1__359_ vdd gnd FILL
XFILL_5__337_ vdd gnd FILL
XFILL_5__406_ vdd gnd FILL
XFILL_3__390_ vdd gnd FILL
XFILL_8__617_ vdd gnd FILL
XFILL_8__548_ vdd gnd FILL
XFILL_8__479_ vdd gnd FILL
XFILL_0__515_ vdd gnd FILL
XFILL_0__446_ vdd gnd FILL
XFILL_9__315_ vdd gnd FILL
XFILL_0__377_ vdd gnd FILL
XFILL_4__424_ vdd gnd FILL
XFILL_4__286_ vdd gnd FILL
XFILL_4__355_ vdd gnd FILL
XFILL_7__497_ vdd gnd FILL
XFILL_8__402_ vdd gnd FILL
XFILL_0__300_ vdd gnd FILL
XFILL_8__333_ vdd gnd FILL
XFILL_3__511_ vdd gnd FILL
XFILL_3__442_ vdd gnd FILL
XFILL_3__373_ vdd gnd FILL
XFILL_0__429_ vdd gnd FILL
XFILL_7__282_ vdd gnd FILL
XFILL_7__420_ vdd gnd FILL
XFILL_7__351_ vdd gnd FILL
XFILL_2__460_ vdd gnd FILL
XFILL_4__407_ vdd gnd FILL
XFILL_2__391_ vdd gnd FILL
XFILL_4__338_ vdd gnd FILL
XFILL_7__618_ vdd gnd FILL
XFILL_7__549_ vdd gnd FILL
XFILL73950x10950 vdd gnd FILL
XFILL_8__316_ vdd gnd FILL
X_595_ _595_/D _595_/CLK _595_/Q vdd gnd DFFPOSX1
XFILL_6_BUFX2_insert15 vdd gnd FILL
XFILL_3__287_ vdd gnd FILL
XFILL_3__425_ vdd gnd FILL
XFILL_3__356_ vdd gnd FILL
XFILL72750x72150 vdd gnd FILL
XFILL_6__498_ vdd gnd FILL
XFILL_7__403_ vdd gnd FILL
XFILL_7__334_ vdd gnd FILL
XFILL_2__512_ vdd gnd FILL
XFILL_2__443_ vdd gnd FILL
XFILL_2__374_ vdd gnd FILL
XFILL73650x57750 vdd gnd FILL
X_380_ _412_/A _414_/B _383_/B vdd gnd NAND2X1
XFILL_6__283_ vdd gnd FILL
XFILL_6__421_ vdd gnd FILL
XFILL_6__352_ vdd gnd FILL
X_578_ _578_/D _581_/CLK _578_/Q vdd gnd DFFPOSX1
XFILL_1__461_ vdd gnd FILL
XFILL_3__408_ vdd gnd FILL
XFILL_1__530_ vdd gnd FILL
XFILL_6__619_ vdd gnd FILL
XFILL_1__392_ vdd gnd FILL
XFILL_3__339_ vdd gnd FILL
XFILL_2_BUFX2_insert24 vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
.ends

