magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -120 -120 2520 320
<< psubstratepdiff >>
rect 0 0 2400 200
<< metal1 >>
rect 0 0 2400 200
use CONT$3  CONT$3_0
timestamp 1569533753
transform 1 0 164 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_1
timestamp 1569533753
transform 1 0 128 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_2
timestamp 1569533753
transform 1 0 92 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_3
timestamp 1569533753
transform 1 0 236 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_4
timestamp 1569533753
transform 1 0 200 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_5
timestamp 1569533753
transform 1 0 164 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_6
timestamp 1569533753
transform 1 0 524 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_7
timestamp 1569533753
transform 1 0 488 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_8
timestamp 1569533753
transform 1 0 452 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_9
timestamp 1569533753
transform 1 0 416 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_10
timestamp 1569533753
transform 1 0 380 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_11
timestamp 1569533753
transform 1 0 344 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_12
timestamp 1569533753
transform 1 0 308 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_13
timestamp 1569533753
transform 1 0 272 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_14
timestamp 1569533753
transform 1 0 596 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_15
timestamp 1569533753
transform 1 0 560 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_16
timestamp 1569533753
transform 1 0 524 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_17
timestamp 1569533753
transform 1 0 488 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_18
timestamp 1569533753
transform 1 0 452 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_19
timestamp 1569533753
transform 1 0 416 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_20
timestamp 1569533753
transform 1 0 380 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_21
timestamp 1569533753
transform 1 0 344 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_22
timestamp 1569533753
transform 1 0 308 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_23
timestamp 1569533753
transform 1 0 272 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_24
timestamp 1569533753
transform 1 0 236 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_25
timestamp 1569533753
transform 1 0 200 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_26
timestamp 1569533753
transform 1 0 164 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_27
timestamp 1569533753
transform 1 0 128 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_28
timestamp 1569533753
transform 1 0 236 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_29
timestamp 1569533753
transform 1 0 200 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_30
timestamp 1569533753
transform 1 0 596 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_31
timestamp 1569533753
transform 1 0 596 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_32
timestamp 1569533753
transform 1 0 560 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_33
timestamp 1569533753
transform 1 0 524 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_34
timestamp 1569533753
transform 1 0 488 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_35
timestamp 1569533753
transform 1 0 452 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_36
timestamp 1569533753
transform 1 0 416 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_37
timestamp 1569533753
transform 1 0 380 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_38
timestamp 1569533753
transform 1 0 344 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_39
timestamp 1569533753
transform 1 0 596 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_40
timestamp 1569533753
transform 1 0 560 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_41
timestamp 1569533753
transform 1 0 524 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_42
timestamp 1569533753
transform 1 0 488 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_43
timestamp 1569533753
transform 1 0 452 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_44
timestamp 1569533753
transform 1 0 416 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_45
timestamp 1569533753
transform 1 0 380 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_46
timestamp 1569533753
transform 1 0 344 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_47
timestamp 1569533753
transform 1 0 308 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_48
timestamp 1569533753
transform 1 0 272 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_49
timestamp 1569533753
transform 1 0 236 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_50
timestamp 1569533753
transform 1 0 200 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_51
timestamp 1569533753
transform 1 0 164 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_52
timestamp 1569533753
transform 1 0 128 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_53
timestamp 1569533753
transform 1 0 92 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_54
timestamp 1569533753
transform 1 0 56 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_55
timestamp 1569533753
transform 1 0 92 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_56
timestamp 1569533753
transform 1 0 56 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_57
timestamp 1569533753
transform 1 0 56 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_58
timestamp 1569533753
transform 1 0 56 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_59
timestamp 1569533753
transform 1 0 308 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_60
timestamp 1569533753
transform 1 0 272 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_61
timestamp 1569533753
transform 1 0 236 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_62
timestamp 1569533753
transform 1 0 200 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_63
timestamp 1569533753
transform 1 0 164 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_64
timestamp 1569533753
transform 1 0 128 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_65
timestamp 1569533753
transform 1 0 92 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_66
timestamp 1569533753
transform 1 0 56 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_67
timestamp 1569533753
transform 1 0 128 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_68
timestamp 1569533753
transform 1 0 92 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_69
timestamp 1569533753
transform 1 0 560 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_70
timestamp 1569533753
transform 1 0 596 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_71
timestamp 1569533753
transform 1 0 560 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_72
timestamp 1569533753
transform 1 0 524 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_73
timestamp 1569533753
transform 1 0 488 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_74
timestamp 1569533753
transform 1 0 452 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_75
timestamp 1569533753
transform 1 0 416 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_76
timestamp 1569533753
transform 1 0 380 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_77
timestamp 1569533753
transform 1 0 344 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_78
timestamp 1569533753
transform 1 0 308 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_79
timestamp 1569533753
transform 1 0 272 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_80
timestamp 1569533753
transform 1 0 1172 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_81
timestamp 1569533753
transform 1 0 1136 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_82
timestamp 1569533753
transform 1 0 920 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_83
timestamp 1569533753
transform 1 0 884 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_84
timestamp 1569533753
transform 1 0 848 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_85
timestamp 1569533753
transform 1 0 812 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_86
timestamp 1569533753
transform 1 0 776 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_87
timestamp 1569533753
transform 1 0 740 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_88
timestamp 1569533753
transform 1 0 704 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_89
timestamp 1569533753
transform 1 0 668 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_90
timestamp 1569533753
transform 1 0 776 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_91
timestamp 1569533753
transform 1 0 1172 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_92
timestamp 1569533753
transform 1 0 1136 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_93
timestamp 1569533753
transform 1 0 920 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_94
timestamp 1569533753
transform 1 0 884 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_95
timestamp 1569533753
transform 1 0 848 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_96
timestamp 1569533753
transform 1 0 812 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_97
timestamp 1569533753
transform 1 0 776 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_98
timestamp 1569533753
transform 1 0 740 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_99
timestamp 1569533753
transform 1 0 704 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_100
timestamp 1569533753
transform 1 0 668 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_101
timestamp 1569533753
transform 1 0 740 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_102
timestamp 1569533753
transform 1 0 1172 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_103
timestamp 1569533753
transform 1 0 1136 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_104
timestamp 1569533753
transform 1 0 920 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_105
timestamp 1569533753
transform 1 0 884 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_106
timestamp 1569533753
transform 1 0 848 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_107
timestamp 1569533753
transform 1 0 812 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_108
timestamp 1569533753
transform 1 0 776 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_109
timestamp 1569533753
transform 1 0 740 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_110
timestamp 1569533753
transform 1 0 704 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_111
timestamp 1569533753
transform 1 0 668 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_112
timestamp 1569533753
transform 1 0 704 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_113
timestamp 1569533753
transform 1 0 1172 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_114
timestamp 1569533753
transform 1 0 1136 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_115
timestamp 1569533753
transform 1 0 920 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_116
timestamp 1569533753
transform 1 0 884 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_117
timestamp 1569533753
transform 1 0 848 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_118
timestamp 1569533753
transform 1 0 812 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_119
timestamp 1569533753
transform 1 0 776 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_120
timestamp 1569533753
transform 1 0 740 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_121
timestamp 1569533753
transform 1 0 704 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_122
timestamp 1569533753
transform 1 0 668 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_123
timestamp 1569533753
transform 1 0 668 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_124
timestamp 1569533753
transform 1 0 1172 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_125
timestamp 1569533753
transform 1 0 1136 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_126
timestamp 1569533753
transform 1 0 920 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_127
timestamp 1569533753
transform 1 0 884 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_128
timestamp 1569533753
transform 1 0 848 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_129
timestamp 1569533753
transform 1 0 812 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_130
timestamp 1569533753
transform 1 0 632 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_131
timestamp 1569533753
transform 1 0 632 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_132
timestamp 1569533753
transform 1 0 632 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_133
timestamp 1569533753
transform 1 0 632 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_134
timestamp 1569533753
transform 1 0 632 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_135
timestamp 1569533753
transform 1 0 1388 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_136
timestamp 1569533753
transform 1 0 1352 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_137
timestamp 1569533753
transform 1 0 1316 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_138
timestamp 1569533753
transform 1 0 1280 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_139
timestamp 1569533753
transform 1 0 1244 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_140
timestamp 1569533753
transform 1 0 1316 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_141
timestamp 1569533753
transform 1 0 1748 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_142
timestamp 1569533753
transform 1 0 1532 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_143
timestamp 1569533753
transform 1 0 1496 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_144
timestamp 1569533753
transform 1 0 1460 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_145
timestamp 1569533753
transform 1 0 1424 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_146
timestamp 1569533753
transform 1 0 1388 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_147
timestamp 1569533753
transform 1 0 1352 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_148
timestamp 1569533753
transform 1 0 1316 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_149
timestamp 1569533753
transform 1 0 1280 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_150
timestamp 1569533753
transform 1 0 1244 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_151
timestamp 1569533753
transform 1 0 1244 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_152
timestamp 1569533753
transform 1 0 1748 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_153
timestamp 1569533753
transform 1 0 1532 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_154
timestamp 1569533753
transform 1 0 1496 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_155
timestamp 1569533753
transform 1 0 1460 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_156
timestamp 1569533753
transform 1 0 1424 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_157
timestamp 1569533753
transform 1 0 1388 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_158
timestamp 1569533753
transform 1 0 1352 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_159
timestamp 1569533753
transform 1 0 1316 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_160
timestamp 1569533753
transform 1 0 1280 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_161
timestamp 1569533753
transform 1 0 1244 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_162
timestamp 1569533753
transform 1 0 1352 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_163
timestamp 1569533753
transform 1 0 1532 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_164
timestamp 1569533753
transform 1 0 1496 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_165
timestamp 1569533753
transform 1 0 1460 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_166
timestamp 1569533753
transform 1 0 1424 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_167
timestamp 1569533753
transform 1 0 1388 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_168
timestamp 1569533753
transform 1 0 1748 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_169
timestamp 1569533753
transform 1 0 1748 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_170
timestamp 1569533753
transform 1 0 1532 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_171
timestamp 1569533753
transform 1 0 1496 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_172
timestamp 1569533753
transform 1 0 1460 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_173
timestamp 1569533753
transform 1 0 1424 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_174
timestamp 1569533753
transform 1 0 1388 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_175
timestamp 1569533753
transform 1 0 1352 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_176
timestamp 1569533753
transform 1 0 1316 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_177
timestamp 1569533753
transform 1 0 1280 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_178
timestamp 1569533753
transform 1 0 1244 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_179
timestamp 1569533753
transform 1 0 1280 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_180
timestamp 1569533753
transform 1 0 1748 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_181
timestamp 1569533753
transform 1 0 1532 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_182
timestamp 1569533753
transform 1 0 1496 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_183
timestamp 1569533753
transform 1 0 1460 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_184
timestamp 1569533753
transform 1 0 1424 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_185
timestamp 1569533753
transform 1 0 2360 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_186
timestamp 1569533753
transform 1 0 2324 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_187
timestamp 1569533753
transform 1 0 2288 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_188
timestamp 1569533753
transform 1 0 2252 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_189
timestamp 1569533753
transform 1 0 2216 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_190
timestamp 1569533753
transform 1 0 2180 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_191
timestamp 1569533753
transform 1 0 2144 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_192
timestamp 1569533753
transform 1 0 2108 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_193
timestamp 1569533753
transform 1 0 2072 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_194
timestamp 1569533753
transform 1 0 2036 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_195
timestamp 1569533753
transform 1 0 2000 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_196
timestamp 1569533753
transform 1 0 1964 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_197
timestamp 1569533753
transform 1 0 1928 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_198
timestamp 1569533753
transform 1 0 1892 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_199
timestamp 1569533753
transform 1 0 1856 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_200
timestamp 1569533753
transform 1 0 1820 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_201
timestamp 1569533753
transform 1 0 1928 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_202
timestamp 1569533753
transform 1 0 2360 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_203
timestamp 1569533753
transform 1 0 2324 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_204
timestamp 1569533753
transform 1 0 2288 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_205
timestamp 1569533753
transform 1 0 2252 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_206
timestamp 1569533753
transform 1 0 2216 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_207
timestamp 1569533753
transform 1 0 2180 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_208
timestamp 1569533753
transform 1 0 2144 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_209
timestamp 1569533753
transform 1 0 2108 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_210
timestamp 1569533753
transform 1 0 2072 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_211
timestamp 1569533753
transform 1 0 2036 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_212
timestamp 1569533753
transform 1 0 2000 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_213
timestamp 1569533753
transform 1 0 1964 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_214
timestamp 1569533753
transform 1 0 1928 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_215
timestamp 1569533753
transform 1 0 1892 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_216
timestamp 1569533753
transform 1 0 1856 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_217
timestamp 1569533753
transform 1 0 1820 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_218
timestamp 1569533753
transform 1 0 1892 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_219
timestamp 1569533753
transform 1 0 2360 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_220
timestamp 1569533753
transform 1 0 2324 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_221
timestamp 1569533753
transform 1 0 2288 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_222
timestamp 1569533753
transform 1 0 2252 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_223
timestamp 1569533753
transform 1 0 2216 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_224
timestamp 1569533753
transform 1 0 2180 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_225
timestamp 1569533753
transform 1 0 2144 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_226
timestamp 1569533753
transform 1 0 2108 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_227
timestamp 1569533753
transform 1 0 2072 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_228
timestamp 1569533753
transform 1 0 2036 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_229
timestamp 1569533753
transform 1 0 2000 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_230
timestamp 1569533753
transform 1 0 1964 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_231
timestamp 1569533753
transform 1 0 1928 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_232
timestamp 1569533753
transform 1 0 1892 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_233
timestamp 1569533753
transform 1 0 1856 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_234
timestamp 1569533753
transform 1 0 1820 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_235
timestamp 1569533753
transform 1 0 1856 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_236
timestamp 1569533753
transform 1 0 2360 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_237
timestamp 1569533753
transform 1 0 2324 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_238
timestamp 1569533753
transform 1 0 2288 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_239
timestamp 1569533753
transform 1 0 2252 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_240
timestamp 1569533753
transform 1 0 2216 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_241
timestamp 1569533753
transform 1 0 2180 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_242
timestamp 1569533753
transform 1 0 2144 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_243
timestamp 1569533753
transform 1 0 2108 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_244
timestamp 1569533753
transform 1 0 2072 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_245
timestamp 1569533753
transform 1 0 2036 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_246
timestamp 1569533753
transform 1 0 2000 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_247
timestamp 1569533753
transform 1 0 1964 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_248
timestamp 1569533753
transform 1 0 1928 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_249
timestamp 1569533753
transform 1 0 1892 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_250
timestamp 1569533753
transform 1 0 1856 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_251
timestamp 1569533753
transform 1 0 1820 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_252
timestamp 1569533753
transform 1 0 1820 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_253
timestamp 1569533753
transform 1 0 2360 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_254
timestamp 1569533753
transform 1 0 2324 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_255
timestamp 1569533753
transform 1 0 2288 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_256
timestamp 1569533753
transform 1 0 2252 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_257
timestamp 1569533753
transform 1 0 2216 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_258
timestamp 1569533753
transform 1 0 2180 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_259
timestamp 1569533753
transform 1 0 2144 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_260
timestamp 1569533753
transform 1 0 2108 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_261
timestamp 1569533753
transform 1 0 2072 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_262
timestamp 1569533753
transform 1 0 2036 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_263
timestamp 1569533753
transform 1 0 2000 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_264
timestamp 1569533753
transform 1 0 1964 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_265
timestamp 1569533753
transform 1 0 1784 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_266
timestamp 1569533753
transform 1 0 1784 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_267
timestamp 1569533753
transform 1 0 1784 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_268
timestamp 1569533753
transform 1 0 1784 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_269
timestamp 1569533753
transform 1 0 1784 0 1 27
box -6 -6 6 6
use CONT$3  CONT$3_270
timestamp 1569533753
transform 1 0 1208 0 1 171
box -6 -6 6 6
use CONT$3  CONT$3_271
timestamp 1569533753
transform 1 0 1208 0 1 135
box -6 -6 6 6
use CONT$3  CONT$3_272
timestamp 1569533753
transform 1 0 1208 0 1 99
box -6 -6 6 6
use CONT$3  CONT$3_273
timestamp 1569533753
transform 1 0 1208 0 1 63
box -6 -6 6 6
use CONT$3  CONT$3_274
timestamp 1569533753
transform 1 0 1208 0 1 27
box -6 -6 6 6
<< end >>
