magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -127 -120 327 5132
<< nwell >>
rect -7 4201 207 4571
rect -7 2241 207 3839
<< psubstratepdiff >>
rect 20 4680 180 5012
rect 20 0 180 1560
<< nsubstratendiff >>
rect 20 4220 180 4552
rect 20 2260 180 3820
<< metal1 >>
rect 24 4680 176 5012
rect 24 4220 176 4552
rect 24 2260 176 3820
rect 24 0 176 1560
<< metal2 >>
rect 24 4680 176 5012
rect 24 4220 176 4552
rect 24 2260 176 3820
rect 24 0 176 1560
<< metal3 >>
rect 0 4680 200 5012
rect 0 4220 200 4552
rect 0 2260 200 3820
rect 0 0 200 1560
use CONT$1  CONT$1_0
array 0 1 64 0 23 64
timestamp 1569533753
transform 1 0 54 0 1 22
box -6 -6 6 6
use CONT$1  CONT$1_1
array 0 1 64 0 23 64
timestamp 1569533753
transform 1 0 48 0 1 2300
box -6 -6 6 6
use CONT$1  CONT$1_2
array 0 1 64 0 3 64
timestamp 1569533753
transform 1 0 48 0 1 4264
box -6 -6 6 6
use CONT$1  CONT$1_3
array 0 1 64 0 3 64
timestamp 1569533753
transform 1 0 48 0 1 4740
box -6 -6 6 6
use VIA1$1  VIA1$1_0
array 0 1 64 0 22 64
timestamp 1569533753
transform 1 0 80 0 1 2332
box -8 -8 8 8
use VIA1$1  VIA1$1_1
array 0 1 64 0 22 64
timestamp 1569533753
transform 1 0 86 0 1 54
box -8 -8 8 8
use VIA1$1  VIA1$1_2
array 0 1 64 0 2 64
timestamp 1569533753
transform 1 0 80 0 1 4296
box -8 -8 8 8
use VIA1$1  VIA1$1_3
array 0 1 64 0 2 64
timestamp 1569533753
transform 1 0 80 0 1 4772
box -8 -8 8 8
use VIA2$1  VIA2$1_0
array 0 1 64 0 23 64
timestamp 1569533753
transform 1 0 54 0 1 22
box -8 -8 8 8
use VIA2$1  VIA2$1_1
array 0 1 64 0 23 64
timestamp 1569533753
transform 1 0 48 0 1 2300
box -8 -8 8 8
use VIA2$1  VIA2$1_2
array 0 1 64 0 3 64
timestamp 1569533753
transform 1 0 48 0 1 4264
box -8 -8 8 8
use VIA2$1  VIA2$1_3
array 0 1 64 0 3 64
timestamp 1569533753
transform 1 0 48 0 1 4740
box -8 -8 8 8
<< end >>
