magic
tech scmos
magscale 1 30
timestamp 1740940952
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 59200 141200 134100 143600
rect 49100 138700 51000 138900
rect 49100 138600 51200 138700
rect 49100 138400 51400 138600
rect 49100 138200 51600 138400
rect 49100 138000 51800 138200
rect 49100 137800 52000 138000
rect 49100 137600 52200 137800
rect 49100 137400 52400 137600
rect 49100 137200 52600 137400
rect 49100 137000 52800 137200
rect 49100 136800 53000 137000
rect 49100 136600 53200 136800
rect 49100 136400 53400 136600
rect 49100 136200 53600 136400
rect 49100 136000 53800 136200
rect 49100 135800 54000 136000
rect 49100 135600 54200 135800
rect 49100 135400 54400 135600
rect 49100 135200 54600 135400
rect 49100 135000 54800 135200
rect 49100 134800 55000 135000
rect 49100 134600 55200 134800
rect 49100 134500 55400 134600
rect 49100 134300 55600 134500
rect 49100 134100 55800 134300
rect 49100 133900 56000 134100
rect 49100 133700 56200 133900
rect 49100 133500 56400 133700
rect 49100 132100 56600 133500
rect 133200 132600 134100 141200
<< m2contact >>
rect 49800 141200 59200 143600
rect 46600 132100 49100 138900
<< metal2 >>
rect 49800 143600 59200 146000
rect 44100 132100 46600 138900
rect 62400 134300 62900 145900
rect 75900 135300 76400 145900
rect 89400 136300 89900 145900
rect 102900 137300 103400 145900
rect 116400 138300 116900 145900
rect 129900 139300 130400 145900
rect 129900 138800 132500 139300
rect 116400 137800 128800 138300
rect 102900 136800 127800 137300
rect 89400 135800 124300 136300
rect 75900 134800 123300 135300
rect 62400 133800 109600 134300
rect 122800 133700 123300 134800
rect 123800 133700 124300 135800
rect 127300 133700 127800 136800
rect 128300 133700 128800 137800
rect 132000 133700 132500 138800
rect 145400 129900 145900 130400
rect 44100 116300 53100 116800
rect 145400 116400 145900 116900
rect 44100 102800 44600 103300
rect 145400 102900 145900 103400
rect 145400 89400 145900 89900
rect 145400 75900 145900 76400
rect 145400 62400 145900 62900
rect 102100 50400 102600 57200
rect 59700 49900 102600 50400
rect 44100 48600 45000 49500
rect 59700 44100 60200 49900
rect 103000 49400 103500 57200
rect 73200 48900 103500 49400
rect 73200 44100 73700 48900
rect 109900 48400 110400 57200
rect 86700 47900 110400 48400
rect 86700 44100 87200 47900
rect 110800 47400 111300 57200
rect 100200 46900 111300 47400
rect 100200 44100 100700 46900
rect 126300 46400 126800 57100
rect 113700 45900 126800 46400
rect 113700 44100 114200 45900
rect 131000 45400 131500 57100
rect 145400 48900 145900 49400
rect 127200 44900 131500 45400
rect 127200 44100 127700 44900
<< m3contact >>
rect 143900 129900 145400 130400
rect 53100 116300 54600 116800
rect 143900 116400 145400 116900
rect 44600 102800 46100 103300
rect 143900 102900 145400 103400
rect 143900 89400 145400 89900
rect 143900 75900 145400 76400
rect 143900 62400 145400 62900
rect 45000 48600 48600 49500
rect 143900 48900 145400 49400
<< metal3 >>
rect 45600 130900 56600 131400
rect 45600 103300 46100 130900
rect 143900 120500 144400 129900
rect 133600 120000 144400 120500
rect 133600 116900 140100 117000
rect 133600 116500 143900 116900
rect 139600 116400 143900 116500
rect 54100 104000 54600 116300
rect 133600 112800 139100 113300
rect 133600 109300 138100 109800
rect 133400 106900 137100 107300
rect 133400 106100 136100 106500
rect 133400 105300 135100 105700
rect 54100 103500 56800 104000
rect 56500 103300 56800 103500
rect 47700 102400 56700 102800
rect 47700 101700 55300 102400
rect 47700 49500 48600 101700
rect 134600 49400 135100 105300
rect 135600 62900 136100 106100
rect 136600 76400 137100 106900
rect 137600 89900 138100 109300
rect 138600 103400 139100 112800
rect 138600 102900 143900 103400
rect 137600 89400 143900 89900
rect 136600 75900 143900 76400
rect 135600 62400 143900 62900
rect 134600 48900 143900 49400
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0
timestamp 1569525083
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569525083
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569525083
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569525083
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569525083
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569525083
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569525083
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569525083
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use output_terminal_Core  output_terminal_Core_0
timestamp 1740696072
transform 1 0 56910 0 1 57390
box -930 -360 77130 76545
use PVDD  PAD_1_VDD
timestamp 1569525083
transform 0 1 18900 -1 0 141500
box 0 -9150 12000 25300
use PIC  PAD_2_Rdy
timestamp 1569525083
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  PAD_3_ISin
timestamp 1569525083
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  PAD_4_none
timestamp 1569525083
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  PAD_5_none
timestamp 1569525083
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  PAD_6_none
timestamp 1569525083
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PIC  PAD_7_clk
timestamp 1569525083
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PIC  PAD_8_Xin1
timestamp 1569525083
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_9_Xin0
timestamp 1569525083
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_10_Yin1
timestamp 1569525083
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_11_Yin0
timestamp 1569525083
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_12_selXY
timestamp 1569525083
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_13_selSign
timestamp 1569525083
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  PAD_14_none
timestamp 1569525083
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use POB8  PAD_15_Dout0
timestamp 1569525083
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use POB8  PAD_16_Dout1
timestamp 1569525083
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use POB8  PAD_17_Dout2
timestamp 1569525083
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  PAD_18_Dout3
timestamp 1569525083
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use POB8  PAD_19_Dout4
timestamp 1569525083
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  PAD_20_Dout5
timestamp 1569525083
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  PAD_21_Dout6
timestamp 1569525083
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB8  PAD_22_Dout7
timestamp 1569525083
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use POB8  PAD_23_Dout8
timestamp 1569525083
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use POB8  PAD_24_Dout9
timestamp 1569525083
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB8  PAD_25_Dout10
timestamp 1569525083
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  PAD_26_Dout11
timestamp 1569525083
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8  PAD_27_Vld
timestamp 1569525083
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PVSS  PAD_28_VSS
timestamp 1569525083
transform 1 0 48500 0 -1 171100
box 0 -9150 12000 25300
use PCORNER  PCORNER_0
timestamp 1569525083
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569525083
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569525083
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569525083
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
<< end >>
