magic
tech scmos
magscale 1 3
timestamp 1569543463
<< checkpaint >>
rect -60 -60 910 910
<< metal1 >>
rect 0 825 850 850
rect 0 25 25 825
rect 825 25 850 825
rect 0 0 850 25
<< metal2 >>
rect 0 825 850 850
rect 0 25 25 825
rect 825 25 850 825
rect 0 0 850 25
<< metal3 >>
rect 0 825 850 850
rect 0 25 25 825
rect 825 25 850 825
rect 0 0 850 25
<< pad >>
rect 25 25 825 825
use via1_array_CDNS_704676826051$1  via1_array_CDNS_704676826051$1_0
array 0 19 40 0 19 40
timestamp 1569543463
transform 1 0 35 0 1 35
box 0 0 20 20
use via2_array_CDNS_704676826052$1  via2_array_CDNS_704676826052$1_0
array 0 18 40 0 18 40
timestamp 1569543463
transform 1 0 55 0 1 55
box 0 0 20 20
<< end >>
