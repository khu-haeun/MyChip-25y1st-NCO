magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -140 -140 2539 620
<< nwell >>
rect -20 -20 2419 220
<< psubstratepdiff >>
rect 0 300 2400 500
<< nsubstratendiff >>
rect 0 0 2400 200
<< metal1 >>
rect 0 300 2400 500
rect 0 0 2400 200
use CONT$3  CONT$3_0
array 0 61 36 0 4 36
timestamp 1569543463
transform 1 0 164 0 1 325
box -6 -6 6 6
use CONT$3  CONT$3_1
array 0 61 36 0 4 36
timestamp 1569543463
transform 1 0 56 0 1 31
box -6 -6 6 6
<< end >>
