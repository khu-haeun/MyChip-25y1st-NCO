magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -120 -1950 2520 5180
<< metal2 >>
rect 516 5032 1884 5060
use METAL_RING$2  METAL_RING$2_0
timestamp 1569543463
transform 1 0 0 0 1 0
box 0 0 2400 5012
use NDRV$1  NDRV$1_0
timestamp 1569543463
transform 1 0 0 0 1 0
box 0 0 2400 1560
use NDRV1$2  NDRV1$2_0
timestamp 1569543463
transform 1 0 252 0 1 3120
box 0 0 1896 1560
use NDRV1$2  NDRV1$2_1
timestamp 1569543463
transform 1 0 252 0 1 1560
box 0 0 1896 1560
use PAD_80$2  PAD_80$2_0
timestamp 1569543463
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_PVDD$1  PAD_METAL_PVDD$1_0
timestamp 1569543463
transform 1 0 0 0 1 0
box 0 0 2400 5060
<< labels >>
flabel m2p s 1175 5060 1175 5060 0 FreeSans 1000 0 0 0 VDD
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 700 0 700 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 4755 0 4755 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 4400 0 4400 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 3000 0 3000 0 FreeSans 1000 0 0 0 VDD
<< end >>
