/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module output_terminal(
    output [11:0] Dout,
    input ISin,
    input Rdy,
    output Vld,
    input [1:0] Xin,
    input [1:0] Yin,
    input clk,
    input selSign,
    input selXY
);

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire [6:0] LoadCtl ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire ISin ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _256_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _48_ ;
wire _121_ ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire _118_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire _212_ ;
wire _250_ ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire ISreg_bF$buf0 ;
wire ISreg_bF$buf1 ;
wire ISreg_bF$buf2 ;
wire ISreg_bF$buf3 ;
wire ISreg_bF$buf4 ;
wire _80_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _147_ ;
wire _185_ ;
wire selXY ;
wire selSign ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire [11:0] Ycalc ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _96__bF$buf0 ;
wire _96__bF$buf1 ;
wire _96__bF$buf2 ;
wire _96__bF$buf3 ;
wire _96__bF$buf4 ;
wire _138_ ;
wire _30_ ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire ISreg ;
wire _264_ ;
wire [11:0] Dout ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire [11:0] Xin12b ;
wire [1:0] Yin ;
wire _255_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire [11:0] Xcalc ;
wire [1:0] Yin0 ;
wire [1:0] Yin1 ;
wire _214_ ;
wire _252_ ;
wire _117_ ;
wire _155_ ;
wire _193_ ;
wire _249_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire [1:0] Xin0 ;
wire [1:0] Xin1 ;
wire _114_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire _146_ ;
wire _184_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire [11:0] _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire LoadCtl_6_bF$buf0 ;
wire LoadCtl_6_bF$buf1 ;
wire LoadCtl_6_bF$buf2 ;
wire LoadCtl_6_bF$buf3 ;
wire LoadCtl_6_bF$buf4 ;
wire _119_ ;
wire _11_ ;
wire [11:0] Yin12b ;
wire _157_ ;
wire _195_ ;
wire _5_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _116_ ;
wire _154_ ;
wire _192_ ;
wire _248_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire [1:0] Xin ;
wire _245_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

BUFX2 BUFX2_insert25 (
    .A(_96_),
    .Y(_96__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .A(_96_),
    .Y(_96__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .A(_96_),
    .Y(_96__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .A(_96_),
    .Y(_96__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .A(_96_),
    .Y(_96__bF$buf4)
);

BUFX2 BUFX2_insert20 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf4)
);

BUFX2 BUFX2_insert15 (
    .A(ISreg),
    .Y(ISreg_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(ISreg),
    .Y(ISreg_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(ISreg),
    .Y(ISreg_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(ISreg),
    .Y(ISreg_bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(ISreg),
    .Y(ISreg_bF$buf4)
);

BUFX2 BUFX2_insert10 (
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .A(selXY),
    .Y(selXY_bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .A(selXY),
    .Y(selXY_bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .A(selXY),
    .Y(selXY_bF$buf3)
);

CLKBUF1 CLKBUF1_insert6 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf6)
);

INVX1 _273_ (
    .A(Ycalc[0]),
    .Y(_49_)
);

NAND2X1 _274_ (
    .A(Xcalc[0]),
    .B(selXY_bF$buf3),
    .Y(_50_)
);

OAI21X1 _275_ (
    .A(selXY_bF$buf2),
    .B(_49_),
    .C(_50_),
    .Y(_272_[0])
);

INVX1 _276_ (
    .A(Ycalc[1]),
    .Y(_51_)
);

NAND2X1 _277_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[1]),
    .Y(_52_)
);

OAI21X1 _278_ (
    .A(selXY_bF$buf0),
    .B(_51_),
    .C(_52_),
    .Y(_272_[1])
);

INVX1 _279_ (
    .A(Ycalc[2]),
    .Y(_53_)
);

NAND2X1 _280_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[2]),
    .Y(_54_)
);

OAI21X1 _281_ (
    .A(selXY_bF$buf2),
    .B(_53_),
    .C(_54_),
    .Y(_272_[2])
);

INVX1 _282_ (
    .A(Ycalc[3]),
    .Y(_55_)
);

NAND2X1 _283_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[3]),
    .Y(_56_)
);

OAI21X1 _284_ (
    .A(selXY_bF$buf0),
    .B(_55_),
    .C(_56_),
    .Y(_272_[3])
);

INVX1 _285_ (
    .A(Ycalc[4]),
    .Y(_57_)
);

NAND2X1 _286_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[4]),
    .Y(_58_)
);

OAI21X1 _287_ (
    .A(selXY_bF$buf2),
    .B(_57_),
    .C(_58_),
    .Y(_272_[4])
);

INVX1 _288_ (
    .A(Ycalc[5]),
    .Y(_59_)
);

NAND2X1 _289_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[5]),
    .Y(_60_)
);

OAI21X1 _290_ (
    .A(selXY_bF$buf0),
    .B(_59_),
    .C(_60_),
    .Y(_272_[5])
);

INVX1 _291_ (
    .A(Ycalc[6]),
    .Y(_61_)
);

NAND2X1 _292_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[6]),
    .Y(_62_)
);

OAI21X1 _293_ (
    .A(selXY_bF$buf2),
    .B(_61_),
    .C(_62_),
    .Y(_272_[6])
);

INVX1 _294_ (
    .A(Ycalc[7]),
    .Y(_63_)
);

NAND2X1 _295_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[7]),
    .Y(_64_)
);

OAI21X1 _296_ (
    .A(selXY_bF$buf0),
    .B(_63_),
    .C(_64_),
    .Y(_272_[7])
);

INVX1 _297_ (
    .A(Ycalc[8]),
    .Y(_65_)
);

NAND2X1 _298_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[8]),
    .Y(_66_)
);

OAI21X1 _299_ (
    .A(selXY_bF$buf2),
    .B(_65_),
    .C(_66_),
    .Y(_272_[8])
);

INVX1 _300_ (
    .A(Ycalc[9]),
    .Y(_67_)
);

NAND2X1 _301_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[9]),
    .Y(_68_)
);

OAI21X1 _302_ (
    .A(selXY_bF$buf0),
    .B(_67_),
    .C(_68_),
    .Y(_272_[9])
);

INVX1 _303_ (
    .A(Ycalc[10]),
    .Y(_69_)
);

NAND2X1 _304_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[10]),
    .Y(_70_)
);

OAI21X1 _305_ (
    .A(selXY_bF$buf2),
    .B(_69_),
    .C(_70_),
    .Y(_272_[10])
);

INVX1 _306_ (
    .A(Ycalc[11]),
    .Y(_71_)
);

NAND2X1 _307_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[11]),
    .Y(_72_)
);

OAI21X1 _308_ (
    .A(selXY_bF$buf0),
    .B(_71_),
    .C(_72_),
    .Y(_272_[11])
);

INVX1 _309_ (
    .A(Yin[1]),
    .Y(_73_)
);

INVX1 _310_ (
    .A(LoadCtl[2]),
    .Y(_74_)
);

NOR2X1 _311_ (
    .A(LoadCtl[0]),
    .B(LoadCtl[1]),
    .Y(_75_)
);

NAND3X1 _312_ (
    .A(_74_),
    .B(LoadCtl[3]),
    .C(_75_),
    .Y(_76_)
);

NAND2X1 _313_ (
    .A(Yin12b[7]),
    .B(_76_),
    .Y(_77_)
);

OAI21X1 _314_ (
    .A(_73_),
    .B(_76_),
    .C(_77_),
    .Y(_1_)
);

INVX1 _315_ (
    .A(Yin12b[4]),
    .Y(_78_)
);

INVX1 _316_ (
    .A(_75_),
    .Y(_79_)
);

NOR2X1 _317_ (
    .A(_74_),
    .B(_79_),
    .Y(_80_)
);

NAND2X1 _318_ (
    .A(Yin[0]),
    .B(_80_),
    .Y(_81_)
);

OAI21X1 _319_ (
    .A(_78_),
    .B(_80_),
    .C(_81_),
    .Y(_2_)
);

INVX1 _320_ (
    .A(Yin12b[5]),
    .Y(_82_)
);

NAND2X1 _321_ (
    .A(Yin[1]),
    .B(_80_),
    .Y(_83_)
);

OAI21X1 _322_ (
    .A(_82_),
    .B(_80_),
    .C(_83_),
    .Y(_3_)
);

INVX1 _323_ (
    .A(Yin[0]),
    .Y(_84_)
);

INVX2 _324_ (
    .A(LoadCtl[1]),
    .Y(_85_)
);

OR2X2 _325_ (
    .A(_85_),
    .B(LoadCtl[0]),
    .Y(_86_)
);

OAI21X1 _326_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[0]),
    .Y(_87_)
);

OAI21X1 _327_ (
    .A(_84_),
    .B(_86_),
    .C(_87_),
    .Y(_4_)
);

OAI21X1 _328_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[1]),
    .Y(_88_)
);

OAI21X1 _329_ (
    .A(_73_),
    .B(_86_),
    .C(_88_),
    .Y(_5_)
);

INVX1 _330_ (
    .A(Yin0[0]),
    .Y(_89_)
);

NAND2X1 _331_ (
    .A(LoadCtl[0]),
    .B(Yin[0]),
    .Y(_90_)
);

OAI21X1 _332_ (
    .A(LoadCtl[0]),
    .B(_89_),
    .C(_90_),
    .Y(_6_)
);

INVX1 _333_ (
    .A(Yin0[1]),
    .Y(_91_)
);

NAND2X1 _334_ (
    .A(LoadCtl[0]),
    .B(Yin[1]),
    .Y(_92_)
);

OAI21X1 _335_ (
    .A(LoadCtl[0]),
    .B(_91_),
    .C(_92_),
    .Y(_7_)
);

INVX4 _336_ (
    .A(ISreg_bF$buf4),
    .Y(_93_)
);

NAND2X1 _337_ (
    .A(ISin),
    .B(LoadCtl_6_bF$buf4),
    .Y(_94_)
);

OAI21X1 _338_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_93_),
    .C(_94_),
    .Y(_8_)
);

INVX1 _339_ (
    .A(Xin0[0]),
    .Y(_95_)
);

INVX8 _340_ (
    .A(LoadCtl_6_bF$buf2),
    .Y(_96_)
);

NAND2X1 _341_ (
    .A(Xcalc[0]),
    .B(_96__bF$buf4),
    .Y(_97_)
);

OAI21X1 _342_ (
    .A(_95_),
    .B(_96__bF$buf3),
    .C(_97_),
    .Y(_9_)
);

NAND3X1 _343_ (
    .A(ISreg_bF$buf3),
    .B(Xin0[0]),
    .C(Xin0[1]),
    .Y(_98_)
);

INVX1 _344_ (
    .A(Xin0[1]),
    .Y(_99_)
);

OAI21X1 _345_ (
    .A(_93_),
    .B(_95_),
    .C(_99_),
    .Y(_100_)
);

NAND2X1 _346_ (
    .A(_98_),
    .B(_100_),
    .Y(_101_)
);

NAND2X1 _347_ (
    .A(Xcalc[1]),
    .B(_96__bF$buf2),
    .Y(_102_)
);

OAI21X1 _348_ (
    .A(_96__bF$buf1),
    .B(_101_),
    .C(_102_),
    .Y(_10_)
);

INVX1 _349_ (
    .A(Xin1[0]),
    .Y(_103_)
);

OAI21X1 _350_ (
    .A(Xin0[0]),
    .B(Xin0[1]),
    .C(ISreg_bF$buf2),
    .Y(_104_)
);

OR2X2 _351_ (
    .A(_104_),
    .B(_103_),
    .Y(_105_)
);

NOR2X1 _352_ (
    .A(Xin0[0]),
    .B(Xin0[1]),
    .Y(_106_)
);

OAI21X1 _353_ (
    .A(_93_),
    .B(_106_),
    .C(_103_),
    .Y(_107_)
);

NAND2X1 _354_ (
    .A(_107_),
    .B(_105_),
    .Y(_108_)
);

NAND2X1 _355_ (
    .A(Xcalc[2]),
    .B(_96__bF$buf0),
    .Y(_109_)
);

OAI21X1 _356_ (
    .A(_96__bF$buf4),
    .B(_108_),
    .C(_109_),
    .Y(_11_)
);

OAI21X1 _357_ (
    .A(_93_),
    .B(_103_),
    .C(_104_),
    .Y(_110_)
);

NAND2X1 _358_ (
    .A(Xin1[1]),
    .B(_110_),
    .Y(_111_)
);

OR2X2 _359_ (
    .A(_110_),
    .B(Xin1[1]),
    .Y(_112_)
);

NAND2X1 _360_ (
    .A(_111_),
    .B(_112_),
    .Y(_113_)
);

NAND2X1 _361_ (
    .A(Xcalc[3]),
    .B(_96__bF$buf3),
    .Y(_114_)
);

OAI21X1 _362_ (
    .A(_96__bF$buf2),
    .B(_113_),
    .C(_114_),
    .Y(_12_)
);

NOR2X1 _363_ (
    .A(Xin1[0]),
    .B(Xin1[1]),
    .Y(_115_)
);

NAND2X1 _364_ (
    .A(_106_),
    .B(_115_),
    .Y(_116_)
);

NAND3X1 _365_ (
    .A(ISreg_bF$buf1),
    .B(Xin12b[4]),
    .C(_116_),
    .Y(_117_)
);

INVX1 _366_ (
    .A(Xin12b[4]),
    .Y(_118_)
);

AND2X2 _367_ (
    .A(_106_),
    .B(_115_),
    .Y(_119_)
);

OAI21X1 _368_ (
    .A(_93_),
    .B(_119_),
    .C(_118_),
    .Y(_120_)
);

NAND2X1 _369_ (
    .A(_117_),
    .B(_120_),
    .Y(_121_)
);

NAND2X1 _370_ (
    .A(Xcalc[4]),
    .B(_96__bF$buf1),
    .Y(_122_)
);

OAI21X1 _371_ (
    .A(_96__bF$buf0),
    .B(_121_),
    .C(_122_),
    .Y(_13_)
);

INVX1 _372_ (
    .A(Xin12b[5]),
    .Y(_123_)
);

OAI21X1 _373_ (
    .A(Xin12b[4]),
    .B(_116_),
    .C(ISreg_bF$buf0),
    .Y(_124_)
);

OR2X2 _374_ (
    .A(_124_),
    .B(_123_),
    .Y(_125_)
);

NAND2X1 _375_ (
    .A(_123_),
    .B(_124_),
    .Y(_126_)
);

NAND2X1 _376_ (
    .A(_126_),
    .B(_125_),
    .Y(_127_)
);

NAND2X1 _377_ (
    .A(Xcalc[5]),
    .B(_96__bF$buf4),
    .Y(_128_)
);

OAI21X1 _378_ (
    .A(_96__bF$buf3),
    .B(_127_),
    .C(_128_),
    .Y(_14_)
);

NOR2X1 _379_ (
    .A(Xin12b[4]),
    .B(Xin12b[5]),
    .Y(_129_)
);

NAND2X1 _380_ (
    .A(_129_),
    .B(_119_),
    .Y(_130_)
);

NAND3X1 _381_ (
    .A(ISreg_bF$buf4),
    .B(Xin12b[6]),
    .C(_130_),
    .Y(_131_)
);

INVX1 _382_ (
    .A(Xin12b[6]),
    .Y(_132_)
);

NAND2X1 _383_ (
    .A(ISreg_bF$buf3),
    .B(_130_),
    .Y(_133_)
);

NAND2X1 _384_ (
    .A(_132_),
    .B(_133_),
    .Y(_134_)
);

NAND2X1 _385_ (
    .A(_131_),
    .B(_134_),
    .Y(_135_)
);

NAND2X1 _386_ (
    .A(Xcalc[6]),
    .B(_96__bF$buf2),
    .Y(_136_)
);

OAI21X1 _387_ (
    .A(_96__bF$buf1),
    .B(_135_),
    .C(_136_),
    .Y(_15_)
);

INVX1 _388_ (
    .A(Xcalc[7]),
    .Y(_137_)
);

NAND3X1 _389_ (
    .A(_132_),
    .B(_129_),
    .C(_119_),
    .Y(_138_)
);

NAND3X1 _390_ (
    .A(ISreg_bF$buf2),
    .B(Xin12b[7]),
    .C(_138_),
    .Y(_139_)
);

INVX1 _391_ (
    .A(Xin12b[7]),
    .Y(_140_)
);

NAND2X1 _392_ (
    .A(ISreg_bF$buf1),
    .B(Xin12b[6]),
    .Y(_141_)
);

NAND3X1 _393_ (
    .A(_140_),
    .B(_141_),
    .C(_133_),
    .Y(_142_)
);

NAND3X1 _394_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_139_),
    .C(_142_),
    .Y(_143_)
);

OAI21X1 _395_ (
    .A(_137_),
    .B(LoadCtl_6_bF$buf0),
    .C(_143_),
    .Y(_16_)
);

INVX1 _396_ (
    .A(Xin12b[8]),
    .Y(_144_)
);

NOR2X1 _397_ (
    .A(Xin12b[6]),
    .B(Xin12b[7]),
    .Y(_145_)
);

NAND2X1 _398_ (
    .A(_129_),
    .B(_145_),
    .Y(_146_)
);

OAI21X1 _399_ (
    .A(_116_),
    .B(_146_),
    .C(ISreg_bF$buf0),
    .Y(_147_)
);

OR2X2 _400_ (
    .A(_147_),
    .B(_144_),
    .Y(_148_)
);

NAND2X1 _401_ (
    .A(_144_),
    .B(_147_),
    .Y(_149_)
);

NAND2X1 _402_ (
    .A(_149_),
    .B(_148_),
    .Y(_150_)
);

NAND2X1 _403_ (
    .A(Xcalc[8]),
    .B(_96__bF$buf0),
    .Y(_151_)
);

OAI21X1 _404_ (
    .A(_96__bF$buf4),
    .B(_150_),
    .C(_151_),
    .Y(_17_)
);

INVX1 _405_ (
    .A(Xcalc[9]),
    .Y(_152_)
);

INVX1 _406_ (
    .A(Xin12b[9]),
    .Y(_153_)
);

OAI21X1 _407_ (
    .A(_93_),
    .B(_144_),
    .C(_147_),
    .Y(_154_)
);

OR2X2 _408_ (
    .A(_154_),
    .B(_153_),
    .Y(_155_)
);

AOI21X1 _409_ (
    .A(_154_),
    .B(_153_),
    .C(_96__bF$buf3),
    .Y(_156_)
);

AOI22X1 _410_ (
    .A(_152_),
    .B(_96__bF$buf2),
    .C(_155_),
    .D(_156_),
    .Y(_18_)
);

INVX1 _411_ (
    .A(Xcalc[10]),
    .Y(_157_)
);

AND2X2 _412_ (
    .A(_129_),
    .B(_145_),
    .Y(_158_)
);

NOR2X1 _413_ (
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .Y(_159_)
);

NAND3X1 _414_ (
    .A(_159_),
    .B(_119_),
    .C(_158_),
    .Y(_160_)
);

NAND3X1 _415_ (
    .A(ISreg_bF$buf4),
    .B(Xin12b[10]),
    .C(_160_),
    .Y(_161_)
);

INVX1 _416_ (
    .A(Xin12b[10]),
    .Y(_162_)
);

NAND2X1 _417_ (
    .A(ISreg_bF$buf3),
    .B(_160_),
    .Y(_163_)
);

NAND2X1 _418_ (
    .A(_162_),
    .B(_163_),
    .Y(_164_)
);

NAND3X1 _419_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_161_),
    .C(_164_),
    .Y(_165_)
);

OAI21X1 _420_ (
    .A(_157_),
    .B(LoadCtl_6_bF$buf3),
    .C(_165_),
    .Y(_19_)
);

NAND2X1 _421_ (
    .A(Xcalc[11]),
    .B(_96__bF$buf1),
    .Y(_166_)
);

INVX1 _422_ (
    .A(Xin12b[11]),
    .Y(_167_)
);

NAND2X1 _423_ (
    .A(selSign),
    .B(_167_),
    .Y(_168_)
);

INVX1 _424_ (
    .A(selSign),
    .Y(_169_)
);

NAND2X1 _425_ (
    .A(Xin12b[11]),
    .B(_169_),
    .Y(_170_)
);

NAND2X1 _426_ (
    .A(_168_),
    .B(_170_),
    .Y(_171_)
);

INVX1 _427_ (
    .A(_171_),
    .Y(_172_)
);

NAND2X1 _428_ (
    .A(ISreg_bF$buf2),
    .B(Xin12b[10]),
    .Y(_173_)
);

NAND3X1 _429_ (
    .A(_172_),
    .B(_173_),
    .C(_163_),
    .Y(_174_)
);

OAI21X1 _430_ (
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .C(ISreg_bF$buf1),
    .Y(_175_)
);

NAND3X1 _431_ (
    .A(_175_),
    .B(_173_),
    .C(_147_),
    .Y(_176_)
);

NAND2X1 _432_ (
    .A(_171_),
    .B(_176_),
    .Y(_177_)
);

NAND3X1 _433_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_177_),
    .C(_174_),
    .Y(_178_)
);

NAND2X1 _434_ (
    .A(_166_),
    .B(_178_),
    .Y(_20_)
);

NAND2X1 _435_ (
    .A(Yin0[0]),
    .B(LoadCtl_6_bF$buf1),
    .Y(_179_)
);

OAI21X1 _436_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_49_),
    .C(_179_),
    .Y(_21_)
);

NAND3X1 _437_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf0),
    .Y(_180_)
);

OAI21X1 _438_ (
    .A(_89_),
    .B(_93_),
    .C(_91_),
    .Y(_181_)
);

NAND3X1 _439_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_180_),
    .C(_181_),
    .Y(_182_)
);

OAI21X1 _440_ (
    .A(_51_),
    .B(LoadCtl_6_bF$buf3),
    .C(_182_),
    .Y(_22_)
);

INVX1 _441_ (
    .A(Yin1[0]),
    .Y(_183_)
);

OAI21X1 _442_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf4),
    .Y(_184_)
);

OR2X2 _443_ (
    .A(_184_),
    .B(_183_),
    .Y(_185_)
);

NOR2X1 _444_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .Y(_186_)
);

OAI21X1 _445_ (
    .A(_93_),
    .B(_186_),
    .C(_183_),
    .Y(_187_)
);

NAND3X1 _446_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_187_),
    .C(_185_),
    .Y(_188_)
);

OAI21X1 _447_ (
    .A(_53_),
    .B(LoadCtl_6_bF$buf1),
    .C(_188_),
    .Y(_23_)
);

OAI21X1 _448_ (
    .A(_93_),
    .B(_183_),
    .C(_184_),
    .Y(_189_)
);

NAND2X1 _449_ (
    .A(Yin1[1]),
    .B(_189_),
    .Y(_190_)
);

OR2X2 _450_ (
    .A(_189_),
    .B(Yin1[1]),
    .Y(_191_)
);

NAND3X1 _451_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_190_),
    .C(_191_),
    .Y(_192_)
);

OAI21X1 _452_ (
    .A(_55_),
    .B(LoadCtl_6_bF$buf4),
    .C(_192_),
    .Y(_24_)
);

NOR2X1 _453_ (
    .A(Yin1[0]),
    .B(Yin1[1]),
    .Y(_193_)
);

NAND2X1 _454_ (
    .A(_186_),
    .B(_193_),
    .Y(_194_)
);

NAND2X1 _455_ (
    .A(ISreg_bF$buf3),
    .B(_194_),
    .Y(_195_)
);

OR2X2 _456_ (
    .A(_195_),
    .B(_78_),
    .Y(_196_)
);

AND2X2 _457_ (
    .A(_186_),
    .B(_193_),
    .Y(_197_)
);

OAI21X1 _458_ (
    .A(_93_),
    .B(_197_),
    .C(_78_),
    .Y(_198_)
);

NAND3X1 _459_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_198_),
    .C(_196_),
    .Y(_199_)
);

OAI21X1 _460_ (
    .A(_57_),
    .B(LoadCtl_6_bF$buf2),
    .C(_199_),
    .Y(_25_)
);

OAI21X1 _461_ (
    .A(_93_),
    .B(_78_),
    .C(_195_),
    .Y(_200_)
);

OR2X2 _462_ (
    .A(_200_),
    .B(_82_),
    .Y(_201_)
);

AOI21X1 _463_ (
    .A(_200_),
    .B(_82_),
    .C(_96__bF$buf0),
    .Y(_202_)
);

AOI22X1 _464_ (
    .A(_59_),
    .B(_96__bF$buf4),
    .C(_201_),
    .D(_202_),
    .Y(_26_)
);

NOR2X1 _465_ (
    .A(Yin12b[4]),
    .B(Yin12b[5]),
    .Y(_203_)
);

NAND2X1 _466_ (
    .A(_203_),
    .B(_197_),
    .Y(_204_)
);

NAND3X1 _467_ (
    .A(ISreg_bF$buf2),
    .B(Yin12b[6]),
    .C(_204_),
    .Y(_205_)
);

INVX1 _468_ (
    .A(Yin12b[6]),
    .Y(_206_)
);

NAND2X1 _469_ (
    .A(ISreg_bF$buf1),
    .B(_204_),
    .Y(_207_)
);

NAND2X1 _470_ (
    .A(_206_),
    .B(_207_),
    .Y(_208_)
);

NAND3X1 _471_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_205_),
    .C(_208_),
    .Y(_209_)
);

OAI21X1 _472_ (
    .A(_61_),
    .B(LoadCtl_6_bF$buf0),
    .C(_209_),
    .Y(_27_)
);

NAND3X1 _473_ (
    .A(_206_),
    .B(_203_),
    .C(_197_),
    .Y(_210_)
);

NAND3X1 _474_ (
    .A(ISreg_bF$buf0),
    .B(Yin12b[7]),
    .C(_210_),
    .Y(_211_)
);

INVX1 _475_ (
    .A(Yin12b[7]),
    .Y(_212_)
);

NAND2X1 _476_ (
    .A(ISreg_bF$buf4),
    .B(Yin12b[6]),
    .Y(_213_)
);

NAND3X1 _477_ (
    .A(_212_),
    .B(_213_),
    .C(_207_),
    .Y(_214_)
);

NAND3X1 _478_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_211_),
    .C(_214_),
    .Y(_215_)
);

OAI21X1 _479_ (
    .A(_63_),
    .B(LoadCtl_6_bF$buf3),
    .C(_215_),
    .Y(_28_)
);

INVX1 _480_ (
    .A(Yin12b[8]),
    .Y(_216_)
);

NOR2X1 _481_ (
    .A(Yin12b[6]),
    .B(Yin12b[7]),
    .Y(_217_)
);

NAND2X1 _482_ (
    .A(_203_),
    .B(_217_),
    .Y(_218_)
);

OAI21X1 _483_ (
    .A(_194_),
    .B(_218_),
    .C(ISreg_bF$buf3),
    .Y(_219_)
);

OR2X2 _484_ (
    .A(_219_),
    .B(_216_),
    .Y(_220_)
);

NAND2X1 _485_ (
    .A(_216_),
    .B(_219_),
    .Y(_221_)
);

NAND2X1 _486_ (
    .A(_221_),
    .B(_220_),
    .Y(_222_)
);

NAND2X1 _487_ (
    .A(Ycalc[8]),
    .B(_96__bF$buf3),
    .Y(_223_)
);

OAI21X1 _488_ (
    .A(_96__bF$buf2),
    .B(_222_),
    .C(_223_),
    .Y(_29_)
);

INVX1 _489_ (
    .A(Yin12b[9]),
    .Y(_224_)
);

OAI21X1 _490_ (
    .A(_93_),
    .B(_216_),
    .C(_219_),
    .Y(_225_)
);

OR2X2 _491_ (
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

AOI21X1 _492_ (
    .A(_225_),
    .B(_224_),
    .C(_96__bF$buf1),
    .Y(_227_)
);

AOI22X1 _493_ (
    .A(_67_),
    .B(_96__bF$buf0),
    .C(_226_),
    .D(_227_),
    .Y(_30_)
);

AND2X2 _494_ (
    .A(_203_),
    .B(_217_),
    .Y(_228_)
);

NOR2X1 _495_ (
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .Y(_229_)
);

NAND3X1 _496_ (
    .A(_229_),
    .B(_197_),
    .C(_228_),
    .Y(_230_)
);

NAND3X1 _497_ (
    .A(ISreg_bF$buf2),
    .B(Yin12b[10]),
    .C(_230_),
    .Y(_231_)
);

INVX1 _498_ (
    .A(Yin12b[10]),
    .Y(_232_)
);

NAND2X1 _499_ (
    .A(ISreg_bF$buf1),
    .B(_230_),
    .Y(_233_)
);

NAND2X1 _500_ (
    .A(_232_),
    .B(_233_),
    .Y(_234_)
);

NAND3X1 _501_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_231_),
    .C(_234_),
    .Y(_235_)
);

OAI21X1 _502_ (
    .A(_69_),
    .B(LoadCtl_6_bF$buf1),
    .C(_235_),
    .Y(_31_)
);

NAND2X1 _503_ (
    .A(Ycalc[11]),
    .B(_96__bF$buf4),
    .Y(_236_)
);

INVX1 _504_ (
    .A(Yin12b[11]),
    .Y(_237_)
);

NAND2X1 _505_ (
    .A(selSign),
    .B(_237_),
    .Y(_238_)
);

NAND2X1 _506_ (
    .A(Yin12b[11]),
    .B(_169_),
    .Y(_239_)
);

NAND2X1 _507_ (
    .A(_238_),
    .B(_239_),
    .Y(_240_)
);

INVX1 _508_ (
    .A(_240_),
    .Y(_241_)
);

NAND2X1 _509_ (
    .A(ISreg_bF$buf0),
    .B(Yin12b[10]),
    .Y(_242_)
);

NAND3X1 _510_ (
    .A(_241_),
    .B(_242_),
    .C(_233_),
    .Y(_243_)
);

OAI21X1 _511_ (
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .C(ISreg_bF$buf4),
    .Y(_244_)
);

NAND3X1 _512_ (
    .A(_244_),
    .B(_242_),
    .C(_219_),
    .Y(_245_)
);

NAND2X1 _513_ (
    .A(_240_),
    .B(_245_),
    .Y(_246_)
);

NAND3X1 _514_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_246_),
    .C(_243_),
    .Y(_247_)
);

NAND2X1 _515_ (
    .A(_236_),
    .B(_247_),
    .Y(_32_)
);

NOR2X1 _516_ (
    .A(LoadCtl[2]),
    .B(LoadCtl[3]),
    .Y(_248_)
);

AND2X2 _517_ (
    .A(_75_),
    .B(_248_),
    .Y(_249_)
);

NAND2X1 _518_ (
    .A(LoadCtl[5]),
    .B(_249_),
    .Y(_250_)
);

NOR2X1 _519_ (
    .A(LoadCtl[4]),
    .B(_250_),
    .Y(_251_)
);

NAND2X1 _520_ (
    .A(Xin[0]),
    .B(_251_),
    .Y(_252_)
);

OAI21X1 _521_ (
    .A(_162_),
    .B(_251_),
    .C(_252_),
    .Y(_33_)
);

NAND2X1 _522_ (
    .A(Xin[1]),
    .B(_251_),
    .Y(_253_)
);

OAI21X1 _523_ (
    .A(_167_),
    .B(_251_),
    .C(_253_),
    .Y(_34_)
);

INVX1 _524_ (
    .A(Xin[0]),
    .Y(_254_)
);

NAND2X1 _525_ (
    .A(LoadCtl[4]),
    .B(_249_),
    .Y(_255_)
);

NAND2X1 _526_ (
    .A(Xin12b[8]),
    .B(_255_),
    .Y(_256_)
);

OAI21X1 _527_ (
    .A(_254_),
    .B(_255_),
    .C(_256_),
    .Y(_35_)
);

INVX1 _528_ (
    .A(Xin[1]),
    .Y(_257_)
);

NAND2X1 _529_ (
    .A(Xin12b[9]),
    .B(_255_),
    .Y(_258_)
);

OAI21X1 _530_ (
    .A(_257_),
    .B(_255_),
    .C(_258_),
    .Y(_36_)
);

NAND2X1 _531_ (
    .A(Xin12b[6]),
    .B(_76_),
    .Y(_259_)
);

OAI21X1 _532_ (
    .A(_254_),
    .B(_76_),
    .C(_259_),
    .Y(_37_)
);

NAND2X1 _533_ (
    .A(Xin12b[7]),
    .B(_76_),
    .Y(_260_)
);

OAI21X1 _534_ (
    .A(_257_),
    .B(_76_),
    .C(_260_),
    .Y(_38_)
);

NAND2X1 _535_ (
    .A(Xin[0]),
    .B(_80_),
    .Y(_261_)
);

OAI21X1 _536_ (
    .A(_118_),
    .B(_80_),
    .C(_261_),
    .Y(_39_)
);

NAND2X1 _537_ (
    .A(Xin[1]),
    .B(_80_),
    .Y(_262_)
);

OAI21X1 _538_ (
    .A(_123_),
    .B(_80_),
    .C(_262_),
    .Y(_40_)
);

OAI21X1 _539_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[0]),
    .Y(_263_)
);

OAI21X1 _540_ (
    .A(_254_),
    .B(_86_),
    .C(_263_),
    .Y(_41_)
);

OAI21X1 _541_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[1]),
    .Y(_264_)
);

OAI21X1 _542_ (
    .A(_257_),
    .B(_86_),
    .C(_264_),
    .Y(_42_)
);

NAND2X1 _543_ (
    .A(LoadCtl[0]),
    .B(Xin[0]),
    .Y(_265_)
);

OAI21X1 _544_ (
    .A(LoadCtl[0]),
    .B(_95_),
    .C(_265_),
    .Y(_43_)
);

NAND2X1 _545_ (
    .A(LoadCtl[0]),
    .B(Xin[1]),
    .Y(_266_)
);

OAI21X1 _546_ (
    .A(LoadCtl[0]),
    .B(_99_),
    .C(_266_),
    .Y(_44_)
);

NAND2X1 _547_ (
    .A(Yin[0]),
    .B(_251_),
    .Y(_267_)
);

OAI21X1 _548_ (
    .A(_232_),
    .B(_251_),
    .C(_267_),
    .Y(_45_)
);

NAND2X1 _549_ (
    .A(Yin[1]),
    .B(_251_),
    .Y(_268_)
);

OAI21X1 _550_ (
    .A(_237_),
    .B(_251_),
    .C(_268_),
    .Y(_46_)
);

NAND2X1 _551_ (
    .A(Yin12b[8]),
    .B(_255_),
    .Y(_269_)
);

OAI21X1 _552_ (
    .A(_84_),
    .B(_255_),
    .C(_269_),
    .Y(_47_)
);

NAND2X1 _553_ (
    .A(Yin12b[9]),
    .B(_255_),
    .Y(_270_)
);

OAI21X1 _554_ (
    .A(_73_),
    .B(_255_),
    .C(_270_),
    .Y(_48_)
);

NAND2X1 _555_ (
    .A(Yin12b[6]),
    .B(_76_),
    .Y(_271_)
);

OAI21X1 _556_ (
    .A(_84_),
    .B(_76_),
    .C(_271_),
    .Y(_0_)
);

DFFPOSX1 _557_ (
    .CLK(clk_bF$buf6),
    .D(_8_),
    .Q(ISreg)
);

DFFPOSX1 _558_ (
    .CLK(clk_bF$buf5),
    .D(_9_),
    .Q(Xcalc[0])
);

DFFPOSX1 _559_ (
    .CLK(clk_bF$buf4),
    .D(_10_),
    .Q(Xcalc[1])
);

DFFPOSX1 _560_ (
    .CLK(clk_bF$buf3),
    .D(_11_),
    .Q(Xcalc[2])
);

DFFPOSX1 _561_ (
    .CLK(clk_bF$buf2),
    .D(_12_),
    .Q(Xcalc[3])
);

DFFPOSX1 _562_ (
    .CLK(clk_bF$buf1),
    .D(_13_),
    .Q(Xcalc[4])
);

DFFPOSX1 _563_ (
    .CLK(clk_bF$buf0),
    .D(_14_),
    .Q(Xcalc[5])
);

DFFPOSX1 _564_ (
    .CLK(clk_bF$buf6),
    .D(_15_),
    .Q(Xcalc[6])
);

DFFPOSX1 _565_ (
    .CLK(clk_bF$buf5),
    .D(_16_),
    .Q(Xcalc[7])
);

DFFPOSX1 _566_ (
    .CLK(clk_bF$buf4),
    .D(_17_),
    .Q(Xcalc[8])
);

DFFPOSX1 _567_ (
    .CLK(clk_bF$buf3),
    .D(_18_),
    .Q(Xcalc[9])
);

DFFPOSX1 _568_ (
    .CLK(clk_bF$buf2),
    .D(_19_),
    .Q(Xcalc[10])
);

DFFPOSX1 _569_ (
    .CLK(clk_bF$buf1),
    .D(_20_),
    .Q(Xcalc[11])
);

DFFPOSX1 _570_ (
    .CLK(clk_bF$buf0),
    .D(_21_),
    .Q(Ycalc[0])
);

DFFPOSX1 _571_ (
    .CLK(clk_bF$buf6),
    .D(_22_),
    .Q(Ycalc[1])
);

DFFPOSX1 _572_ (
    .CLK(clk_bF$buf5),
    .D(_23_),
    .Q(Ycalc[2])
);

DFFPOSX1 _573_ (
    .CLK(clk_bF$buf4),
    .D(_24_),
    .Q(Ycalc[3])
);

DFFPOSX1 _574_ (
    .CLK(clk_bF$buf3),
    .D(_25_),
    .Q(Ycalc[4])
);

DFFPOSX1 _575_ (
    .CLK(clk_bF$buf2),
    .D(_26_),
    .Q(Ycalc[5])
);

DFFPOSX1 _576_ (
    .CLK(clk_bF$buf1),
    .D(_27_),
    .Q(Ycalc[6])
);

DFFPOSX1 _577_ (
    .CLK(clk_bF$buf0),
    .D(_28_),
    .Q(Ycalc[7])
);

DFFPOSX1 _578_ (
    .CLK(clk_bF$buf6),
    .D(_29_),
    .Q(Ycalc[8])
);

DFFPOSX1 _579_ (
    .CLK(clk_bF$buf5),
    .D(_30_),
    .Q(Ycalc[9])
);

DFFPOSX1 _580_ (
    .CLK(clk_bF$buf4),
    .D(_31_),
    .Q(Ycalc[10])
);

DFFPOSX1 _581_ (
    .CLK(clk_bF$buf3),
    .D(_32_),
    .Q(Ycalc[11])
);

DFFPOSX1 _582_ (
    .CLK(clk_bF$buf2),
    .D(_33_),
    .Q(Xin12b[10])
);

DFFPOSX1 _583_ (
    .CLK(clk_bF$buf1),
    .D(_34_),
    .Q(Xin12b[11])
);

DFFPOSX1 _584_ (
    .CLK(clk_bF$buf0),
    .D(_35_),
    .Q(Xin12b[8])
);

DFFPOSX1 _585_ (
    .CLK(clk_bF$buf6),
    .D(_36_),
    .Q(Xin12b[9])
);

DFFPOSX1 _586_ (
    .CLK(clk_bF$buf5),
    .D(_37_),
    .Q(Xin12b[6])
);

DFFPOSX1 _587_ (
    .CLK(clk_bF$buf4),
    .D(_38_),
    .Q(Xin12b[7])
);

DFFPOSX1 _588_ (
    .CLK(clk_bF$buf3),
    .D(_39_),
    .Q(Xin12b[4])
);

DFFPOSX1 _589_ (
    .CLK(clk_bF$buf2),
    .D(_40_),
    .Q(Xin12b[5])
);

DFFPOSX1 _590_ (
    .CLK(clk_bF$buf1),
    .D(_41_),
    .Q(Xin1[0])
);

DFFPOSX1 _591_ (
    .CLK(clk_bF$buf0),
    .D(_42_),
    .Q(Xin1[1])
);

DFFPOSX1 _592_ (
    .CLK(clk_bF$buf6),
    .D(_43_),
    .Q(Xin0[0])
);

DFFPOSX1 _593_ (
    .CLK(clk_bF$buf5),
    .D(_44_),
    .Q(Xin0[1])
);

DFFPOSX1 _594_ (
    .CLK(clk_bF$buf4),
    .D(_45_),
    .Q(Yin12b[10])
);

DFFPOSX1 _595_ (
    .CLK(clk_bF$buf3),
    .D(_46_),
    .Q(Yin12b[11])
);

DFFPOSX1 _596_ (
    .CLK(clk_bF$buf2),
    .D(_47_),
    .Q(Yin12b[8])
);

DFFPOSX1 _597_ (
    .CLK(clk_bF$buf1),
    .D(_48_),
    .Q(Yin12b[9])
);

DFFPOSX1 _598_ (
    .CLK(clk_bF$buf0),
    .D(_0_),
    .Q(Yin12b[6])
);

DFFPOSX1 _599_ (
    .CLK(clk_bF$buf6),
    .D(_1_),
    .Q(Yin12b[7])
);

DFFPOSX1 _600_ (
    .CLK(clk_bF$buf5),
    .D(_2_),
    .Q(Yin12b[4])
);

DFFPOSX1 _601_ (
    .CLK(clk_bF$buf4),
    .D(_3_),
    .Q(Yin12b[5])
);

DFFPOSX1 _602_ (
    .CLK(clk_bF$buf3),
    .D(_4_),
    .Q(Yin1[0])
);

DFFPOSX1 _603_ (
    .CLK(clk_bF$buf2),
    .D(_5_),
    .Q(Yin1[1])
);

DFFPOSX1 _604_ (
    .CLK(clk_bF$buf1),
    .D(_6_),
    .Q(Yin0[0])
);

DFFPOSX1 _605_ (
    .CLK(clk_bF$buf0),
    .D(_7_),
    .Q(Yin0[1])
);

DFFPOSX1 _606_ (
    .CLK(clk_bF$buf6),
    .D(Rdy),
    .Q(LoadCtl[0])
);

DFFPOSX1 _607_ (
    .CLK(clk_bF$buf5),
    .D(LoadCtl[0]),
    .Q(LoadCtl[1])
);

DFFPOSX1 _608_ (
    .CLK(clk_bF$buf4),
    .D(LoadCtl[1]),
    .Q(LoadCtl[2])
);

DFFPOSX1 _609_ (
    .CLK(clk_bF$buf3),
    .D(LoadCtl[2]),
    .Q(LoadCtl[3])
);

DFFPOSX1 _610_ (
    .CLK(clk_bF$buf2),
    .D(LoadCtl[3]),
    .Q(LoadCtl[4])
);

DFFPOSX1 _611_ (
    .CLK(clk_bF$buf1),
    .D(LoadCtl[4]),
    .Q(LoadCtl[5])
);

DFFPOSX1 _612_ (
    .CLK(clk_bF$buf0),
    .D(LoadCtl[5]),
    .Q(LoadCtl[6])
);

BUFX2 _613_ (
    .A(_272_[0]),
    .Y(Dout[0])
);

BUFX2 _614_ (
    .A(_272_[1]),
    .Y(Dout[1])
);

BUFX2 _615_ (
    .A(_272_[10]),
    .Y(Dout[10])
);

BUFX2 _616_ (
    .A(_272_[11]),
    .Y(Dout[11])
);

BUFX2 _617_ (
    .A(_272_[2]),
    .Y(Dout[2])
);

BUFX2 _618_ (
    .A(_272_[3]),
    .Y(Dout[3])
);

BUFX2 _619_ (
    .A(_272_[4]),
    .Y(Dout[4])
);

BUFX2 _620_ (
    .A(_272_[5]),
    .Y(Dout[5])
);

BUFX2 _621_ (
    .A(_272_[6]),
    .Y(Dout[6])
);

BUFX2 _622_ (
    .A(_272_[7]),
    .Y(Dout[7])
);

BUFX2 _623_ (
    .A(_272_[8]),
    .Y(Dout[8])
);

BUFX2 _624_ (
    .A(_272_[9]),
    .Y(Dout[9])
);

BUFX2 _625_ (
    .A(LoadCtl_6_bF$buf4),
    .Y(Vld)
);

endmodule
