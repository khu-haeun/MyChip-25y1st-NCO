magic
tech scmos
magscale 1 2
timestamp 1740654108
<< metal1 >>
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 1327 4677 1353 4683
rect 1307 4657 1473 4663
rect 5102 4578 5162 4818
rect 5070 4562 5162 4578
rect 2777 4477 2793 4483
rect 1287 4437 1453 4443
rect 2777 4403 2783 4477
rect 2777 4397 2793 4403
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 5102 4098 5162 4562
rect 5070 4082 5162 4098
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 5102 3618 5162 4082
rect 5070 3602 5162 3618
rect 4337 3537 4353 3543
rect 4337 3467 4343 3537
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 5102 3138 5162 3602
rect 5070 3122 5162 3138
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 567 2817 713 2823
rect 2727 2757 2893 2763
rect 5102 2658 5162 3122
rect 5070 2642 5162 2658
rect 3827 2577 3893 2583
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 5102 2178 5162 2642
rect 5070 2162 5162 2178
rect 4147 2097 4163 2103
rect 4157 2023 4163 2097
rect 4147 2017 4163 2023
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 5102 1698 5162 2162
rect 5070 1682 5162 1698
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 5102 1218 5162 1682
rect 5070 1202 5162 1218
rect -62 962 30 978
rect -62 498 -2 962
rect 1727 797 1753 803
rect 5102 738 5162 1202
rect 5070 722 5162 738
rect 4887 657 4913 663
rect -62 482 30 498
rect -62 18 -2 482
rect 4847 337 4893 343
rect 5102 258 5162 722
rect 5070 242 5162 258
rect -62 2 30 18
rect 5102 2 5162 242
<< m2contact >>
rect 1313 4673 1327 4687
rect 1353 4673 1367 4687
rect 1293 4653 1307 4667
rect 1473 4653 1487 4667
rect 1273 4433 1287 4447
rect 1453 4433 1467 4447
rect 2793 4473 2807 4487
rect 2793 4393 2807 4407
rect 4353 3533 4367 3547
rect 4333 3453 4347 3467
rect 553 2813 567 2827
rect 713 2813 727 2827
rect 2713 2753 2727 2767
rect 2893 2753 2907 2767
rect 3813 2573 3827 2587
rect 3893 2573 3907 2587
rect 4133 2093 4147 2107
rect 4133 2013 4147 2027
rect 1713 793 1727 807
rect 1753 793 1767 807
rect 4873 653 4887 667
rect 4913 653 4927 667
rect 4833 333 4847 347
rect 4893 333 4907 347
<< metal2 >>
rect 956 4696 983 4703
rect 216 4647 223 4663
rect 16 4007 23 4493
rect 36 3267 43 4533
rect 176 4447 183 4633
rect 256 4627 263 4663
rect 256 4443 263 4613
rect 436 4507 443 4673
rect 476 4547 483 4683
rect 756 4676 763 4693
rect 956 4667 963 4696
rect 996 4667 1003 4683
rect 1296 4676 1313 4683
rect 1476 4676 1503 4683
rect 536 4647 543 4663
rect 236 4436 263 4443
rect 216 4196 223 4333
rect 276 4167 283 4453
rect 436 4347 443 4493
rect 496 4483 503 4633
rect 696 4507 703 4533
rect 736 4496 743 4643
rect 1236 4627 1243 4663
rect 1276 4623 1283 4663
rect 1336 4663 1343 4673
rect 1316 4656 1343 4663
rect 1296 4647 1303 4653
rect 1316 4623 1323 4656
rect 1276 4616 1323 4623
rect 1356 4607 1363 4673
rect 1476 4667 1483 4676
rect 1436 4647 1443 4653
rect 476 4476 503 4483
rect 476 4223 483 4476
rect 476 4216 503 4223
rect 456 4167 463 4203
rect 496 4196 503 4216
rect 236 3736 243 3973
rect 296 3767 303 3993
rect 296 3703 303 3753
rect 336 3707 343 4013
rect 376 3996 383 4013
rect 476 3747 483 4183
rect 636 4027 643 4413
rect 696 4187 703 4493
rect 756 4476 763 4493
rect 796 4223 803 4483
rect 876 4476 903 4483
rect 896 4427 903 4476
rect 1296 4467 1303 4493
rect 1276 4447 1283 4463
rect 776 4216 803 4223
rect 756 4187 763 4203
rect 796 4167 803 4216
rect 976 4196 983 4273
rect 1256 4223 1263 4433
rect 1276 4287 1283 4433
rect 1236 4216 1263 4223
rect 636 3996 643 4013
rect 736 4003 743 4013
rect 716 3996 743 4003
rect 216 3687 223 3703
rect 276 3696 303 3703
rect 176 3516 203 3523
rect 176 3247 183 3516
rect 256 3516 263 3533
rect 436 3527 443 3733
rect 536 3707 543 3993
rect 956 3967 963 3983
rect 1016 3736 1023 3753
rect 1076 3743 1083 4013
rect 1236 3967 1243 3983
rect 1056 3736 1083 3743
rect 816 3716 843 3723
rect 516 3687 523 3703
rect 496 3547 503 3683
rect 236 3483 243 3513
rect 436 3496 443 3513
rect 456 3487 463 3533
rect 216 3476 243 3483
rect 496 3287 503 3483
rect 516 3267 523 3673
rect 836 3667 843 3716
rect 756 3516 763 3653
rect 227 3256 243 3263
rect 196 3047 203 3223
rect 216 3083 223 3253
rect 216 3076 243 3083
rect 236 3036 243 3076
rect 476 3067 483 3223
rect 516 3047 523 3213
rect 536 3207 543 3493
rect 736 3487 743 3503
rect 776 3496 783 3533
rect 256 2767 263 3033
rect 556 2827 563 3273
rect 716 3207 723 3253
rect 736 3227 743 3243
rect 716 3056 723 3193
rect 756 3087 763 3223
rect 796 3207 803 3223
rect 756 3036 783 3043
rect 16 2147 23 2333
rect 136 2107 143 2743
rect 216 2736 223 2753
rect 216 2556 223 2693
rect 256 2556 263 2753
rect 316 2707 323 2753
rect 176 2536 203 2543
rect 176 2227 183 2536
rect 236 2487 243 2543
rect 476 2507 483 2523
rect 556 2507 563 2813
rect 576 2487 583 2713
rect 696 2527 703 2793
rect 716 2556 723 2813
rect 776 2807 783 3036
rect 796 2783 803 3073
rect 836 3027 843 3053
rect 776 2776 803 2783
rect 856 2607 863 3713
rect 1036 3687 1043 3723
rect 1076 3523 1083 3736
rect 1256 3687 1263 4216
rect 1296 4207 1303 4453
rect 1396 4427 1403 4493
rect 1436 4447 1443 4633
rect 1456 4476 1483 4483
rect 1456 4447 1463 4476
rect 1536 4467 1543 4593
rect 1556 4487 1563 4663
rect 1576 4483 1583 4613
rect 1576 4476 1603 4483
rect 1676 4476 1683 4493
rect 1396 4003 1403 4413
rect 1416 4027 1423 4193
rect 1476 4187 1483 4203
rect 1556 4183 1563 4213
rect 1596 4187 1603 4453
rect 1736 4216 1743 4693
rect 1756 4647 1763 4673
rect 1776 4487 1783 4653
rect 1776 4227 1783 4473
rect 1816 4467 1823 4663
rect 1836 4607 1843 4683
rect 2056 4663 2063 4863
rect 2036 4647 2043 4663
rect 2056 4656 2083 4663
rect 2036 4507 2043 4633
rect 2356 4507 2363 4663
rect 2636 4663 2643 4693
rect 2616 4656 2643 4663
rect 2596 4503 2603 4643
rect 2636 4627 2643 4656
rect 2896 4663 2903 4793
rect 3936 4707 3943 4713
rect 3336 4696 3363 4703
rect 2876 4656 2903 4663
rect 3096 4676 3123 4683
rect 2596 4496 2623 4503
rect 1916 4476 1923 4493
rect 1996 4203 2003 4333
rect 1376 3996 1403 4003
rect 1296 3716 1323 3723
rect 1316 3687 1323 3716
rect 996 3516 1023 3523
rect 1056 3516 1083 3523
rect 996 3247 1003 3516
rect 1076 3387 1083 3516
rect 1296 3516 1303 3673
rect 1056 3207 1063 3223
rect 876 2787 883 3053
rect 1016 3036 1023 3053
rect 1036 3016 1043 3203
rect 976 2727 983 2743
rect 1016 2707 1023 2743
rect 1116 2647 1123 2743
rect 1016 2556 1023 2593
rect 196 2307 203 2313
rect 196 2276 203 2293
rect 576 2287 583 2473
rect 336 2276 363 2283
rect 356 2267 363 2276
rect 356 2107 363 2253
rect 96 2076 123 2083
rect 136 2076 143 2093
rect 116 1787 123 2076
rect 216 1967 223 2083
rect 276 2067 283 2083
rect 356 2076 363 2093
rect 276 1867 283 2053
rect 236 1796 243 1813
rect 296 1787 303 1953
rect 236 1756 263 1763
rect 236 1576 243 1756
rect 216 1547 223 1563
rect 196 1087 203 1303
rect 216 1116 223 1253
rect 276 1116 283 1293
rect 156 -24 163 1073
rect 296 983 303 1773
rect 316 1307 323 1853
rect 496 1827 503 2273
rect 556 2067 563 2263
rect 596 2067 603 2263
rect 616 2227 623 2283
rect 496 1796 503 1813
rect 616 1807 623 2213
rect 716 2103 723 2273
rect 736 2127 743 2263
rect 716 2096 743 2103
rect 736 2056 763 2063
rect 496 1616 503 1753
rect 436 1547 443 1593
rect 536 1567 543 1593
rect 736 1576 743 2056
rect 756 1767 763 1783
rect 796 1767 803 1783
rect 776 1747 783 1763
rect 776 1563 783 1573
rect 436 1247 443 1533
rect 716 1387 723 1563
rect 756 1556 783 1563
rect 816 1387 823 2553
rect 1036 2347 1043 2543
rect 856 2256 883 2263
rect 876 2247 883 2256
rect 956 1847 963 2253
rect 976 2227 983 2333
rect 976 2076 983 2213
rect 1016 2076 1023 2133
rect 896 1747 903 1783
rect 956 1783 963 1833
rect 936 1776 963 1783
rect 456 1267 463 1303
rect 496 1287 503 1303
rect 656 1287 663 1313
rect 676 1307 683 1373
rect 776 1323 783 1373
rect 756 1316 783 1323
rect 456 1107 463 1253
rect 476 1147 483 1283
rect 696 1267 703 1303
rect 496 1116 503 1233
rect 796 1167 803 1353
rect 536 1147 543 1153
rect 576 1103 583 1133
rect 756 1116 763 1153
rect 816 1116 823 1153
rect 556 1096 583 1103
rect 276 976 303 983
rect 196 816 223 823
rect 196 667 203 816
rect 236 787 243 803
rect 196 636 203 653
rect 276 643 283 976
rect 456 807 463 1093
rect 736 836 763 843
rect 456 656 463 793
rect 256 636 283 643
rect 216 383 223 603
rect 196 376 223 383
rect 196 343 203 376
rect 276 343 283 636
rect 436 607 443 623
rect 476 356 483 593
rect 196 336 223 343
rect 256 336 283 343
rect 196 -24 203 336
rect 676 327 683 813
rect 756 623 763 836
rect 796 787 803 1073
rect 836 827 843 873
rect 736 616 763 623
rect 696 356 703 373
rect 276 123 283 293
rect 536 156 543 193
rect 216 107 223 123
rect 256 116 283 123
rect 216 -17 223 93
rect 216 -24 243 -17
rect 496 -24 503 113
rect 736 107 743 343
rect 756 307 763 323
rect 916 307 923 1773
rect 936 1347 943 1593
rect 1096 1567 1103 2533
rect 1156 2267 1163 2743
rect 1256 2703 1263 3223
rect 1296 3207 1303 3223
rect 1316 3027 1323 3673
rect 1236 2696 1263 2703
rect 1216 2267 1223 2273
rect 1216 2067 1223 2253
rect 1236 2147 1243 2696
rect 1256 2556 1263 2593
rect 1276 2576 1283 2633
rect 1316 2327 1323 3013
rect 1356 2587 1363 3953
rect 1396 3887 1403 3996
rect 1436 3716 1443 3873
rect 1456 3667 1463 4003
rect 1476 3647 1483 4173
rect 1496 3987 1503 4183
rect 1536 4176 1563 4183
rect 1756 4047 1763 4203
rect 1976 4196 2003 4203
rect 1716 3976 1743 3983
rect 1527 3516 1543 3523
rect 1556 3516 1563 3713
rect 1656 3667 1663 3703
rect 1716 3647 1723 3723
rect 1736 3707 1743 3976
rect 1756 3967 1763 3983
rect 1996 3976 2003 4196
rect 2056 4163 2063 4193
rect 2036 4156 2063 4163
rect 2256 4047 2263 4203
rect 2276 4047 2283 4183
rect 2036 3976 2043 4033
rect 2236 3996 2243 4013
rect 2316 3983 2323 4033
rect 1936 3716 1963 3723
rect 2096 3716 2103 3793
rect 1936 3687 1943 3716
rect 1536 3487 1543 3516
rect 1716 3507 1723 3633
rect 1856 3527 1863 3653
rect 1716 3267 1723 3493
rect 1776 3263 1783 3513
rect 1836 3387 1843 3503
rect 1776 3256 1803 3263
rect 1456 3047 1463 3223
rect 1536 3216 1563 3223
rect 1556 3187 1563 3216
rect 1636 3056 1643 3173
rect 1456 3027 1463 3033
rect 1676 3023 1683 3233
rect 1716 3207 1723 3253
rect 1796 3236 1803 3256
rect 1656 3016 1683 3023
rect 1476 2756 1483 2773
rect 1536 2536 1543 2613
rect 1316 2276 1323 2293
rect 1516 2267 1523 2523
rect 1576 2287 1583 2333
rect 1676 2307 1683 2773
rect 1696 2756 1723 2763
rect 1696 2567 1703 2756
rect 1736 2647 1743 2723
rect 1736 2556 1743 2573
rect 1696 2547 1703 2553
rect 1796 2536 1803 2613
rect 1696 2527 1703 2533
rect 1587 2276 1603 2283
rect 1676 2263 1683 2293
rect 1656 2256 1683 2263
rect 1236 2076 1243 2113
rect 1256 2047 1263 2063
rect 1216 1647 1223 1813
rect 1256 1796 1263 1813
rect 1316 1803 1323 2213
rect 1336 2047 1343 2073
rect 1356 2067 1363 2093
rect 1516 2056 1523 2213
rect 1576 2076 1603 2083
rect 1596 2027 1603 2076
rect 1296 1796 1323 1803
rect 1436 1783 1443 1833
rect 1656 1787 1663 2093
rect 1736 2063 1743 2273
rect 1836 2263 1843 2633
rect 1856 2547 1863 3233
rect 1916 3207 1923 3373
rect 1876 3036 1903 3043
rect 1916 3036 1923 3193
rect 1896 2307 1903 3036
rect 1956 2787 1963 3273
rect 2076 3256 2083 3273
rect 2056 3063 2063 3243
rect 2036 3056 2063 3063
rect 2116 3223 2123 3473
rect 2256 3287 2263 3983
rect 2296 3976 2323 3983
rect 2296 3736 2323 3743
rect 2356 3736 2383 3743
rect 2296 3527 2303 3736
rect 2376 3667 2383 3736
rect 2316 3547 2323 3633
rect 2376 3527 2383 3653
rect 2476 3547 2483 4493
rect 2596 4443 2603 4473
rect 2616 4467 2623 4496
rect 2796 4487 2803 4653
rect 2856 4476 2863 4493
rect 2776 4456 2803 4463
rect 2536 4347 2543 4443
rect 2576 4436 2603 4443
rect 2516 4176 2543 4183
rect 2516 4027 2523 4176
rect 2596 4183 2603 4353
rect 2776 4207 2783 4456
rect 2796 4227 2803 4393
rect 2956 4207 2963 4513
rect 3076 4367 3083 4463
rect 3096 4447 3103 4676
rect 3136 4663 3143 4693
rect 3136 4656 3163 4663
rect 3336 4647 3343 4696
rect 4156 4696 4163 4733
rect 3136 4507 3143 4533
rect 2856 4196 2883 4203
rect 2587 4176 2603 4183
rect 2776 4183 2783 4193
rect 2776 4176 2803 4183
rect 2876 4167 2883 4196
rect 2516 3976 2523 4013
rect 2556 4007 2563 4163
rect 2836 4147 2843 4163
rect 2776 3963 2783 4133
rect 2816 3996 2843 4003
rect 2496 3727 2503 3963
rect 2496 3507 2503 3553
rect 2516 3223 2523 3913
rect 2536 3567 2543 3963
rect 2776 3956 2803 3963
rect 2556 3647 2563 3703
rect 2596 3647 2603 3703
rect 2756 3687 2763 3733
rect 2616 3507 2623 3633
rect 2116 3216 2143 3223
rect 2036 3036 2043 3056
rect 1976 2347 1983 2763
rect 2096 2743 2103 3033
rect 2116 2923 2123 3216
rect 2216 3087 2223 3223
rect 2256 3207 2263 3223
rect 2516 3216 2543 3223
rect 2176 3043 2183 3053
rect 2216 3047 2223 3073
rect 2156 3036 2183 3043
rect 2116 2916 2143 2923
rect 2016 2736 2043 2743
rect 2096 2736 2113 2743
rect 2016 2647 2023 2736
rect 2136 2723 2143 2916
rect 2116 2716 2143 2723
rect 2116 2707 2123 2716
rect 2036 2576 2043 2633
rect 1996 2527 2003 2553
rect 1836 2256 1863 2263
rect 1736 2056 1783 2063
rect 1236 1596 1243 1733
rect 1276 1663 1283 1783
rect 1416 1747 1423 1783
rect 1436 1776 1463 1783
rect 1716 1767 1723 2053
rect 1756 1796 1763 2056
rect 1816 1747 1823 1783
rect 1256 1656 1283 1663
rect 1256 1627 1263 1656
rect 1276 1616 1283 1633
rect 1536 1596 1543 1713
rect 956 1367 963 1563
rect 976 1336 983 1353
rect 936 1087 943 1333
rect 996 1307 1003 1323
rect 956 847 963 1273
rect 1056 1116 1063 1193
rect 1096 1147 1103 1553
rect 1296 1307 1303 1583
rect 1276 1287 1283 1303
rect 1256 1107 1263 1283
rect 1336 1167 1343 1333
rect 1456 1327 1463 1593
rect 1516 1387 1523 1583
rect 1556 1576 1583 1583
rect 1476 1336 1483 1353
rect 1336 1136 1343 1153
rect 1076 827 1083 1103
rect 1296 1103 1303 1133
rect 1376 1116 1383 1133
rect 1296 1096 1323 1103
rect 1356 887 1363 1103
rect 936 647 943 823
rect 1316 807 1323 853
rect 1356 807 1363 873
rect 1496 836 1503 853
rect 1536 847 1543 1353
rect 1536 807 1543 833
rect 1576 827 1583 1576
rect 1716 1336 1743 1343
rect 1616 1116 1643 1123
rect 1636 827 1643 1116
rect 1676 1103 1683 1333
rect 1656 1096 1683 1103
rect 956 383 963 793
rect 1196 656 1223 663
rect 996 616 1003 633
rect 1196 607 1203 656
rect 976 407 983 593
rect 1016 507 1023 603
rect 956 376 983 383
rect 996 287 1003 363
rect 776 176 783 273
rect 796 156 803 173
rect 976 156 983 193
rect 1016 183 1023 353
rect 1036 347 1043 363
rect 1056 347 1063 493
rect 1316 347 1323 793
rect 1456 643 1463 653
rect 1436 636 1463 643
rect 1496 636 1503 673
rect 1636 647 1643 813
rect 1436 627 1443 636
rect 1516 616 1543 623
rect 1536 507 1543 616
rect 1496 376 1523 383
rect 1007 176 1023 183
rect 816 127 823 153
rect 1036 147 1043 333
rect 1236 307 1243 333
rect 1236 187 1243 193
rect 1316 143 1323 313
rect 1336 187 1343 373
rect 1336 163 1343 173
rect 1336 156 1363 163
rect 1436 156 1443 173
rect 1476 156 1483 213
rect 1496 167 1503 376
rect 1696 187 1703 853
rect 1716 807 1723 1336
rect 1756 1307 1763 1323
rect 1796 1187 1803 1583
rect 1736 627 1743 1133
rect 1796 867 1803 1173
rect 1896 1147 1903 2073
rect 1956 1587 1963 2313
rect 1996 2127 2003 2293
rect 2036 2287 2043 2533
rect 2056 2187 2063 2543
rect 1996 2087 2003 2113
rect 2076 2067 2083 2073
rect 2076 1847 2083 2053
rect 1936 1576 1953 1583
rect 1896 1116 1903 1133
rect 2016 1127 2023 1303
rect 2036 1267 2043 1803
rect 2076 1796 2083 1833
rect 2096 1707 2103 1783
rect 2056 1287 2063 1303
rect 2116 1287 2123 2693
rect 2156 2667 2163 2743
rect 2136 2267 2143 2283
rect 2176 2276 2183 2753
rect 2296 2576 2303 2653
rect 2316 2607 2323 3153
rect 2456 2787 2463 3033
rect 2516 3027 2523 3216
rect 2576 3167 2583 3223
rect 2536 3036 2543 3073
rect 2576 3036 2583 3073
rect 2707 2756 2713 2763
rect 2336 2727 2343 2743
rect 2456 2736 2483 2743
rect 2476 2727 2483 2736
rect 2316 2556 2323 2593
rect 2336 2507 2343 2553
rect 2336 2267 2343 2493
rect 2156 2047 2163 2263
rect 2216 2256 2243 2263
rect 2296 2256 2323 2263
rect 2196 2067 2203 2253
rect 2216 2187 2223 2256
rect 2256 2096 2263 2173
rect 2296 1587 2303 2256
rect 2416 2147 2423 2553
rect 2676 2296 2683 2553
rect 2776 2503 2783 3933
rect 2836 3787 2843 3996
rect 2856 3947 2863 4153
rect 3096 4147 3103 4163
rect 3096 3983 3103 4133
rect 3116 4127 3123 4183
rect 3076 3976 3103 3983
rect 2836 3716 2863 3723
rect 2796 3683 2803 3713
rect 2796 3676 2823 3683
rect 2856 3647 2863 3716
rect 2816 3487 2823 3513
rect 2816 3027 2823 3243
rect 2856 3236 2863 3273
rect 2876 3263 2883 3693
rect 2896 3516 2903 3733
rect 3036 3727 3043 3953
rect 3056 3767 3063 3963
rect 2876 3256 2903 3263
rect 2816 2567 2823 3013
rect 2836 2767 2843 3223
rect 2896 3036 2903 3256
rect 2916 3227 2923 3673
rect 3056 3467 3063 3733
rect 3156 3723 3163 4193
rect 3176 3987 3183 4493
rect 3376 4476 3383 4533
rect 3296 3983 3303 4193
rect 3356 4187 3363 4453
rect 3367 4176 3383 4183
rect 3376 4147 3383 4176
rect 3416 4163 3423 4193
rect 3396 4156 3423 4163
rect 3336 4016 3343 4033
rect 3556 4007 3563 4633
rect 3576 4443 3583 4673
rect 3936 4663 3943 4693
rect 3636 4527 3643 4663
rect 3676 4567 3683 4663
rect 3876 4647 3883 4663
rect 3916 4656 3943 4663
rect 3836 4476 3863 4483
rect 3576 4436 3603 4443
rect 3516 3996 3543 4003
rect 3296 3976 3323 3983
rect 3176 3747 3183 3973
rect 3356 3967 3363 3983
rect 3136 3716 3163 3723
rect 3136 3467 3143 3483
rect 3116 3056 3123 3073
rect 3096 3036 3103 3053
rect 3136 3036 3143 3053
rect 2907 2756 2923 2763
rect 3156 2567 3163 3233
rect 3176 2763 3183 3513
rect 3256 3267 3263 3493
rect 3276 3063 3283 3753
rect 3296 3507 3303 3713
rect 3316 3703 3323 3953
rect 3516 3807 3523 3996
rect 3316 3696 3363 3703
rect 3396 3687 3403 3703
rect 3416 3527 3423 3733
rect 3536 3527 3543 3793
rect 3556 3687 3563 3993
rect 3576 3883 3583 4213
rect 3636 4196 3643 4213
rect 3676 4207 3683 4473
rect 3836 4227 3843 4476
rect 3916 4467 3923 4553
rect 4076 4507 4083 4693
rect 3876 4443 3883 4463
rect 3876 4436 3903 4443
rect 3616 4047 3623 4183
rect 3656 4147 3663 4163
rect 3836 4127 3843 4213
rect 3896 4196 3903 4436
rect 3836 3996 3843 4113
rect 3916 4007 3923 4153
rect 3996 3996 4003 4033
rect 4016 3996 4043 4003
rect 3576 3876 3603 3883
rect 3596 3743 3603 3876
rect 3596 3736 3623 3743
rect 3576 3516 3583 3533
rect 3336 3243 3343 3513
rect 3396 3487 3403 3503
rect 3396 3287 3403 3473
rect 3336 3236 3363 3243
rect 3396 3203 3403 3273
rect 3496 3223 3503 3513
rect 3596 3487 3603 3736
rect 3636 3687 3643 3723
rect 3776 3487 3783 3493
rect 3416 3216 3443 3223
rect 3496 3216 3523 3223
rect 3416 3207 3423 3216
rect 3336 3187 3343 3203
rect 3376 3196 3403 3203
rect 3276 3056 3303 3063
rect 3176 2756 3203 2763
rect 2836 2507 2843 2523
rect 2776 2496 2803 2503
rect 2716 2247 2723 2263
rect 2376 1796 2383 1813
rect 2316 1627 2323 1783
rect 2396 1767 2403 1833
rect 2336 1567 2343 1753
rect 2416 1307 2423 2133
rect 2496 2076 2503 2233
rect 2516 2047 2523 2063
rect 2536 1807 2543 2033
rect 2576 1816 2583 2233
rect 2796 2076 2803 2496
rect 2976 2276 2983 2553
rect 3216 2547 3223 2743
rect 3096 2507 3103 2543
rect 2996 2247 3003 2263
rect 2996 2043 3003 2233
rect 3036 2056 3043 2273
rect 3196 2247 3203 2263
rect 3196 2087 3203 2233
rect 2996 2036 3023 2043
rect 2436 1596 2443 1613
rect 2476 1603 2483 1613
rect 2576 1603 2583 1633
rect 2456 1596 2483 1603
rect 2556 1596 2583 1603
rect 2456 1587 2463 1596
rect 2296 1267 2303 1303
rect 2156 1116 2163 1133
rect 1916 823 1923 853
rect 1756 636 1763 793
rect 1796 667 1803 823
rect 1896 767 1903 823
rect 1916 816 1943 823
rect 2176 807 2183 1113
rect 2276 807 2283 823
rect 1996 656 2003 673
rect 1776 356 1783 593
rect 1756 307 1763 323
rect 1816 227 1823 633
rect 1936 307 1943 373
rect 1976 367 1983 653
rect 2016 636 2023 653
rect 2056 607 2063 623
rect 2036 376 2063 383
rect 2056 327 2063 376
rect 2176 367 2183 793
rect 2256 687 2263 803
rect 2236 623 2243 673
rect 2316 636 2323 653
rect 2336 627 2343 1113
rect 2436 1103 2443 1153
rect 2456 1116 2463 1553
rect 2496 1116 2503 1333
rect 2556 1167 2563 1303
rect 2416 1096 2443 1103
rect 2416 847 2423 1096
rect 2516 887 2523 1113
rect 2536 1107 2543 1133
rect 2416 747 2423 833
rect 2476 823 2483 873
rect 2536 836 2543 1093
rect 2696 827 2703 1553
rect 2736 1136 2743 1593
rect 2796 1576 2803 2033
rect 2996 1847 3003 2036
rect 2856 1796 2863 1813
rect 2916 1776 2923 1833
rect 2876 1647 2883 1763
rect 2996 1627 3003 1783
rect 3056 1747 3063 2043
rect 3196 1767 3203 2073
rect 2976 1596 2983 1613
rect 3056 1567 3063 1603
rect 2776 1547 2783 1563
rect 3196 1327 3203 1733
rect 3256 1687 3263 2283
rect 3276 2127 3283 3033
rect 3296 2747 3303 3056
rect 3376 3036 3383 3196
rect 3396 3007 3403 3196
rect 3396 2727 3403 2993
rect 3336 2576 3343 2653
rect 3376 2556 3403 2563
rect 3296 2536 3323 2543
rect 3276 2076 3283 2113
rect 3296 1727 3303 2536
rect 3316 2076 3323 2493
rect 3396 2287 3403 2556
rect 3416 2507 3423 3173
rect 3496 2667 3503 2723
rect 3516 2607 3523 2743
rect 3536 2263 3543 3453
rect 3636 3036 3643 3053
rect 3676 3047 3683 3213
rect 3776 3027 3783 3473
rect 3656 3007 3663 3023
rect 3796 2987 3803 3993
rect 3816 3167 3823 3713
rect 3836 3236 3843 3773
rect 3936 3716 3963 3723
rect 3956 3707 3963 3716
rect 3876 3547 3883 3703
rect 3936 3283 3943 3673
rect 4016 3527 4023 3996
rect 4076 3747 4083 4493
rect 4136 4483 4143 4683
rect 4116 4476 4143 4483
rect 4096 4227 4103 4473
rect 4116 4467 4123 4476
rect 4156 4456 4163 4473
rect 4116 4443 4123 4453
rect 4196 4443 4203 4453
rect 4116 4436 4143 4443
rect 4176 4436 4203 4443
rect 4096 4167 4103 4183
rect 4136 3823 4143 4013
rect 4116 3816 4143 3823
rect 4116 3703 4123 3816
rect 4156 3716 4163 4183
rect 4116 3696 4143 3703
rect 3956 3487 3963 3523
rect 4076 3516 4103 3523
rect 3936 3276 3963 3283
rect 3876 3236 3883 3253
rect 3556 2547 3563 2753
rect 3636 2556 3643 2973
rect 3756 2756 3763 2773
rect 3696 2607 3703 2723
rect 3676 2556 3683 2593
rect 3816 2587 3823 3153
rect 3516 2256 3543 2263
rect 3556 2076 3563 2533
rect 3656 2403 3663 2533
rect 3636 2396 3663 2403
rect 3396 1767 3403 1783
rect 3436 1776 3443 2013
rect 3576 2007 3583 2043
rect 3296 1576 3303 1673
rect 3396 1567 3403 1753
rect 3516 1747 3523 1783
rect 3516 1627 3523 1733
rect 3536 1583 3543 1813
rect 3556 1767 3563 1783
rect 3616 1603 3623 2013
rect 3596 1596 3623 1603
rect 3516 1576 3543 1583
rect 2776 1287 2783 1303
rect 2756 1116 2763 1153
rect 2816 863 2823 1303
rect 2956 1087 2963 1103
rect 3056 1003 3063 1303
rect 3076 1167 3083 1283
rect 3176 1116 3183 1173
rect 3196 1087 3203 1313
rect 3276 1307 3283 1553
rect 3316 1547 3323 1553
rect 3516 1327 3523 1576
rect 3576 1563 3583 1583
rect 3576 1556 3603 1563
rect 3596 1327 3603 1556
rect 3056 996 3083 1003
rect 2836 863 2843 873
rect 2816 856 2843 863
rect 2476 816 2523 823
rect 2556 787 2563 823
rect 2236 616 2263 623
rect 2296 347 2303 363
rect 2236 207 2243 343
rect 1696 156 1703 173
rect 1796 163 1803 193
rect 2276 183 2283 343
rect 2256 176 2283 183
rect 1776 156 1803 163
rect 1296 136 1323 143
rect 2096 127 2103 173
rect 2116 147 2123 173
rect 2256 167 2263 176
rect 2316 156 2323 173
rect 2336 167 2343 613
rect 2416 347 2423 733
rect 2756 667 2763 823
rect 2836 807 2843 856
rect 2996 856 3023 863
rect 2996 787 3003 856
rect 2816 636 2823 673
rect 2836 656 2843 753
rect 2536 607 2543 623
rect 2536 367 2543 573
rect 2616 367 2623 613
rect 2576 356 2603 363
rect 2416 167 2423 333
rect 2516 307 2523 343
rect 2536 156 2543 193
rect 2576 156 2583 333
rect 2596 167 2603 356
rect 2796 347 2803 633
rect 2876 383 2883 773
rect 3076 587 3083 996
rect 3096 616 3103 733
rect 3116 636 3123 813
rect 3216 727 3223 1173
rect 3296 1123 3303 1283
rect 3516 1267 3523 1313
rect 3576 1287 3583 1303
rect 3256 1116 3303 1123
rect 3276 836 3283 853
rect 3316 743 3323 823
rect 3356 803 3363 1193
rect 3436 1116 3463 1123
rect 3436 827 3443 1116
rect 3516 1107 3523 1253
rect 3636 1207 3643 2396
rect 3716 2263 3723 2573
rect 3656 1747 3663 2263
rect 3696 2256 3723 2263
rect 3856 2056 3863 3203
rect 3896 3087 3903 3223
rect 3936 3187 3943 3253
rect 3956 3227 3963 3276
rect 4016 3223 4023 3513
rect 4096 3227 4103 3516
rect 4016 3216 4043 3223
rect 4076 3187 4083 3223
rect 3916 3036 3923 3053
rect 3976 2763 3983 3073
rect 4016 3027 4023 3073
rect 4136 3027 4143 3053
rect 4156 3036 4163 3173
rect 4196 3087 4203 3713
rect 4296 3467 4303 4813
rect 4316 4667 4323 4863
rect 4356 4827 4363 4863
rect 4396 4807 4403 4863
rect 4636 4856 4663 4863
rect 4896 4856 4923 4863
rect 4656 4707 4663 4856
rect 4676 4747 4683 4753
rect 4596 4696 4623 4703
rect 4436 4647 4443 4663
rect 4596 4647 4603 4696
rect 4396 4447 4403 4633
rect 4436 4456 4443 4473
rect 4416 4427 4423 4443
rect 4336 4187 4343 4413
rect 4336 3927 4343 4173
rect 4356 4163 4363 4193
rect 4356 4156 4383 4163
rect 4376 3976 4383 4156
rect 4416 4047 4423 4183
rect 4456 4007 4463 4433
rect 4476 4207 4483 4473
rect 4636 4447 4643 4683
rect 4676 4476 4683 4733
rect 4856 4667 4863 4693
rect 4867 4636 4883 4643
rect 4596 3963 4603 4193
rect 4596 3956 4623 3963
rect 4396 3736 4423 3743
rect 4316 3287 4323 3493
rect 4336 3487 4343 3733
rect 4396 3687 4403 3736
rect 4476 3727 4483 3953
rect 4676 3747 4683 4153
rect 4696 3716 4703 3953
rect 4736 3547 4743 4453
rect 4856 4167 4863 4633
rect 4916 4423 4923 4856
rect 4996 4443 5003 4673
rect 4976 4436 5003 4443
rect 4916 4416 4943 4423
rect 4876 4196 4903 4203
rect 4796 3547 4803 4013
rect 4816 3996 4843 4003
rect 4876 3996 4883 4196
rect 4936 4163 4943 4416
rect 4916 4156 4943 4163
rect 4816 3967 4823 3996
rect 4916 3743 4923 4156
rect 4896 3736 4923 3743
rect 4896 3707 4903 3736
rect 4916 3687 4923 3703
rect 4367 3536 4383 3543
rect 4376 3496 4383 3536
rect 4416 3487 4423 3533
rect 4336 3247 4343 3453
rect 4396 3427 4403 3483
rect 4376 3236 4383 3273
rect 4196 3056 4203 3073
rect 4256 2776 4263 3053
rect 3976 2756 4003 2763
rect 4036 2756 4043 2773
rect 3896 2556 3903 2573
rect 3936 2556 3963 2563
rect 3936 2287 3943 2513
rect 3956 2507 3963 2556
rect 3916 2047 3923 2073
rect 3876 2007 3883 2043
rect 3716 1707 3723 1773
rect 3756 1747 3763 1783
rect 3656 1347 3663 1633
rect 3656 1296 3663 1333
rect 3696 1327 3703 1613
rect 3716 1327 3723 1693
rect 3796 1667 3803 1783
rect 3816 1596 3823 1753
rect 3876 1727 3883 1993
rect 3896 1583 3903 1673
rect 3876 1576 3903 1583
rect 3476 1087 3483 1103
rect 3536 843 3543 1093
rect 3696 887 3703 1313
rect 3736 1187 3743 1303
rect 3776 1267 3783 1303
rect 3796 1116 3803 1333
rect 3776 887 3783 1103
rect 3916 1067 3923 2033
rect 3956 1807 3963 2493
rect 3536 836 3563 843
rect 3596 836 3603 873
rect 3776 827 3783 873
rect 3576 807 3583 823
rect 3336 796 3363 803
rect 3316 736 3343 743
rect 3276 636 3283 713
rect 3316 636 3323 653
rect 3136 587 3143 623
rect 2856 376 2883 383
rect 2876 327 2883 376
rect 2936 347 2943 373
rect 3116 356 3123 373
rect 2836 156 2843 213
rect 2336 147 2343 153
rect 2596 136 2603 153
rect 2996 -24 3003 333
rect 3196 327 3203 633
rect 3336 347 3343 736
rect 3356 723 3363 796
rect 3356 716 3383 723
rect 3376 607 3383 716
rect 3616 616 3623 773
rect 3376 347 3383 363
rect 3596 347 3603 603
rect 3656 387 3663 593
rect 3676 587 3683 813
rect 3796 807 3803 833
rect 3796 636 3803 713
rect 3816 647 3823 823
rect 3876 587 3883 643
rect 3976 607 3983 2593
rect 4056 2547 4063 2743
rect 4016 1827 4023 2263
rect 4056 2247 4063 2263
rect 4076 2043 4083 2733
rect 4356 2547 4363 3223
rect 4416 2903 4423 3003
rect 4396 2896 4423 2903
rect 4396 2767 4403 2896
rect 4416 2767 4423 2773
rect 4416 2556 4423 2753
rect 4476 2727 4483 3053
rect 4536 2756 4543 3033
rect 4576 2743 4583 3233
rect 4636 3207 4643 3503
rect 4696 3236 4703 3253
rect 4736 3036 4743 3213
rect 4756 3207 4763 3413
rect 4876 3267 4883 3503
rect 4856 3087 4863 3233
rect 4896 3227 4903 3273
rect 4756 3007 4763 3053
rect 4756 2756 4783 2763
rect 4556 2736 4583 2743
rect 4476 2563 4483 2573
rect 4456 2556 4483 2563
rect 4396 2536 4403 2553
rect 4436 2527 4443 2543
rect 4276 2247 4283 2263
rect 4116 2096 4133 2103
rect 4116 2056 4123 2096
rect 4076 2036 4093 2043
rect 4156 2043 4163 2093
rect 4276 2067 4283 2233
rect 4296 2107 4303 2243
rect 4356 2107 4363 2293
rect 4476 2287 4483 2556
rect 4696 2543 4703 2713
rect 4736 2547 4743 2753
rect 4756 2747 4763 2756
rect 4856 2743 4863 3073
rect 4896 3027 4903 3213
rect 4916 3063 4923 3533
rect 4936 3287 4943 3683
rect 4976 3667 4983 3713
rect 4976 3207 4983 3223
rect 4916 3056 4943 3063
rect 4916 3047 4923 3056
rect 4936 3036 4943 3056
rect 4976 3036 4983 3053
rect 4996 3016 5003 3073
rect 4836 2736 4863 2743
rect 4856 2576 4883 2583
rect 4856 2567 4863 2576
rect 4676 2536 4703 2543
rect 4516 2296 4523 2313
rect 4736 2283 4743 2313
rect 4736 2276 4763 2283
rect 4636 2096 4643 2253
rect 4396 2076 4423 2083
rect 4336 2047 4343 2063
rect 4136 2036 4163 2043
rect 4136 1823 4143 2013
rect 4116 1816 4143 1823
rect 4096 1687 4103 1803
rect 4416 1803 4423 2076
rect 4596 2076 4623 2083
rect 4596 2027 4603 2076
rect 4416 1796 4443 1803
rect 4096 1596 4103 1653
rect 4076 1316 4103 1323
rect 4016 1116 4023 1253
rect 4096 1167 4103 1316
rect 4116 1307 4123 1583
rect 4076 856 4083 1053
rect 4096 827 4103 843
rect 3656 356 3663 373
rect 3076 123 3083 213
rect 3216 167 3223 313
rect 3396 163 3403 193
rect 3616 183 3623 353
rect 3636 227 3643 343
rect 4036 327 4043 633
rect 3596 176 3623 183
rect 3396 156 3423 163
rect 3216 127 3223 153
rect 3416 127 3423 156
rect 3576 147 3583 173
rect 3596 156 3603 176
rect 3636 156 3643 173
rect 3816 167 3823 193
rect 4056 187 4063 773
rect 4116 687 4123 863
rect 4136 787 4143 843
rect 4156 827 4163 1273
rect 4256 1087 4263 1793
rect 4356 1627 4363 1783
rect 4396 1747 4403 1763
rect 4416 1596 4423 1733
rect 4436 1616 4443 1796
rect 4616 1743 4623 1783
rect 4616 1736 4643 1743
rect 4336 1303 4343 1333
rect 4316 1296 4343 1303
rect 4536 1303 4543 1713
rect 4636 1647 4643 1736
rect 4636 1596 4643 1633
rect 4576 1347 4583 1593
rect 4576 1316 4583 1333
rect 4616 1316 4623 1353
rect 4656 1307 4663 1753
rect 4736 1747 4743 2276
rect 4856 2267 4863 2553
rect 4836 2076 4863 2083
rect 4836 2027 4843 2076
rect 4876 2043 4883 2273
rect 4916 2076 4923 2233
rect 4856 2036 4883 2043
rect 4856 1783 4863 2036
rect 5016 1787 5023 4793
rect 5096 4627 5103 4673
rect 5036 2276 5063 2283
rect 4856 1776 4883 1783
rect 4916 1776 4943 1783
rect 4756 1567 4763 1773
rect 4836 1327 4843 1593
rect 4856 1336 4863 1553
rect 4876 1347 4883 1776
rect 4896 1747 4903 1763
rect 4936 1616 4943 1776
rect 4956 1596 4983 1603
rect 4976 1567 4983 1596
rect 5036 1367 5043 2276
rect 5076 1767 5083 2243
rect 4536 1296 4563 1303
rect 4836 1303 4843 1313
rect 4816 1296 4843 1303
rect 4336 1136 4343 1153
rect 4536 1136 4563 1143
rect 4296 1116 4303 1133
rect 4536 1107 4543 1136
rect 4576 1116 4583 1153
rect 4316 1087 4323 1103
rect 4336 856 4343 873
rect 4076 636 4103 643
rect 4076 347 4083 636
rect 4356 616 4363 673
rect 4376 596 4383 813
rect 4396 616 4403 653
rect 4436 627 4443 853
rect 4536 847 4543 1093
rect 4616 1087 4623 1103
rect 4636 863 4643 873
rect 4636 856 4663 863
rect 4656 823 4663 856
rect 4636 816 4663 823
rect 4396 356 4403 373
rect 4636 367 4643 816
rect 4676 383 4683 653
rect 4696 636 4703 673
rect 4736 383 4743 673
rect 4816 647 4823 1273
rect 4836 1116 4863 1123
rect 4896 1116 4903 1273
rect 4856 863 4863 1116
rect 4876 883 4883 1083
rect 4876 876 4903 883
rect 4836 856 4863 863
rect 4896 863 4903 876
rect 4896 856 4923 863
rect 4836 587 4843 856
rect 4916 667 4923 856
rect 4936 656 4943 673
rect 4656 376 4683 383
rect 4716 376 4743 383
rect 4656 347 4663 376
rect 4836 347 4843 573
rect 4876 347 4883 653
rect 4956 636 4983 643
rect 4907 336 4923 343
rect 3076 116 3103 123
rect 3816 27 3823 153
rect 4156 136 4163 313
rect 4176 187 4183 323
rect 4396 176 4403 193
rect 3896 27 3903 123
rect 4116 123 4123 133
rect 4196 123 4203 133
rect 4256 127 4263 173
rect 4416 127 4423 143
rect 4896 127 4903 143
rect 4116 116 4143 123
rect 4176 116 4203 123
rect 4956 27 4963 333
rect 4976 327 4983 636
rect 3816 -24 3823 13
rect 4876 -24 4883 13
<< m3contact >>
rect 753 4693 767 4707
rect 433 4673 447 4687
rect 173 4633 187 4647
rect 213 4633 227 4647
rect 233 4633 247 4647
rect 33 4533 47 4547
rect 13 4493 27 4507
rect 13 3993 27 4007
rect 253 4613 267 4627
rect 213 4453 227 4467
rect 173 4433 187 4447
rect 193 4433 207 4447
rect 513 4673 527 4687
rect 1013 4693 1027 4707
rect 1733 4693 1747 4707
rect 1253 4673 1267 4687
rect 1333 4673 1347 4687
rect 493 4653 507 4667
rect 953 4653 967 4667
rect 993 4653 1007 4667
rect 493 4633 507 4647
rect 533 4633 547 4647
rect 473 4533 487 4547
rect 433 4493 447 4507
rect 273 4453 287 4467
rect 213 4333 227 4347
rect 693 4533 707 4547
rect 513 4493 527 4507
rect 693 4493 707 4507
rect 1233 4613 1247 4627
rect 1293 4633 1307 4647
rect 1533 4673 1547 4687
rect 1433 4653 1447 4667
rect 1433 4633 1447 4647
rect 1513 4633 1527 4647
rect 1353 4593 1367 4607
rect 753 4493 767 4507
rect 1253 4493 1267 4507
rect 1293 4493 1307 4507
rect 1393 4493 1407 4507
rect 453 4453 467 4467
rect 433 4333 447 4347
rect 633 4413 647 4427
rect 233 4153 247 4167
rect 273 4153 287 4167
rect 453 4153 467 4167
rect 233 4013 247 4027
rect 333 4013 347 4027
rect 373 4013 387 4027
rect 213 3993 227 4007
rect 253 3993 267 4007
rect 293 3993 307 4007
rect 233 3973 247 3987
rect 293 3753 307 3767
rect 413 3993 427 4007
rect 513 4173 527 4187
rect 713 4473 727 4487
rect 733 4213 747 4227
rect 913 4473 927 4487
rect 1213 4473 1227 4487
rect 1233 4453 1247 4467
rect 1293 4453 1307 4467
rect 1253 4433 1267 4447
rect 893 4413 907 4427
rect 973 4273 987 4287
rect 693 4173 707 4187
rect 753 4173 767 4187
rect 1193 4213 1207 4227
rect 1273 4273 1287 4287
rect 1213 4193 1227 4207
rect 793 4153 807 4167
rect 953 4153 967 4167
rect 633 4013 647 4027
rect 733 4013 747 4027
rect 933 4013 947 4027
rect 1073 4013 1087 4027
rect 1213 4013 1227 4027
rect 533 3993 547 4007
rect 593 3993 607 4007
rect 433 3733 447 3747
rect 473 3733 487 3747
rect 333 3693 347 3707
rect 213 3673 227 3687
rect 253 3533 267 3547
rect 33 3253 47 3267
rect 233 3513 247 3527
rect 953 3953 967 3967
rect 1013 3753 1027 3767
rect 1173 3993 1187 4007
rect 1193 3973 1207 3987
rect 1233 3953 1247 3967
rect 773 3713 787 3727
rect 473 3693 487 3707
rect 533 3693 547 3707
rect 753 3693 767 3707
rect 513 3673 527 3687
rect 793 3673 807 3687
rect 453 3533 467 3547
rect 493 3533 507 3547
rect 433 3513 447 3527
rect 473 3493 487 3507
rect 453 3473 467 3487
rect 493 3273 507 3287
rect 853 3713 867 3727
rect 753 3653 767 3667
rect 833 3653 847 3667
rect 713 3513 727 3527
rect 773 3533 787 3547
rect 533 3493 547 3507
rect 213 3253 227 3267
rect 513 3253 527 3267
rect 173 3233 187 3247
rect 253 3213 267 3227
rect 213 3053 227 3067
rect 193 3033 207 3047
rect 513 3213 527 3227
rect 493 3193 507 3207
rect 473 3053 487 3067
rect 493 3053 507 3067
rect 733 3473 747 3487
rect 553 3273 567 3287
rect 533 3193 547 3207
rect 253 3033 267 3047
rect 513 3033 527 3047
rect 473 3013 487 3027
rect 713 3253 727 3267
rect 773 3233 787 3247
rect 733 3213 747 3227
rect 713 3193 727 3207
rect 793 3193 807 3207
rect 753 3073 767 3087
rect 793 3073 807 3087
rect 693 3013 707 3027
rect 733 3013 747 3027
rect 213 2753 227 2767
rect 253 2753 267 2767
rect 313 2753 327 2767
rect 473 2753 487 2767
rect 513 2753 527 2767
rect 93 2733 107 2747
rect 13 2333 27 2347
rect 13 2133 27 2147
rect 213 2693 227 2707
rect 453 2733 467 2747
rect 493 2713 507 2727
rect 313 2693 327 2707
rect 493 2533 507 2547
rect 513 2513 527 2527
rect 693 2793 707 2807
rect 573 2713 587 2727
rect 473 2493 487 2507
rect 553 2493 567 2507
rect 773 2793 787 2807
rect 733 2773 747 2787
rect 833 3053 847 3067
rect 833 3013 847 3027
rect 753 2753 767 2767
rect 1033 3673 1047 3687
rect 1033 3533 1047 3547
rect 1533 4593 1547 4607
rect 1513 4473 1527 4487
rect 1573 4613 1587 4627
rect 1553 4473 1567 4487
rect 1673 4493 1687 4507
rect 1713 4473 1727 4487
rect 1493 4453 1507 4467
rect 1533 4453 1547 4467
rect 1593 4453 1607 4467
rect 1433 4433 1447 4447
rect 1393 4413 1407 4427
rect 1293 4193 1307 4207
rect 1333 3993 1347 4007
rect 1553 4213 1567 4227
rect 1413 4193 1427 4207
rect 1513 4193 1527 4207
rect 1473 4173 1487 4187
rect 1753 4673 1767 4687
rect 1793 4673 1807 4687
rect 1773 4653 1787 4667
rect 1753 4633 1767 4647
rect 1773 4473 1787 4487
rect 4293 4813 4307 4827
rect 2893 4793 2907 4807
rect 2333 4693 2347 4707
rect 2633 4693 2647 4707
rect 2293 4653 2307 4667
rect 2033 4633 2047 4647
rect 1833 4593 1847 4607
rect 2573 4653 2587 4667
rect 1913 4493 1927 4507
rect 2033 4493 2047 4507
rect 2293 4493 2307 4507
rect 2353 4493 2367 4507
rect 2473 4493 2487 4507
rect 2793 4653 2807 4667
rect 2833 4653 2847 4667
rect 4153 4733 4167 4747
rect 3933 4713 3947 4727
rect 3133 4693 3147 4707
rect 2633 4613 2647 4627
rect 1833 4473 1847 4487
rect 1953 4473 1967 4487
rect 2253 4473 2267 4487
rect 1813 4453 1827 4467
rect 2273 4453 2287 4467
rect 2313 4453 2327 4467
rect 1993 4333 2007 4347
rect 1773 4213 1787 4227
rect 1413 4013 1427 4027
rect 1353 3953 1367 3967
rect 1253 3673 1267 3687
rect 1293 3673 1307 3687
rect 1313 3673 1327 3687
rect 1253 3513 1267 3527
rect 1073 3373 1087 3387
rect 993 3233 1007 3247
rect 1013 3213 1027 3227
rect 873 3053 887 3067
rect 1013 3053 1027 3067
rect 973 3033 987 3047
rect 993 3013 1007 3027
rect 1053 3193 1067 3207
rect 873 2773 887 2787
rect 973 2713 987 2727
rect 1013 2693 1027 2707
rect 1113 2633 1127 2647
rect 853 2593 867 2607
rect 1013 2593 1027 2607
rect 773 2553 787 2567
rect 813 2553 827 2567
rect 693 2513 707 2527
rect 753 2513 767 2527
rect 233 2473 247 2487
rect 573 2473 587 2487
rect 193 2313 207 2327
rect 193 2293 207 2307
rect 493 2273 507 2287
rect 573 2273 587 2287
rect 353 2253 367 2267
rect 173 2213 187 2227
rect 133 2093 147 2107
rect 353 2093 367 2107
rect 393 2073 407 2087
rect 273 2053 287 2067
rect 213 1953 227 1967
rect 293 1953 307 1967
rect 273 1853 287 1867
rect 233 1813 247 1827
rect 273 1793 287 1807
rect 313 1853 327 1867
rect 113 1773 127 1787
rect 213 1773 227 1787
rect 293 1773 307 1787
rect 253 1553 267 1567
rect 213 1533 227 1547
rect 233 1293 247 1307
rect 273 1293 287 1307
rect 213 1273 227 1287
rect 213 1253 227 1267
rect 153 1073 167 1087
rect 193 1073 207 1087
rect 233 1073 247 1087
rect 713 2273 727 2287
rect 613 2213 627 2227
rect 553 2053 567 2067
rect 593 2053 607 2067
rect 493 1813 507 1827
rect 773 2253 787 2267
rect 733 2113 747 2127
rect 693 2073 707 2087
rect 713 2053 727 2067
rect 533 1793 547 1807
rect 613 1793 627 1807
rect 473 1773 487 1787
rect 513 1773 527 1787
rect 493 1753 507 1767
rect 433 1593 447 1607
rect 473 1593 487 1607
rect 513 1593 527 1607
rect 533 1593 547 1607
rect 753 1753 767 1767
rect 793 1753 807 1767
rect 773 1733 787 1747
rect 773 1573 787 1587
rect 533 1553 547 1567
rect 433 1533 447 1547
rect 313 1293 327 1307
rect 1093 2533 1107 2547
rect 973 2333 987 2347
rect 1033 2333 1047 2347
rect 953 2253 967 2267
rect 873 2233 887 2247
rect 1073 2273 1087 2287
rect 1053 2233 1067 2247
rect 973 2213 987 2227
rect 1013 2133 1027 2147
rect 953 1833 967 1847
rect 913 1773 927 1787
rect 1013 1773 1027 1787
rect 893 1733 907 1747
rect 673 1373 687 1387
rect 713 1373 727 1387
rect 773 1373 787 1387
rect 813 1373 827 1387
rect 653 1313 667 1327
rect 713 1313 727 1327
rect 793 1353 807 1367
rect 673 1293 687 1307
rect 453 1253 467 1267
rect 433 1233 447 1247
rect 493 1273 507 1287
rect 653 1273 667 1287
rect 733 1293 747 1307
rect 693 1253 707 1267
rect 493 1233 507 1247
rect 473 1133 487 1147
rect 533 1153 547 1167
rect 753 1153 767 1167
rect 793 1153 807 1167
rect 813 1153 827 1167
rect 533 1133 547 1147
rect 573 1133 587 1147
rect 453 1093 467 1107
rect 513 1093 527 1107
rect 253 813 267 827
rect 233 773 247 787
rect 193 653 207 667
rect 793 1073 807 1087
rect 473 833 487 847
rect 693 833 707 847
rect 673 813 687 827
rect 713 813 727 827
rect 453 793 467 807
rect 493 793 507 807
rect 493 633 507 647
rect 473 613 487 627
rect 433 593 447 607
rect 473 593 487 607
rect 713 653 727 667
rect 833 873 847 887
rect 833 813 847 827
rect 793 773 807 787
rect 693 373 707 387
rect 233 313 247 327
rect 453 313 467 327
rect 673 313 687 327
rect 273 293 287 307
rect 233 133 247 147
rect 533 193 547 207
rect 473 153 487 167
rect 493 113 507 127
rect 213 93 227 107
rect 933 1593 947 1607
rect 973 1573 987 1587
rect 1233 2733 1247 2747
rect 1293 3193 1307 3207
rect 1273 3013 1287 3027
rect 1313 3013 1327 3027
rect 1213 2273 1227 2287
rect 1153 2253 1167 2267
rect 1213 2253 1227 2267
rect 1273 2633 1287 2647
rect 1253 2593 1267 2607
rect 1293 2553 1307 2567
rect 1393 3873 1407 3887
rect 1433 3873 1447 3887
rect 1453 3653 1467 3667
rect 1593 4173 1607 4187
rect 1753 4033 1767 4047
rect 1733 4013 1747 4027
rect 1693 3993 1707 4007
rect 1493 3973 1507 3987
rect 1553 3713 1567 3727
rect 1673 3713 1687 3727
rect 1473 3633 1487 3647
rect 1513 3513 1527 3527
rect 1693 3693 1707 3707
rect 1653 3653 1667 3667
rect 2053 4193 2067 4207
rect 2013 4173 2027 4187
rect 2293 4193 2307 4207
rect 2313 4173 2327 4187
rect 2033 4033 2047 4047
rect 2253 4033 2267 4047
rect 2273 4033 2287 4047
rect 2313 4033 2327 4047
rect 2233 4013 2247 4027
rect 2273 4013 2287 4027
rect 1753 3953 1767 3967
rect 1973 3953 1987 3967
rect 2013 3953 2027 3967
rect 2093 3793 2107 3807
rect 1733 3693 1747 3707
rect 1933 3673 1947 3687
rect 1853 3653 1867 3667
rect 1713 3633 1727 3647
rect 2093 3533 2107 3547
rect 1773 3513 1787 3527
rect 1813 3513 1827 3527
rect 1853 3513 1867 3527
rect 1713 3493 1727 3507
rect 1533 3473 1547 3487
rect 1713 3253 1727 3267
rect 1793 3493 1807 3507
rect 2073 3493 2087 3507
rect 2113 3473 2127 3487
rect 1833 3373 1847 3387
rect 1913 3373 1927 3387
rect 1673 3233 1687 3247
rect 1413 3213 1427 3227
rect 1553 3173 1567 3187
rect 1633 3173 1647 3187
rect 1453 3033 1467 3047
rect 1413 3013 1427 3027
rect 1453 3013 1467 3027
rect 1833 3233 1847 3247
rect 1853 3233 1867 3247
rect 1773 3213 1787 3227
rect 1713 3193 1727 3207
rect 1813 3193 1827 3207
rect 1473 2773 1487 2787
rect 1673 2773 1687 2787
rect 1453 2713 1467 2727
rect 1533 2613 1547 2627
rect 1353 2573 1367 2587
rect 1313 2313 1327 2327
rect 1313 2293 1327 2307
rect 1353 2273 1367 2287
rect 1553 2513 1567 2527
rect 1573 2333 1587 2347
rect 1733 2633 1747 2647
rect 1833 2633 1847 2647
rect 1793 2613 1807 2627
rect 1733 2573 1747 2587
rect 1693 2553 1707 2567
rect 1773 2553 1787 2567
rect 1693 2533 1707 2547
rect 1753 2533 1767 2547
rect 1693 2513 1707 2527
rect 1673 2293 1687 2307
rect 1573 2273 1587 2287
rect 1633 2273 1647 2287
rect 1293 2253 1307 2267
rect 1333 2253 1347 2267
rect 1513 2253 1527 2267
rect 1613 2253 1627 2267
rect 1733 2273 1747 2287
rect 1313 2213 1327 2227
rect 1513 2213 1527 2227
rect 1233 2133 1247 2147
rect 1233 2113 1247 2127
rect 1273 2093 1287 2107
rect 1213 2053 1227 2067
rect 1293 2053 1307 2067
rect 1253 2033 1267 2047
rect 1213 1813 1227 1827
rect 1253 1813 1267 1827
rect 1353 2093 1367 2107
rect 1333 2073 1347 2087
rect 1353 2053 1367 2067
rect 1653 2093 1667 2107
rect 1533 2073 1547 2087
rect 1553 2053 1567 2067
rect 1333 2033 1347 2047
rect 1593 2013 1607 2027
rect 1433 1833 1447 1847
rect 1233 1773 1247 1787
rect 1713 2053 1727 2067
rect 1953 3273 1967 3287
rect 2073 3273 2087 3287
rect 1913 3193 1927 3207
rect 1853 2533 1867 2547
rect 2033 3253 2047 3267
rect 2333 3713 2347 3727
rect 2373 3653 2387 3667
rect 2313 3633 2327 3647
rect 2313 3533 2327 3547
rect 2593 4473 2607 4487
rect 2553 4453 2567 4467
rect 2953 4513 2967 4527
rect 2853 4493 2867 4507
rect 2813 4473 2827 4487
rect 2613 4453 2627 4467
rect 2593 4353 2607 4367
rect 2533 4333 2547 4347
rect 2573 4173 2587 4187
rect 2833 4453 2847 4467
rect 2793 4213 2807 4227
rect 3393 4693 3407 4707
rect 3933 4693 3947 4707
rect 4073 4693 4087 4707
rect 4113 4693 4127 4707
rect 3373 4673 3387 4687
rect 3573 4673 3587 4687
rect 3613 4673 3627 4687
rect 3653 4673 3667 4687
rect 3173 4633 3187 4647
rect 3333 4633 3347 4647
rect 3553 4633 3567 4647
rect 3133 4533 3147 4547
rect 3373 4533 3387 4547
rect 3133 4493 3147 4507
rect 3173 4493 3187 4507
rect 3353 4493 3367 4507
rect 3113 4473 3127 4487
rect 3093 4433 3107 4447
rect 3073 4353 3087 4367
rect 2773 4193 2787 4207
rect 2813 4193 2827 4207
rect 2953 4193 2967 4207
rect 3153 4193 3167 4207
rect 3073 4173 3087 4187
rect 2513 4013 2527 4027
rect 2853 4153 2867 4167
rect 2873 4153 2887 4167
rect 2773 4133 2787 4147
rect 2833 4133 2847 4147
rect 2553 3993 2567 4007
rect 2753 3993 2767 4007
rect 2513 3913 2527 3927
rect 2493 3713 2507 3727
rect 2493 3553 2507 3567
rect 2473 3533 2487 3547
rect 2293 3513 2307 3527
rect 2333 3513 2347 3527
rect 2373 3513 2387 3527
rect 2493 3493 2507 3507
rect 2253 3273 2267 3287
rect 2773 3933 2787 3947
rect 2753 3733 2767 3747
rect 2573 3673 2587 3687
rect 2753 3673 2767 3687
rect 2553 3633 2567 3647
rect 2593 3633 2607 3647
rect 2613 3633 2627 3647
rect 2533 3553 2547 3567
rect 2553 3533 2567 3547
rect 2593 3513 2607 3527
rect 2533 3493 2547 3507
rect 2573 3493 2587 3507
rect 2613 3493 2627 3507
rect 2073 3033 2087 3047
rect 2093 3033 2107 3047
rect 1953 2773 1967 2787
rect 1993 2773 2007 2787
rect 2253 3193 2267 3207
rect 2313 3153 2327 3167
rect 2213 3073 2227 3087
rect 2173 3053 2187 3067
rect 2213 3033 2227 3047
rect 2113 2733 2127 2747
rect 2173 2753 2187 2767
rect 2113 2693 2127 2707
rect 2013 2633 2027 2647
rect 2033 2633 2047 2647
rect 1993 2553 2007 2567
rect 2073 2553 2087 2567
rect 2013 2533 2027 2547
rect 2033 2533 2047 2547
rect 1993 2513 2007 2527
rect 1973 2333 1987 2347
rect 1953 2313 1967 2327
rect 1893 2293 1907 2307
rect 1873 2273 1887 2287
rect 1913 2273 1927 2287
rect 1893 2253 1907 2267
rect 1753 2093 1767 2107
rect 1893 2073 1907 2087
rect 1233 1733 1247 1747
rect 1213 1633 1227 1647
rect 1533 1773 1547 1787
rect 1653 1773 1667 1787
rect 1793 1793 1807 1807
rect 1713 1753 1727 1767
rect 1773 1753 1787 1767
rect 1413 1733 1427 1747
rect 1813 1733 1827 1747
rect 1533 1713 1547 1727
rect 1273 1633 1287 1647
rect 1253 1613 1267 1627
rect 1453 1593 1467 1607
rect 1493 1593 1507 1607
rect 1253 1573 1267 1587
rect 993 1553 1007 1567
rect 1093 1553 1107 1567
rect 953 1353 967 1367
rect 973 1353 987 1367
rect 933 1333 947 1347
rect 1013 1333 1027 1347
rect 993 1293 1007 1307
rect 953 1273 967 1287
rect 933 1073 947 1087
rect 1053 1193 1067 1207
rect 1333 1333 1347 1347
rect 1233 1293 1247 1307
rect 1293 1293 1307 1307
rect 1093 1133 1107 1147
rect 1273 1273 1287 1287
rect 1513 1373 1527 1387
rect 1473 1353 1487 1367
rect 1533 1353 1547 1367
rect 1513 1333 1527 1347
rect 1453 1313 1467 1327
rect 1493 1313 1507 1327
rect 1333 1153 1347 1167
rect 1293 1133 1307 1147
rect 1373 1133 1387 1147
rect 953 833 967 847
rect 993 833 1007 847
rect 1113 1093 1127 1107
rect 1253 1093 1267 1107
rect 1353 873 1367 887
rect 1313 853 1327 867
rect 1233 833 1247 847
rect 973 813 987 827
rect 1073 813 1087 827
rect 1493 853 1507 867
rect 1453 833 1467 847
rect 1533 833 1547 847
rect 1513 813 1527 827
rect 1673 1333 1687 1347
rect 1593 1133 1607 1147
rect 1693 853 1707 867
rect 1573 813 1587 827
rect 1633 813 1647 827
rect 953 793 967 807
rect 1253 793 1267 807
rect 1313 793 1327 807
rect 1353 793 1367 807
rect 1473 793 1487 807
rect 1533 793 1547 807
rect 933 633 947 647
rect 993 633 1007 647
rect 1233 613 1247 627
rect 973 593 987 607
rect 1193 593 1207 607
rect 1013 493 1027 507
rect 1053 493 1067 507
rect 973 393 987 407
rect 1013 373 1027 387
rect 753 293 767 307
rect 913 293 927 307
rect 1013 353 1027 367
rect 773 273 787 287
rect 993 273 1007 287
rect 973 193 987 207
rect 793 173 807 187
rect 753 153 767 167
rect 813 153 827 167
rect 993 173 1007 187
rect 1253 353 1267 367
rect 1293 353 1307 367
rect 1493 673 1507 687
rect 1453 653 1467 667
rect 1633 633 1647 647
rect 1433 613 1447 627
rect 1473 613 1487 627
rect 1533 493 1547 507
rect 1333 373 1347 387
rect 1033 333 1047 347
rect 1053 333 1067 347
rect 1233 333 1247 347
rect 1273 333 1287 347
rect 1313 333 1327 347
rect 1013 153 1027 167
rect 1313 313 1327 327
rect 1233 293 1247 307
rect 1233 193 1247 207
rect 1233 173 1247 187
rect 1253 153 1267 167
rect 1033 133 1047 147
rect 1473 213 1487 227
rect 1333 173 1347 187
rect 1433 173 1447 187
rect 1553 373 1567 387
rect 1533 353 1547 367
rect 1773 1333 1787 1347
rect 1753 1293 1767 1307
rect 1793 1173 1807 1187
rect 1733 1133 1747 1147
rect 1993 2293 2007 2307
rect 2033 2273 2047 2287
rect 2053 2173 2067 2187
rect 1993 2113 2007 2127
rect 1993 2073 2007 2087
rect 2033 2073 2047 2087
rect 2073 2073 2087 2087
rect 2073 2053 2087 2067
rect 2073 1833 2087 1847
rect 1953 1573 1967 1587
rect 1893 1133 1907 1147
rect 2053 1773 2067 1787
rect 2093 1693 2107 1707
rect 2153 2653 2167 2667
rect 2293 2653 2307 2667
rect 2373 3053 2387 3067
rect 2453 3033 2467 3047
rect 2393 3013 2407 3027
rect 2553 3193 2567 3207
rect 2573 3153 2587 3167
rect 2533 3073 2547 3087
rect 2573 3073 2587 3087
rect 2513 3013 2527 3027
rect 2453 2773 2467 2787
rect 2693 2753 2707 2767
rect 2373 2733 2387 2747
rect 2333 2713 2347 2727
rect 2473 2713 2487 2727
rect 2673 2713 2687 2727
rect 2313 2593 2327 2607
rect 2273 2553 2287 2567
rect 2333 2553 2347 2567
rect 2413 2553 2427 2567
rect 2513 2553 2527 2567
rect 2553 2553 2567 2567
rect 2673 2553 2687 2567
rect 2333 2493 2347 2507
rect 2133 2253 2147 2267
rect 2193 2253 2207 2267
rect 2213 2173 2227 2187
rect 2253 2173 2267 2187
rect 2193 2053 2207 2067
rect 2273 2053 2287 2067
rect 2153 2033 2167 2047
rect 2333 2253 2347 2267
rect 2353 2253 2367 2267
rect 3093 4133 3107 4147
rect 3113 4113 3127 4127
rect 3113 3973 3127 3987
rect 3033 3953 3047 3967
rect 2853 3933 2867 3947
rect 2833 3773 2847 3787
rect 2893 3733 2907 3747
rect 2793 3713 2807 3727
rect 2873 3693 2887 3707
rect 2853 3633 2867 3647
rect 2813 3513 2827 3527
rect 2833 3513 2847 3527
rect 2813 3473 2827 3487
rect 2853 3473 2867 3487
rect 2853 3273 2867 3287
rect 3093 3953 3107 3967
rect 3053 3753 3067 3767
rect 3053 3733 3067 3747
rect 3073 3733 3087 3747
rect 3113 3733 3127 3747
rect 3033 3713 3047 3727
rect 2913 3673 2927 3687
rect 2813 3013 2827 3027
rect 2873 3213 2887 3227
rect 2873 3053 2887 3067
rect 2853 3033 2867 3047
rect 3093 3713 3107 3727
rect 3333 4473 3347 4487
rect 3353 4453 3367 4467
rect 3293 4193 3307 4207
rect 3333 4193 3347 4207
rect 3173 3973 3187 3987
rect 3413 4193 3427 4207
rect 3353 4173 3367 4187
rect 3373 4133 3387 4147
rect 3333 4033 3347 4047
rect 3873 4633 3887 4647
rect 3893 4633 3907 4647
rect 3673 4553 3687 4567
rect 3913 4553 3927 4567
rect 3633 4513 3647 4527
rect 3673 4473 3687 4487
rect 3613 4453 3627 4467
rect 3633 4433 3647 4447
rect 3573 4213 3587 4227
rect 3633 4213 3647 4227
rect 3373 3993 3387 4007
rect 3493 3993 3507 4007
rect 3313 3953 3327 3967
rect 3353 3953 3367 3967
rect 3273 3753 3287 3767
rect 3173 3733 3187 3747
rect 3173 3513 3187 3527
rect 3113 3493 3127 3507
rect 3093 3473 3107 3487
rect 3053 3453 3067 3467
rect 3133 3453 3147 3467
rect 3093 3233 3107 3247
rect 3153 3233 3167 3247
rect 2913 3213 2927 3227
rect 3073 3193 3087 3207
rect 3113 3073 3127 3087
rect 3093 3053 3107 3067
rect 3133 3053 3147 3067
rect 2833 2753 2847 2767
rect 2953 2753 2967 2767
rect 2973 2733 2987 2747
rect 2933 2713 2947 2727
rect 3253 3493 3267 3507
rect 3253 3253 3267 3267
rect 3293 3713 3307 3727
rect 3553 3993 3567 4007
rect 3513 3793 3527 3807
rect 3533 3793 3547 3807
rect 3413 3733 3427 3747
rect 3333 3713 3347 3727
rect 3373 3713 3387 3727
rect 3393 3673 3407 3687
rect 3893 4473 3907 4487
rect 4073 4493 4087 4507
rect 3913 4453 3927 4467
rect 3833 4213 3847 4227
rect 3673 4193 3687 4207
rect 3653 4133 3667 4147
rect 3913 4153 3927 4167
rect 3833 4113 3847 4127
rect 3613 4033 3627 4047
rect 3613 3993 3627 4007
rect 3793 3993 3807 4007
rect 3853 4013 3867 4027
rect 3993 4033 4007 4047
rect 3873 3993 3887 4007
rect 3913 3993 3927 4007
rect 3553 3673 3567 3687
rect 3573 3533 3587 3547
rect 3333 3513 3347 3527
rect 3373 3513 3387 3527
rect 3413 3513 3427 3527
rect 3453 3513 3467 3527
rect 3493 3513 3507 3527
rect 3533 3513 3547 3527
rect 3293 3493 3307 3507
rect 3313 3233 3327 3247
rect 3353 3493 3367 3507
rect 3393 3473 3407 3487
rect 3393 3273 3407 3287
rect 3373 3213 3387 3227
rect 3653 3733 3667 3747
rect 3633 3673 3647 3687
rect 3773 3493 3787 3507
rect 3593 3473 3607 3487
rect 3773 3473 3787 3487
rect 3533 3453 3547 3467
rect 3333 3173 3347 3187
rect 3273 3033 3287 3047
rect 3233 2753 3247 2767
rect 2813 2553 2827 2567
rect 2973 2553 2987 2567
rect 3073 2553 3087 2567
rect 3113 2553 3127 2567
rect 3153 2553 3167 2567
rect 2813 2533 2827 2547
rect 2793 2513 2807 2527
rect 2653 2253 2667 2267
rect 2493 2233 2507 2247
rect 2573 2233 2587 2247
rect 2713 2233 2727 2247
rect 2413 2133 2427 2147
rect 2393 1833 2407 1847
rect 2373 1813 2387 1827
rect 2333 1793 2347 1807
rect 2333 1753 2347 1767
rect 2353 1753 2367 1767
rect 2393 1753 2407 1767
rect 2313 1613 2327 1627
rect 2173 1573 2187 1587
rect 2293 1573 2307 1587
rect 2313 1573 2327 1587
rect 2333 1553 2347 1567
rect 2533 2073 2547 2087
rect 2553 2053 2567 2067
rect 2513 2033 2527 2047
rect 2533 2033 2547 2047
rect 2833 2493 2847 2507
rect 2933 2273 2947 2287
rect 3253 2733 3267 2747
rect 3053 2533 3067 2547
rect 3213 2533 3227 2547
rect 3093 2493 3107 2507
rect 3033 2273 3047 2287
rect 3213 2273 3227 2287
rect 2953 2253 2967 2267
rect 2993 2233 3007 2247
rect 2833 2073 2847 2087
rect 2773 2053 2787 2067
rect 2813 2053 2827 2067
rect 2793 2033 2807 2047
rect 3233 2253 3247 2267
rect 3193 2233 3207 2247
rect 3193 2073 3207 2087
rect 2613 1813 2627 1827
rect 2533 1793 2547 1807
rect 2593 1793 2607 1807
rect 2573 1633 2587 1647
rect 2433 1613 2447 1627
rect 2473 1613 2487 1627
rect 2733 1593 2747 1607
rect 2453 1573 2467 1587
rect 2453 1553 2467 1567
rect 2693 1553 2707 1567
rect 2253 1293 2267 1307
rect 2053 1273 2067 1287
rect 2113 1273 2127 1287
rect 2413 1293 2427 1307
rect 2033 1253 2047 1267
rect 2293 1253 2307 1267
rect 2433 1153 2447 1167
rect 2153 1133 2167 1147
rect 1933 1113 1947 1127
rect 2013 1113 2027 1127
rect 2173 1113 2187 1127
rect 2193 1113 2207 1127
rect 2333 1113 2347 1127
rect 1793 853 1807 867
rect 1913 853 1927 867
rect 1753 813 1767 827
rect 1773 793 1787 807
rect 2013 813 2027 827
rect 2233 813 2247 827
rect 2173 793 2187 807
rect 1893 753 1907 767
rect 1993 673 2007 687
rect 1793 653 1807 667
rect 1973 653 1987 667
rect 2013 653 2027 667
rect 1793 633 1807 647
rect 1813 633 1827 647
rect 1733 613 1747 627
rect 1773 613 1787 627
rect 1773 593 1787 607
rect 1753 293 1767 307
rect 1933 373 1947 387
rect 2053 593 2067 607
rect 1993 373 2007 387
rect 1973 353 1987 367
rect 2013 353 2027 367
rect 2273 793 2287 807
rect 2233 673 2247 687
rect 2253 673 2267 687
rect 2273 653 2287 667
rect 2313 653 2327 667
rect 2493 1333 2507 1347
rect 2513 1293 2527 1307
rect 2553 1153 2567 1167
rect 2533 1133 2547 1147
rect 2513 1113 2527 1127
rect 2473 1093 2487 1107
rect 2533 1093 2547 1107
rect 2473 873 2487 887
rect 2513 873 2527 887
rect 2413 833 2427 847
rect 2493 833 2507 847
rect 2913 1833 2927 1847
rect 2993 1833 3007 1847
rect 2853 1813 2867 1827
rect 2873 1633 2887 1647
rect 3033 1773 3047 1787
rect 3193 1753 3207 1767
rect 3053 1733 3067 1747
rect 3193 1733 3207 1747
rect 2973 1613 2987 1627
rect 2993 1613 3007 1627
rect 2933 1593 2947 1607
rect 2813 1553 2827 1567
rect 3053 1553 3067 1567
rect 2773 1533 2787 1547
rect 3333 3033 3347 3047
rect 3413 3193 3427 3207
rect 3413 3173 3427 3187
rect 3393 2993 3407 3007
rect 3293 2733 3307 2747
rect 3393 2713 3407 2727
rect 3333 2653 3347 2667
rect 3273 2113 3287 2127
rect 3353 2533 3367 2547
rect 3313 2493 3327 2507
rect 3473 2733 3487 2747
rect 3493 2653 3507 2667
rect 3513 2593 3527 2607
rect 3413 2493 3427 2507
rect 3393 2273 3407 2287
rect 3473 2253 3487 2267
rect 3553 3213 3567 3227
rect 3673 3213 3687 3227
rect 3633 3053 3647 3067
rect 3673 3033 3687 3047
rect 3613 3013 3627 3027
rect 3773 3013 3787 3027
rect 3653 2993 3667 3007
rect 3833 3773 3847 3787
rect 3813 3713 3827 3727
rect 3893 3713 3907 3727
rect 3953 3693 3967 3707
rect 3913 3673 3927 3687
rect 3933 3673 3947 3687
rect 3873 3533 3887 3547
rect 3893 3493 3907 3507
rect 3873 3473 3887 3487
rect 3913 3473 3927 3487
rect 4093 4473 4107 4487
rect 4153 4473 4167 4487
rect 4113 4453 4127 4467
rect 4193 4453 4207 4467
rect 4093 4213 4107 4227
rect 4133 4213 4147 4227
rect 4093 4153 4107 4167
rect 4133 4013 4147 4027
rect 4113 3993 4127 4007
rect 4073 3733 4087 3747
rect 4193 3713 4207 3727
rect 4173 3693 4187 3707
rect 4013 3513 4027 3527
rect 4033 3513 4047 3527
rect 3953 3473 3967 3487
rect 3873 3253 3887 3267
rect 3933 3253 3947 3267
rect 3813 3153 3827 3167
rect 3633 2973 3647 2987
rect 3793 2973 3807 2987
rect 3553 2753 3567 2767
rect 3753 2773 3767 2787
rect 3713 2733 3727 2747
rect 3673 2593 3687 2607
rect 3693 2593 3707 2607
rect 3713 2573 3727 2587
rect 3553 2533 3567 2547
rect 3613 2533 3627 2547
rect 3653 2533 3667 2547
rect 3573 2253 3587 2267
rect 3613 2073 3627 2087
rect 3433 2013 3447 2027
rect 3353 1813 3367 1827
rect 3333 1773 3347 1787
rect 3613 2013 3627 2027
rect 3573 1993 3587 2007
rect 3533 1813 3547 1827
rect 3393 1753 3407 1767
rect 3293 1713 3307 1727
rect 3253 1673 3267 1687
rect 3293 1673 3307 1687
rect 3513 1733 3527 1747
rect 3513 1613 3527 1627
rect 3553 1753 3567 1767
rect 3553 1593 3567 1607
rect 3273 1553 3287 1567
rect 3313 1553 3327 1567
rect 3393 1553 3407 1567
rect 3193 1313 3207 1327
rect 2773 1273 2787 1287
rect 2753 1153 2767 1167
rect 2713 1113 2727 1127
rect 2973 1133 2987 1147
rect 3013 1113 3027 1127
rect 2993 1093 3007 1107
rect 2953 1073 2967 1087
rect 3093 1293 3107 1307
rect 3173 1173 3187 1187
rect 3073 1153 3087 1167
rect 3133 1113 3147 1127
rect 3313 1533 3327 1547
rect 3313 1313 3327 1327
rect 3513 1313 3527 1327
rect 3553 1313 3567 1327
rect 3593 1313 3607 1327
rect 3273 1293 3287 1307
rect 3213 1173 3227 1187
rect 3193 1073 3207 1087
rect 2833 873 2847 887
rect 2773 833 2787 847
rect 2813 833 2827 847
rect 2693 813 2707 827
rect 2553 773 2567 787
rect 2413 733 2427 747
rect 2293 613 2307 627
rect 2333 613 2347 627
rect 2173 353 2187 367
rect 2253 353 2267 367
rect 2053 313 2067 327
rect 1933 293 1947 307
rect 1813 213 1827 227
rect 1793 193 1807 207
rect 2233 193 2247 207
rect 1693 173 1707 187
rect 1493 153 1507 167
rect 1653 153 1667 167
rect 2053 173 2067 187
rect 2093 173 2107 187
rect 2113 173 2127 187
rect 2293 333 2307 347
rect 2013 153 2027 167
rect 2033 133 2047 147
rect 2073 133 2087 147
rect 2293 173 2307 187
rect 2313 173 2327 187
rect 2253 153 2267 167
rect 2273 153 2287 167
rect 2793 793 2807 807
rect 2833 793 2847 807
rect 3053 853 3067 867
rect 3033 833 3047 847
rect 2873 773 2887 787
rect 2993 773 3007 787
rect 2833 753 2847 767
rect 2813 673 2827 687
rect 2553 653 2567 667
rect 2753 653 2767 667
rect 2593 633 2607 647
rect 2793 633 2807 647
rect 2853 633 2867 647
rect 2573 613 2587 627
rect 2613 613 2627 627
rect 2533 593 2547 607
rect 2533 573 2547 587
rect 2533 353 2547 367
rect 2413 333 2427 347
rect 2553 333 2567 347
rect 2573 333 2587 347
rect 2513 293 2527 307
rect 2533 193 2547 207
rect 2333 153 2347 167
rect 2413 153 2427 167
rect 2613 353 2627 367
rect 2813 373 2827 387
rect 3113 813 3127 827
rect 3093 733 3107 747
rect 3613 1293 3627 1307
rect 3573 1273 3587 1287
rect 3513 1253 3527 1267
rect 3353 1193 3367 1207
rect 3273 853 3287 867
rect 3493 1113 3507 1127
rect 3953 3213 3967 3227
rect 4093 3213 4107 3227
rect 3933 3173 3947 3187
rect 4073 3173 4087 3187
rect 4153 3173 4167 3187
rect 3893 3073 3907 3087
rect 3973 3073 3987 3087
rect 4013 3073 4027 3087
rect 3913 3053 3927 3067
rect 3953 3033 3967 3047
rect 3893 3013 3907 3027
rect 3933 3013 3947 3027
rect 4133 3053 4147 3067
rect 4353 4813 4367 4827
rect 4393 4793 4407 4807
rect 4673 4753 4687 4767
rect 4673 4733 4687 4747
rect 4313 4653 4327 4667
rect 4393 4653 4407 4667
rect 4653 4693 4667 4707
rect 4393 4633 4407 4647
rect 4433 4633 4447 4647
rect 4593 4633 4607 4647
rect 4433 4473 4447 4487
rect 4473 4473 4487 4487
rect 4393 4433 4407 4447
rect 4453 4433 4467 4447
rect 4333 4413 4347 4427
rect 4413 4413 4427 4427
rect 4353 4193 4367 4207
rect 4393 4193 4407 4207
rect 4433 4193 4447 4207
rect 4333 4173 4347 4187
rect 4373 4173 4387 4187
rect 4413 4033 4427 4047
rect 4653 4493 4667 4507
rect 4853 4693 4867 4707
rect 4853 4653 4867 4667
rect 4893 4653 4907 4667
rect 4853 4633 4867 4647
rect 4713 4453 4727 4467
rect 4733 4453 4747 4467
rect 4633 4433 4647 4447
rect 4473 4193 4487 4207
rect 4593 4193 4607 4207
rect 4653 4193 4667 4207
rect 4453 3993 4467 4007
rect 4353 3953 4367 3967
rect 4393 3953 4407 3967
rect 4473 3953 4487 3967
rect 4673 4153 4687 4167
rect 4633 3973 4647 3987
rect 4653 3953 4667 3967
rect 4333 3913 4347 3927
rect 4333 3733 4347 3747
rect 4313 3493 4327 3507
rect 4293 3453 4307 3467
rect 4453 3733 4467 3747
rect 4693 3953 4707 3967
rect 4673 3733 4687 3747
rect 4433 3713 4447 3727
rect 4473 3713 4487 3727
rect 4393 3673 4407 3687
rect 4713 3673 4727 3687
rect 5013 4793 5027 4807
rect 4933 4673 4947 4687
rect 4993 4673 5007 4687
rect 4953 4453 4967 4467
rect 4933 4433 4947 4447
rect 4853 4153 4867 4167
rect 4793 4013 4807 4027
rect 4853 4013 4867 4027
rect 4813 3953 4827 3967
rect 4973 3713 4987 3727
rect 4893 3693 4907 3707
rect 4953 3693 4967 3707
rect 4913 3673 4927 3687
rect 4413 3533 4427 3547
rect 4613 3533 4627 3547
rect 4733 3533 4747 3547
rect 4793 3533 4807 3547
rect 4893 3533 4907 3547
rect 4913 3533 4927 3547
rect 4333 3473 4347 3487
rect 4353 3473 4367 3487
rect 4313 3273 4327 3287
rect 4413 3473 4427 3487
rect 4393 3413 4407 3427
rect 4373 3273 4387 3287
rect 4333 3233 4347 3247
rect 4413 3233 4427 3247
rect 4573 3233 4587 3247
rect 4193 3073 4207 3087
rect 4253 3053 4267 3067
rect 4013 3013 4027 3027
rect 4133 3013 4147 3027
rect 4173 3013 4187 3027
rect 4213 3013 4227 3027
rect 4033 2773 4047 2787
rect 4293 2773 4307 2787
rect 4273 2753 4287 2767
rect 4013 2733 4027 2747
rect 3973 2593 3987 2607
rect 3913 2573 3927 2587
rect 3933 2513 3947 2527
rect 3953 2493 3967 2507
rect 3933 2273 3947 2287
rect 3913 2073 3927 2087
rect 3833 2033 3847 2047
rect 3913 2033 3927 2047
rect 3873 1993 3887 2007
rect 3673 1773 3687 1787
rect 3713 1773 3727 1787
rect 3653 1733 3667 1747
rect 3753 1733 3767 1747
rect 3713 1693 3727 1707
rect 3653 1633 3667 1647
rect 3693 1613 3707 1627
rect 3653 1333 3667 1347
rect 3813 1753 3827 1767
rect 3793 1653 3807 1667
rect 3873 1713 3887 1727
rect 3893 1673 3907 1687
rect 3853 1613 3867 1627
rect 3833 1573 3847 1587
rect 3793 1333 3807 1347
rect 3693 1313 3707 1327
rect 3713 1313 3727 1327
rect 3633 1193 3647 1207
rect 3513 1093 3527 1107
rect 3533 1093 3547 1107
rect 3473 1073 3487 1087
rect 3773 1253 3787 1267
rect 3733 1173 3747 1187
rect 3753 1113 3767 1127
rect 3733 1093 3747 1107
rect 3953 1793 3967 1807
rect 3913 1053 3927 1067
rect 3593 873 3607 887
rect 3693 873 3707 887
rect 3773 873 3787 887
rect 3793 833 3807 847
rect 3833 833 3847 847
rect 3873 833 3887 847
rect 3433 813 3447 827
rect 3613 813 3627 827
rect 3673 813 3687 827
rect 3773 813 3787 827
rect 3213 713 3227 727
rect 3273 713 3287 727
rect 3153 633 3167 647
rect 3193 633 3207 647
rect 3313 653 3327 667
rect 3073 573 3087 587
rect 3133 573 3147 587
rect 2833 353 2847 367
rect 2793 333 2807 347
rect 2933 373 2947 387
rect 3113 373 3127 387
rect 2933 333 2947 347
rect 2993 333 3007 347
rect 3073 333 3087 347
rect 2873 313 2887 327
rect 2833 213 2847 227
rect 2593 153 2607 167
rect 2853 173 2867 187
rect 2873 153 2887 167
rect 2113 133 2127 147
rect 2333 133 2347 147
rect 2553 133 2567 147
rect 813 113 827 127
rect 2093 113 2107 127
rect 733 93 747 107
rect 3573 793 3587 807
rect 3613 773 3627 787
rect 3373 593 3387 607
rect 3353 373 3367 387
rect 3393 373 3407 387
rect 3633 593 3647 607
rect 3653 593 3667 607
rect 3793 793 3807 807
rect 3793 713 3807 727
rect 3753 633 3767 647
rect 3853 793 3867 807
rect 3813 633 3827 647
rect 4073 2733 4087 2747
rect 4053 2533 4067 2547
rect 3993 2273 4007 2287
rect 4033 2273 4047 2287
rect 4053 2233 4067 2247
rect 4133 2573 4147 2587
rect 4393 3213 4407 3227
rect 4433 3213 4447 3227
rect 4473 3053 4487 3067
rect 4433 3013 4447 3027
rect 4453 2993 4467 3007
rect 4413 2773 4427 2787
rect 4393 2753 4407 2767
rect 4413 2753 4427 2767
rect 4393 2553 4407 2567
rect 4533 3033 4547 3047
rect 4493 2753 4507 2767
rect 4753 3413 4767 3427
rect 4693 3253 4707 3267
rect 4653 3233 4667 3247
rect 4713 3213 4727 3227
rect 4733 3213 4747 3227
rect 4633 3193 4647 3207
rect 4673 3193 4687 3207
rect 4713 3053 4727 3067
rect 4693 3033 4707 3047
rect 4893 3273 4907 3287
rect 4873 3253 4887 3267
rect 4853 3233 4867 3247
rect 4753 3193 4767 3207
rect 4893 3213 4907 3227
rect 4853 3073 4867 3087
rect 4753 3053 4767 3067
rect 4753 2993 4767 3007
rect 4733 2753 4747 2767
rect 4473 2713 4487 2727
rect 4513 2713 4527 2727
rect 4693 2713 4707 2727
rect 4473 2573 4487 2587
rect 4653 2573 4667 2587
rect 4153 2533 4167 2547
rect 4353 2533 4367 2547
rect 4433 2513 4447 2527
rect 4353 2293 4367 2307
rect 4313 2253 4327 2267
rect 4273 2233 4287 2247
rect 4153 2093 4167 2107
rect 4093 2033 4107 2047
rect 4813 2753 4827 2767
rect 4753 2733 4767 2747
rect 4973 3653 4987 3667
rect 4933 3273 4947 3287
rect 4953 3233 4967 3247
rect 4993 3233 5007 3247
rect 4933 3213 4947 3227
rect 4973 3193 4987 3207
rect 4993 3073 5007 3087
rect 4913 3033 4927 3047
rect 4973 3053 4987 3067
rect 4893 3013 4907 3027
rect 4953 3013 4967 3027
rect 4793 2713 4807 2727
rect 4853 2553 4867 2567
rect 4733 2533 4747 2547
rect 4513 2313 4527 2327
rect 4733 2313 4747 2327
rect 4553 2293 4567 2307
rect 4473 2273 4487 2287
rect 4533 2273 4547 2287
rect 4633 2253 4647 2267
rect 4293 2093 4307 2107
rect 4353 2093 4367 2107
rect 4273 2053 4287 2067
rect 4373 2053 4387 2067
rect 4333 2033 4347 2047
rect 4013 1813 4027 1827
rect 4073 1813 4087 1827
rect 4253 1793 4267 1807
rect 4373 1793 4387 1807
rect 4653 2073 4667 2087
rect 4593 2013 4607 2027
rect 4093 1673 4107 1687
rect 4093 1653 4107 1667
rect 4133 1613 4147 1627
rect 4053 1273 4067 1287
rect 4013 1253 4027 1267
rect 4153 1573 4167 1587
rect 4113 1293 4127 1307
rect 4153 1273 4167 1287
rect 4093 1153 4107 1167
rect 4053 1133 4067 1147
rect 4033 1093 4047 1107
rect 4073 1093 4087 1107
rect 4073 1053 4087 1067
rect 4093 813 4107 827
rect 4053 773 4067 787
rect 4033 633 4047 647
rect 3973 593 3987 607
rect 3673 573 3687 587
rect 3873 573 3887 587
rect 3653 373 3667 387
rect 3613 353 3627 367
rect 3933 353 3947 367
rect 3333 333 3347 347
rect 3373 333 3387 347
rect 3593 333 3607 347
rect 3053 313 3067 327
rect 3193 313 3207 327
rect 3213 313 3227 327
rect 3073 213 3087 227
rect 3393 193 3407 207
rect 3373 173 3387 187
rect 3213 153 3227 167
rect 3353 153 3367 167
rect 3573 173 3587 187
rect 3673 333 3687 347
rect 3893 333 3907 347
rect 3873 313 3887 327
rect 4033 313 4047 327
rect 3633 213 3647 227
rect 3813 193 3827 207
rect 3113 133 3127 147
rect 3633 173 3647 187
rect 4393 1733 4407 1747
rect 4413 1733 4427 1747
rect 4353 1613 4367 1627
rect 4653 1773 4667 1787
rect 4633 1753 4647 1767
rect 4653 1753 4667 1767
rect 4533 1713 4547 1727
rect 4373 1573 4387 1587
rect 4333 1333 4347 1347
rect 4273 1293 4287 1307
rect 4633 1633 4647 1647
rect 4573 1593 4587 1607
rect 4613 1353 4627 1367
rect 4573 1333 4587 1347
rect 4793 2273 4807 2287
rect 4893 2533 4907 2547
rect 4873 2273 4887 2287
rect 4813 2253 4827 2267
rect 4853 2253 4867 2267
rect 4773 2233 4787 2247
rect 4913 2233 4927 2247
rect 4833 2013 4847 2027
rect 4753 1773 4767 1787
rect 4893 2033 4907 2047
rect 5093 4673 5107 4687
rect 5093 4613 5107 4627
rect 4733 1733 4747 1747
rect 4693 1593 4707 1607
rect 4833 1593 4847 1607
rect 4673 1553 4687 1567
rect 4753 1553 4767 1567
rect 4853 1553 4867 1567
rect 4893 1733 4907 1747
rect 5013 1773 5027 1787
rect 4913 1593 4927 1607
rect 4973 1553 4987 1567
rect 5073 1753 5087 1767
rect 5033 1353 5047 1367
rect 4873 1333 4887 1347
rect 4833 1313 4847 1327
rect 4653 1293 4667 1307
rect 4873 1293 4887 1307
rect 4293 1273 4307 1287
rect 4593 1273 4607 1287
rect 4813 1273 4827 1287
rect 4893 1273 4907 1287
rect 4333 1153 4347 1167
rect 4573 1153 4587 1167
rect 4293 1133 4307 1147
rect 4353 1093 4367 1107
rect 4533 1093 4547 1107
rect 4253 1073 4267 1087
rect 4313 1073 4327 1087
rect 4333 873 4347 887
rect 4373 853 4387 867
rect 4433 853 4447 867
rect 4353 833 4367 847
rect 4153 813 4167 827
rect 4373 813 4387 827
rect 4133 773 4147 787
rect 4113 673 4127 687
rect 4353 673 4367 687
rect 4113 653 4127 667
rect 4133 633 4147 647
rect 4393 653 4407 667
rect 4613 1073 4627 1087
rect 4633 873 4647 887
rect 4593 853 4607 867
rect 4533 833 4547 847
rect 4613 833 4627 847
rect 4433 613 4447 627
rect 4413 593 4427 607
rect 4393 373 4407 387
rect 4153 353 4167 367
rect 4693 673 4707 687
rect 4733 673 4747 687
rect 4673 653 4687 667
rect 4653 613 4667 627
rect 4713 653 4727 667
rect 4813 633 4827 647
rect 4873 833 4887 847
rect 4933 673 4947 687
rect 4833 573 4847 587
rect 4433 353 4447 367
rect 4633 353 4647 367
rect 4693 353 4707 367
rect 4913 633 4927 647
rect 4073 333 4087 347
rect 4373 333 4387 347
rect 4413 333 4427 347
rect 4653 333 4667 347
rect 4873 333 4887 347
rect 4953 333 4967 347
rect 4153 313 4167 327
rect 4053 173 4067 187
rect 3813 153 3827 167
rect 3573 133 3587 147
rect 3613 133 3627 147
rect 3653 133 3667 147
rect 3133 113 3147 127
rect 3213 113 3227 127
rect 3413 113 3427 127
rect 3913 133 3927 147
rect 4113 133 4127 147
rect 4933 313 4947 327
rect 4393 193 4407 207
rect 4173 173 4187 187
rect 4253 173 4267 187
rect 4873 173 4887 187
rect 4193 133 4207 147
rect 3933 113 3947 127
rect 4653 133 4667 147
rect 4253 113 4267 127
rect 4413 113 4427 127
rect 4633 113 4647 127
rect 4673 113 4687 127
rect 4893 113 4907 127
rect 4973 313 4987 327
rect 3813 13 3827 27
rect 3893 13 3907 27
rect 4873 13 4887 27
rect 4953 13 4967 27
<< metal3 >>
rect 4307 4816 4353 4824
rect 2907 4796 4393 4804
rect 5027 4796 5144 4804
rect 4687 4756 5144 4764
rect 4167 4736 4673 4744
rect 3947 4716 5144 4724
rect 767 4696 1013 4704
rect 1747 4696 2333 4704
rect 2347 4696 2633 4704
rect 3147 4696 3393 4704
rect 3407 4696 3933 4704
rect 4087 4696 4113 4704
rect 4667 4696 4853 4704
rect 447 4676 513 4684
rect 1267 4676 1324 4684
rect 507 4656 953 4664
rect 1316 4664 1324 4676
rect 1347 4676 1533 4684
rect 1767 4676 1793 4684
rect 3387 4676 3573 4684
rect 3587 4676 3613 4684
rect 4947 4676 4993 4684
rect 5107 4676 5144 4684
rect 1007 4656 1304 4664
rect 1316 4656 1433 4664
rect 1296 4647 1304 4656
rect 1787 4656 2293 4664
rect 2307 4656 2573 4664
rect 2807 4656 2833 4664
rect 3656 4664 3664 4673
rect 3656 4656 3904 4664
rect 3896 4647 3904 4656
rect 4327 4656 4393 4664
rect 4867 4656 4893 4664
rect 187 4636 213 4644
rect 247 4636 493 4644
rect 507 4636 533 4644
rect 1447 4636 1513 4644
rect 1527 4636 1753 4644
rect 1767 4636 2033 4644
rect 3187 4636 3333 4644
rect 3347 4636 3553 4644
rect 3567 4636 3873 4644
rect 4407 4636 4433 4644
rect 4607 4636 4853 4644
rect 267 4616 1233 4624
rect 1247 4616 1573 4624
rect 2647 4616 5093 4624
rect 1367 4596 1533 4604
rect 1547 4596 1833 4604
rect 3687 4556 3913 4564
rect -24 4536 33 4544
rect 487 4536 693 4544
rect 3147 4536 3373 4544
rect 2967 4516 3633 4524
rect -24 4496 13 4504
rect 447 4496 513 4504
rect 707 4496 753 4504
rect 1267 4496 1293 4504
rect 1407 4496 1673 4504
rect 1687 4496 1913 4504
rect 2047 4496 2293 4504
rect 2367 4496 2473 4504
rect 2487 4496 2853 4504
rect 2867 4496 3133 4504
rect 3187 4496 3353 4504
rect 4087 4496 4653 4504
rect 927 4476 1213 4484
rect 1236 4476 1513 4484
rect -24 4444 -16 4464
rect 227 4456 273 4464
rect 716 4464 724 4473
rect 1236 4467 1244 4476
rect 1567 4476 1713 4484
rect 1787 4476 1833 4484
rect 1967 4476 2253 4484
rect 2607 4476 2813 4484
rect 3127 4476 3333 4484
rect 3687 4476 3893 4484
rect 4107 4476 4153 4484
rect 4447 4476 4473 4484
rect 467 4456 724 4464
rect 1307 4456 1493 4464
rect 1547 4456 1593 4464
rect 1827 4456 2273 4464
rect 2327 4456 2553 4464
rect 2627 4456 2833 4464
rect 3116 4464 3124 4473
rect 2847 4456 3124 4464
rect 3367 4456 3613 4464
rect 3927 4456 4113 4464
rect 4207 4456 4713 4464
rect 4747 4456 4953 4464
rect -24 4436 173 4444
rect 187 4436 193 4444
rect 1267 4436 1433 4444
rect 3107 4436 3633 4444
rect 4407 4436 4453 4444
rect 4647 4436 4933 4444
rect 647 4416 893 4424
rect 907 4416 1393 4424
rect 4347 4416 4413 4424
rect 2607 4356 3073 4364
rect 227 4336 433 4344
rect 2007 4336 2533 4344
rect 987 4276 1273 4284
rect -24 4216 733 4224
rect -24 4196 -16 4216
rect 747 4216 1193 4224
rect 1567 4216 1773 4224
rect 3587 4216 3633 4224
rect 3847 4216 4093 4224
rect 4107 4216 4133 4224
rect 1227 4196 1293 4204
rect 1427 4196 1513 4204
rect 2067 4196 2293 4204
rect 2307 4196 2773 4204
rect 527 4176 693 4184
rect 707 4176 753 4184
rect 1487 4176 1593 4184
rect 2027 4176 2313 4184
rect 2327 4176 2573 4184
rect 247 4156 273 4164
rect 287 4156 453 4164
rect 807 4156 953 4164
rect 2796 4164 2804 4213
rect 2827 4196 2953 4204
rect 2967 4196 3153 4204
rect 3307 4196 3333 4204
rect 3427 4196 3673 4204
rect 4367 4196 4393 4204
rect 4447 4196 4473 4204
rect 4607 4196 4653 4204
rect 3087 4176 3353 4184
rect 4347 4176 4373 4184
rect 2796 4156 2853 4164
rect 2887 4156 3913 4164
rect 3927 4156 4093 4164
rect 4687 4156 4853 4164
rect 2787 4136 2833 4144
rect 2847 4136 3093 4144
rect 3387 4136 3653 4144
rect 3127 4116 3833 4124
rect 1767 4036 2033 4044
rect 2047 4036 2253 4044
rect 2287 4036 2313 4044
rect 3347 4036 3613 4044
rect 4007 4036 4413 4044
rect 247 4016 333 4024
rect 387 4016 633 4024
rect 747 4016 933 4024
rect 1087 4016 1213 4024
rect 1227 4016 1413 4024
rect 1747 4016 2233 4024
rect 2287 4016 2513 4024
rect 3867 4016 4133 4024
rect 4807 4016 4853 4024
rect 27 3996 213 4004
rect 267 3996 293 4004
rect 427 3996 533 4004
rect 607 3996 1173 4004
rect 1347 3996 1693 4004
rect 2567 3996 2753 4004
rect 3387 3996 3493 4004
rect 3567 3996 3613 4004
rect 3807 3996 3873 4004
rect 3887 3996 3913 4004
rect 4127 3996 4453 4004
rect 216 3984 224 3993
rect 216 3976 233 3984
rect 1207 3976 1493 3984
rect 3127 3976 3173 3984
rect 4356 3976 4633 3984
rect 4356 3967 4364 3976
rect 967 3956 1233 3964
rect 1247 3956 1353 3964
rect 1767 3956 1973 3964
rect 2027 3956 3033 3964
rect 3047 3956 3093 3964
rect 3327 3956 3353 3964
rect 4407 3956 4473 3964
rect 4667 3956 4693 3964
rect 4707 3956 4813 3964
rect 2787 3936 2853 3944
rect 2527 3916 4333 3924
rect 1407 3876 1433 3884
rect 2107 3796 3513 3804
rect 3527 3796 3533 3804
rect 2847 3776 3833 3784
rect 307 3756 1013 3764
rect 3067 3756 3273 3764
rect 447 3736 473 3744
rect 2767 3736 2884 3744
rect 787 3716 853 3724
rect 1567 3716 1673 3724
rect 1687 3716 2244 3724
rect 347 3696 473 3704
rect 547 3696 753 3704
rect 1707 3696 1733 3704
rect 2236 3704 2244 3716
rect 2347 3716 2493 3724
rect 2507 3716 2793 3724
rect 2876 3724 2884 3736
rect 2907 3736 3053 3744
rect 3067 3736 3073 3744
rect 3127 3736 3173 3744
rect 3427 3736 3653 3744
rect 3667 3736 4073 3744
rect 4347 3736 4453 3744
rect 4467 3736 4673 3744
rect 2876 3716 3033 3724
rect 3047 3716 3093 3724
rect 3307 3716 3333 3724
rect 3827 3716 3893 3724
rect 3936 3716 4193 3724
rect 2236 3696 2873 3704
rect 3376 3704 3384 3713
rect 3936 3704 3944 3716
rect 4447 3716 4473 3724
rect 4987 3716 5144 3724
rect 2887 3696 3944 3704
rect 3967 3696 4173 3704
rect 4907 3696 4953 3704
rect 227 3676 513 3684
rect 807 3676 1033 3684
rect 1267 3676 1293 3684
rect 1327 3676 1933 3684
rect 2587 3676 2753 3684
rect 2927 3676 3393 3684
rect 3407 3676 3553 3684
rect 3647 3676 3913 3684
rect 3947 3676 4393 3684
rect 4407 3676 4713 3684
rect 4727 3676 4913 3684
rect 767 3656 833 3664
rect 1467 3656 1653 3664
rect 1667 3656 1853 3664
rect 2387 3656 4973 3664
rect 1487 3636 1713 3644
rect 2327 3636 2553 3644
rect 2607 3636 2613 3644
rect 2627 3636 2853 3644
rect 2507 3556 2533 3564
rect 267 3536 453 3544
rect 467 3536 493 3544
rect 787 3536 1033 3544
rect 2107 3536 2313 3544
rect 2487 3536 2553 3544
rect 3587 3536 3873 3544
rect 4427 3536 4613 3544
rect 4627 3536 4733 3544
rect 4807 3536 4893 3544
rect 4907 3536 4913 3544
rect 247 3516 433 3524
rect 447 3516 713 3524
rect 1267 3516 1513 3524
rect 1787 3516 1813 3524
rect 1867 3516 2293 3524
rect 2347 3516 2373 3524
rect 2607 3516 2813 3524
rect 2847 3516 3173 3524
rect 3347 3516 3373 3524
rect 3427 3516 3453 3524
rect 3507 3516 3533 3524
rect 3547 3516 4013 3524
rect 4027 3516 4033 3524
rect 487 3496 533 3504
rect 1727 3496 1793 3504
rect 2087 3496 2493 3504
rect 2507 3496 2533 3504
rect 2587 3496 2613 3504
rect 3127 3496 3253 3504
rect 3307 3496 3353 3504
rect 3367 3496 3773 3504
rect 3907 3496 4313 3504
rect 467 3476 733 3484
rect 1547 3476 2113 3484
rect 2827 3476 2853 3484
rect 2867 3476 3093 3484
rect 3407 3476 3593 3484
rect 3787 3476 3873 3484
rect 3927 3476 3953 3484
rect 3967 3476 4333 3484
rect 4367 3476 4413 3484
rect 3067 3456 3133 3464
rect 3547 3456 4293 3464
rect 4407 3416 4753 3424
rect 1087 3376 1833 3384
rect 1847 3376 1913 3384
rect 507 3276 553 3284
rect 1967 3276 2073 3284
rect 2267 3276 2853 3284
rect 2867 3276 3393 3284
rect 4327 3276 4373 3284
rect 4907 3276 4933 3284
rect 47 3256 213 3264
rect 527 3256 713 3264
rect 1727 3256 2033 3264
rect 3267 3256 3873 3264
rect 3947 3256 4693 3264
rect 4887 3256 5004 3264
rect 4996 3247 5004 3256
rect 187 3236 773 3244
rect 787 3236 993 3244
rect 1007 3236 1024 3244
rect 1016 3227 1024 3236
rect 1687 3236 1833 3244
rect 1847 3236 1853 3244
rect 3107 3236 3153 3244
rect 3167 3236 3313 3244
rect 4347 3236 4413 3244
rect 4587 3236 4653 3244
rect 4867 3236 4953 3244
rect 267 3216 513 3224
rect 676 3216 733 3224
rect 507 3196 533 3204
rect 676 3204 684 3216
rect 1427 3216 1773 3224
rect 2887 3216 2913 3224
rect 3387 3216 3553 3224
rect 3687 3216 3953 3224
rect 4107 3216 4393 3224
rect 4447 3216 4713 3224
rect 4747 3216 4893 3224
rect 4907 3216 4933 3224
rect 547 3196 684 3204
rect 727 3196 793 3204
rect 807 3196 1053 3204
rect 1307 3196 1713 3204
rect 1827 3196 1913 3204
rect 2267 3196 2553 3204
rect 3087 3196 3413 3204
rect 4647 3196 4673 3204
rect 4767 3196 4973 3204
rect 1567 3176 1633 3184
rect 3347 3176 3413 3184
rect 3427 3176 3933 3184
rect 4087 3176 4153 3184
rect 2327 3156 2573 3164
rect 2587 3156 3813 3164
rect 767 3076 793 3084
rect 2227 3076 2533 3084
rect 2587 3076 3113 3084
rect 3907 3076 3973 3084
rect 4027 3076 4193 3084
rect 4867 3076 4993 3084
rect 227 3056 473 3064
rect 487 3056 493 3064
rect 507 3056 833 3064
rect 887 3056 1013 3064
rect 2187 3056 2373 3064
rect 2887 3056 3093 3064
rect 3147 3056 3633 3064
rect 3927 3056 4133 3064
rect 4267 3056 4473 3064
rect 4487 3056 4713 3064
rect 4767 3056 4973 3064
rect 207 3036 253 3044
rect 527 3036 973 3044
rect 736 3027 744 3036
rect 1467 3036 2073 3044
rect 2087 3036 2093 3044
rect 2107 3036 2213 3044
rect 2467 3036 2853 3044
rect 3287 3036 3333 3044
rect 3687 3036 3953 3044
rect 4547 3036 4693 3044
rect 4707 3036 4913 3044
rect 487 3016 693 3024
rect 847 3016 993 3024
rect 1287 3016 1313 3024
rect 1427 3016 1453 3024
rect 2407 3016 2513 3024
rect 2827 3016 3613 3024
rect 3627 3016 3773 3024
rect 3787 3016 3893 3024
rect 3947 3016 4013 3024
rect 4147 3016 4173 3024
rect 4227 3016 4433 3024
rect 4907 3016 4953 3024
rect 3407 2996 3653 3004
rect 4467 2996 4753 3004
rect 3647 2976 3793 2984
rect 707 2796 773 2804
rect 747 2776 873 2784
rect 1487 2776 1673 2784
rect 1687 2776 1953 2784
rect 2007 2776 2453 2784
rect 3767 2776 4033 2784
rect 4307 2776 4413 2784
rect 227 2756 253 2764
rect 327 2756 473 2764
rect 527 2756 753 2764
rect 2187 2756 2693 2764
rect 2847 2756 2953 2764
rect 3247 2756 3553 2764
rect 4287 2756 4393 2764
rect 4427 2756 4493 2764
rect 4747 2756 4813 2764
rect 107 2736 453 2744
rect 2127 2736 2373 2744
rect 2396 2736 2973 2744
rect 507 2716 573 2724
rect 587 2716 973 2724
rect 1236 2724 1244 2733
rect 1236 2716 1453 2724
rect 2396 2724 2404 2736
rect 3267 2736 3293 2744
rect 3307 2736 3473 2744
rect 3487 2736 3713 2744
rect 4027 2736 4073 2744
rect 4087 2736 4753 2744
rect 2347 2716 2404 2724
rect 2487 2716 2673 2724
rect 2947 2716 3393 2724
rect 4487 2716 4513 2724
rect 4707 2716 4793 2724
rect 227 2696 313 2704
rect 1027 2696 2113 2704
rect 2167 2656 2293 2664
rect 3347 2656 3493 2664
rect 1127 2636 1273 2644
rect 1747 2636 1833 2644
rect 1847 2636 2013 2644
rect 2027 2636 2033 2644
rect 1547 2616 1793 2624
rect 867 2596 1013 2604
rect 1027 2596 1253 2604
rect 1267 2596 2313 2604
rect 3527 2596 3673 2604
rect 3687 2596 3693 2604
rect 3707 2596 3973 2604
rect 1367 2576 1733 2584
rect 3727 2576 3913 2584
rect 3927 2576 4133 2584
rect 4487 2576 4653 2584
rect 787 2556 813 2564
rect 1307 2556 1693 2564
rect 1787 2556 1993 2564
rect 2036 2556 2073 2564
rect 2036 2547 2044 2556
rect 2287 2556 2333 2564
rect 2427 2556 2513 2564
rect 2567 2556 2673 2564
rect 2687 2556 2813 2564
rect 2987 2556 3073 2564
rect 3127 2556 3153 2564
rect 4407 2556 4853 2564
rect 507 2536 1093 2544
rect 1707 2536 1753 2544
rect 1867 2536 2013 2544
rect 2827 2536 3053 2544
rect 3227 2536 3353 2544
rect 3567 2536 3613 2544
rect 3667 2536 4053 2544
rect 4167 2536 4353 2544
rect 4747 2536 4893 2544
rect 527 2516 693 2524
rect 707 2516 753 2524
rect 1567 2516 1693 2524
rect 2007 2516 2793 2524
rect 3947 2516 4433 2524
rect 487 2496 553 2504
rect 2347 2496 2833 2504
rect 2847 2496 3093 2504
rect 3327 2496 3413 2504
rect 3427 2496 3953 2504
rect 247 2476 573 2484
rect -24 2336 13 2344
rect 987 2336 1033 2344
rect 1587 2336 1973 2344
rect 207 2316 1313 2324
rect 1327 2316 1953 2324
rect 4527 2316 4733 2324
rect -24 2296 193 2304
rect 1327 2296 1673 2304
rect 1907 2296 1993 2304
rect 4367 2296 4553 2304
rect 507 2276 573 2284
rect 587 2276 713 2284
rect 1087 2276 1213 2284
rect 1367 2276 1573 2284
rect 1647 2276 1733 2284
rect 1927 2276 2033 2284
rect 2947 2276 3033 2284
rect 3407 2276 3933 2284
rect 3947 2276 3993 2284
rect 4487 2276 4533 2284
rect 4807 2276 4873 2284
rect 367 2256 773 2264
rect 787 2256 953 2264
rect 967 2256 1153 2264
rect 1227 2256 1293 2264
rect 1347 2256 1513 2264
rect 1876 2264 1884 2273
rect 1627 2256 1884 2264
rect 1907 2256 2133 2264
rect 2207 2256 2333 2264
rect 2367 2256 2653 2264
rect 3216 2264 3224 2273
rect 2967 2256 3224 2264
rect 3247 2256 3473 2264
rect 3536 2256 3573 2264
rect 887 2236 1053 2244
rect 2507 2236 2573 2244
rect 2587 2236 2713 2244
rect 2727 2236 2993 2244
rect 3536 2244 3544 2256
rect 4036 2264 4044 2273
rect 4036 2256 4313 2264
rect 4327 2256 4633 2264
rect 4827 2256 4853 2264
rect 3207 2236 3544 2244
rect 4067 2236 4273 2244
rect 4287 2236 4773 2244
rect 4787 2236 4913 2244
rect 187 2216 613 2224
rect 627 2216 973 2224
rect 987 2216 1313 2224
rect 1327 2216 1513 2224
rect 2067 2176 2213 2184
rect 2227 2176 2253 2184
rect 27 2136 1013 2144
rect 1027 2136 1233 2144
rect 1247 2136 2413 2144
rect 747 2116 1233 2124
rect 2007 2116 3273 2124
rect 147 2096 353 2104
rect 1287 2096 1353 2104
rect 1667 2096 1753 2104
rect 4167 2096 4293 2104
rect 4307 2096 4353 2104
rect 407 2076 693 2084
rect 1347 2076 1533 2084
rect 1907 2076 1993 2084
rect 2047 2076 2073 2084
rect 2547 2076 2824 2084
rect 2816 2067 2824 2076
rect 2847 2076 3193 2084
rect 3627 2076 3913 2084
rect 287 2056 553 2064
rect 607 2056 713 2064
rect 1227 2056 1293 2064
rect 1367 2056 1553 2064
rect 1567 2056 1713 2064
rect 1727 2056 2073 2064
rect 2207 2056 2273 2064
rect 4287 2056 4373 2064
rect 1267 2036 1333 2044
rect 2167 2036 2513 2044
rect 2556 2044 2564 2053
rect 2547 2036 2564 2044
rect 2776 2044 2784 2053
rect 2776 2036 2793 2044
rect 3847 2036 3913 2044
rect 4107 2036 4333 2044
rect 4656 2044 4664 2073
rect 4656 2036 4893 2044
rect 4907 2036 5144 2044
rect 1607 2016 3433 2024
rect 3447 2016 3613 2024
rect 3627 2016 4593 2024
rect 4607 2016 4833 2024
rect 3587 1996 3873 2004
rect 227 1956 293 1964
rect 287 1856 313 1864
rect 967 1836 1433 1844
rect 2087 1836 2393 1844
rect 2927 1836 2993 1844
rect 247 1816 304 1824
rect 296 1804 304 1816
rect 507 1816 1213 1824
rect 1227 1816 1253 1824
rect 2387 1816 2613 1824
rect 2627 1816 2853 1824
rect 3367 1816 3533 1824
rect 4027 1816 4073 1824
rect 296 1796 504 1804
rect 127 1776 213 1784
rect 276 1744 284 1793
rect 307 1776 473 1784
rect 496 1784 504 1796
rect 547 1796 613 1804
rect 2547 1796 2593 1804
rect 3967 1796 4253 1804
rect 4267 1796 4373 1804
rect 496 1776 513 1784
rect 927 1776 1013 1784
rect 1027 1776 1233 1784
rect 1547 1776 1653 1784
rect 1796 1784 1804 1793
rect 1796 1776 2053 1784
rect 2336 1767 2344 1793
rect 3047 1776 3333 1784
rect 3687 1776 3713 1784
rect 4667 1776 4753 1784
rect 4767 1776 5013 1784
rect 507 1756 753 1764
rect 807 1756 1713 1764
rect 1727 1756 1773 1764
rect 2367 1756 2393 1764
rect 3207 1756 3393 1764
rect 3567 1756 3813 1764
rect 4647 1756 4653 1764
rect 4667 1756 5073 1764
rect 276 1736 773 1744
rect 907 1736 1233 1744
rect 1427 1736 1813 1744
rect 3067 1736 3193 1744
rect 3527 1736 3653 1744
rect 3667 1736 3753 1744
rect 4407 1736 4413 1744
rect 4427 1736 4733 1744
rect 4747 1736 4893 1744
rect 1547 1716 3293 1724
rect 3887 1716 4533 1724
rect 2107 1696 3713 1704
rect 3267 1676 3293 1684
rect 3907 1676 4093 1684
rect 3807 1656 4093 1664
rect 1227 1636 1273 1644
rect 2587 1636 2873 1644
rect 3667 1636 4633 1644
rect 2327 1616 2433 1624
rect 2487 1616 2973 1624
rect 2987 1616 2993 1624
rect 3007 1616 3513 1624
rect 3707 1616 3853 1624
rect 4147 1616 4353 1624
rect 447 1596 473 1604
rect 527 1596 533 1604
rect 547 1596 933 1604
rect 1256 1587 1264 1613
rect 1467 1596 1493 1604
rect 2747 1596 2933 1604
rect 3567 1596 3844 1604
rect 3836 1587 3844 1596
rect 4587 1596 4693 1604
rect 4847 1596 4913 1604
rect 787 1576 973 1584
rect 1967 1576 2173 1584
rect 2307 1576 2313 1584
rect 2327 1576 2453 1584
rect 4167 1576 4373 1584
rect 267 1556 533 1564
rect 1007 1556 1093 1564
rect 2347 1556 2453 1564
rect 2707 1556 2813 1564
rect 3067 1556 3273 1564
rect 3327 1556 3393 1564
rect 4687 1556 4753 1564
rect 4867 1556 4973 1564
rect 4987 1556 5144 1564
rect 227 1536 433 1544
rect 2787 1536 3313 1544
rect 687 1376 713 1384
rect 787 1376 813 1384
rect 827 1376 1513 1384
rect 807 1356 953 1364
rect 967 1356 973 1364
rect 1487 1356 1533 1364
rect 4627 1356 5033 1364
rect 947 1336 1013 1344
rect 1347 1336 1513 1344
rect 1687 1336 1773 1344
rect 2507 1336 3653 1344
rect 3667 1336 3793 1344
rect 4347 1336 4573 1344
rect 667 1316 713 1324
rect 1467 1316 1493 1324
rect 3207 1316 3313 1324
rect 3527 1316 3553 1324
rect 3607 1316 3693 1324
rect 3727 1316 4833 1324
rect 247 1296 273 1304
rect 287 1296 313 1304
rect 687 1296 733 1304
rect 1007 1296 1233 1304
rect 1307 1296 1753 1304
rect 2267 1296 2413 1304
rect 2427 1296 2513 1304
rect 3107 1296 3273 1304
rect 3716 1304 3724 1313
rect 4876 1307 4884 1333
rect 3627 1296 3724 1304
rect 4036 1296 4113 1304
rect 227 1276 493 1284
rect 507 1276 653 1284
rect 967 1276 1273 1284
rect 2067 1276 2113 1284
rect 2127 1276 2773 1284
rect 4036 1284 4044 1296
rect 4287 1296 4653 1304
rect 3587 1276 4044 1284
rect 4067 1276 4153 1284
rect 4167 1276 4293 1284
rect 4607 1276 4813 1284
rect 4827 1276 4893 1284
rect 227 1256 453 1264
rect 467 1256 693 1264
rect 2047 1256 2293 1264
rect 2307 1256 3513 1264
rect 3787 1256 4013 1264
rect 447 1236 493 1244
rect 1067 1196 3353 1204
rect 3367 1196 3633 1204
rect 1807 1176 3173 1184
rect 3187 1176 3213 1184
rect 3227 1176 3733 1184
rect 547 1156 753 1164
rect 767 1156 793 1164
rect 827 1156 1333 1164
rect 2447 1156 2553 1164
rect 2767 1156 3073 1164
rect 4107 1156 4333 1164
rect 4347 1156 4573 1164
rect 487 1136 533 1144
rect 587 1136 1093 1144
rect 1107 1136 1293 1144
rect 1387 1136 1593 1144
rect 1607 1136 1733 1144
rect 1907 1136 2153 1144
rect 2547 1136 2973 1144
rect 4067 1136 4293 1144
rect 1947 1116 2013 1124
rect 2027 1116 2173 1124
rect 2207 1116 2333 1124
rect 2347 1116 2484 1124
rect 2476 1107 2484 1116
rect 2527 1116 2713 1124
rect 3027 1116 3133 1124
rect 3156 1116 3493 1124
rect 467 1096 513 1104
rect 1127 1096 1253 1104
rect 2487 1096 2533 1104
rect 3156 1104 3164 1116
rect 3767 1116 4044 1124
rect 4036 1107 4044 1116
rect 3007 1096 3164 1104
rect 3527 1096 3533 1104
rect 3547 1096 3733 1104
rect 4087 1096 4344 1104
rect 167 1076 193 1084
rect 207 1076 233 1084
rect 807 1076 933 1084
rect 2967 1076 3193 1084
rect 3487 1076 4253 1084
rect 4267 1076 4313 1084
rect 4336 1084 4344 1096
rect 4367 1096 4533 1104
rect 4336 1076 4613 1084
rect 3927 1056 4073 1064
rect 847 876 1353 884
rect 2487 876 2513 884
rect 2847 876 3593 884
rect 3607 876 3693 884
rect 3707 876 3773 884
rect 4347 876 4633 884
rect 1327 856 1493 864
rect 1707 856 1793 864
rect 1807 856 1913 864
rect 3067 856 3273 864
rect 4387 856 4433 864
rect 4607 856 4644 864
rect 487 836 693 844
rect 1007 836 1233 844
rect 1467 836 1533 844
rect 2427 836 2493 844
rect 2827 836 3033 844
rect 3807 836 3833 844
rect 3887 836 4353 844
rect 4547 836 4613 844
rect 4636 844 4644 856
rect 4636 836 4873 844
rect 267 816 673 824
rect 727 816 833 824
rect 956 807 964 833
rect 987 816 1073 824
rect 1527 816 1573 824
rect 1647 816 1753 824
rect 2027 816 2233 824
rect 2247 816 2693 824
rect 2776 824 2784 833
rect 2776 816 3113 824
rect 3447 816 3613 824
rect 3627 816 3673 824
rect 3787 816 3864 824
rect 3856 807 3864 816
rect 4107 816 4153 824
rect 4167 816 4373 824
rect 467 796 493 804
rect 1267 796 1313 804
rect 1367 796 1473 804
rect 1547 796 1773 804
rect 2187 796 2273 804
rect 2807 796 2833 804
rect 3587 796 3793 804
rect 247 776 793 784
rect 2567 776 2873 784
rect 3007 776 3613 784
rect 4067 776 4133 784
rect 1907 756 2833 764
rect 2427 736 3093 744
rect 3227 716 3273 724
rect 3287 716 3793 724
rect 1507 676 1993 684
rect 2007 676 2233 684
rect 2267 676 2813 684
rect 4127 676 4353 684
rect 4367 676 4693 684
rect 4707 676 4733 684
rect 4747 676 4933 684
rect 207 656 713 664
rect 476 627 484 656
rect 1467 656 1784 664
rect 507 636 933 644
rect 1007 636 1633 644
rect 1776 627 1784 656
rect 1807 656 1973 664
rect 1987 656 2013 664
rect 2027 656 2273 664
rect 2327 656 2553 664
rect 2767 656 3313 664
rect 4127 656 4393 664
rect 4687 656 4713 664
rect 1827 636 2593 644
rect 2807 636 2853 644
rect 3167 636 3193 644
rect 3767 636 3813 644
rect 4047 636 4133 644
rect 4827 636 4913 644
rect 1247 616 1433 624
rect 1487 616 1733 624
rect 447 596 473 604
rect 987 596 1193 604
rect 1796 604 1804 633
rect 2307 616 2333 624
rect 2587 616 2613 624
rect 4447 616 4653 624
rect 1787 596 1804 604
rect 2067 596 2533 604
rect 3387 596 3633 604
rect 3647 596 3653 604
rect 3987 596 4413 604
rect 2547 576 3073 584
rect 3087 576 3133 584
rect 3687 576 3873 584
rect 3887 576 4833 584
rect 1027 496 1053 504
rect 1067 496 1533 504
rect 976 384 984 393
rect 707 376 1013 384
rect 1347 376 1553 384
rect 1567 376 1933 384
rect 1956 376 1993 384
rect 1027 356 1253 364
rect 1307 356 1533 364
rect 1956 364 1964 376
rect 2827 376 2933 384
rect 3127 376 3353 384
rect 3667 376 4393 384
rect 1547 356 1964 364
rect 1987 356 2013 364
rect 2187 356 2253 364
rect 2267 356 2533 364
rect 2556 356 2613 364
rect 2556 347 2564 356
rect 3396 364 3404 373
rect 2847 356 3613 364
rect 3947 356 4144 364
rect 1047 336 1053 344
rect 1067 336 1233 344
rect 1287 336 1313 344
rect 2307 336 2413 344
rect 2587 336 2793 344
rect 2947 336 2993 344
rect 3007 336 3073 344
rect 3347 336 3373 344
rect 3387 336 3593 344
rect 3607 336 3673 344
rect 3687 336 3893 344
rect 3907 336 4073 344
rect 4136 344 4144 356
rect 4167 356 4433 364
rect 4647 356 4693 364
rect 4136 336 4373 344
rect 4427 336 4653 344
rect 4887 336 4953 344
rect 247 316 453 324
rect 467 316 673 324
rect 1327 316 2053 324
rect 2887 316 3053 324
rect 3067 316 3193 324
rect 3227 316 3873 324
rect 3887 316 4033 324
rect 4047 316 4153 324
rect 4947 316 4973 324
rect 287 296 753 304
rect 767 296 913 304
rect 1247 296 1753 304
rect 1947 296 2513 304
rect 787 276 993 284
rect 1487 216 1813 224
rect 2847 216 3073 224
rect 3087 216 3633 224
rect 547 196 973 204
rect 987 196 1233 204
rect 1807 196 2233 204
rect 2247 196 2533 204
rect 2547 196 3393 204
rect 3827 196 4393 204
rect 807 176 993 184
rect 1247 176 1333 184
rect 1447 176 1693 184
rect 2067 176 2093 184
rect 2127 176 2293 184
rect 2327 176 2853 184
rect 3387 176 3573 184
rect 3647 176 4053 184
rect 4067 176 4173 184
rect 4267 176 4873 184
rect 487 156 753 164
rect 827 156 1013 164
rect 1027 156 1253 164
rect 1267 156 1493 164
rect 1667 156 2013 164
rect 2036 156 2253 164
rect 2036 147 2044 156
rect 2287 156 2333 164
rect 2427 156 2593 164
rect 2887 156 3213 164
rect 3367 156 3813 164
rect 247 136 1033 144
rect 2087 136 2113 144
rect 2347 136 2553 144
rect 2576 136 3113 144
rect 507 116 813 124
rect 2576 124 2584 136
rect 3587 136 3613 144
rect 3667 136 3913 144
rect 3927 136 4113 144
rect 4207 136 4653 144
rect 2107 116 2584 124
rect 3147 116 3213 124
rect 3427 116 3933 124
rect 3947 116 4253 124
rect 4427 116 4633 124
rect 4687 116 4893 124
rect 227 96 733 104
rect 3827 16 3893 24
rect 4887 16 4953 24
use OAI21X1  _313_
timestamp 0
transform 1 0 1230 0 1 250
box -6 -8 106 248
use INVX1  _314_
timestamp 0
transform -1 0 1270 0 1 730
box -6 -8 66 248
use OAI21X1  _315_
timestamp 0
transform 1 0 930 0 1 730
box -6 -8 106 248
use AOI21X1  _316_
timestamp 0
transform -1 0 1130 0 -1 1210
box -6 -8 106 248
use NAND2X1  _317_
timestamp 0
transform -1 0 2870 0 1 250
box -6 -8 86 248
use OR2X2  _318_
timestamp 0
transform 1 0 3050 0 1 250
box -6 -8 106 248
use NAND2X1  _319_
timestamp 0
transform -1 0 3410 0 1 250
box -6 -8 86 248
use OR2X2  _320_
timestamp 0
transform -1 0 3350 0 1 730
box -6 -8 106 248
use NAND2X1  _321_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 86 248
use NAND2X1  _322_
timestamp 0
transform 1 0 3010 0 1 730
box -6 -8 86 248
use OAI21X1  _323_
timestamp 0
transform -1 0 3170 0 -1 730
box -6 -8 106 248
use AOI21X1  _324_
timestamp 0
transform -1 0 2830 0 1 730
box -6 -8 106 248
use OAI21X1  _325_
timestamp 0
transform -1 0 3690 0 1 250
box -6 -8 106 248
use NAND2X1  _326_
timestamp 0
transform -1 0 3950 0 -1 250
box -6 -8 86 248
use INVX1  _327_
timestamp 0
transform 1 0 4870 0 -1 250
box -6 -8 66 248
use INVX1  _328_
timestamp 0
transform 1 0 4390 0 -1 250
box -6 -8 66 248
use NAND2X1  _329_
timestamp 0
transform -1 0 4690 0 -1 250
box -6 -8 86 248
use NAND2X1  _330_
timestamp 0
transform 1 0 4130 0 -1 250
box -6 -8 86 248
use NAND2X1  _331_
timestamp 0
transform -1 0 3150 0 -1 250
box -6 -8 86 248
use NOR2X1  _332_
timestamp 0
transform -1 0 2890 0 -1 250
box -6 -8 86 248
use NOR2X1  _333_
timestamp 0
transform 1 0 2270 0 -1 250
box -6 -8 86 248
use OAI21X1  _334_
timestamp 0
transform 1 0 2230 0 1 250
box -6 -8 106 248
use AOI21X1  _335_
timestamp 0
transform -1 0 2090 0 -1 250
box -6 -8 106 248
use NOR2X1  _336_
timestamp 0
transform -1 0 3410 0 -1 250
box -6 -8 86 248
use OAI21X1  _337_
timestamp 0
transform 1 0 3590 0 -1 250
box -6 -8 106 248
use INVX1  _338_
timestamp 0
transform -1 0 4190 0 1 250
box -6 -8 66 248
use OR2X2  _339_
timestamp 0
transform 1 0 3870 0 1 250
box -6 -8 106 248
use OAI21X1  _340_
timestamp 0
transform 1 0 4370 0 1 250
box -6 -8 106 248
use AND2X2  _341_
timestamp 0
transform 1 0 4830 0 -1 1210
box -6 -8 106 248
use NOR2X1  _342_
timestamp 0
transform 1 0 4910 0 1 250
box -6 -8 86 248
use NOR2X1  _343_
timestamp 0
transform -1 0 4970 0 -1 730
box -6 -8 86 248
use NAND2X1  _344_
timestamp 0
transform -1 0 4730 0 1 250
box -6 -8 86 248
use OR2X2  _345_
timestamp 0
transform -1 0 4730 0 -1 730
box -6 -8 106 248
use NAND2X1  _346_
timestamp 0
transform 1 0 4330 0 1 730
box -6 -8 86 248
use OAI21X1  _347_
timestamp 0
transform -1 0 3630 0 1 730
box -6 -8 106 248
use AOI21X1  _348_
timestamp 0
transform -1 0 3890 0 1 730
box -6 -8 106 248
use NAND2X1  _349_
timestamp 0
transform 1 0 4850 0 1 730
box -6 -8 86 248
use NAND2X1  _350_
timestamp 0
transform 1 0 4590 0 1 730
box -6 -8 86 248
use AND2X2  _351_
timestamp 0
transform 1 0 4630 0 -1 1690
box -6 -8 106 248
use NOR2X1  _352_
timestamp 0
transform 1 0 4610 0 1 1690
box -6 -8 86 248
use NOR2X1  _353_
timestamp 0
transform 1 0 4270 0 1 1210
box -6 -8 86 248
use INVX1  _354_
timestamp 0
transform 1 0 4050 0 1 1210
box -6 -8 66 248
use OR2X2  _355_
timestamp 0
transform 1 0 4550 0 -1 1210
box -6 -8 106 248
use AOI21X1  _356_
timestamp 0
transform -1 0 4370 0 -1 1210
box -6 -8 106 248
use OAI21X1  _357_
timestamp 0
transform -1 0 3810 0 -1 1210
box -6 -8 106 248
use AOI21X1  _358_
timestamp 0
transform -1 0 4090 0 -1 1210
box -6 -8 106 248
use NAND2X1  _359_
timestamp 0
transform -1 0 3670 0 1 3610
box -6 -8 86 248
use NOR2X1  _360_
timestamp 0
transform 1 0 4090 0 -1 730
box -6 -8 86 248
use NAND3X1  _361_
timestamp 0
transform 1 0 4350 0 -1 730
box -6 -8 106 248
use NAND3X1  _362_
timestamp 0
transform -1 0 4150 0 1 730
box -6 -8 106 248
use INVX1  _363_
timestamp 0
transform -1 0 5090 0 1 2170
box -6 -8 66 248
use AOI21X1  _364_
timestamp 0
transform -1 0 4630 0 1 1210
box -6 -8 106 248
use AND2X2  _365_
timestamp 0
transform -1 0 3630 0 -1 2170
box -6 -8 106 248
use OAI21X1  _366_
timestamp 0
transform -1 0 3690 0 -1 2650
box -6 -8 106 248
use NAND2X1  _367_
timestamp 0
transform 1 0 4110 0 1 4570
box -6 -8 86 248
use OR2X2  _368_
timestamp 0
transform 1 0 4650 0 -1 4570
box -6 -8 106 248
use NAND2X1  _369_
timestamp 0
transform 1 0 4130 0 -1 4570
box -6 -8 86 248
use NOR2X1  _370_
timestamp 0
transform 1 0 3830 0 -1 4090
box -6 -8 86 248
use AND2X2  _371_
timestamp 0
transform 1 0 4090 0 1 4090
box -6 -8 106 248
use OAI21X1  _372_
timestamp 0
transform 1 0 4130 0 1 3610
box -6 -8 106 248
use AOI21X1  _373_
timestamp 0
transform -1 0 3950 0 1 3610
box -6 -8 106 248
use INVX1  _374_
timestamp 0
transform -1 0 3930 0 1 4090
box -6 -8 66 248
use OAI21X1  _375_
timestamp 0
transform 1 0 3850 0 -1 4570
box -6 -8 106 248
use NAND2X1  _376_
timestamp 0
transform 1 0 3350 0 1 4570
box -6 -8 86 248
use OR2X2  _377_
timestamp 0
transform -1 0 3190 0 1 4570
box -6 -8 106 248
use NAND2X1  _378_
timestamp 0
transform 1 0 3590 0 -1 4570
box -6 -8 86 248
use OR2X2  _379_
timestamp 0
transform -1 0 3410 0 1 4090
box -6 -8 106 248
use AOI21X1  _380_
timestamp 0
transform -1 0 3690 0 1 4090
box -6 -8 106 248
use OAI21X1  _381_
timestamp 0
transform -1 0 3410 0 1 3610
box -6 -8 106 248
use AOI21X1  _382_
timestamp 0
transform 1 0 3310 0 -1 4090
box -6 -8 106 248
use NOR2X1  _383_
timestamp 0
transform -1 0 3130 0 1 4090
box -6 -8 86 248
use NOR2X1  _384_
timestamp 0
transform 1 0 3870 0 1 4570
box -6 -8 86 248
use OAI21X1  _385_
timestamp 0
transform -1 0 3690 0 1 4570
box -6 -8 106 248
use AOI21X1  _386_
timestamp 0
transform -1 0 2870 0 1 4090
box -6 -8 106 248
use AND2X2  _387_
timestamp 0
transform 1 0 2290 0 1 4570
box -6 -8 106 248
use NOR2X1  _388_
timestamp 0
transform 1 0 2570 0 1 4570
box -6 -8 86 248
use OR2X2  _389_
timestamp 0
transform -1 0 3150 0 -1 4570
box -6 -8 106 248
use OR2X2  _390_
timestamp 0
transform -1 0 2050 0 1 4090
box -6 -8 106 248
use OAI21X1  _391_
timestamp 0
transform -1 0 2870 0 -1 4570
box -6 -8 106 248
use NAND2X1  _392_
timestamp 0
transform -1 0 2590 0 -1 4570
box -6 -8 86 248
use OAI21X1  _393_
timestamp 0
transform 1 0 1770 0 1 4570
box -6 -8 106 248
use AOI21X1  _394_
timestamp 0
transform -1 0 2330 0 -1 4570
box -6 -8 106 248
use NAND2X1  _395_
timestamp 0
transform -1 0 1790 0 1 4090
box -6 -8 86 248
use NAND2X1  _396_
timestamp 0
transform 1 0 2310 0 1 3610
box -6 -8 86 248
use INVX1  _397_
timestamp 0
transform 1 0 2810 0 1 3610
box -6 -8 66 248
use NOR2X1  _398_
timestamp 0
transform 1 0 2290 0 -1 3610
box -6 -8 86 248
use NOR2X1  _399_
timestamp 0
transform 1 0 2550 0 1 3610
box -6 -8 86 248
use NAND3X1  _400_
timestamp 0
transform -1 0 2050 0 -1 4090
box -6 -8 106 248
use OAI21X1  _401_
timestamp 0
transform -1 0 2330 0 1 4090
box -6 -8 106 248
use INVX1  _402_
timestamp 0
transform -1 0 2110 0 -1 3610
box -6 -8 66 248
use NAND2X1  _403_
timestamp 0
transform 1 0 2490 0 -1 4090
box -6 -8 86 248
use AOI21X1  _404_
timestamp 0
transform -1 0 2310 0 -1 4090
box -6 -8 106 248
use OAI21X1  _405_
timestamp 0
transform 1 0 1650 0 1 3610
box -6 -8 106 248
use AOI21X1  _406_
timestamp 0
transform -1 0 1770 0 -1 4090
box -6 -8 106 248
use NOR2X1  _407_
timestamp 0
transform 1 0 3330 0 -1 4570
box -6 -8 86 248
use NAND3X1  _408_
timestamp 0
transform -1 0 3130 0 -1 4090
box -6 -8 106 248
use OR2X2  _409_
timestamp 0
transform 1 0 3690 0 1 2650
box -6 -8 106 248
use NAND2X1  _410_
timestamp 0
transform -1 0 3890 0 -1 2170
box -6 -8 86 248
use NOR2X1  _411_
timestamp 0
transform -1 0 2590 0 1 4090
box -6 -8 86 248
use AND2X2  _412_
timestamp 0
transform 1 0 2750 0 -1 4090
box -6 -8 106 248
use NAND3X1  _413_
timestamp 0
transform -1 0 3150 0 1 3610
box -6 -8 106 248
use AOI21X1  _414_
timestamp 0
transform 1 0 2530 0 -1 3610
box -6 -8 106 248
use NAND2X1  _415_
timestamp 0
transform 1 0 3090 0 -1 3610
box -6 -8 86 248
use AOI21X1  _416_
timestamp 0
transform 1 0 3830 0 1 3130
box -6 -8 106 248
use OAI21X1  _417_
timestamp 0
transform -1 0 4070 0 1 2650
box -6 -8 106 248
use AND2X2  _418_
timestamp 0
transform 1 0 4850 0 -1 2170
box -6 -8 106 248
use NOR2X1  _419_
timestamp 0
transform 1 0 4610 0 -1 2170
box -6 -8 86 248
use NOR2X1  _420_
timestamp 0
transform -1 0 4330 0 1 2170
box -6 -8 86 248
use NAND2X1  _421_
timestamp 0
transform -1 0 4150 0 -1 2170
box -6 -8 86 248
use NOR2X1  _422_
timestamp 0
transform -1 0 1810 0 1 730
box -6 -8 86 248
use NAND2X1  _423_
timestamp 0
transform 1 0 1470 0 1 1210
box -6 -8 86 248
use AOI21X1  _424_
timestamp 0
transform 1 0 1450 0 1 730
box -6 -8 106 248
use OAI21X1  _425_
timestamp 0
transform 1 0 1490 0 -1 1690
box -6 -8 106 248
use NOR2X1  _426_
timestamp 0
transform -1 0 3530 0 1 2650
box -6 -8 86 248
use AND2X2  _427_
timestamp 0
transform -1 0 2910 0 -1 3610
box -6 -8 106 248
use OAI21X1  _428_
timestamp 0
transform -1 0 3270 0 1 2650
box -6 -8 106 248
use AOI21X1  _429_
timestamp 0
transform 1 0 3310 0 -1 2650
box -6 -8 106 248
use OAI21X1  _430_
timestamp 0
transform -1 0 4070 0 1 2170
box -6 -8 106 248
use NAND2X1  _431_
timestamp 0
transform 1 0 4070 0 1 1690
box -6 -8 86 248
use OAI21X1  _432_
timestamp 0
transform -1 0 3610 0 -1 1690
box -6 -8 106 248
use AOI21X1  _433_
timestamp 0
transform -1 0 3890 0 -1 1690
box -6 -8 106 248
use AOI21X1  _434_
timestamp 0
transform 1 0 4330 0 -1 2170
box -6 -8 106 248
use AND2X2  _435_
timestamp 0
transform 1 0 4810 0 1 1210
box -6 -8 106 248
use NOR2X1  _436_
timestamp 0
transform 1 0 4910 0 -1 1690
box -6 -8 86 248
use NOR2X1  _437_
timestamp 0
transform -1 0 4930 0 1 1690
box -6 -8 86 248
use OR2X2  _438_
timestamp 0
transform -1 0 4450 0 -1 1690
box -6 -8 106 248
use AOI21X1  _439_
timestamp 0
transform -1 0 4430 0 1 1690
box -6 -8 106 248
use OAI21X1  _440_
timestamp 0
transform -1 0 3630 0 1 1210
box -6 -8 106 248
use AOI21X1  _441_
timestamp 0
transform -1 0 4170 0 -1 1690
box -6 -8 106 248
use NAND2X1  _442_
timestamp 0
transform -1 0 4570 0 1 2170
box -6 -8 86 248
use AOI21X1  _443_
timestamp 0
transform 1 0 4750 0 1 2170
box -6 -8 106 248
use OAI21X1  _444_
timestamp 0
transform -1 0 4470 0 -1 2650
box -6 -8 106 248
use INVX1  _445_
timestamp 0
transform -1 0 4930 0 1 4090
box -6 -8 66 248
use NOR2X1  _446_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 86 248
use NOR2X1  _447_
timestamp 0
transform 1 0 4910 0 1 3610
box -6 -8 86 248
use NOR2X1  _448_
timestamp 0
transform -1 0 4750 0 -1 3130
box -6 -8 86 248
use NAND2X1  _449_
timestamp 0
transform 1 0 4250 0 1 2650
box -6 -8 86 248
use INVX1  _450_
timestamp 0
transform 1 0 4650 0 -1 2650
box -6 -8 66 248
use INVX1  _451_
timestamp 0
transform 1 0 4870 0 -1 2650
box -6 -8 66 248
use AOI21X1  _452_
timestamp 0
transform 1 0 4770 0 1 2650
box -6 -8 106 248
use OAI21X1  _453_
timestamp 0
transform 1 0 4930 0 -1 3130
box -6 -8 106 248
use NAND2X1  _454_
timestamp 0
transform 1 0 4410 0 -1 3130
box -6 -8 86 248
use OAI21X1  _455_
timestamp 0
transform -1 0 3970 0 -1 3130
box -6 -8 106 248
use AOI21X1  _456_
timestamp 0
transform -1 0 4230 0 -1 3130
box -6 -8 106 248
use INVX1  _457_
timestamp 0
transform 1 0 4130 0 -1 2650
box -6 -8 66 248
use NAND2X1  _458_
timestamp 0
transform -1 0 3930 0 -1 3610
box -6 -8 86 248
use INVX1  _459_
timestamp 0
transform -1 0 4910 0 -1 3610
box -6 -8 66 248
use OAI21X1  _460_
timestamp 0
transform 1 0 4930 0 1 3130
box -6 -8 106 248
use NAND2X1  _461_
timestamp 0
transform 1 0 4610 0 1 4570
box -6 -8 86 248
use OR2X2  _462_
timestamp 0
transform 1 0 4870 0 1 4570
box -6 -8 106 248
use NAND2X1  _463_
timestamp 0
transform 1 0 4930 0 -1 4570
box -6 -8 86 248
use NAND2X1  _464_
timestamp 0
transform 1 0 4350 0 -1 3610
box -6 -8 86 248
use AOI21X1  _465_
timestamp 0
transform 1 0 4490 0 1 2650
box -6 -8 106 248
use INVX1  _466_
timestamp 0
transform 1 0 4610 0 -1 3610
box -6 -8 66 248
use AOI21X1  _467_
timestamp 0
transform 1 0 4650 0 1 3130
box -6 -8 106 248
use AOI22X1  _468_
timestamp 0
transform 1 0 4350 0 1 3130
box -6 -8 126 248
use NOR2X1  _469_
timestamp 0
transform -1 0 3110 0 1 1210
box -6 -8 86 248
use OAI21X1  _470_
timestamp 0
transform -1 0 2570 0 1 730
box -6 -8 106 248
use NOR2X1  _471_
timestamp 0
transform -1 0 2770 0 -1 1210
box -6 -8 86 248
use NOR2X1  _472_
timestamp 0
transform 1 0 2230 0 1 730
box -6 -8 86 248
use OAI21X1  _473_
timestamp 0
transform 1 0 2530 0 -1 250
box -6 -8 106 248
use NOR2X1  _474_
timestamp 0
transform 1 0 2810 0 -1 730
box -6 -8 86 248
use OAI21X1  _475_
timestamp 0
transform 1 0 3450 0 -1 1210
box -6 -8 106 248
use AOI21X1  _476_
timestamp 0
transform 1 0 2950 0 -1 1210
box -6 -8 106 248
use OAI21X1  _477_
timestamp 0
transform -1 0 2510 0 -1 1210
box -6 -8 106 248
use AOI21X1  _478_
timestamp 0
transform -1 0 2390 0 1 1690
box -6 -8 106 248
use OAI21X1  _479_
timestamp 0
transform -1 0 3430 0 -1 3610
box -6 -8 106 248
use AOI21X1  _480_
timestamp 0
transform 1 0 3310 0 1 3130
box -6 -8 106 248
use OAI21X1  _481_
timestamp 0
transform -1 0 2890 0 1 3130
box -6 -8 106 248
use AOI21X1  _482_
timestamp 0
transform 1 0 2910 0 1 2650
box -6 -8 106 248
use OAI21X1  _483_
timestamp 0
transform -1 0 1550 0 1 4090
box -6 -8 106 248
use AOI21X1  _484_
timestamp 0
transform -1 0 1250 0 -1 4090
box -6 -8 106 248
use OAI21X1  _485_
timestamp 0
transform -1 0 1870 0 -1 3610
box -6 -8 106 248
use AOI21X1  _486_
timestamp 0
transform -1 0 1850 0 1 3130
box -6 -8 106 248
use OAI21X1  _487_
timestamp 0
transform -1 0 1590 0 -1 2170
box -6 -8 106 248
use AOI21X1  _488_
timestamp 0
transform -1 0 1310 0 -1 2170
box -6 -8 106 248
use OAI21X1  _489_
timestamp 0
transform -1 0 2110 0 1 1690
box -6 -8 106 248
use AOI21X1  _490_
timestamp 0
transform 1 0 1750 0 1 1690
box -6 -8 106 248
use NOR2X1  _491_
timestamp 0
transform 1 0 2850 0 -1 3130
box -6 -8 86 248
use OAI21X1  _492_
timestamp 0
transform -1 0 3690 0 -1 3130
box -6 -8 106 248
use NOR2X1  _493_
timestamp 0
transform 1 0 3090 0 -1 3130
box -6 -8 86 248
use INVX1  _494_
timestamp 0
transform 1 0 3070 0 1 3130
box -6 -8 66 248
use INVX1  _495_
timestamp 0
transform 1 0 2250 0 -1 2170
box -6 -8 66 248
use INVX1  _496_
timestamp 0
transform 1 0 930 0 -1 4090
box -6 -8 66 248
use INVX1  _497_
timestamp 0
transform -1 0 1750 0 1 2650
box -6 -8 66 248
use INVX1  _498_
timestamp 0
transform 1 0 1050 0 1 2170
box -6 -8 66 248
use INVX1  _499_
timestamp 0
transform 1 0 1450 0 1 2650
box -6 -8 66 248
use NAND2X1  _500_
timestamp 0
transform -1 0 2010 0 1 2650
box -6 -8 86 248
use OAI21X1  _501_
timestamp 0
transform 1 0 1290 0 1 2170
box -6 -8 106 248
use NAND2X1  _502_
timestamp 0
transform -1 0 1570 0 -1 2650
box -6 -8 86 248
use OAI21X1  _503_
timestamp 0
transform 1 0 1730 0 -1 2650
box -6 -8 106 248
use NAND2X1  _504_
timestamp 0
transform -1 0 2850 0 -1 2650
box -6 -8 86 248
use OAI21X1  _505_
timestamp 0
transform -1 0 3130 0 -1 2650
box -6 -8 106 248
use INVX1  _506_
timestamp 0
transform 1 0 3290 0 1 1210
box -6 -8 66 248
use NAND2X1  _507_
timestamp 0
transform 1 0 3010 0 -1 2170
box -6 -8 86 248
use OAI21X1  _508_
timestamp 0
transform -1 0 3010 0 1 2170
box -6 -8 106 248
use NAND2X1  _509_
timestamp 0
transform 1 0 3270 0 -1 1690
box -6 -8 86 248
use OAI21X1  _510_
timestamp 0
transform 1 0 3190 0 1 2170
box -6 -8 106 248
use INVX1  _511_
timestamp 0
transform 1 0 2670 0 1 2650
box -6 -8 66 248
use INVX1  _512_
timestamp 0
transform 1 0 1750 0 -1 2170
box -6 -8 66 248
use OAI21X1  _513_
timestamp 0
transform -1 0 1670 0 1 2170
box -6 -8 106 248
use INVX1  _514_
timestamp 0
transform 1 0 1630 0 -1 3130
box -6 -8 66 248
use AOI21X1  _515_
timestamp 0
transform 1 0 2010 0 -1 2650
box -6 -8 106 248
use OAI21X1  _516_
timestamp 0
transform 1 0 1850 0 1 2170
box -6 -8 106 248
use OAI21X1  _517_
timestamp 0
transform -1 0 2210 0 1 2170
box -6 -8 106 248
use INVX1  _518_
timestamp 0
transform -1 0 2890 0 1 1690
box -6 -8 66 248
use NAND2X1  _519_
timestamp 0
transform 1 0 2570 0 1 1690
box -6 -8 86 248
use OAI21X1  _520_
timestamp 0
transform 1 0 2490 0 -1 2170
box -6 -8 106 248
use NAND2X1  _521_
timestamp 0
transform 1 0 2770 0 -1 1690
box -6 -8 86 248
use OAI21X1  _522_
timestamp 0
transform -1 0 2850 0 -1 2170
box -6 -8 106 248
use INVX1  _523_
timestamp 0
transform 1 0 2370 0 -1 3130
box -6 -8 66 248
use NAND2X1  _524_
timestamp 0
transform 1 0 4410 0 1 3610
box -6 -8 86 248
use INVX1  _525_
timestamp 0
transform -1 0 4730 0 1 3610
box -6 -8 66 248
use INVX1  _526_
timestamp 0
transform -1 0 4690 0 1 4090
box -6 -8 66 248
use NAND2X1  _527_
timestamp 0
transform -1 0 4670 0 -1 4090
box -6 -8 86 248
use NAND2X1  _528_
timestamp 0
transform -1 0 4410 0 -1 4090
box -6 -8 86 248
use NAND2X1  _529_
timestamp 0
transform -1 0 4470 0 -1 4570
box -6 -8 86 248
use OAI21X1  _530_
timestamp 0
transform 1 0 4370 0 1 4090
box -6 -8 106 248
use INVX8  _531_
timestamp 0
transform -1 0 1970 0 -1 1210
box -6 -8 126 248
use INVX2  _532_
timestamp 0
transform -1 0 1050 0 -1 2650
box -6 -8 66 248
use NOR2X1  _533_
timestamp 0
transform -1 0 3950 0 -1 2650
box -6 -8 86 248
use AND2X2  _534_
timestamp 0
transform -1 0 3410 0 1 1690
box -6 -8 106 248
use AND2X2  _535_
timestamp 0
transform -1 0 2730 0 1 2170
box -6 -8 106 248
use NOR2X1  _536_
timestamp 0
transform 1 0 2270 0 -1 2650
box -6 -8 86 248
use NOR2X1  _537_
timestamp 0
transform -1 0 1310 0 -1 2650
box -6 -8 86 248
use NAND2X1  _538_
timestamp 0
transform 1 0 2030 0 1 3130
box -6 -8 86 248
use NOR2X1  _539_
timestamp 0
transform 1 0 2530 0 1 3130
box -6 -8 86 248
use INVX1  _540_
timestamp 0
transform 1 0 950 0 1 4090
box -6 -8 66 248
use NAND2X1  _541_
timestamp 0
transform 1 0 1190 0 1 4090
box -6 -8 86 248
use OAI21X1  _542_
timestamp 0
transform 1 0 1470 0 -1 4570
box -6 -8 106 248
use AOI21X1  _543_
timestamp 0
transform -1 0 1290 0 -1 4570
box -6 -8 106 248
use NAND2X1  _544_
timestamp 0
transform -1 0 790 0 1 4090
box -6 -8 86 248
use NAND2X1  _545_
timestamp 0
transform -1 0 250 0 -1 4570
box -6 -8 86 248
use INVX1  _546_
timestamp 0
transform -1 0 250 0 1 4090
box -6 -8 66 248
use NOR2X1  _547_
timestamp 0
transform -1 0 270 0 1 4570
box -6 -8 86 248
use OAI21X1  _548_
timestamp 0
transform -1 0 550 0 1 4570
box -6 -8 106 248
use OR2X2  _549_
timestamp 0
transform -1 0 530 0 -1 4570
box -6 -8 106 248
use NOR2X1  _550_
timestamp 0
transform -1 0 770 0 -1 4570
box -6 -8 86 248
use INVX1  _551_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 66 248
use NAND2X1  _552_
timestamp 0
transform 1 0 970 0 1 4570
box -6 -8 86 248
use OAI21X1  _553_
timestamp 0
transform 1 0 1230 0 1 4570
box -6 -8 106 248
use AOI21X1  _554_
timestamp 0
transform 1 0 1490 0 1 4570
box -6 -8 106 248
use OAI21X1  _555_
timestamp 0
transform -1 0 530 0 1 4090
box -6 -8 106 248
use AND2X2  _556_
timestamp 0
transform -1 0 290 0 1 3610
box -6 -8 106 248
use NOR2X1  _557_
timestamp 0
transform -1 0 270 0 -1 4090
box -6 -8 86 248
use NOR2X1  _558_
timestamp 0
transform 1 0 470 0 1 3610
box -6 -8 86 248
use AND2X2  _559_
timestamp 0
transform -1 0 270 0 -1 3610
box -6 -8 106 248
use NOR2X1  _560_
timestamp 0
transform -1 0 1070 0 -1 3610
box -6 -8 86 248
use OAI21X1  _561_
timestamp 0
transform 1 0 710 0 -1 3610
box -6 -8 106 248
use NAND2X1  _562_
timestamp 0
transform 1 0 1010 0 1 3610
box -6 -8 86 248
use AOI21X1  _563_
timestamp 0
transform -1 0 830 0 1 3610
box -6 -8 106 248
use OAI21X1  _564_
timestamp 0
transform -1 0 270 0 -1 2650
box -6 -8 106 248
use AND2X2  _565_
timestamp 0
transform 1 0 190 0 1 3130
box -6 -8 106 248
use NOR2X1  _566_
timestamp 0
transform 1 0 190 0 -1 3130
box -6 -8 86 248
use NOR2X1  _567_
timestamp 0
transform 1 0 470 0 1 3130
box -6 -8 86 248
use OAI21X1  _568_
timestamp 0
transform -1 0 810 0 1 3130
box -6 -8 106 248
use NOR2X1  _569_
timestamp 0
transform -1 0 1070 0 1 3130
box -6 -8 86 248
use OAI21X1  _570_
timestamp 0
transform 1 0 970 0 -1 3130
box -6 -8 106 248
use NAND2X1  _571_
timestamp 0
transform -1 0 790 0 1 2650
box -6 -8 86 248
use AOI21X1  _572_
timestamp 0
transform -1 0 530 0 1 2650
box -6 -8 106 248
use NAND3X1  _573_
timestamp 0
transform 1 0 430 0 -1 3610
box -6 -8 106 248
use INVX1  _574_
timestamp 0
transform -1 0 510 0 -1 3130
box -6 -8 66 248
use AOI21X1  _575_
timestamp 0
transform 1 0 690 0 -1 3130
box -6 -8 106 248
use AND2X2  _576_
timestamp 0
transform 1 0 710 0 -1 2650
box -6 -8 106 248
use AND2X2  _577_
timestamp 0
transform -1 0 290 0 -1 1210
box -6 -8 106 248
use NOR2X1  _578_
timestamp 0
transform -1 0 250 0 1 1210
box -6 -8 86 248
use OAI21X1  _579_
timestamp 0
transform 1 0 690 0 1 1210
box -6 -8 106 248
use NAND2X1  _580_
timestamp 0
transform -1 0 530 0 -1 2650
box -6 -8 86 248
use NOR2X1  _581_
timestamp 0
transform -1 0 510 0 1 1210
box -6 -8 86 248
use NAND2X1  _582_
timestamp 0
transform 1 0 950 0 -1 1690
box -6 -8 86 248
use NAND2X1  _583_
timestamp 0
transform -1 0 770 0 -1 1690
box -6 -8 86 248
use OAI21X1  _584_
timestamp 0
transform 1 0 550 0 1 2170
box -6 -8 106 248
use AOI21X1  _585_
timestamp 0
transform -1 0 770 0 -1 2170
box -6 -8 106 248
use AOI21X1  _586_
timestamp 0
transform -1 0 570 0 -1 1210
box -6 -8 106 248
use AND2X2  _587_
timestamp 0
transform -1 0 270 0 -1 730
box -6 -8 106 248
use NOR2X1  _588_
timestamp 0
transform -1 0 270 0 1 250
box -6 -8 86 248
use NOR2X1  _589_
timestamp 0
transform -1 0 270 0 1 730
box -6 -8 86 248
use NAND2X1  _590_
timestamp 0
transform -1 0 270 0 -1 1690
box -6 -8 86 248
use NOR2X1  _591_
timestamp 0
transform -1 0 530 0 -1 1690
box -6 -8 86 248
use NOR2X1  _592_
timestamp 0
transform -1 0 810 0 1 1690
box -6 -8 86 248
use OAI21X1  _593_
timestamp 0
transform 1 0 470 0 1 1690
box -6 -8 106 248
use AOI21X1  _594_
timestamp 0
transform -1 0 290 0 1 1690
box -6 -8 106 248
use INVX1  _595_
timestamp 0
transform -1 0 510 0 1 730
box -6 -8 66 248
use INVX1  _596_
timestamp 0
transform 1 0 710 0 -1 730
box -6 -8 66 248
use OAI21X1  _597_
timestamp 0
transform 1 0 670 0 1 730
box -6 -8 106 248
use AND2X2  _598_
timestamp 0
transform 1 0 750 0 -1 1210
box -6 -8 106 248
use AOI21X1  _599_
timestamp 0
transform 1 0 1310 0 -1 1210
box -6 -8 106 248
use NAND2X1  _600_
timestamp 0
transform -1 0 270 0 -1 250
box -6 -8 86 248
use OR2X2  _601_
timestamp 0
transform -1 0 770 0 1 250
box -6 -8 106 248
use NAND2X1  _602_
timestamp 0
transform -1 0 1030 0 -1 730
box -6 -8 86 248
use OR2X2  _603_
timestamp 0
transform 1 0 1590 0 -1 1210
box -6 -8 106 248
use INVX1  _604_
timestamp 0
transform 1 0 1750 0 1 250
box -6 -8 66 248
use INVX1  _605_
timestamp 0
transform 1 0 1210 0 -1 730
box -6 -8 66 248
use OAI21X1  _606_
timestamp 0
transform -1 0 1810 0 -1 730
box -6 -8 106 248
use NAND2X1  _607_
timestamp 0
transform 1 0 1730 0 1 1210
box -6 -8 86 248
use OAI21X1  _608_
timestamp 0
transform 1 0 1230 0 1 1690
box -6 -8 106 248
use AOI21X1  _609_
timestamp 0
transform -1 0 1310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _610_
timestamp 0
transform 1 0 1450 0 -1 730
box -6 -8 106 248
use NAND2X1  _611_
timestamp 0
transform -1 0 1570 0 1 250
box -6 -8 86 248
use OR2X2  _612_
timestamp 0
transform 1 0 1230 0 -1 250
box -6 -8 106 248
use NAND2X1  _613_
timestamp 0
transform 1 0 1990 0 1 250
box -6 -8 86 248
use OR2X2  _614_
timestamp 0
transform 1 0 1990 0 -1 730
box -6 -8 106 248
use AOI21X1  _615_
timestamp 0
transform 1 0 2250 0 -1 730
box -6 -8 106 248
use OAI21X1  _616_
timestamp 0
transform 1 0 2510 0 1 250
box -6 -8 106 248
use AOI21X1  _617_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 106 248
use NAND2X1  _618_
timestamp 0
transform 1 0 970 0 1 1210
box -6 -8 86 248
use AND2X2  _619_
timestamp 0
transform -1 0 550 0 -1 250
box -6 -8 106 248
use NOR2X1  _620_
timestamp 0
transform 1 0 970 0 -1 250
box -6 -8 86 248
use NOR2X1  _621_
timestamp 0
transform -1 0 810 0 -1 250
box -6 -8 86 248
use NAND3X1  _622_
timestamp 0
transform -1 0 1050 0 1 250
box -6 -8 106 248
use NOR2X1  _623_
timestamp 0
transform 1 0 1230 0 1 1210
box -6 -8 86 248
use INVX1  _624_
timestamp 0
transform 1 0 450 0 1 250
box -6 -8 66 248
use AOI21X1  _625_
timestamp 0
transform 1 0 430 0 -1 730
box -6 -8 106 248
use DFFPOSX1  _626_
timestamp 0
transform -1 0 3790 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _627_
timestamp 0
transform -1 0 3130 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _628_
timestamp 0
transform -1 0 2450 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _629_
timestamp 0
transform -1 0 2250 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _630_
timestamp 0
transform 1 0 1030 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _631_
timestamp 0
transform 1 0 1950 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _632_
timestamp 0
transform -1 0 2350 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _633_
timestamp 0
transform -1 0 1010 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _634_
timestamp 0
transform -1 0 1810 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _635_
timestamp 0
transform -1 0 510 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _636_
timestamp 0
transform 1 0 10 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _637_
timestamp 0
transform -1 0 490 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _638_
timestamp 0
transform 1 0 10 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _639_
timestamp 0
transform 1 0 810 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _640_
timestamp 0
transform -1 0 1570 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _641_
timestamp 0
transform -1 0 3410 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _642_
timestamp 0
transform 1 0 1570 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _643_
timestamp 0
transform 1 0 3670 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _644_
timestamp 0
transform -1 0 3870 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _645_
timestamp 0
transform -1 0 3670 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _646_
timestamp 0
transform 1 0 3410 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _647_
timestamp 0
transform -1 0 2050 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _648_
timestamp 0
transform 1 0 1250 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _649_
timestamp 0
transform -1 0 3650 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _650_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _651_
timestamp 0
transform -1 0 4170 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _652_
timestamp 0
transform -1 0 4170 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _653_
timestamp 0
transform 1 0 2850 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _654_
timestamp 0
transform 1 0 1810 0 1 730
box -6 -8 246 248
use DFFPOSX1  _655_
timestamp 0
transform 1 0 3050 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _656_
timestamp 0
transform 1 0 2350 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _657_
timestamp 0
transform -1 0 3650 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _658_
timestamp 0
transform 1 0 2250 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _659_
timestamp 0
transform 1 0 510 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _660_
timestamp 0
transform 1 0 1330 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _661_
timestamp 0
transform 1 0 650 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _662_
timestamp 0
transform 1 0 1330 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _663_
timestamp 0
transform -1 0 2670 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _664_
timestamp 0
transform 1 0 3910 0 -1 4090
box -6 -8 246 248
use BUFX2  _665_
timestamp 0
transform 1 0 3470 0 1 2170
box -6 -8 86 248
use BUFX2  _666_
timestamp 0
transform 1 0 2830 0 1 4570
box -6 -8 86 248
use BUFX2  _667_
timestamp 0
transform -1 0 4450 0 1 4570
box -6 -8 86 248
use BUFX2  _668_
timestamp 0
transform 1 0 2030 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 1030 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 2770 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform 1 0 1510 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 1250 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform -1 0 2070 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 2510 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 1250 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 2250 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert14
timestamp 0
transform -1 0 1030 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 2510 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 3330 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 1990 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform 1 0 3270 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform 1 0 2150 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 1870 0 -1 3130
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert0
timestamp 0
transform 1 0 2150 0 -1 1690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert1
timestamp 0
transform -1 0 1970 0 -1 1690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert2
timestamp 0
transform 1 0 170 0 1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert3
timestamp 0
transform 1 0 1930 0 1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert4
timestamp 0
transform 1 0 1250 0 -1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert5
timestamp 0
transform 1 0 1270 0 1 3610
box -6 -8 206 248
use FILL  FILL73050x39750
timestamp 0
transform 1 0 4870 0 1 2650
box -6 -8 26 248
use FILL  FILL73350x39750
timestamp 0
transform 1 0 4890 0 1 2650
box -6 -8 26 248
use FILL  FILL73650x18150
timestamp 0
transform 1 0 4910 0 1 1210
box -6 -8 26 248
use FILL  FILL73650x39750
timestamp 0
transform 1 0 4910 0 1 2650
box -6 -8 26 248
use FILL  FILL73650x50550
timestamp 0
transform -1 0 4930 0 -1 3610
box -6 -8 26 248
use FILL  FILL73650x57750
timestamp 0
transform -1 0 4930 0 -1 4090
box -6 -8 26 248
use FILL  FILL73950x150
timestamp 0
transform -1 0 4950 0 -1 250
box -6 -8 26 248
use FILL  FILL73950x10950
timestamp 0
transform 1 0 4930 0 1 730
box -6 -8 26 248
use FILL  FILL73950x14550
timestamp 0
transform -1 0 4950 0 -1 1210
box -6 -8 26 248
use FILL  FILL73950x18150
timestamp 0
transform 1 0 4930 0 1 1210
box -6 -8 26 248
use FILL  FILL73950x25350
timestamp 0
transform 1 0 4930 0 1 1690
box -6 -8 26 248
use FILL  FILL73950x36150
timestamp 0
transform -1 0 4950 0 -1 2650
box -6 -8 26 248
use FILL  FILL73950x39750
timestamp 0
transform 1 0 4930 0 1 2650
box -6 -8 26 248
use FILL  FILL73950x50550
timestamp 0
transform -1 0 4950 0 -1 3610
box -6 -8 26 248
use FILL  FILL73950x57750
timestamp 0
transform -1 0 4950 0 -1 4090
box -6 -8 26 248
use FILL  FILL73950x61350
timestamp 0
transform 1 0 4930 0 1 4090
box -6 -8 26 248
use FILL  FILL74250x150
timestamp 0
transform -1 0 4970 0 -1 250
box -6 -8 26 248
use FILL  FILL74250x10950
timestamp 0
transform 1 0 4950 0 1 730
box -6 -8 26 248
use FILL  FILL74250x14550
timestamp 0
transform -1 0 4970 0 -1 1210
box -6 -8 26 248
use FILL  FILL74250x18150
timestamp 0
transform 1 0 4950 0 1 1210
box -6 -8 26 248
use FILL  FILL74250x25350
timestamp 0
transform 1 0 4950 0 1 1690
box -6 -8 26 248
use FILL  FILL74250x28950
timestamp 0
transform -1 0 4970 0 -1 2170
box -6 -8 26 248
use FILL  FILL74250x36150
timestamp 0
transform -1 0 4970 0 -1 2650
box -6 -8 26 248
use FILL  FILL74250x39750
timestamp 0
transform 1 0 4950 0 1 2650
box -6 -8 26 248
use FILL  FILL74250x50550
timestamp 0
transform -1 0 4970 0 -1 3610
box -6 -8 26 248
use FILL  FILL74250x57750
timestamp 0
transform -1 0 4970 0 -1 4090
box -6 -8 26 248
use FILL  FILL74250x61350
timestamp 0
transform 1 0 4950 0 1 4090
box -6 -8 26 248
use FILL  FILL74550x150
timestamp 0
transform -1 0 4990 0 -1 250
box -6 -8 26 248
use FILL  FILL74550x7350
timestamp 0
transform -1 0 4990 0 -1 730
box -6 -8 26 248
use FILL  FILL74550x10950
timestamp 0
transform 1 0 4970 0 1 730
box -6 -8 26 248
use FILL  FILL74550x14550
timestamp 0
transform -1 0 4990 0 -1 1210
box -6 -8 26 248
use FILL  FILL74550x18150
timestamp 0
transform 1 0 4970 0 1 1210
box -6 -8 26 248
use FILL  FILL74550x25350
timestamp 0
transform 1 0 4970 0 1 1690
box -6 -8 26 248
use FILL  FILL74550x28950
timestamp 0
transform -1 0 4990 0 -1 2170
box -6 -8 26 248
use FILL  FILL74550x36150
timestamp 0
transform -1 0 4990 0 -1 2650
box -6 -8 26 248
use FILL  FILL74550x39750
timestamp 0
transform 1 0 4970 0 1 2650
box -6 -8 26 248
use FILL  FILL74550x50550
timestamp 0
transform -1 0 4990 0 -1 3610
box -6 -8 26 248
use FILL  FILL74550x57750
timestamp 0
transform -1 0 4990 0 -1 4090
box -6 -8 26 248
use FILL  FILL74550x61350
timestamp 0
transform 1 0 4970 0 1 4090
box -6 -8 26 248
use FILL  FILL74550x68550
timestamp 0
transform 1 0 4970 0 1 4570
box -6 -8 26 248
use FILL  FILL74850x150
timestamp 0
transform -1 0 5010 0 -1 250
box -6 -8 26 248
use FILL  FILL74850x3750
timestamp 0
transform 1 0 4990 0 1 250
box -6 -8 26 248
use FILL  FILL74850x7350
timestamp 0
transform -1 0 5010 0 -1 730
box -6 -8 26 248
use FILL  FILL74850x10950
timestamp 0
transform 1 0 4990 0 1 730
box -6 -8 26 248
use FILL  FILL74850x14550
timestamp 0
transform -1 0 5010 0 -1 1210
box -6 -8 26 248
use FILL  FILL74850x18150
timestamp 0
transform 1 0 4990 0 1 1210
box -6 -8 26 248
use FILL  FILL74850x21750
timestamp 0
transform -1 0 5010 0 -1 1690
box -6 -8 26 248
use FILL  FILL74850x25350
timestamp 0
transform 1 0 4990 0 1 1690
box -6 -8 26 248
use FILL  FILL74850x28950
timestamp 0
transform -1 0 5010 0 -1 2170
box -6 -8 26 248
use FILL  FILL74850x36150
timestamp 0
transform -1 0 5010 0 -1 2650
box -6 -8 26 248
use FILL  FILL74850x39750
timestamp 0
transform 1 0 4990 0 1 2650
box -6 -8 26 248
use FILL  FILL74850x50550
timestamp 0
transform -1 0 5010 0 -1 3610
box -6 -8 26 248
use FILL  FILL74850x54150
timestamp 0
transform 1 0 4990 0 1 3610
box -6 -8 26 248
use FILL  FILL74850x57750
timestamp 0
transform -1 0 5010 0 -1 4090
box -6 -8 26 248
use FILL  FILL74850x61350
timestamp 0
transform 1 0 4990 0 1 4090
box -6 -8 26 248
use FILL  FILL74850x68550
timestamp 0
transform 1 0 4990 0 1 4570
box -6 -8 26 248
use FILL  FILL75150x150
timestamp 0
transform -1 0 5030 0 -1 250
box -6 -8 26 248
use FILL  FILL75150x3750
timestamp 0
transform 1 0 5010 0 1 250
box -6 -8 26 248
use FILL  FILL75150x7350
timestamp 0
transform -1 0 5030 0 -1 730
box -6 -8 26 248
use FILL  FILL75150x10950
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 26 248
use FILL  FILL75150x14550
timestamp 0
transform -1 0 5030 0 -1 1210
box -6 -8 26 248
use FILL  FILL75150x18150
timestamp 0
transform 1 0 5010 0 1 1210
box -6 -8 26 248
use FILL  FILL75150x21750
timestamp 0
transform -1 0 5030 0 -1 1690
box -6 -8 26 248
use FILL  FILL75150x25350
timestamp 0
transform 1 0 5010 0 1 1690
box -6 -8 26 248
use FILL  FILL75150x28950
timestamp 0
transform -1 0 5030 0 -1 2170
box -6 -8 26 248
use FILL  FILL75150x36150
timestamp 0
transform -1 0 5030 0 -1 2650
box -6 -8 26 248
use FILL  FILL75150x39750
timestamp 0
transform 1 0 5010 0 1 2650
box -6 -8 26 248
use FILL  FILL75150x50550
timestamp 0
transform -1 0 5030 0 -1 3610
box -6 -8 26 248
use FILL  FILL75150x54150
timestamp 0
transform 1 0 5010 0 1 3610
box -6 -8 26 248
use FILL  FILL75150x57750
timestamp 0
transform -1 0 5030 0 -1 4090
box -6 -8 26 248
use FILL  FILL75150x61350
timestamp 0
transform 1 0 5010 0 1 4090
box -6 -8 26 248
use FILL  FILL75150x64950
timestamp 0
transform -1 0 5030 0 -1 4570
box -6 -8 26 248
use FILL  FILL75150x68550
timestamp 0
transform 1 0 5010 0 1 4570
box -6 -8 26 248
use FILL  FILL75450x150
timestamp 0
transform -1 0 5050 0 -1 250
box -6 -8 26 248
use FILL  FILL75450x3750
timestamp 0
transform 1 0 5030 0 1 250
box -6 -8 26 248
use FILL  FILL75450x7350
timestamp 0
transform -1 0 5050 0 -1 730
box -6 -8 26 248
use FILL  FILL75450x10950
timestamp 0
transform 1 0 5030 0 1 730
box -6 -8 26 248
use FILL  FILL75450x14550
timestamp 0
transform -1 0 5050 0 -1 1210
box -6 -8 26 248
use FILL  FILL75450x18150
timestamp 0
transform 1 0 5030 0 1 1210
box -6 -8 26 248
use FILL  FILL75450x21750
timestamp 0
transform -1 0 5050 0 -1 1690
box -6 -8 26 248
use FILL  FILL75450x25350
timestamp 0
transform 1 0 5030 0 1 1690
box -6 -8 26 248
use FILL  FILL75450x28950
timestamp 0
transform -1 0 5050 0 -1 2170
box -6 -8 26 248
use FILL  FILL75450x36150
timestamp 0
transform -1 0 5050 0 -1 2650
box -6 -8 26 248
use FILL  FILL75450x39750
timestamp 0
transform 1 0 5030 0 1 2650
box -6 -8 26 248
use FILL  FILL75450x43350
timestamp 0
transform -1 0 5050 0 -1 3130
box -6 -8 26 248
use FILL  FILL75450x46950
timestamp 0
transform 1 0 5030 0 1 3130
box -6 -8 26 248
use FILL  FILL75450x50550
timestamp 0
transform -1 0 5050 0 -1 3610
box -6 -8 26 248
use FILL  FILL75450x54150
timestamp 0
transform 1 0 5030 0 1 3610
box -6 -8 26 248
use FILL  FILL75450x57750
timestamp 0
transform -1 0 5050 0 -1 4090
box -6 -8 26 248
use FILL  FILL75450x61350
timestamp 0
transform 1 0 5030 0 1 4090
box -6 -8 26 248
use FILL  FILL75450x64950
timestamp 0
transform -1 0 5050 0 -1 4570
box -6 -8 26 248
use FILL  FILL75450x68550
timestamp 0
transform 1 0 5030 0 1 4570
box -6 -8 26 248
use FILL  FILL75750x150
timestamp 0
transform -1 0 5070 0 -1 250
box -6 -8 26 248
use FILL  FILL75750x3750
timestamp 0
transform 1 0 5050 0 1 250
box -6 -8 26 248
use FILL  FILL75750x7350
timestamp 0
transform -1 0 5070 0 -1 730
box -6 -8 26 248
use FILL  FILL75750x10950
timestamp 0
transform 1 0 5050 0 1 730
box -6 -8 26 248
use FILL  FILL75750x14550
timestamp 0
transform -1 0 5070 0 -1 1210
box -6 -8 26 248
use FILL  FILL75750x18150
timestamp 0
transform 1 0 5050 0 1 1210
box -6 -8 26 248
use FILL  FILL75750x21750
timestamp 0
transform -1 0 5070 0 -1 1690
box -6 -8 26 248
use FILL  FILL75750x25350
timestamp 0
transform 1 0 5050 0 1 1690
box -6 -8 26 248
use FILL  FILL75750x28950
timestamp 0
transform -1 0 5070 0 -1 2170
box -6 -8 26 248
use FILL  FILL75750x36150
timestamp 0
transform -1 0 5070 0 -1 2650
box -6 -8 26 248
use FILL  FILL75750x39750
timestamp 0
transform 1 0 5050 0 1 2650
box -6 -8 26 248
use FILL  FILL75750x43350
timestamp 0
transform -1 0 5070 0 -1 3130
box -6 -8 26 248
use FILL  FILL75750x46950
timestamp 0
transform 1 0 5050 0 1 3130
box -6 -8 26 248
use FILL  FILL75750x50550
timestamp 0
transform -1 0 5070 0 -1 3610
box -6 -8 26 248
use FILL  FILL75750x54150
timestamp 0
transform 1 0 5050 0 1 3610
box -6 -8 26 248
use FILL  FILL75750x57750
timestamp 0
transform -1 0 5070 0 -1 4090
box -6 -8 26 248
use FILL  FILL75750x61350
timestamp 0
transform 1 0 5050 0 1 4090
box -6 -8 26 248
use FILL  FILL75750x64950
timestamp 0
transform -1 0 5070 0 -1 4570
box -6 -8 26 248
use FILL  FILL75750x68550
timestamp 0
transform 1 0 5050 0 1 4570
box -6 -8 26 248
use FILL  FILL76050x150
timestamp 0
transform -1 0 5090 0 -1 250
box -6 -8 26 248
use FILL  FILL76050x3750
timestamp 0
transform 1 0 5070 0 1 250
box -6 -8 26 248
use FILL  FILL76050x7350
timestamp 0
transform -1 0 5090 0 -1 730
box -6 -8 26 248
use FILL  FILL76050x10950
timestamp 0
transform 1 0 5070 0 1 730
box -6 -8 26 248
use FILL  FILL76050x14550
timestamp 0
transform -1 0 5090 0 -1 1210
box -6 -8 26 248
use FILL  FILL76050x18150
timestamp 0
transform 1 0 5070 0 1 1210
box -6 -8 26 248
use FILL  FILL76050x21750
timestamp 0
transform -1 0 5090 0 -1 1690
box -6 -8 26 248
use FILL  FILL76050x25350
timestamp 0
transform 1 0 5070 0 1 1690
box -6 -8 26 248
use FILL  FILL76050x28950
timestamp 0
transform -1 0 5090 0 -1 2170
box -6 -8 26 248
use FILL  FILL76050x36150
timestamp 0
transform -1 0 5090 0 -1 2650
box -6 -8 26 248
use FILL  FILL76050x39750
timestamp 0
transform 1 0 5070 0 1 2650
box -6 -8 26 248
use FILL  FILL76050x43350
timestamp 0
transform -1 0 5090 0 -1 3130
box -6 -8 26 248
use FILL  FILL76050x46950
timestamp 0
transform 1 0 5070 0 1 3130
box -6 -8 26 248
use FILL  FILL76050x50550
timestamp 0
transform -1 0 5090 0 -1 3610
box -6 -8 26 248
use FILL  FILL76050x54150
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL76050x57750
timestamp 0
transform -1 0 5090 0 -1 4090
box -6 -8 26 248
use FILL  FILL76050x61350
timestamp 0
transform 1 0 5070 0 1 4090
box -6 -8 26 248
use FILL  FILL76050x64950
timestamp 0
transform -1 0 5090 0 -1 4570
box -6 -8 26 248
use FILL  FILL76050x68550
timestamp 0
transform 1 0 5070 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__313_
timestamp 0
transform 1 0 1050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__314_
timestamp 0
transform -1 0 1050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__315_
timestamp 0
transform 1 0 770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__316_
timestamp 0
transform -1 0 870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__317_
timestamp 0
transform -1 0 2630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__318_
timestamp 0
transform 1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__319_
timestamp 0
transform -1 0 3170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__320_
timestamp 0
transform -1 0 3110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__321_
timestamp 0
transform 1 0 3410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__322_
timestamp 0
transform 1 0 2830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__323_
timestamp 0
transform -1 0 2910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__324_
timestamp 0
transform -1 0 2590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__325_
timestamp 0
transform -1 0 3430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__326_
timestamp 0
transform -1 0 3710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__327_
timestamp 0
transform 1 0 4690 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__328_
timestamp 0
transform 1 0 4210 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__329_
timestamp 0
transform -1 0 4470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__330_
timestamp 0
transform 1 0 3950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__331_
timestamp 0
transform -1 0 2910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__332_
timestamp 0
transform -1 0 2650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__333_
timestamp 0
transform 1 0 2090 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__334_
timestamp 0
transform 1 0 2070 0 1 250
box -6 -8 26 248
use FILL  FILL_0__335_
timestamp 0
transform -1 0 1830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__336_
timestamp 0
transform -1 0 3170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__337_
timestamp 0
transform 1 0 3410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__338_
timestamp 0
transform -1 0 3990 0 1 250
box -6 -8 26 248
use FILL  FILL_0__339_
timestamp 0
transform 1 0 3690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__340_
timestamp 0
transform 1 0 4190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__341_
timestamp 0
transform 1 0 4650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__342_
timestamp 0
transform 1 0 4730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__343_
timestamp 0
transform -1 0 4750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__344_
timestamp 0
transform -1 0 4490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__345_
timestamp 0
transform -1 0 4470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__346_
timestamp 0
transform 1 0 4150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__347_
timestamp 0
transform -1 0 3370 0 1 730
box -6 -8 26 248
use FILL  FILL_0__348_
timestamp 0
transform -1 0 3650 0 1 730
box -6 -8 26 248
use FILL  FILL_0__349_
timestamp 0
transform 1 0 4670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__350_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__351_
timestamp 0
transform 1 0 4450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__352_
timestamp 0
transform 1 0 4430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__353_
timestamp 0
transform 1 0 4110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__354_
timestamp 0
transform 1 0 3870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__355_
timestamp 0
transform 1 0 4370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__356_
timestamp 0
transform -1 0 4110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__357_
timestamp 0
transform -1 0 3570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__358_
timestamp 0
transform -1 0 3830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__359_
timestamp 0
transform -1 0 3430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__360_
timestamp 0
transform 1 0 3910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__361_
timestamp 0
transform 1 0 4170 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__362_
timestamp 0
transform -1 0 3910 0 1 730
box -6 -8 26 248
use FILL  FILL_0__363_
timestamp 0
transform -1 0 4870 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__364_
timestamp 0
transform -1 0 4370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__365_
timestamp 0
transform -1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__366_
timestamp 0
transform -1 0 3430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__367_
timestamp 0
transform 1 0 3950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__368_
timestamp 0
transform 1 0 4470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__369_
timestamp 0
transform 1 0 3950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__370_
timestamp 0
transform 1 0 3650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__371_
timestamp 0
transform 1 0 3930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__372_
timestamp 0
transform 1 0 3950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__373_
timestamp 0
transform -1 0 3690 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__374_
timestamp 0
transform -1 0 3710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__375_
timestamp 0
transform 1 0 3670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__376_
timestamp 0
transform 1 0 3190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__377_
timestamp 0
transform -1 0 2930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__378_
timestamp 0
transform 1 0 3410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__379_
timestamp 0
transform -1 0 3150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__380_
timestamp 0
transform -1 0 3430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__381_
timestamp 0
transform -1 0 3170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__382_
timestamp 0
transform 1 0 3130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__383_
timestamp 0
transform -1 0 2890 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__384_
timestamp 0
transform 1 0 3690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__385_
timestamp 0
transform -1 0 3450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__386_
timestamp 0
transform -1 0 2610 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__387_
timestamp 0
transform 1 0 2110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__388_
timestamp 0
transform 1 0 2390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__389_
timestamp 0
transform -1 0 2890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__390_
timestamp 0
transform -1 0 1810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__391_
timestamp 0
transform -1 0 2610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__392_
timestamp 0
transform -1 0 2350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__393_
timestamp 0
transform 1 0 1590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__394_
timestamp 0
transform -1 0 2070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__395_
timestamp 0
transform -1 0 1570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__396_
timestamp 0
transform 1 0 2130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__397_
timestamp 0
transform 1 0 2630 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__398_
timestamp 0
transform 1 0 2110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__399_
timestamp 0
transform 1 0 2390 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__400_
timestamp 0
transform -1 0 1790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__401_
timestamp 0
transform -1 0 2070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__402_
timestamp 0
transform -1 0 1890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__403_
timestamp 0
transform 1 0 2310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__404_
timestamp 0
transform -1 0 2070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__405_
timestamp 0
transform 1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__406_
timestamp 0
transform -1 0 1510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__407_
timestamp 0
transform 1 0 3150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__408_
timestamp 0
transform -1 0 2870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__409_
timestamp 0
transform 1 0 3530 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__410_
timestamp 0
transform -1 0 3650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__411_
timestamp 0
transform -1 0 2350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__412_
timestamp 0
transform 1 0 2570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__413_
timestamp 0
transform -1 0 2890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__414_
timestamp 0
transform 1 0 2370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__415_
timestamp 0
transform 1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__416_
timestamp 0
transform 1 0 3650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__417_
timestamp 0
transform -1 0 3810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__418_
timestamp 0
transform 1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__419_
timestamp 0
transform 1 0 4430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__420_
timestamp 0
transform -1 0 4090 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__421_
timestamp 0
transform -1 0 3910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__422_
timestamp 0
transform -1 0 1570 0 1 730
box -6 -8 26 248
use FILL  FILL_0__423_
timestamp 0
transform 1 0 1310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__424_
timestamp 0
transform 1 0 1270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__425_
timestamp 0
transform 1 0 1310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__426_
timestamp 0
transform -1 0 3290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__427_
timestamp 0
transform -1 0 2650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__428_
timestamp 0
transform -1 0 3030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__429_
timestamp 0
transform 1 0 3130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__430_
timestamp 0
transform -1 0 3810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__431_
timestamp 0
transform 1 0 3890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__432_
timestamp 0
transform -1 0 3370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__433_
timestamp 0
transform -1 0 3630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__434_
timestamp 0
transform 1 0 4150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__435_
timestamp 0
transform 1 0 4630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__436_
timestamp 0
transform 1 0 4730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__437_
timestamp 0
transform -1 0 4710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__438_
timestamp 0
transform -1 0 4190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__439_
timestamp 0
transform -1 0 4170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__440_
timestamp 0
transform -1 0 3370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__441_
timestamp 0
transform -1 0 3910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__442_
timestamp 0
transform -1 0 4350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__443_
timestamp 0
transform 1 0 4570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__444_
timestamp 0
transform -1 0 4210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__445_
timestamp 0
transform -1 0 4710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__446_
timestamp 0
transform 1 0 4670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__447_
timestamp 0
transform 1 0 4730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__448_
timestamp 0
transform -1 0 4510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__449_
timestamp 0
transform 1 0 4070 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__450_
timestamp 0
transform 1 0 4470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__451_
timestamp 0
transform 1 0 4710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__452_
timestamp 0
transform 1 0 4590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__453_
timestamp 0
transform 1 0 4750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__454_
timestamp 0
transform 1 0 4230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__455_
timestamp 0
transform -1 0 3710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__456_
timestamp 0
transform -1 0 3990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__457_
timestamp 0
transform 1 0 3950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__458_
timestamp 0
transform -1 0 3690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__459_
timestamp 0
transform -1 0 4690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__460_
timestamp 0
transform 1 0 4750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__461_
timestamp 0
transform 1 0 4450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__462_
timestamp 0
transform 1 0 4690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__463_
timestamp 0
transform 1 0 4750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__464_
timestamp 0
transform 1 0 4170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__465_
timestamp 0
transform 1 0 4330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__466_
timestamp 0
transform 1 0 4430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__467_
timestamp 0
transform 1 0 4470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__468_
timestamp 0
transform 1 0 4170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__469_
timestamp 0
transform -1 0 2870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__470_
timestamp 0
transform -1 0 2330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__471_
timestamp 0
transform -1 0 2530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__472_
timestamp 0
transform 1 0 2050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__473_
timestamp 0
transform 1 0 2350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__474_
timestamp 0
transform 1 0 2630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__475_
timestamp 0
transform 1 0 3290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__476_
timestamp 0
transform 1 0 2770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__477_
timestamp 0
transform -1 0 2250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__478_
timestamp 0
transform -1 0 2130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__479_
timestamp 0
transform -1 0 3190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__480_
timestamp 0
transform 1 0 3130 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__481_
timestamp 0
transform -1 0 2630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__482_
timestamp 0
transform 1 0 2730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__483_
timestamp 0
transform -1 0 1290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__484_
timestamp 0
transform -1 0 1010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__485_
timestamp 0
transform -1 0 1610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__486_
timestamp 0
transform -1 0 1590 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__487_
timestamp 0
transform -1 0 1330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__488_
timestamp 0
transform -1 0 1050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__489_
timestamp 0
transform -1 0 1870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__490_
timestamp 0
transform 1 0 1570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__491_
timestamp 0
transform 1 0 2670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__492_
timestamp 0
transform -1 0 3430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__493_
timestamp 0
transform 1 0 2930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__494_
timestamp 0
transform 1 0 2890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__495_
timestamp 0
transform 1 0 2070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__496_
timestamp 0
transform 1 0 750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__497_
timestamp 0
transform -1 0 1530 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__498_
timestamp 0
transform 1 0 890 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__499_
timestamp 0
transform 1 0 1270 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__500_
timestamp 0
transform -1 0 1770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__501_
timestamp 0
transform 1 0 1110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__502_
timestamp 0
transform -1 0 1330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__503_
timestamp 0
transform 1 0 1570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__504_
timestamp 0
transform -1 0 2610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__505_
timestamp 0
transform -1 0 2870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__506_
timestamp 0
transform 1 0 3110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__507_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__508_
timestamp 0
transform -1 0 2750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__509_
timestamp 0
transform 1 0 3090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__510_
timestamp 0
transform 1 0 3010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__511_
timestamp 0
transform 1 0 2490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__512_
timestamp 0
transform 1 0 1590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__513_
timestamp 0
transform -1 0 1410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__514_
timestamp 0
transform 1 0 1450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__515_
timestamp 0
transform 1 0 1830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__516_
timestamp 0
transform 1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__517_
timestamp 0
transform -1 0 1970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__518_
timestamp 0
transform -1 0 2670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__519_
timestamp 0
transform 1 0 2390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__520_
timestamp 0
transform 1 0 2310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__521_
timestamp 0
transform 1 0 2590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__522_
timestamp 0
transform -1 0 2610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__523_
timestamp 0
transform 1 0 2190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__524_
timestamp 0
transform 1 0 4230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__525_
timestamp 0
transform -1 0 4510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__526_
timestamp 0
transform -1 0 4490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__527_
timestamp 0
transform -1 0 4430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__528_
timestamp 0
transform -1 0 4170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__529_
timestamp 0
transform -1 0 4230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__530_
timestamp 0
transform 1 0 4190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__531_
timestamp 0
transform -1 0 1710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__532_
timestamp 0
transform -1 0 830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__533_
timestamp 0
transform -1 0 3710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__534_
timestamp 0
transform -1 0 3150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__535_
timestamp 0
transform -1 0 2470 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__536_
timestamp 0
transform 1 0 2110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__537_
timestamp 0
transform -1 0 1070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__538_
timestamp 0
transform 1 0 1850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__539_
timestamp 0
transform 1 0 2350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__540_
timestamp 0
transform 1 0 790 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__541_
timestamp 0
transform 1 0 1010 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__542_
timestamp 0
transform 1 0 1290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__543_
timestamp 0
transform -1 0 1030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__544_
timestamp 0
transform -1 0 550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__545_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__546_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__547_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__548_
timestamp 0
transform -1 0 290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__549_
timestamp 0
transform -1 0 270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__550_
timestamp 0
transform -1 0 550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__551_
timestamp 0
transform 1 0 550 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__552_
timestamp 0
transform 1 0 790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__553_
timestamp 0
transform 1 0 1050 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__554_
timestamp 0
transform 1 0 1330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__555_
timestamp 0
transform -1 0 270 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__556_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__557_
timestamp 0
transform -1 0 30 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__558_
timestamp 0
transform 1 0 290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__559_
timestamp 0
transform -1 0 30 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__560_
timestamp 0
transform -1 0 830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__561_
timestamp 0
transform 1 0 530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__562_
timestamp 0
transform 1 0 830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__563_
timestamp 0
transform -1 0 570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__564_
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__565_
timestamp 0
transform 1 0 10 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__566_
timestamp 0
transform 1 0 10 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__567_
timestamp 0
transform 1 0 290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__568_
timestamp 0
transform -1 0 570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__569_
timestamp 0
transform -1 0 830 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__570_
timestamp 0
transform 1 0 790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__571_
timestamp 0
transform -1 0 550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__572_
timestamp 0
transform -1 0 270 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__573_
timestamp 0
transform 1 0 270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__574_
timestamp 0
transform -1 0 290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__575_
timestamp 0
transform 1 0 510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__576_
timestamp 0
transform 1 0 530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__577_
timestamp 0
transform -1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__578_
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__579_
timestamp 0
transform 1 0 510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__580_
timestamp 0
transform -1 0 290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__581_
timestamp 0
transform -1 0 270 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__582_
timestamp 0
transform 1 0 770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__583_
timestamp 0
transform -1 0 550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__584_
timestamp 0
transform 1 0 370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__585_
timestamp 0
transform -1 0 510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__586_
timestamp 0
transform -1 0 310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__587_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__588_
timestamp 0
transform -1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_0__589_
timestamp 0
transform -1 0 30 0 1 730
box -6 -8 26 248
use FILL  FILL_0__590_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__591_
timestamp 0
transform -1 0 290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__592_
timestamp 0
transform -1 0 590 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__593_
timestamp 0
transform 1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__594_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__595_
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__596_
timestamp 0
transform 1 0 530 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__597_
timestamp 0
transform 1 0 510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__598_
timestamp 0
transform 1 0 570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__599_
timestamp 0
transform 1 0 1130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__600_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__601_
timestamp 0
transform -1 0 530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__602_
timestamp 0
transform -1 0 790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__603_
timestamp 0
transform 1 0 1410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__604_
timestamp 0
transform 1 0 1570 0 1 250
box -6 -8 26 248
use FILL  FILL_0__605_
timestamp 0
transform 1 0 1030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__606_
timestamp 0
transform -1 0 1570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__607_
timestamp 0
transform 1 0 1550 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__608_
timestamp 0
transform 1 0 1050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__609_
timestamp 0
transform -1 0 1050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__610_
timestamp 0
transform 1 0 1270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__611_
timestamp 0
transform -1 0 1350 0 1 250
box -6 -8 26 248
use FILL  FILL_0__612_
timestamp 0
transform 1 0 1050 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__613_
timestamp 0
transform 1 0 1810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__614_
timestamp 0
transform 1 0 1810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__615_
timestamp 0
transform 1 0 2090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__616_
timestamp 0
transform 1 0 2330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__617_
timestamp 0
transform 1 0 2350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__618_
timestamp 0
transform 1 0 790 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__619_
timestamp 0
transform -1 0 290 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__620_
timestamp 0
transform 1 0 810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__621_
timestamp 0
transform -1 0 570 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__622_
timestamp 0
transform -1 0 790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__623_
timestamp 0
transform 1 0 1050 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__624_
timestamp 0
transform 1 0 270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__625_
timestamp 0
transform 1 0 270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__665_
timestamp 0
transform 1 0 3290 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__666_
timestamp 0
transform 1 0 2650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__667_
timestamp 0
transform -1 0 4210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__668_
timestamp 0
transform 1 0 1870 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 2590 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform 1 0 1330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 1070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform -1 0 1830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 1070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 2070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform -1 0 790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 2330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 3170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 1810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform 1 0 3090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform 1 0 1970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 1690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert0
timestamp 0
transform 1 0 1970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert1
timestamp 0
transform -1 0 1610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert2
timestamp 0
transform 1 0 10 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert3
timestamp 0
transform 1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert4
timestamp 0
transform 1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert5
timestamp 0
transform 1 0 1090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__313_
timestamp 0
transform 1 0 1070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__314_
timestamp 0
transform -1 0 1070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__315_
timestamp 0
transform 1 0 790 0 1 730
box -6 -8 26 248
use FILL  FILL_1__316_
timestamp 0
transform -1 0 890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__317_
timestamp 0
transform -1 0 2650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__318_
timestamp 0
transform 1 0 2890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__319_
timestamp 0
transform -1 0 3190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__320_
timestamp 0
transform -1 0 3130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__321_
timestamp 0
transform 1 0 3430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__322_
timestamp 0
transform 1 0 2850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__323_
timestamp 0
transform -1 0 2930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__324_
timestamp 0
transform -1 0 2610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__325_
timestamp 0
transform -1 0 3450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__326_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__327_
timestamp 0
transform 1 0 4710 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__328_
timestamp 0
transform 1 0 4230 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__329_
timestamp 0
transform -1 0 4490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__330_
timestamp 0
transform 1 0 3970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__331_
timestamp 0
transform -1 0 2930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__332_
timestamp 0
transform -1 0 2670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__333_
timestamp 0
transform 1 0 2110 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__334_
timestamp 0
transform 1 0 2090 0 1 250
box -6 -8 26 248
use FILL  FILL_1__335_
timestamp 0
transform -1 0 1850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__336_
timestamp 0
transform -1 0 3190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__337_
timestamp 0
transform 1 0 3430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__338_
timestamp 0
transform -1 0 4010 0 1 250
box -6 -8 26 248
use FILL  FILL_1__339_
timestamp 0
transform 1 0 3710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__340_
timestamp 0
transform 1 0 4210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__341_
timestamp 0
transform 1 0 4670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__342_
timestamp 0
transform 1 0 4750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__343_
timestamp 0
transform -1 0 4770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__344_
timestamp 0
transform -1 0 4510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__345_
timestamp 0
transform -1 0 4490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__346_
timestamp 0
transform 1 0 4170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__347_
timestamp 0
transform -1 0 3390 0 1 730
box -6 -8 26 248
use FILL  FILL_1__348_
timestamp 0
transform -1 0 3670 0 1 730
box -6 -8 26 248
use FILL  FILL_1__349_
timestamp 0
transform 1 0 4690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__350_
timestamp 0
transform 1 0 4430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__351_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__352_
timestamp 0
transform 1 0 4450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__353_
timestamp 0
transform 1 0 4130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__354_
timestamp 0
transform 1 0 3890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__355_
timestamp 0
transform 1 0 4390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__356_
timestamp 0
transform -1 0 4130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__357_
timestamp 0
transform -1 0 3590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__358_
timestamp 0
transform -1 0 3850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__359_
timestamp 0
transform -1 0 3450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__360_
timestamp 0
transform 1 0 3930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__361_
timestamp 0
transform 1 0 4190 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__362_
timestamp 0
transform -1 0 3930 0 1 730
box -6 -8 26 248
use FILL  FILL_1__363_
timestamp 0
transform -1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__364_
timestamp 0
transform -1 0 4390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__365_
timestamp 0
transform -1 0 3390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__366_
timestamp 0
transform -1 0 3450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__367_
timestamp 0
transform 1 0 3970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__368_
timestamp 0
transform 1 0 4490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__369_
timestamp 0
transform 1 0 3970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__370_
timestamp 0
transform 1 0 3670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__371_
timestamp 0
transform 1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__372_
timestamp 0
transform 1 0 3970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__373_
timestamp 0
transform -1 0 3710 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__374_
timestamp 0
transform -1 0 3730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__375_
timestamp 0
transform 1 0 3690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__376_
timestamp 0
transform 1 0 3210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__377_
timestamp 0
transform -1 0 2950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__378_
timestamp 0
transform 1 0 3430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__379_
timestamp 0
transform -1 0 3170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__380_
timestamp 0
transform -1 0 3450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__381_
timestamp 0
transform -1 0 3190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__382_
timestamp 0
transform 1 0 3150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__383_
timestamp 0
transform -1 0 2910 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__384_
timestamp 0
transform 1 0 3710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__385_
timestamp 0
transform -1 0 3470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__386_
timestamp 0
transform -1 0 2630 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__387_
timestamp 0
transform 1 0 2130 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__388_
timestamp 0
transform 1 0 2410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__389_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__390_
timestamp 0
transform -1 0 1830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__391_
timestamp 0
transform -1 0 2630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__392_
timestamp 0
transform -1 0 2370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__393_
timestamp 0
transform 1 0 1610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__394_
timestamp 0
transform -1 0 2090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__395_
timestamp 0
transform -1 0 1590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__396_
timestamp 0
transform 1 0 2150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__397_
timestamp 0
transform 1 0 2650 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__398_
timestamp 0
transform 1 0 2130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__399_
timestamp 0
transform 1 0 2410 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__400_
timestamp 0
transform -1 0 1810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__401_
timestamp 0
transform -1 0 2090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__402_
timestamp 0
transform -1 0 1910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__403_
timestamp 0
transform 1 0 2330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__404_
timestamp 0
transform -1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__405_
timestamp 0
transform 1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__406_
timestamp 0
transform -1 0 1530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__407_
timestamp 0
transform 1 0 3170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__408_
timestamp 0
transform -1 0 2890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__409_
timestamp 0
transform 1 0 3550 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__410_
timestamp 0
transform -1 0 3670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__411_
timestamp 0
transform -1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__412_
timestamp 0
transform 1 0 2590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__413_
timestamp 0
transform -1 0 2910 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__414_
timestamp 0
transform 1 0 2390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__415_
timestamp 0
transform 1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__416_
timestamp 0
transform 1 0 3670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__417_
timestamp 0
transform -1 0 3830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__418_
timestamp 0
transform 1 0 4710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__419_
timestamp 0
transform 1 0 4450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__420_
timestamp 0
transform -1 0 4110 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__421_
timestamp 0
transform -1 0 3930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__422_
timestamp 0
transform -1 0 1590 0 1 730
box -6 -8 26 248
use FILL  FILL_1__423_
timestamp 0
transform 1 0 1330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__424_
timestamp 0
transform 1 0 1290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__425_
timestamp 0
transform 1 0 1330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__426_
timestamp 0
transform -1 0 3310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__427_
timestamp 0
transform -1 0 2670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__428_
timestamp 0
transform -1 0 3050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__429_
timestamp 0
transform 1 0 3150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__430_
timestamp 0
transform -1 0 3830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__431_
timestamp 0
transform 1 0 3910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__432_
timestamp 0
transform -1 0 3390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__433_
timestamp 0
transform -1 0 3650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__434_
timestamp 0
transform 1 0 4170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__435_
timestamp 0
transform 1 0 4650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__436_
timestamp 0
transform 1 0 4750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__437_
timestamp 0
transform -1 0 4730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__438_
timestamp 0
transform -1 0 4210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__439_
timestamp 0
transform -1 0 4190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__440_
timestamp 0
transform -1 0 3390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__441_
timestamp 0
transform -1 0 3930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__442_
timestamp 0
transform -1 0 4370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__443_
timestamp 0
transform 1 0 4590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__444_
timestamp 0
transform -1 0 4230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__445_
timestamp 0
transform -1 0 4730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__446_
timestamp 0
transform 1 0 4690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__447_
timestamp 0
transform 1 0 4750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__448_
timestamp 0
transform -1 0 4530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__449_
timestamp 0
transform 1 0 4090 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__450_
timestamp 0
transform 1 0 4490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__451_
timestamp 0
transform 1 0 4730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__452_
timestamp 0
transform 1 0 4610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__453_
timestamp 0
transform 1 0 4770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__454_
timestamp 0
transform 1 0 4250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__455_
timestamp 0
transform -1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__456_
timestamp 0
transform -1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__457_
timestamp 0
transform 1 0 3970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__458_
timestamp 0
transform -1 0 3710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__459_
timestamp 0
transform -1 0 4710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__460_
timestamp 0
transform 1 0 4770 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__461_
timestamp 0
transform 1 0 4470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__462_
timestamp 0
transform 1 0 4710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__463_
timestamp 0
transform 1 0 4770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__464_
timestamp 0
transform 1 0 4190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__465_
timestamp 0
transform 1 0 4350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__466_
timestamp 0
transform 1 0 4450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__467_
timestamp 0
transform 1 0 4490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__468_
timestamp 0
transform 1 0 4190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__469_
timestamp 0
transform -1 0 2890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__470_
timestamp 0
transform -1 0 2350 0 1 730
box -6 -8 26 248
use FILL  FILL_1__471_
timestamp 0
transform -1 0 2550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__472_
timestamp 0
transform 1 0 2070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__473_
timestamp 0
transform 1 0 2370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__474_
timestamp 0
transform 1 0 2650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__475_
timestamp 0
transform 1 0 3310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__476_
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__477_
timestamp 0
transform -1 0 2270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__478_
timestamp 0
transform -1 0 2150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__479_
timestamp 0
transform -1 0 3210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__480_
timestamp 0
transform 1 0 3150 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__481_
timestamp 0
transform -1 0 2650 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__482_
timestamp 0
transform 1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__483_
timestamp 0
transform -1 0 1310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__484_
timestamp 0
transform -1 0 1030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__485_
timestamp 0
transform -1 0 1630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__486_
timestamp 0
transform -1 0 1610 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__487_
timestamp 0
transform -1 0 1350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__488_
timestamp 0
transform -1 0 1070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__489_
timestamp 0
transform -1 0 1890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__490_
timestamp 0
transform 1 0 1590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__491_
timestamp 0
transform 1 0 2690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__492_
timestamp 0
transform -1 0 3450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__493_
timestamp 0
transform 1 0 2950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__494_
timestamp 0
transform 1 0 2910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__495_
timestamp 0
transform 1 0 2090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__496_
timestamp 0
transform 1 0 770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__497_
timestamp 0
transform -1 0 1550 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__498_
timestamp 0
transform 1 0 910 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__499_
timestamp 0
transform 1 0 1290 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__500_
timestamp 0
transform -1 0 1790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__501_
timestamp 0
transform 1 0 1130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__502_
timestamp 0
transform -1 0 1350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__503_
timestamp 0
transform 1 0 1590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__504_
timestamp 0
transform -1 0 2630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__505_
timestamp 0
transform -1 0 2890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__506_
timestamp 0
transform 1 0 3130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__507_
timestamp 0
transform 1 0 2870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__508_
timestamp 0
transform -1 0 2770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__509_
timestamp 0
transform 1 0 3110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__510_
timestamp 0
transform 1 0 3030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__511_
timestamp 0
transform 1 0 2510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__512_
timestamp 0
transform 1 0 1610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__513_
timestamp 0
transform -1 0 1430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__514_
timestamp 0
transform 1 0 1470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__515_
timestamp 0
transform 1 0 1850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__516_
timestamp 0
transform 1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__517_
timestamp 0
transform -1 0 1990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__518_
timestamp 0
transform -1 0 2690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__519_
timestamp 0
transform 1 0 2410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__520_
timestamp 0
transform 1 0 2330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__521_
timestamp 0
transform 1 0 2610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__522_
timestamp 0
transform -1 0 2630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__523_
timestamp 0
transform 1 0 2210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__524_
timestamp 0
transform 1 0 4250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__525_
timestamp 0
transform -1 0 4530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__526_
timestamp 0
transform -1 0 4510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__527_
timestamp 0
transform -1 0 4450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__528_
timestamp 0
transform -1 0 4190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__529_
timestamp 0
transform -1 0 4250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__530_
timestamp 0
transform 1 0 4210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__531_
timestamp 0
transform -1 0 1730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__532_
timestamp 0
transform -1 0 850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__533_
timestamp 0
transform -1 0 3730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__534_
timestamp 0
transform -1 0 3170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__535_
timestamp 0
transform -1 0 2490 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__536_
timestamp 0
transform 1 0 2130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__537_
timestamp 0
transform -1 0 1090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__538_
timestamp 0
transform 1 0 1870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__539_
timestamp 0
transform 1 0 2370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__540_
timestamp 0
transform 1 0 810 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__541_
timestamp 0
transform 1 0 1030 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__542_
timestamp 0
transform 1 0 1310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__543_
timestamp 0
transform -1 0 1050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__544_
timestamp 0
transform -1 0 570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__545_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__546_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__547_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__548_
timestamp 0
transform -1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__549_
timestamp 0
transform -1 0 290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__550_
timestamp 0
transform -1 0 570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__551_
timestamp 0
transform 1 0 570 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__552_
timestamp 0
transform 1 0 810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__553_
timestamp 0
transform 1 0 1070 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__554_
timestamp 0
transform 1 0 1350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__555_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__556_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__557_
timestamp 0
transform -1 0 50 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__558_
timestamp 0
transform 1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__559_
timestamp 0
transform -1 0 50 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__560_
timestamp 0
transform -1 0 850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__561_
timestamp 0
transform 1 0 550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__562_
timestamp 0
transform 1 0 850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__563_
timestamp 0
transform -1 0 590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__564_
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__565_
timestamp 0
transform 1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__566_
timestamp 0
transform 1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__567_
timestamp 0
transform 1 0 310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__568_
timestamp 0
transform -1 0 590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__569_
timestamp 0
transform -1 0 850 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__570_
timestamp 0
transform 1 0 810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__571_
timestamp 0
transform -1 0 570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__572_
timestamp 0
transform -1 0 290 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__573_
timestamp 0
transform 1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__574_
timestamp 0
transform -1 0 310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__575_
timestamp 0
transform 1 0 530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__576_
timestamp 0
transform 1 0 550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__577_
timestamp 0
transform -1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__578_
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__579_
timestamp 0
transform 1 0 530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__580_
timestamp 0
transform -1 0 310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__581_
timestamp 0
transform -1 0 290 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__582_
timestamp 0
transform 1 0 790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__583_
timestamp 0
transform -1 0 570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__584_
timestamp 0
transform 1 0 390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__585_
timestamp 0
transform -1 0 530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__586_
timestamp 0
transform -1 0 330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__587_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__588_
timestamp 0
transform -1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_1__589_
timestamp 0
transform -1 0 50 0 1 730
box -6 -8 26 248
use FILL  FILL_1__590_
timestamp 0
transform -1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__591_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__592_
timestamp 0
transform -1 0 610 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__593_
timestamp 0
transform 1 0 310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__594_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__595_
timestamp 0
transform -1 0 310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__596_
timestamp 0
transform 1 0 550 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__597_
timestamp 0
transform 1 0 530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__598_
timestamp 0
transform 1 0 590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__599_
timestamp 0
transform 1 0 1150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__600_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__601_
timestamp 0
transform -1 0 550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__602_
timestamp 0
transform -1 0 810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__603_
timestamp 0
transform 1 0 1430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__604_
timestamp 0
transform 1 0 1590 0 1 250
box -6 -8 26 248
use FILL  FILL_1__605_
timestamp 0
transform 1 0 1050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__606_
timestamp 0
transform -1 0 1590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__607_
timestamp 0
transform 1 0 1570 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__608_
timestamp 0
transform 1 0 1070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__609_
timestamp 0
transform -1 0 1070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__610_
timestamp 0
transform 1 0 1290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__611_
timestamp 0
transform -1 0 1370 0 1 250
box -6 -8 26 248
use FILL  FILL_1__612_
timestamp 0
transform 1 0 1070 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__613_
timestamp 0
transform 1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__614_
timestamp 0
transform 1 0 1830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__615_
timestamp 0
transform 1 0 2110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__616_
timestamp 0
transform 1 0 2350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__617_
timestamp 0
transform 1 0 2370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__618_
timestamp 0
transform 1 0 810 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__619_
timestamp 0
transform -1 0 310 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__620_
timestamp 0
transform 1 0 830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__621_
timestamp 0
transform -1 0 590 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__622_
timestamp 0
transform -1 0 810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__623_
timestamp 0
transform 1 0 1070 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__624_
timestamp 0
transform 1 0 290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__625_
timestamp 0
transform 1 0 290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__665_
timestamp 0
transform 1 0 3310 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__666_
timestamp 0
transform 1 0 2670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__667_
timestamp 0
transform -1 0 4230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__668_
timestamp 0
transform 1 0 1890 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 2610 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform 1 0 1350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 1090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform -1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 1090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 2090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform -1 0 810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 2350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 3190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 1830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform 1 0 3110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform 1 0 1990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 1710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert0
timestamp 0
transform 1 0 1990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert1
timestamp 0
transform -1 0 1630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert2
timestamp 0
transform 1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert3
timestamp 0
transform 1 0 1770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert4
timestamp 0
transform 1 0 1090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert5
timestamp 0
transform 1 0 1110 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__313_
timestamp 0
transform 1 0 1090 0 1 250
box -6 -8 26 248
use FILL  FILL_2__314_
timestamp 0
transform -1 0 1090 0 1 730
box -6 -8 26 248
use FILL  FILL_2__315_
timestamp 0
transform 1 0 810 0 1 730
box -6 -8 26 248
use FILL  FILL_2__316_
timestamp 0
transform -1 0 910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__317_
timestamp 0
transform -1 0 2670 0 1 250
box -6 -8 26 248
use FILL  FILL_2__318_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 26 248
use FILL  FILL_2__319_
timestamp 0
transform -1 0 3210 0 1 250
box -6 -8 26 248
use FILL  FILL_2__320_
timestamp 0
transform -1 0 3150 0 1 730
box -6 -8 26 248
use FILL  FILL_2__321_
timestamp 0
transform 1 0 3450 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__322_
timestamp 0
transform 1 0 2870 0 1 730
box -6 -8 26 248
use FILL  FILL_2__323_
timestamp 0
transform -1 0 2950 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__324_
timestamp 0
transform -1 0 2630 0 1 730
box -6 -8 26 248
use FILL  FILL_2__325_
timestamp 0
transform -1 0 3470 0 1 250
box -6 -8 26 248
use FILL  FILL_2__326_
timestamp 0
transform -1 0 3750 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__327_
timestamp 0
transform 1 0 4730 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__328_
timestamp 0
transform 1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__329_
timestamp 0
transform -1 0 4510 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__330_
timestamp 0
transform 1 0 3990 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__331_
timestamp 0
transform -1 0 2950 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__332_
timestamp 0
transform -1 0 2690 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__333_
timestamp 0
transform 1 0 2130 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__334_
timestamp 0
transform 1 0 2110 0 1 250
box -6 -8 26 248
use FILL  FILL_2__335_
timestamp 0
transform -1 0 1870 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__336_
timestamp 0
transform -1 0 3210 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__337_
timestamp 0
transform 1 0 3450 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__338_
timestamp 0
transform -1 0 4030 0 1 250
box -6 -8 26 248
use FILL  FILL_2__339_
timestamp 0
transform 1 0 3730 0 1 250
box -6 -8 26 248
use FILL  FILL_2__340_
timestamp 0
transform 1 0 4230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__341_
timestamp 0
transform 1 0 4690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__342_
timestamp 0
transform 1 0 4770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__343_
timestamp 0
transform -1 0 4790 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__344_
timestamp 0
transform -1 0 4530 0 1 250
box -6 -8 26 248
use FILL  FILL_2__345_
timestamp 0
transform -1 0 4510 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__346_
timestamp 0
transform 1 0 4190 0 1 730
box -6 -8 26 248
use FILL  FILL_2__347_
timestamp 0
transform -1 0 3410 0 1 730
box -6 -8 26 248
use FILL  FILL_2__348_
timestamp 0
transform -1 0 3690 0 1 730
box -6 -8 26 248
use FILL  FILL_2__349_
timestamp 0
transform 1 0 4710 0 1 730
box -6 -8 26 248
use FILL  FILL_2__350_
timestamp 0
transform 1 0 4450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__351_
timestamp 0
transform 1 0 4490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__352_
timestamp 0
transform 1 0 4470 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__353_
timestamp 0
transform 1 0 4150 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__354_
timestamp 0
transform 1 0 3910 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__355_
timestamp 0
transform 1 0 4410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__356_
timestamp 0
transform -1 0 4150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__357_
timestamp 0
transform -1 0 3610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__358_
timestamp 0
transform -1 0 3870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__359_
timestamp 0
transform -1 0 3470 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__360_
timestamp 0
transform 1 0 3950 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__361_
timestamp 0
transform 1 0 4210 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__362_
timestamp 0
transform -1 0 3950 0 1 730
box -6 -8 26 248
use FILL  FILL_2__363_
timestamp 0
transform -1 0 4910 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__364_
timestamp 0
transform -1 0 4410 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__365_
timestamp 0
transform -1 0 3410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__366_
timestamp 0
transform -1 0 3470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__367_
timestamp 0
transform 1 0 3990 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__368_
timestamp 0
transform 1 0 4510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__369_
timestamp 0
transform 1 0 3990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__370_
timestamp 0
transform 1 0 3690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__371_
timestamp 0
transform 1 0 3970 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__372_
timestamp 0
transform 1 0 3990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__373_
timestamp 0
transform -1 0 3730 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__374_
timestamp 0
transform -1 0 3750 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__375_
timestamp 0
transform 1 0 3710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__376_
timestamp 0
transform 1 0 3230 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__377_
timestamp 0
transform -1 0 2970 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__378_
timestamp 0
transform 1 0 3450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__379_
timestamp 0
transform -1 0 3190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__380_
timestamp 0
transform -1 0 3470 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__381_
timestamp 0
transform -1 0 3210 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__382_
timestamp 0
transform 1 0 3170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__383_
timestamp 0
transform -1 0 2930 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__384_
timestamp 0
transform 1 0 3730 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__385_
timestamp 0
transform -1 0 3490 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__386_
timestamp 0
transform -1 0 2650 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__387_
timestamp 0
transform 1 0 2150 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__388_
timestamp 0
transform 1 0 2430 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__389_
timestamp 0
transform -1 0 2930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__390_
timestamp 0
transform -1 0 1850 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__391_
timestamp 0
transform -1 0 2650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__392_
timestamp 0
transform -1 0 2390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__393_
timestamp 0
transform 1 0 1630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__394_
timestamp 0
transform -1 0 2110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__395_
timestamp 0
transform -1 0 1610 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__396_
timestamp 0
transform 1 0 2170 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__397_
timestamp 0
transform 1 0 2670 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__398_
timestamp 0
transform 1 0 2150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__399_
timestamp 0
transform 1 0 2430 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__400_
timestamp 0
transform -1 0 1830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__401_
timestamp 0
transform -1 0 2110 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__402_
timestamp 0
transform -1 0 1930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__403_
timestamp 0
transform 1 0 2350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__404_
timestamp 0
transform -1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__405_
timestamp 0
transform 1 0 1510 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__406_
timestamp 0
transform -1 0 1550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__407_
timestamp 0
transform 1 0 3190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__408_
timestamp 0
transform -1 0 2910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__409_
timestamp 0
transform 1 0 3570 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__410_
timestamp 0
transform -1 0 3690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__411_
timestamp 0
transform -1 0 2390 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__412_
timestamp 0
transform 1 0 2610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__413_
timestamp 0
transform -1 0 2930 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__414_
timestamp 0
transform 1 0 2410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__415_
timestamp 0
transform 1 0 2950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__416_
timestamp 0
transform 1 0 3690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__417_
timestamp 0
transform -1 0 3850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__418_
timestamp 0
transform 1 0 4730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__419_
timestamp 0
transform 1 0 4470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__420_
timestamp 0
transform -1 0 4130 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__421_
timestamp 0
transform -1 0 3950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__422_
timestamp 0
transform -1 0 1610 0 1 730
box -6 -8 26 248
use FILL  FILL_2__423_
timestamp 0
transform 1 0 1350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__424_
timestamp 0
transform 1 0 1310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__425_
timestamp 0
transform 1 0 1350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__426_
timestamp 0
transform -1 0 3330 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__427_
timestamp 0
transform -1 0 2690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__428_
timestamp 0
transform -1 0 3070 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__429_
timestamp 0
transform 1 0 3170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__430_
timestamp 0
transform -1 0 3850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__431_
timestamp 0
transform 1 0 3930 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__432_
timestamp 0
transform -1 0 3410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__433_
timestamp 0
transform -1 0 3670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__434_
timestamp 0
transform 1 0 4190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__435_
timestamp 0
transform 1 0 4670 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__436_
timestamp 0
transform 1 0 4770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__437_
timestamp 0
transform -1 0 4750 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__438_
timestamp 0
transform -1 0 4230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__439_
timestamp 0
transform -1 0 4210 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__440_
timestamp 0
transform -1 0 3410 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__441_
timestamp 0
transform -1 0 3950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__442_
timestamp 0
transform -1 0 4390 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__443_
timestamp 0
transform 1 0 4610 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__444_
timestamp 0
transform -1 0 4250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__445_
timestamp 0
transform -1 0 4750 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__446_
timestamp 0
transform 1 0 4710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__447_
timestamp 0
transform 1 0 4770 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__448_
timestamp 0
transform -1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__449_
timestamp 0
transform 1 0 4110 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__450_
timestamp 0
transform 1 0 4510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__451_
timestamp 0
transform 1 0 4750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__452_
timestamp 0
transform 1 0 4630 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__453_
timestamp 0
transform 1 0 4790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__454_
timestamp 0
transform 1 0 4270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__455_
timestamp 0
transform -1 0 3750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__456_
timestamp 0
transform -1 0 4030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__457_
timestamp 0
transform 1 0 3990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__458_
timestamp 0
transform -1 0 3730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__459_
timestamp 0
transform -1 0 4730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__460_
timestamp 0
transform 1 0 4790 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__461_
timestamp 0
transform 1 0 4490 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__462_
timestamp 0
transform 1 0 4730 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__463_
timestamp 0
transform 1 0 4790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__464_
timestamp 0
transform 1 0 4210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__465_
timestamp 0
transform 1 0 4370 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__466_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__467_
timestamp 0
transform 1 0 4510 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__468_
timestamp 0
transform 1 0 4210 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__469_
timestamp 0
transform -1 0 2910 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__470_
timestamp 0
transform -1 0 2370 0 1 730
box -6 -8 26 248
use FILL  FILL_2__471_
timestamp 0
transform -1 0 2570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__472_
timestamp 0
transform 1 0 2090 0 1 730
box -6 -8 26 248
use FILL  FILL_2__473_
timestamp 0
transform 1 0 2390 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__474_
timestamp 0
transform 1 0 2670 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__475_
timestamp 0
transform 1 0 3330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__476_
timestamp 0
transform 1 0 2810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__477_
timestamp 0
transform -1 0 2290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__478_
timestamp 0
transform -1 0 2170 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__479_
timestamp 0
transform -1 0 3230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__480_
timestamp 0
transform 1 0 3170 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__481_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__482_
timestamp 0
transform 1 0 2770 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__483_
timestamp 0
transform -1 0 1330 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__484_
timestamp 0
transform -1 0 1050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__485_
timestamp 0
transform -1 0 1650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__486_
timestamp 0
transform -1 0 1630 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__487_
timestamp 0
transform -1 0 1370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__488_
timestamp 0
transform -1 0 1090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__489_
timestamp 0
transform -1 0 1910 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__490_
timestamp 0
transform 1 0 1610 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__491_
timestamp 0
transform 1 0 2710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__492_
timestamp 0
transform -1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__493_
timestamp 0
transform 1 0 2970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__494_
timestamp 0
transform 1 0 2930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__495_
timestamp 0
transform 1 0 2110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__496_
timestamp 0
transform 1 0 790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__497_
timestamp 0
transform -1 0 1570 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__498_
timestamp 0
transform 1 0 930 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__499_
timestamp 0
transform 1 0 1310 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__500_
timestamp 0
transform -1 0 1810 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__501_
timestamp 0
transform 1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__502_
timestamp 0
transform -1 0 1370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__503_
timestamp 0
transform 1 0 1610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__504_
timestamp 0
transform -1 0 2650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__505_
timestamp 0
transform -1 0 2910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__506_
timestamp 0
transform 1 0 3150 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__507_
timestamp 0
transform 1 0 2890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__508_
timestamp 0
transform -1 0 2790 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__509_
timestamp 0
transform 1 0 3130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__510_
timestamp 0
transform 1 0 3050 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__511_
timestamp 0
transform 1 0 2530 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__512_
timestamp 0
transform 1 0 1630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__513_
timestamp 0
transform -1 0 1450 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__514_
timestamp 0
transform 1 0 1490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__515_
timestamp 0
transform 1 0 1870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__516_
timestamp 0
transform 1 0 1710 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__517_
timestamp 0
transform -1 0 2010 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__518_
timestamp 0
transform -1 0 2710 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__519_
timestamp 0
transform 1 0 2430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__520_
timestamp 0
transform 1 0 2350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__521_
timestamp 0
transform 1 0 2630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__522_
timestamp 0
transform -1 0 2650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__523_
timestamp 0
transform 1 0 2230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__524_
timestamp 0
transform 1 0 4270 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__525_
timestamp 0
transform -1 0 4550 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__526_
timestamp 0
transform -1 0 4530 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__527_
timestamp 0
transform -1 0 4470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__528_
timestamp 0
transform -1 0 4210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__529_
timestamp 0
transform -1 0 4270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__530_
timestamp 0
transform 1 0 4230 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__531_
timestamp 0
transform -1 0 1750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__532_
timestamp 0
transform -1 0 870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__533_
timestamp 0
transform -1 0 3750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__534_
timestamp 0
transform -1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__535_
timestamp 0
transform -1 0 2510 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__536_
timestamp 0
transform 1 0 2150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__537_
timestamp 0
transform -1 0 1110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__538_
timestamp 0
transform 1 0 1890 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__539_
timestamp 0
transform 1 0 2390 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__540_
timestamp 0
transform 1 0 830 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__541_
timestamp 0
transform 1 0 1050 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__542_
timestamp 0
transform 1 0 1330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__543_
timestamp 0
transform -1 0 1070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__544_
timestamp 0
transform -1 0 590 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__545_
timestamp 0
transform -1 0 70 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__546_
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__547_
timestamp 0
transform -1 0 70 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__548_
timestamp 0
transform -1 0 330 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__549_
timestamp 0
transform -1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__550_
timestamp 0
transform -1 0 590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__551_
timestamp 0
transform 1 0 590 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__552_
timestamp 0
transform 1 0 830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__553_
timestamp 0
transform 1 0 1090 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__554_
timestamp 0
transform 1 0 1370 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__555_
timestamp 0
transform -1 0 310 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__556_
timestamp 0
transform -1 0 70 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__557_
timestamp 0
transform -1 0 70 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__558_
timestamp 0
transform 1 0 330 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__559_
timestamp 0
transform -1 0 70 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__560_
timestamp 0
transform -1 0 870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__561_
timestamp 0
transform 1 0 570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__562_
timestamp 0
transform 1 0 870 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__563_
timestamp 0
transform -1 0 610 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__564_
timestamp 0
transform -1 0 70 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__565_
timestamp 0
transform 1 0 50 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__566_
timestamp 0
transform 1 0 50 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__567_
timestamp 0
transform 1 0 330 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__568_
timestamp 0
transform -1 0 610 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__569_
timestamp 0
transform -1 0 870 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__570_
timestamp 0
transform 1 0 830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__571_
timestamp 0
transform -1 0 590 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__572_
timestamp 0
transform -1 0 310 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__573_
timestamp 0
transform 1 0 310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__574_
timestamp 0
transform -1 0 330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__575_
timestamp 0
transform 1 0 550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__576_
timestamp 0
transform 1 0 570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__577_
timestamp 0
transform -1 0 70 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__578_
timestamp 0
transform -1 0 70 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__579_
timestamp 0
transform 1 0 550 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__580_
timestamp 0
transform -1 0 330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__581_
timestamp 0
transform -1 0 310 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__582_
timestamp 0
transform 1 0 810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__583_
timestamp 0
transform -1 0 590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__584_
timestamp 0
transform 1 0 410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__585_
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__586_
timestamp 0
transform -1 0 350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__587_
timestamp 0
transform -1 0 70 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__588_
timestamp 0
transform -1 0 70 0 1 250
box -6 -8 26 248
use FILL  FILL_2__589_
timestamp 0
transform -1 0 70 0 1 730
box -6 -8 26 248
use FILL  FILL_2__590_
timestamp 0
transform -1 0 70 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__591_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__592_
timestamp 0
transform -1 0 630 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__593_
timestamp 0
transform 1 0 330 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__594_
timestamp 0
transform -1 0 70 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__595_
timestamp 0
transform -1 0 330 0 1 730
box -6 -8 26 248
use FILL  FILL_2__596_
timestamp 0
transform 1 0 570 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__597_
timestamp 0
transform 1 0 550 0 1 730
box -6 -8 26 248
use FILL  FILL_2__598_
timestamp 0
transform 1 0 610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__599_
timestamp 0
transform 1 0 1170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__600_
timestamp 0
transform -1 0 70 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__601_
timestamp 0
transform -1 0 570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__602_
timestamp 0
transform -1 0 830 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__603_
timestamp 0
transform 1 0 1450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__604_
timestamp 0
transform 1 0 1610 0 1 250
box -6 -8 26 248
use FILL  FILL_2__605_
timestamp 0
transform 1 0 1070 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__606_
timestamp 0
transform -1 0 1610 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__607_
timestamp 0
transform 1 0 1590 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__608_
timestamp 0
transform 1 0 1090 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__609_
timestamp 0
transform -1 0 1090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__610_
timestamp 0
transform 1 0 1310 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__611_
timestamp 0
transform -1 0 1390 0 1 250
box -6 -8 26 248
use FILL  FILL_2__612_
timestamp 0
transform 1 0 1090 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__613_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__614_
timestamp 0
transform 1 0 1850 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__615_
timestamp 0
transform 1 0 2130 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__616_
timestamp 0
transform 1 0 2370 0 1 250
box -6 -8 26 248
use FILL  FILL_2__617_
timestamp 0
transform 1 0 2390 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__618_
timestamp 0
transform 1 0 830 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__619_
timestamp 0
transform -1 0 330 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__620_
timestamp 0
transform 1 0 850 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__621_
timestamp 0
transform -1 0 610 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__622_
timestamp 0
transform -1 0 830 0 1 250
box -6 -8 26 248
use FILL  FILL_2__623_
timestamp 0
transform 1 0 1090 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__624_
timestamp 0
transform 1 0 310 0 1 250
box -6 -8 26 248
use FILL  FILL_2__625_
timestamp 0
transform 1 0 310 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__665_
timestamp 0
transform 1 0 3330 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__666_
timestamp 0
transform 1 0 2690 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__667_
timestamp 0
transform -1 0 4250 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__668_
timestamp 0
transform 1 0 1910 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform -1 0 850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform 1 0 2630 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform 1 0 1370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert9
timestamp 0
transform 1 0 1110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform -1 0 1870 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform 1 0 2390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 1110 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 2110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform -1 0 830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 2370 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 3210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 1850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform 1 0 3130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform 1 0 2010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 1730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert0
timestamp 0
transform 1 0 2010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert1
timestamp 0
transform -1 0 1650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert2
timestamp 0
transform 1 0 50 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert3
timestamp 0
transform 1 0 1790 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert4
timestamp 0
transform 1 0 1110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert5
timestamp 0
transform 1 0 1130 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__313_
timestamp 0
transform 1 0 1110 0 1 250
box -6 -8 26 248
use FILL  FILL_3__314_
timestamp 0
transform -1 0 1110 0 1 730
box -6 -8 26 248
use FILL  FILL_3__315_
timestamp 0
transform 1 0 830 0 1 730
box -6 -8 26 248
use FILL  FILL_3__316_
timestamp 0
transform -1 0 930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__317_
timestamp 0
transform -1 0 2690 0 1 250
box -6 -8 26 248
use FILL  FILL_3__318_
timestamp 0
transform 1 0 2930 0 1 250
box -6 -8 26 248
use FILL  FILL_3__319_
timestamp 0
transform -1 0 3230 0 1 250
box -6 -8 26 248
use FILL  FILL_3__320_
timestamp 0
transform -1 0 3170 0 1 730
box -6 -8 26 248
use FILL  FILL_3__321_
timestamp 0
transform 1 0 3470 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__322_
timestamp 0
transform 1 0 2890 0 1 730
box -6 -8 26 248
use FILL  FILL_3__323_
timestamp 0
transform -1 0 2970 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__324_
timestamp 0
transform -1 0 2650 0 1 730
box -6 -8 26 248
use FILL  FILL_3__325_
timestamp 0
transform -1 0 3490 0 1 250
box -6 -8 26 248
use FILL  FILL_3__326_
timestamp 0
transform -1 0 3770 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__327_
timestamp 0
transform 1 0 4750 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__328_
timestamp 0
transform 1 0 4270 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__329_
timestamp 0
transform -1 0 4530 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__330_
timestamp 0
transform 1 0 4010 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__331_
timestamp 0
transform -1 0 2970 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__332_
timestamp 0
transform -1 0 2710 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__333_
timestamp 0
transform 1 0 2150 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__334_
timestamp 0
transform 1 0 2130 0 1 250
box -6 -8 26 248
use FILL  FILL_3__335_
timestamp 0
transform -1 0 1890 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__336_
timestamp 0
transform -1 0 3230 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__337_
timestamp 0
transform 1 0 3470 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__338_
timestamp 0
transform -1 0 4050 0 1 250
box -6 -8 26 248
use FILL  FILL_3__339_
timestamp 0
transform 1 0 3750 0 1 250
box -6 -8 26 248
use FILL  FILL_3__340_
timestamp 0
transform 1 0 4250 0 1 250
box -6 -8 26 248
use FILL  FILL_3__341_
timestamp 0
transform 1 0 4710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__342_
timestamp 0
transform 1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__343_
timestamp 0
transform -1 0 4810 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__344_
timestamp 0
transform -1 0 4550 0 1 250
box -6 -8 26 248
use FILL  FILL_3__345_
timestamp 0
transform -1 0 4530 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__346_
timestamp 0
transform 1 0 4210 0 1 730
box -6 -8 26 248
use FILL  FILL_3__347_
timestamp 0
transform -1 0 3430 0 1 730
box -6 -8 26 248
use FILL  FILL_3__348_
timestamp 0
transform -1 0 3710 0 1 730
box -6 -8 26 248
use FILL  FILL_3__349_
timestamp 0
transform 1 0 4730 0 1 730
box -6 -8 26 248
use FILL  FILL_3__350_
timestamp 0
transform 1 0 4470 0 1 730
box -6 -8 26 248
use FILL  FILL_3__351_
timestamp 0
transform 1 0 4510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__352_
timestamp 0
transform 1 0 4490 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__353_
timestamp 0
transform 1 0 4170 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__354_
timestamp 0
transform 1 0 3930 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__355_
timestamp 0
transform 1 0 4430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__356_
timestamp 0
transform -1 0 4170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__357_
timestamp 0
transform -1 0 3630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__358_
timestamp 0
transform -1 0 3890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__359_
timestamp 0
transform -1 0 3490 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__360_
timestamp 0
transform 1 0 3970 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__361_
timestamp 0
transform 1 0 4230 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__362_
timestamp 0
transform -1 0 3970 0 1 730
box -6 -8 26 248
use FILL  FILL_3__363_
timestamp 0
transform -1 0 4930 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__364_
timestamp 0
transform -1 0 4430 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__365_
timestamp 0
transform -1 0 3430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__366_
timestamp 0
transform -1 0 3490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__367_
timestamp 0
transform 1 0 4010 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__368_
timestamp 0
transform 1 0 4530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__369_
timestamp 0
transform 1 0 4010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__370_
timestamp 0
transform 1 0 3710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__371_
timestamp 0
transform 1 0 3990 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__372_
timestamp 0
transform 1 0 4010 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__373_
timestamp 0
transform -1 0 3750 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__374_
timestamp 0
transform -1 0 3770 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__375_
timestamp 0
transform 1 0 3730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__376_
timestamp 0
transform 1 0 3250 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__377_
timestamp 0
transform -1 0 2990 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__378_
timestamp 0
transform 1 0 3470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__379_
timestamp 0
transform -1 0 3210 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__380_
timestamp 0
transform -1 0 3490 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__381_
timestamp 0
transform -1 0 3230 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__382_
timestamp 0
transform 1 0 3190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__383_
timestamp 0
transform -1 0 2950 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__384_
timestamp 0
transform 1 0 3750 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__385_
timestamp 0
transform -1 0 3510 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__386_
timestamp 0
transform -1 0 2670 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__387_
timestamp 0
transform 1 0 2170 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__388_
timestamp 0
transform 1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__389_
timestamp 0
transform -1 0 2950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__390_
timestamp 0
transform -1 0 1870 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__391_
timestamp 0
transform -1 0 2670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__392_
timestamp 0
transform -1 0 2410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__393_
timestamp 0
transform 1 0 1650 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__394_
timestamp 0
transform -1 0 2130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__395_
timestamp 0
transform -1 0 1630 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__396_
timestamp 0
transform 1 0 2190 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__397_
timestamp 0
transform 1 0 2690 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__398_
timestamp 0
transform 1 0 2170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__399_
timestamp 0
transform 1 0 2450 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__400_
timestamp 0
transform -1 0 1850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__401_
timestamp 0
transform -1 0 2130 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__402_
timestamp 0
transform -1 0 1950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__403_
timestamp 0
transform 1 0 2370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__404_
timestamp 0
transform -1 0 2130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__405_
timestamp 0
transform 1 0 1530 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__406_
timestamp 0
transform -1 0 1570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__407_
timestamp 0
transform 1 0 3210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__408_
timestamp 0
transform -1 0 2930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__409_
timestamp 0
transform 1 0 3590 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__410_
timestamp 0
transform -1 0 3710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__411_
timestamp 0
transform -1 0 2410 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__412_
timestamp 0
transform 1 0 2630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__413_
timestamp 0
transform -1 0 2950 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__414_
timestamp 0
transform 1 0 2430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__415_
timestamp 0
transform 1 0 2970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__416_
timestamp 0
transform 1 0 3710 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__417_
timestamp 0
transform -1 0 3870 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__418_
timestamp 0
transform 1 0 4750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__419_
timestamp 0
transform 1 0 4490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__420_
timestamp 0
transform -1 0 4150 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__421_
timestamp 0
transform -1 0 3970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__422_
timestamp 0
transform -1 0 1630 0 1 730
box -6 -8 26 248
use FILL  FILL_3__423_
timestamp 0
transform 1 0 1370 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__424_
timestamp 0
transform 1 0 1330 0 1 730
box -6 -8 26 248
use FILL  FILL_3__425_
timestamp 0
transform 1 0 1370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__426_
timestamp 0
transform -1 0 3350 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__427_
timestamp 0
transform -1 0 2710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__428_
timestamp 0
transform -1 0 3090 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__429_
timestamp 0
transform 1 0 3190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__430_
timestamp 0
transform -1 0 3870 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__431_
timestamp 0
transform 1 0 3950 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__432_
timestamp 0
transform -1 0 3430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__433_
timestamp 0
transform -1 0 3690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__434_
timestamp 0
transform 1 0 4210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__435_
timestamp 0
transform 1 0 4690 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__436_
timestamp 0
transform 1 0 4790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__437_
timestamp 0
transform -1 0 4770 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__438_
timestamp 0
transform -1 0 4250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__439_
timestamp 0
transform -1 0 4230 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__440_
timestamp 0
transform -1 0 3430 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__441_
timestamp 0
transform -1 0 3970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__442_
timestamp 0
transform -1 0 4410 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__443_
timestamp 0
transform 1 0 4630 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__444_
timestamp 0
transform -1 0 4270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__445_
timestamp 0
transform -1 0 4770 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__446_
timestamp 0
transform 1 0 4730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__447_
timestamp 0
transform 1 0 4790 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__448_
timestamp 0
transform -1 0 4570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__449_
timestamp 0
transform 1 0 4130 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__450_
timestamp 0
transform 1 0 4530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__451_
timestamp 0
transform 1 0 4770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__452_
timestamp 0
transform 1 0 4650 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__453_
timestamp 0
transform 1 0 4810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__454_
timestamp 0
transform 1 0 4290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__455_
timestamp 0
transform -1 0 3770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__456_
timestamp 0
transform -1 0 4050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__457_
timestamp 0
transform 1 0 4010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__458_
timestamp 0
transform -1 0 3750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__459_
timestamp 0
transform -1 0 4750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__460_
timestamp 0
transform 1 0 4810 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__461_
timestamp 0
transform 1 0 4510 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__462_
timestamp 0
transform 1 0 4750 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__463_
timestamp 0
transform 1 0 4810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__464_
timestamp 0
transform 1 0 4230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__465_
timestamp 0
transform 1 0 4390 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__466_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__467_
timestamp 0
transform 1 0 4530 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__468_
timestamp 0
transform 1 0 4230 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__469_
timestamp 0
transform -1 0 2930 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__470_
timestamp 0
transform -1 0 2390 0 1 730
box -6 -8 26 248
use FILL  FILL_3__471_
timestamp 0
transform -1 0 2590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__472_
timestamp 0
transform 1 0 2110 0 1 730
box -6 -8 26 248
use FILL  FILL_3__473_
timestamp 0
transform 1 0 2410 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__474_
timestamp 0
transform 1 0 2690 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__475_
timestamp 0
transform 1 0 3350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__476_
timestamp 0
transform 1 0 2830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__477_
timestamp 0
transform -1 0 2310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__478_
timestamp 0
transform -1 0 2190 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__479_
timestamp 0
transform -1 0 3250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__480_
timestamp 0
transform 1 0 3190 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__481_
timestamp 0
transform -1 0 2690 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__482_
timestamp 0
transform 1 0 2790 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__483_
timestamp 0
transform -1 0 1350 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__484_
timestamp 0
transform -1 0 1070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__485_
timestamp 0
transform -1 0 1670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__486_
timestamp 0
transform -1 0 1650 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__487_
timestamp 0
transform -1 0 1390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__488_
timestamp 0
transform -1 0 1110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__489_
timestamp 0
transform -1 0 1930 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__490_
timestamp 0
transform 1 0 1630 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__491_
timestamp 0
transform 1 0 2730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__492_
timestamp 0
transform -1 0 3490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__493_
timestamp 0
transform 1 0 2990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__494_
timestamp 0
transform 1 0 2950 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__495_
timestamp 0
transform 1 0 2130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__496_
timestamp 0
transform 1 0 810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__497_
timestamp 0
transform -1 0 1590 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__498_
timestamp 0
transform 1 0 950 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__499_
timestamp 0
transform 1 0 1330 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__500_
timestamp 0
transform -1 0 1830 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__501_
timestamp 0
transform 1 0 1170 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__502_
timestamp 0
transform -1 0 1390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__503_
timestamp 0
transform 1 0 1630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__504_
timestamp 0
transform -1 0 2670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__505_
timestamp 0
transform -1 0 2930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__506_
timestamp 0
transform 1 0 3170 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__507_
timestamp 0
transform 1 0 2910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__508_
timestamp 0
transform -1 0 2810 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__509_
timestamp 0
transform 1 0 3150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__510_
timestamp 0
transform 1 0 3070 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__511_
timestamp 0
transform 1 0 2550 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__512_
timestamp 0
transform 1 0 1650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__513_
timestamp 0
transform -1 0 1470 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__514_
timestamp 0
transform 1 0 1510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__515_
timestamp 0
transform 1 0 1890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__516_
timestamp 0
transform 1 0 1730 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__517_
timestamp 0
transform -1 0 2030 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__518_
timestamp 0
transform -1 0 2730 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__519_
timestamp 0
transform 1 0 2450 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__520_
timestamp 0
transform 1 0 2370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__521_
timestamp 0
transform 1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__522_
timestamp 0
transform -1 0 2670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__523_
timestamp 0
transform 1 0 2250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__524_
timestamp 0
transform 1 0 4290 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__525_
timestamp 0
transform -1 0 4570 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__526_
timestamp 0
transform -1 0 4550 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__527_
timestamp 0
transform -1 0 4490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__528_
timestamp 0
transform -1 0 4230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__529_
timestamp 0
transform -1 0 4290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__530_
timestamp 0
transform 1 0 4250 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__531_
timestamp 0
transform -1 0 1770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__532_
timestamp 0
transform -1 0 890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__533_
timestamp 0
transform -1 0 3770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__534_
timestamp 0
transform -1 0 3210 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__535_
timestamp 0
transform -1 0 2530 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__536_
timestamp 0
transform 1 0 2170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__537_
timestamp 0
transform -1 0 1130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__538_
timestamp 0
transform 1 0 1910 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__539_
timestamp 0
transform 1 0 2410 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__540_
timestamp 0
transform 1 0 850 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__541_
timestamp 0
transform 1 0 1070 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__542_
timestamp 0
transform 1 0 1350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__543_
timestamp 0
transform -1 0 1090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__544_
timestamp 0
transform -1 0 610 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__545_
timestamp 0
transform -1 0 90 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__546_
timestamp 0
transform -1 0 90 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__547_
timestamp 0
transform -1 0 90 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__548_
timestamp 0
transform -1 0 350 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__549_
timestamp 0
transform -1 0 330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__550_
timestamp 0
transform -1 0 610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__551_
timestamp 0
transform 1 0 610 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__552_
timestamp 0
transform 1 0 850 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__553_
timestamp 0
transform 1 0 1110 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__554_
timestamp 0
transform 1 0 1390 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__555_
timestamp 0
transform -1 0 330 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__556_
timestamp 0
transform -1 0 90 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__557_
timestamp 0
transform -1 0 90 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__558_
timestamp 0
transform 1 0 350 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__559_
timestamp 0
transform -1 0 90 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__560_
timestamp 0
transform -1 0 890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__561_
timestamp 0
transform 1 0 590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__562_
timestamp 0
transform 1 0 890 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__563_
timestamp 0
transform -1 0 630 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__564_
timestamp 0
transform -1 0 90 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__565_
timestamp 0
transform 1 0 70 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__566_
timestamp 0
transform 1 0 70 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__567_
timestamp 0
transform 1 0 350 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__568_
timestamp 0
transform -1 0 630 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__569_
timestamp 0
transform -1 0 890 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__570_
timestamp 0
transform 1 0 850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__571_
timestamp 0
transform -1 0 610 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__572_
timestamp 0
transform -1 0 330 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__573_
timestamp 0
transform 1 0 330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__574_
timestamp 0
transform -1 0 350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__575_
timestamp 0
transform 1 0 570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__576_
timestamp 0
transform 1 0 590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__577_
timestamp 0
transform -1 0 90 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__578_
timestamp 0
transform -1 0 90 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__579_
timestamp 0
transform 1 0 570 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__580_
timestamp 0
transform -1 0 350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__581_
timestamp 0
transform -1 0 330 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__582_
timestamp 0
transform 1 0 830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__583_
timestamp 0
transform -1 0 610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__584_
timestamp 0
transform 1 0 430 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__585_
timestamp 0
transform -1 0 570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__586_
timestamp 0
transform -1 0 370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__587_
timestamp 0
transform -1 0 90 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__588_
timestamp 0
transform -1 0 90 0 1 250
box -6 -8 26 248
use FILL  FILL_3__589_
timestamp 0
transform -1 0 90 0 1 730
box -6 -8 26 248
use FILL  FILL_3__590_
timestamp 0
transform -1 0 90 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__591_
timestamp 0
transform -1 0 350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__592_
timestamp 0
transform -1 0 650 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__593_
timestamp 0
transform 1 0 350 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__594_
timestamp 0
transform -1 0 90 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__595_
timestamp 0
transform -1 0 350 0 1 730
box -6 -8 26 248
use FILL  FILL_3__596_
timestamp 0
transform 1 0 590 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__597_
timestamp 0
transform 1 0 570 0 1 730
box -6 -8 26 248
use FILL  FILL_3__598_
timestamp 0
transform 1 0 630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__599_
timestamp 0
transform 1 0 1190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__600_
timestamp 0
transform -1 0 90 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__601_
timestamp 0
transform -1 0 590 0 1 250
box -6 -8 26 248
use FILL  FILL_3__602_
timestamp 0
transform -1 0 850 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__603_
timestamp 0
transform 1 0 1470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__604_
timestamp 0
transform 1 0 1630 0 1 250
box -6 -8 26 248
use FILL  FILL_3__605_
timestamp 0
transform 1 0 1090 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__606_
timestamp 0
transform -1 0 1630 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__607_
timestamp 0
transform 1 0 1610 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__608_
timestamp 0
transform 1 0 1110 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__609_
timestamp 0
transform -1 0 1110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__610_
timestamp 0
transform 1 0 1330 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__611_
timestamp 0
transform -1 0 1410 0 1 250
box -6 -8 26 248
use FILL  FILL_3__612_
timestamp 0
transform 1 0 1110 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__613_
timestamp 0
transform 1 0 1870 0 1 250
box -6 -8 26 248
use FILL  FILL_3__614_
timestamp 0
transform 1 0 1870 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__615_
timestamp 0
transform 1 0 2150 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__616_
timestamp 0
transform 1 0 2390 0 1 250
box -6 -8 26 248
use FILL  FILL_3__617_
timestamp 0
transform 1 0 2410 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__618_
timestamp 0
transform 1 0 850 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__619_
timestamp 0
transform -1 0 350 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__620_
timestamp 0
transform 1 0 870 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__621_
timestamp 0
transform -1 0 630 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__622_
timestamp 0
transform -1 0 850 0 1 250
box -6 -8 26 248
use FILL  FILL_3__623_
timestamp 0
transform 1 0 1110 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__624_
timestamp 0
transform 1 0 330 0 1 250
box -6 -8 26 248
use FILL  FILL_3__625_
timestamp 0
transform 1 0 330 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__665_
timestamp 0
transform 1 0 3350 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__666_
timestamp 0
transform 1 0 2710 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__667_
timestamp 0
transform -1 0 4270 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__668_
timestamp 0
transform 1 0 1930 0 1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert6
timestamp 0
transform -1 0 870 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert7
timestamp 0
transform 1 0 2650 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert8
timestamp 0
transform 1 0 1390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert9
timestamp 0
transform 1 0 1130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert10
timestamp 0
transform -1 0 1890 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform 1 0 2410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 1130 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform 1 0 2130 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform -1 0 850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform 1 0 2390 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 3230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 1870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform 1 0 3150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform 1 0 2030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert20
timestamp 0
transform 1 0 1750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert0
timestamp 0
transform 1 0 2030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert1
timestamp 0
transform -1 0 1670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert2
timestamp 0
transform 1 0 70 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert3
timestamp 0
transform 1 0 1810 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert4
timestamp 0
transform 1 0 1130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert5
timestamp 0
transform 1 0 1150 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__313_
timestamp 0
transform 1 0 1130 0 1 250
box -6 -8 26 248
use FILL  FILL_4__314_
timestamp 0
transform -1 0 1130 0 1 730
box -6 -8 26 248
use FILL  FILL_4__315_
timestamp 0
transform 1 0 850 0 1 730
box -6 -8 26 248
use FILL  FILL_4__316_
timestamp 0
transform -1 0 950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__317_
timestamp 0
transform -1 0 2710 0 1 250
box -6 -8 26 248
use FILL  FILL_4__318_
timestamp 0
transform 1 0 2950 0 1 250
box -6 -8 26 248
use FILL  FILL_4__319_
timestamp 0
transform -1 0 3250 0 1 250
box -6 -8 26 248
use FILL  FILL_4__320_
timestamp 0
transform -1 0 3190 0 1 730
box -6 -8 26 248
use FILL  FILL_4__321_
timestamp 0
transform 1 0 3490 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__322_
timestamp 0
transform 1 0 2910 0 1 730
box -6 -8 26 248
use FILL  FILL_4__323_
timestamp 0
transform -1 0 2990 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__324_
timestamp 0
transform -1 0 2670 0 1 730
box -6 -8 26 248
use FILL  FILL_4__325_
timestamp 0
transform -1 0 3510 0 1 250
box -6 -8 26 248
use FILL  FILL_4__326_
timestamp 0
transform -1 0 3790 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__327_
timestamp 0
transform 1 0 4770 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__328_
timestamp 0
transform 1 0 4290 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__329_
timestamp 0
transform -1 0 4550 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__330_
timestamp 0
transform 1 0 4030 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__331_
timestamp 0
transform -1 0 2990 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__332_
timestamp 0
transform -1 0 2730 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__333_
timestamp 0
transform 1 0 2170 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__334_
timestamp 0
transform 1 0 2150 0 1 250
box -6 -8 26 248
use FILL  FILL_4__335_
timestamp 0
transform -1 0 1910 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__336_
timestamp 0
transform -1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__337_
timestamp 0
transform 1 0 3490 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__338_
timestamp 0
transform -1 0 4070 0 1 250
box -6 -8 26 248
use FILL  FILL_4__339_
timestamp 0
transform 1 0 3770 0 1 250
box -6 -8 26 248
use FILL  FILL_4__340_
timestamp 0
transform 1 0 4270 0 1 250
box -6 -8 26 248
use FILL  FILL_4__341_
timestamp 0
transform 1 0 4730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__342_
timestamp 0
transform 1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__343_
timestamp 0
transform -1 0 4830 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__344_
timestamp 0
transform -1 0 4570 0 1 250
box -6 -8 26 248
use FILL  FILL_4__345_
timestamp 0
transform -1 0 4550 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__346_
timestamp 0
transform 1 0 4230 0 1 730
box -6 -8 26 248
use FILL  FILL_4__347_
timestamp 0
transform -1 0 3450 0 1 730
box -6 -8 26 248
use FILL  FILL_4__348_
timestamp 0
transform -1 0 3730 0 1 730
box -6 -8 26 248
use FILL  FILL_4__349_
timestamp 0
transform 1 0 4750 0 1 730
box -6 -8 26 248
use FILL  FILL_4__350_
timestamp 0
transform 1 0 4490 0 1 730
box -6 -8 26 248
use FILL  FILL_4__351_
timestamp 0
transform 1 0 4530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__352_
timestamp 0
transform 1 0 4510 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__353_
timestamp 0
transform 1 0 4190 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__354_
timestamp 0
transform 1 0 3950 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__355_
timestamp 0
transform 1 0 4450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__356_
timestamp 0
transform -1 0 4190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__357_
timestamp 0
transform -1 0 3650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__358_
timestamp 0
transform -1 0 3910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__359_
timestamp 0
transform -1 0 3510 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__360_
timestamp 0
transform 1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__361_
timestamp 0
transform 1 0 4250 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__362_
timestamp 0
transform -1 0 3990 0 1 730
box -6 -8 26 248
use FILL  FILL_4__363_
timestamp 0
transform -1 0 4950 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__364_
timestamp 0
transform -1 0 4450 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__365_
timestamp 0
transform -1 0 3450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__366_
timestamp 0
transform -1 0 3510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__367_
timestamp 0
transform 1 0 4030 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__368_
timestamp 0
transform 1 0 4550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__369_
timestamp 0
transform 1 0 4030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__370_
timestamp 0
transform 1 0 3730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__371_
timestamp 0
transform 1 0 4010 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__372_
timestamp 0
transform 1 0 4030 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__373_
timestamp 0
transform -1 0 3770 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__374_
timestamp 0
transform -1 0 3790 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__375_
timestamp 0
transform 1 0 3750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__376_
timestamp 0
transform 1 0 3270 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__377_
timestamp 0
transform -1 0 3010 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__378_
timestamp 0
transform 1 0 3490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__379_
timestamp 0
transform -1 0 3230 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__380_
timestamp 0
transform -1 0 3510 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__381_
timestamp 0
transform -1 0 3250 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__382_
timestamp 0
transform 1 0 3210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__383_
timestamp 0
transform -1 0 2970 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__384_
timestamp 0
transform 1 0 3770 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__385_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__386_
timestamp 0
transform -1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__387_
timestamp 0
transform 1 0 2190 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__388_
timestamp 0
transform 1 0 2470 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__389_
timestamp 0
transform -1 0 2970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__390_
timestamp 0
transform -1 0 1890 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__391_
timestamp 0
transform -1 0 2690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__392_
timestamp 0
transform -1 0 2430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__393_
timestamp 0
transform 1 0 1670 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__394_
timestamp 0
transform -1 0 2150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__395_
timestamp 0
transform -1 0 1650 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__396_
timestamp 0
transform 1 0 2210 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__397_
timestamp 0
transform 1 0 2710 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__398_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__399_
timestamp 0
transform 1 0 2470 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__400_
timestamp 0
transform -1 0 1870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__401_
timestamp 0
transform -1 0 2150 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__402_
timestamp 0
transform -1 0 1970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__403_
timestamp 0
transform 1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__404_
timestamp 0
transform -1 0 2150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__405_
timestamp 0
transform 1 0 1550 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__406_
timestamp 0
transform -1 0 1590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__407_
timestamp 0
transform 1 0 3230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__408_
timestamp 0
transform -1 0 2950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__409_
timestamp 0
transform 1 0 3610 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__410_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__411_
timestamp 0
transform -1 0 2430 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__412_
timestamp 0
transform 1 0 2650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__413_
timestamp 0
transform -1 0 2970 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__414_
timestamp 0
transform 1 0 2450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__415_
timestamp 0
transform 1 0 2990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__416_
timestamp 0
transform 1 0 3730 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__417_
timestamp 0
transform -1 0 3890 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__418_
timestamp 0
transform 1 0 4770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__419_
timestamp 0
transform 1 0 4510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__420_
timestamp 0
transform -1 0 4170 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__421_
timestamp 0
transform -1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__422_
timestamp 0
transform -1 0 1650 0 1 730
box -6 -8 26 248
use FILL  FILL_4__423_
timestamp 0
transform 1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__424_
timestamp 0
transform 1 0 1350 0 1 730
box -6 -8 26 248
use FILL  FILL_4__425_
timestamp 0
transform 1 0 1390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__426_
timestamp 0
transform -1 0 3370 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__427_
timestamp 0
transform -1 0 2730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__428_
timestamp 0
transform -1 0 3110 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__429_
timestamp 0
transform 1 0 3210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__430_
timestamp 0
transform -1 0 3890 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__431_
timestamp 0
transform 1 0 3970 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__432_
timestamp 0
transform -1 0 3450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__433_
timestamp 0
transform -1 0 3710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__434_
timestamp 0
transform 1 0 4230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__435_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__436_
timestamp 0
transform 1 0 4810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__437_
timestamp 0
transform -1 0 4790 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__438_
timestamp 0
transform -1 0 4270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__439_
timestamp 0
transform -1 0 4250 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__440_
timestamp 0
transform -1 0 3450 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__441_
timestamp 0
transform -1 0 3990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__442_
timestamp 0
transform -1 0 4430 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__443_
timestamp 0
transform 1 0 4650 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__444_
timestamp 0
transform -1 0 4290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__445_
timestamp 0
transform -1 0 4790 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__446_
timestamp 0
transform 1 0 4750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__447_
timestamp 0
transform 1 0 4810 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__448_
timestamp 0
transform -1 0 4590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__449_
timestamp 0
transform 1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__450_
timestamp 0
transform 1 0 4550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__451_
timestamp 0
transform 1 0 4790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__452_
timestamp 0
transform 1 0 4670 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__453_
timestamp 0
transform 1 0 4830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__454_
timestamp 0
transform 1 0 4310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__455_
timestamp 0
transform -1 0 3790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__456_
timestamp 0
transform -1 0 4070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__457_
timestamp 0
transform 1 0 4030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__458_
timestamp 0
transform -1 0 3770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__459_
timestamp 0
transform -1 0 4770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__460_
timestamp 0
transform 1 0 4830 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__461_
timestamp 0
transform 1 0 4530 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__462_
timestamp 0
transform 1 0 4770 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__463_
timestamp 0
transform 1 0 4830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__464_
timestamp 0
transform 1 0 4250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__465_
timestamp 0
transform 1 0 4410 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__466_
timestamp 0
transform 1 0 4510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__467_
timestamp 0
transform 1 0 4550 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__468_
timestamp 0
transform 1 0 4250 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__469_
timestamp 0
transform -1 0 2950 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__470_
timestamp 0
transform -1 0 2410 0 1 730
box -6 -8 26 248
use FILL  FILL_4__471_
timestamp 0
transform -1 0 2610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__472_
timestamp 0
transform 1 0 2130 0 1 730
box -6 -8 26 248
use FILL  FILL_4__473_
timestamp 0
transform 1 0 2430 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__474_
timestamp 0
transform 1 0 2710 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__475_
timestamp 0
transform 1 0 3370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__476_
timestamp 0
transform 1 0 2850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__477_
timestamp 0
transform -1 0 2330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__478_
timestamp 0
transform -1 0 2210 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__479_
timestamp 0
transform -1 0 3270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__480_
timestamp 0
transform 1 0 3210 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__481_
timestamp 0
transform -1 0 2710 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__482_
timestamp 0
transform 1 0 2810 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__483_
timestamp 0
transform -1 0 1370 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__484_
timestamp 0
transform -1 0 1090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__485_
timestamp 0
transform -1 0 1690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__486_
timestamp 0
transform -1 0 1670 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__487_
timestamp 0
transform -1 0 1410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__488_
timestamp 0
transform -1 0 1130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__489_
timestamp 0
transform -1 0 1950 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__490_
timestamp 0
transform 1 0 1650 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__491_
timestamp 0
transform 1 0 2750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__492_
timestamp 0
transform -1 0 3510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__493_
timestamp 0
transform 1 0 3010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__494_
timestamp 0
transform 1 0 2970 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__495_
timestamp 0
transform 1 0 2150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__496_
timestamp 0
transform 1 0 830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__497_
timestamp 0
transform -1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__498_
timestamp 0
transform 1 0 970 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__499_
timestamp 0
transform 1 0 1350 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__500_
timestamp 0
transform -1 0 1850 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__501_
timestamp 0
transform 1 0 1190 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__502_
timestamp 0
transform -1 0 1410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__503_
timestamp 0
transform 1 0 1650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__504_
timestamp 0
transform -1 0 2690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__505_
timestamp 0
transform -1 0 2950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__506_
timestamp 0
transform 1 0 3190 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__507_
timestamp 0
transform 1 0 2930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__508_
timestamp 0
transform -1 0 2830 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__509_
timestamp 0
transform 1 0 3170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__510_
timestamp 0
transform 1 0 3090 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__511_
timestamp 0
transform 1 0 2570 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__512_
timestamp 0
transform 1 0 1670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__513_
timestamp 0
transform -1 0 1490 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__514_
timestamp 0
transform 1 0 1530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__515_
timestamp 0
transform 1 0 1910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__516_
timestamp 0
transform 1 0 1750 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__517_
timestamp 0
transform -1 0 2050 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__518_
timestamp 0
transform -1 0 2750 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__519_
timestamp 0
transform 1 0 2470 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__520_
timestamp 0
transform 1 0 2390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__521_
timestamp 0
transform 1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__522_
timestamp 0
transform -1 0 2690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__523_
timestamp 0
transform 1 0 2270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__524_
timestamp 0
transform 1 0 4310 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__525_
timestamp 0
transform -1 0 4590 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__526_
timestamp 0
transform -1 0 4570 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__527_
timestamp 0
transform -1 0 4510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__528_
timestamp 0
transform -1 0 4250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__529_
timestamp 0
transform -1 0 4310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__530_
timestamp 0
transform 1 0 4270 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__531_
timestamp 0
transform -1 0 1790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__532_
timestamp 0
transform -1 0 910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__533_
timestamp 0
transform -1 0 3790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__534_
timestamp 0
transform -1 0 3230 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__535_
timestamp 0
transform -1 0 2550 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__536_
timestamp 0
transform 1 0 2190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__537_
timestamp 0
transform -1 0 1150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__538_
timestamp 0
transform 1 0 1930 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__539_
timestamp 0
transform 1 0 2430 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__540_
timestamp 0
transform 1 0 870 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__541_
timestamp 0
transform 1 0 1090 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__542_
timestamp 0
transform 1 0 1370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__543_
timestamp 0
transform -1 0 1110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__544_
timestamp 0
transform -1 0 630 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__545_
timestamp 0
transform -1 0 110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__546_
timestamp 0
transform -1 0 110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__547_
timestamp 0
transform -1 0 110 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__548_
timestamp 0
transform -1 0 370 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__549_
timestamp 0
transform -1 0 350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__550_
timestamp 0
transform -1 0 630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__551_
timestamp 0
transform 1 0 630 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__552_
timestamp 0
transform 1 0 870 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__553_
timestamp 0
transform 1 0 1130 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__554_
timestamp 0
transform 1 0 1410 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__555_
timestamp 0
transform -1 0 350 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__556_
timestamp 0
transform -1 0 110 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__557_
timestamp 0
transform -1 0 110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__558_
timestamp 0
transform 1 0 370 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__559_
timestamp 0
transform -1 0 110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__560_
timestamp 0
transform -1 0 910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__561_
timestamp 0
transform 1 0 610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__562_
timestamp 0
transform 1 0 910 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__563_
timestamp 0
transform -1 0 650 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__564_
timestamp 0
transform -1 0 110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__565_
timestamp 0
transform 1 0 90 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__566_
timestamp 0
transform 1 0 90 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__567_
timestamp 0
transform 1 0 370 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__568_
timestamp 0
transform -1 0 650 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__569_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__570_
timestamp 0
transform 1 0 870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__571_
timestamp 0
transform -1 0 630 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__572_
timestamp 0
transform -1 0 350 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__573_
timestamp 0
transform 1 0 350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__574_
timestamp 0
transform -1 0 370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__575_
timestamp 0
transform 1 0 590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__576_
timestamp 0
transform 1 0 610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__577_
timestamp 0
transform -1 0 110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__578_
timestamp 0
transform -1 0 110 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__579_
timestamp 0
transform 1 0 590 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__580_
timestamp 0
transform -1 0 370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__581_
timestamp 0
transform -1 0 350 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__582_
timestamp 0
transform 1 0 850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__583_
timestamp 0
transform -1 0 630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__584_
timestamp 0
transform 1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__585_
timestamp 0
transform -1 0 590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__586_
timestamp 0
transform -1 0 390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__587_
timestamp 0
transform -1 0 110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__588_
timestamp 0
transform -1 0 110 0 1 250
box -6 -8 26 248
use FILL  FILL_4__589_
timestamp 0
transform -1 0 110 0 1 730
box -6 -8 26 248
use FILL  FILL_4__590_
timestamp 0
transform -1 0 110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__591_
timestamp 0
transform -1 0 370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__592_
timestamp 0
transform -1 0 670 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__593_
timestamp 0
transform 1 0 370 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__594_
timestamp 0
transform -1 0 110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__595_
timestamp 0
transform -1 0 370 0 1 730
box -6 -8 26 248
use FILL  FILL_4__596_
timestamp 0
transform 1 0 610 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__597_
timestamp 0
transform 1 0 590 0 1 730
box -6 -8 26 248
use FILL  FILL_4__598_
timestamp 0
transform 1 0 650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__599_
timestamp 0
transform 1 0 1210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__600_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__601_
timestamp 0
transform -1 0 610 0 1 250
box -6 -8 26 248
use FILL  FILL_4__602_
timestamp 0
transform -1 0 870 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__603_
timestamp 0
transform 1 0 1490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__604_
timestamp 0
transform 1 0 1650 0 1 250
box -6 -8 26 248
use FILL  FILL_4__605_
timestamp 0
transform 1 0 1110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__606_
timestamp 0
transform -1 0 1650 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__607_
timestamp 0
transform 1 0 1630 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__608_
timestamp 0
transform 1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__609_
timestamp 0
transform -1 0 1130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__610_
timestamp 0
transform 1 0 1350 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__611_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 26 248
use FILL  FILL_4__612_
timestamp 0
transform 1 0 1130 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__613_
timestamp 0
transform 1 0 1890 0 1 250
box -6 -8 26 248
use FILL  FILL_4__614_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__615_
timestamp 0
transform 1 0 2170 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__616_
timestamp 0
transform 1 0 2410 0 1 250
box -6 -8 26 248
use FILL  FILL_4__617_
timestamp 0
transform 1 0 2430 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__618_
timestamp 0
transform 1 0 870 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__619_
timestamp 0
transform -1 0 370 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__620_
timestamp 0
transform 1 0 890 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__621_
timestamp 0
transform -1 0 650 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__622_
timestamp 0
transform -1 0 870 0 1 250
box -6 -8 26 248
use FILL  FILL_4__623_
timestamp 0
transform 1 0 1130 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__624_
timestamp 0
transform 1 0 350 0 1 250
box -6 -8 26 248
use FILL  FILL_4__625_
timestamp 0
transform 1 0 350 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__665_
timestamp 0
transform 1 0 3370 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__666_
timestamp 0
transform 1 0 2730 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__667_
timestamp 0
transform -1 0 4290 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__668_
timestamp 0
transform 1 0 1950 0 1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert6
timestamp 0
transform -1 0 890 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert7
timestamp 0
transform 1 0 2670 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert8
timestamp 0
transform 1 0 1410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert9
timestamp 0
transform 1 0 1150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert10
timestamp 0
transform -1 0 1910 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert11
timestamp 0
transform 1 0 2430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert12
timestamp 0
transform 1 0 1150 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform 1 0 2150 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform -1 0 870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert15
timestamp 0
transform 1 0 2410 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert16
timestamp 0
transform 1 0 3250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform 1 0 1890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert18
timestamp 0
transform 1 0 3170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert19
timestamp 0
transform 1 0 2050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert20
timestamp 0
transform 1 0 1770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert0
timestamp 0
transform 1 0 2050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert1
timestamp 0
transform -1 0 1690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert2
timestamp 0
transform 1 0 90 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert3
timestamp 0
transform 1 0 1830 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert4
timestamp 0
transform 1 0 1150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert5
timestamp 0
transform 1 0 1170 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__313_
timestamp 0
transform 1 0 1150 0 1 250
box -6 -8 26 248
use FILL  FILL_5__314_
timestamp 0
transform -1 0 1150 0 1 730
box -6 -8 26 248
use FILL  FILL_5__315_
timestamp 0
transform 1 0 870 0 1 730
box -6 -8 26 248
use FILL  FILL_5__316_
timestamp 0
transform -1 0 970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__317_
timestamp 0
transform -1 0 2730 0 1 250
box -6 -8 26 248
use FILL  FILL_5__318_
timestamp 0
transform 1 0 2970 0 1 250
box -6 -8 26 248
use FILL  FILL_5__319_
timestamp 0
transform -1 0 3270 0 1 250
box -6 -8 26 248
use FILL  FILL_5__320_
timestamp 0
transform -1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_5__321_
timestamp 0
transform 1 0 3510 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__322_
timestamp 0
transform 1 0 2930 0 1 730
box -6 -8 26 248
use FILL  FILL_5__323_
timestamp 0
transform -1 0 3010 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__324_
timestamp 0
transform -1 0 2690 0 1 730
box -6 -8 26 248
use FILL  FILL_5__325_
timestamp 0
transform -1 0 3530 0 1 250
box -6 -8 26 248
use FILL  FILL_5__326_
timestamp 0
transform -1 0 3810 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__327_
timestamp 0
transform 1 0 4790 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__328_
timestamp 0
transform 1 0 4310 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__329_
timestamp 0
transform -1 0 4570 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__330_
timestamp 0
transform 1 0 4050 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__331_
timestamp 0
transform -1 0 3010 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__332_
timestamp 0
transform -1 0 2750 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__333_
timestamp 0
transform 1 0 2190 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__334_
timestamp 0
transform 1 0 2170 0 1 250
box -6 -8 26 248
use FILL  FILL_5__335_
timestamp 0
transform -1 0 1930 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__336_
timestamp 0
transform -1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__337_
timestamp 0
transform 1 0 3510 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__338_
timestamp 0
transform -1 0 4090 0 1 250
box -6 -8 26 248
use FILL  FILL_5__339_
timestamp 0
transform 1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_5__340_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 26 248
use FILL  FILL_5__341_
timestamp 0
transform 1 0 4750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__342_
timestamp 0
transform 1 0 4830 0 1 250
box -6 -8 26 248
use FILL  FILL_5__343_
timestamp 0
transform -1 0 4850 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__344_
timestamp 0
transform -1 0 4590 0 1 250
box -6 -8 26 248
use FILL  FILL_5__345_
timestamp 0
transform -1 0 4570 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__346_
timestamp 0
transform 1 0 4250 0 1 730
box -6 -8 26 248
use FILL  FILL_5__347_
timestamp 0
transform -1 0 3470 0 1 730
box -6 -8 26 248
use FILL  FILL_5__348_
timestamp 0
transform -1 0 3750 0 1 730
box -6 -8 26 248
use FILL  FILL_5__349_
timestamp 0
transform 1 0 4770 0 1 730
box -6 -8 26 248
use FILL  FILL_5__350_
timestamp 0
transform 1 0 4510 0 1 730
box -6 -8 26 248
use FILL  FILL_5__351_
timestamp 0
transform 1 0 4550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__352_
timestamp 0
transform 1 0 4530 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__353_
timestamp 0
transform 1 0 4210 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__354_
timestamp 0
transform 1 0 3970 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__355_
timestamp 0
transform 1 0 4470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__356_
timestamp 0
transform -1 0 4210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__357_
timestamp 0
transform -1 0 3670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__358_
timestamp 0
transform -1 0 3930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__359_
timestamp 0
transform -1 0 3530 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__360_
timestamp 0
transform 1 0 4010 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__361_
timestamp 0
transform 1 0 4270 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__362_
timestamp 0
transform -1 0 4010 0 1 730
box -6 -8 26 248
use FILL  FILL_5__363_
timestamp 0
transform -1 0 4970 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__364_
timestamp 0
transform -1 0 4470 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__365_
timestamp 0
transform -1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__366_
timestamp 0
transform -1 0 3530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__367_
timestamp 0
transform 1 0 4050 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__368_
timestamp 0
transform 1 0 4570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__369_
timestamp 0
transform 1 0 4050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__370_
timestamp 0
transform 1 0 3750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__371_
timestamp 0
transform 1 0 4030 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__372_
timestamp 0
transform 1 0 4050 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__373_
timestamp 0
transform -1 0 3790 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__374_
timestamp 0
transform -1 0 3810 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__375_
timestamp 0
transform 1 0 3770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__376_
timestamp 0
transform 1 0 3290 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__377_
timestamp 0
transform -1 0 3030 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__378_
timestamp 0
transform 1 0 3510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__379_
timestamp 0
transform -1 0 3250 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__380_
timestamp 0
transform -1 0 3530 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__381_
timestamp 0
transform -1 0 3270 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__382_
timestamp 0
transform 1 0 3230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__383_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__384_
timestamp 0
transform 1 0 3790 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__385_
timestamp 0
transform -1 0 3550 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__386_
timestamp 0
transform -1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__387_
timestamp 0
transform 1 0 2210 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__388_
timestamp 0
transform 1 0 2490 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__389_
timestamp 0
transform -1 0 2990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__390_
timestamp 0
transform -1 0 1910 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__391_
timestamp 0
transform -1 0 2710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__392_
timestamp 0
transform -1 0 2450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__393_
timestamp 0
transform 1 0 1690 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__394_
timestamp 0
transform -1 0 2170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__395_
timestamp 0
transform -1 0 1670 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__396_
timestamp 0
transform 1 0 2230 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__397_
timestamp 0
transform 1 0 2730 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__398_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__399_
timestamp 0
transform 1 0 2490 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__400_
timestamp 0
transform -1 0 1890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__401_
timestamp 0
transform -1 0 2170 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__402_
timestamp 0
transform -1 0 1990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__403_
timestamp 0
transform 1 0 2410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__404_
timestamp 0
transform -1 0 2170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__405_
timestamp 0
transform 1 0 1570 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__406_
timestamp 0
transform -1 0 1610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__407_
timestamp 0
transform 1 0 3250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__408_
timestamp 0
transform -1 0 2970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__409_
timestamp 0
transform 1 0 3630 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__410_
timestamp 0
transform -1 0 3750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__411_
timestamp 0
transform -1 0 2450 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__412_
timestamp 0
transform 1 0 2670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__413_
timestamp 0
transform -1 0 2990 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__414_
timestamp 0
transform 1 0 2470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__415_
timestamp 0
transform 1 0 3010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__416_
timestamp 0
transform 1 0 3750 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__417_
timestamp 0
transform -1 0 3910 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__418_
timestamp 0
transform 1 0 4790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__419_
timestamp 0
transform 1 0 4530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__420_
timestamp 0
transform -1 0 4190 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__421_
timestamp 0
transform -1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__422_
timestamp 0
transform -1 0 1670 0 1 730
box -6 -8 26 248
use FILL  FILL_5__423_
timestamp 0
transform 1 0 1410 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__424_
timestamp 0
transform 1 0 1370 0 1 730
box -6 -8 26 248
use FILL  FILL_5__425_
timestamp 0
transform 1 0 1410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__426_
timestamp 0
transform -1 0 3390 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__427_
timestamp 0
transform -1 0 2750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__428_
timestamp 0
transform -1 0 3130 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__429_
timestamp 0
transform 1 0 3230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__430_
timestamp 0
transform -1 0 3910 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__431_
timestamp 0
transform 1 0 3990 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__432_
timestamp 0
transform -1 0 3470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__433_
timestamp 0
transform -1 0 3730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__434_
timestamp 0
transform 1 0 4250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__435_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__436_
timestamp 0
transform 1 0 4830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__437_
timestamp 0
transform -1 0 4810 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__438_
timestamp 0
transform -1 0 4290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__439_
timestamp 0
transform -1 0 4270 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__440_
timestamp 0
transform -1 0 3470 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__441_
timestamp 0
transform -1 0 4010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__442_
timestamp 0
transform -1 0 4450 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__443_
timestamp 0
transform 1 0 4670 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__444_
timestamp 0
transform -1 0 4310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__445_
timestamp 0
transform -1 0 4810 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__446_
timestamp 0
transform 1 0 4770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__447_
timestamp 0
transform 1 0 4830 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__448_
timestamp 0
transform -1 0 4610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__449_
timestamp 0
transform 1 0 4170 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__450_
timestamp 0
transform 1 0 4570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__451_
timestamp 0
transform 1 0 4810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__452_
timestamp 0
transform 1 0 4690 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__453_
timestamp 0
transform 1 0 4850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__454_
timestamp 0
transform 1 0 4330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__455_
timestamp 0
transform -1 0 3810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__456_
timestamp 0
transform -1 0 4090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__457_
timestamp 0
transform 1 0 4050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__458_
timestamp 0
transform -1 0 3790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__459_
timestamp 0
transform -1 0 4790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__460_
timestamp 0
transform 1 0 4850 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__461_
timestamp 0
transform 1 0 4550 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__462_
timestamp 0
transform 1 0 4790 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__463_
timestamp 0
transform 1 0 4850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__464_
timestamp 0
transform 1 0 4270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__465_
timestamp 0
transform 1 0 4430 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__466_
timestamp 0
transform 1 0 4530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__467_
timestamp 0
transform 1 0 4570 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__468_
timestamp 0
transform 1 0 4270 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__469_
timestamp 0
transform -1 0 2970 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__470_
timestamp 0
transform -1 0 2430 0 1 730
box -6 -8 26 248
use FILL  FILL_5__471_
timestamp 0
transform -1 0 2630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__472_
timestamp 0
transform 1 0 2150 0 1 730
box -6 -8 26 248
use FILL  FILL_5__473_
timestamp 0
transform 1 0 2450 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__474_
timestamp 0
transform 1 0 2730 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__475_
timestamp 0
transform 1 0 3390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__476_
timestamp 0
transform 1 0 2870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__477_
timestamp 0
transform -1 0 2350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__478_
timestamp 0
transform -1 0 2230 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__479_
timestamp 0
transform -1 0 3290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__480_
timestamp 0
transform 1 0 3230 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__481_
timestamp 0
transform -1 0 2730 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__482_
timestamp 0
transform 1 0 2830 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__483_
timestamp 0
transform -1 0 1390 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__484_
timestamp 0
transform -1 0 1110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__485_
timestamp 0
transform -1 0 1710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__486_
timestamp 0
transform -1 0 1690 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__487_
timestamp 0
transform -1 0 1430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__488_
timestamp 0
transform -1 0 1150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__489_
timestamp 0
transform -1 0 1970 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__490_
timestamp 0
transform 1 0 1670 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__491_
timestamp 0
transform 1 0 2770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__492_
timestamp 0
transform -1 0 3530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__493_
timestamp 0
transform 1 0 3030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__494_
timestamp 0
transform 1 0 2990 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__495_
timestamp 0
transform 1 0 2170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__496_
timestamp 0
transform 1 0 850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__497_
timestamp 0
transform -1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__498_
timestamp 0
transform 1 0 990 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__499_
timestamp 0
transform 1 0 1370 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__500_
timestamp 0
transform -1 0 1870 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__501_
timestamp 0
transform 1 0 1210 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__502_
timestamp 0
transform -1 0 1430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__503_
timestamp 0
transform 1 0 1670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__504_
timestamp 0
transform -1 0 2710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__505_
timestamp 0
transform -1 0 2970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__506_
timestamp 0
transform 1 0 3210 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__507_
timestamp 0
transform 1 0 2950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__508_
timestamp 0
transform -1 0 2850 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__509_
timestamp 0
transform 1 0 3190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__510_
timestamp 0
transform 1 0 3110 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__511_
timestamp 0
transform 1 0 2590 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__512_
timestamp 0
transform 1 0 1690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__513_
timestamp 0
transform -1 0 1510 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__514_
timestamp 0
transform 1 0 1550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__515_
timestamp 0
transform 1 0 1930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__516_
timestamp 0
transform 1 0 1770 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__517_
timestamp 0
transform -1 0 2070 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__518_
timestamp 0
transform -1 0 2770 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__519_
timestamp 0
transform 1 0 2490 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__520_
timestamp 0
transform 1 0 2410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__521_
timestamp 0
transform 1 0 2690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__522_
timestamp 0
transform -1 0 2710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__523_
timestamp 0
transform 1 0 2290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__524_
timestamp 0
transform 1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__525_
timestamp 0
transform -1 0 4610 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__526_
timestamp 0
transform -1 0 4590 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__527_
timestamp 0
transform -1 0 4530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__528_
timestamp 0
transform -1 0 4270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__529_
timestamp 0
transform -1 0 4330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__530_
timestamp 0
transform 1 0 4290 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__531_
timestamp 0
transform -1 0 1810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__532_
timestamp 0
transform -1 0 930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__533_
timestamp 0
transform -1 0 3810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__534_
timestamp 0
transform -1 0 3250 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__535_
timestamp 0
transform -1 0 2570 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__536_
timestamp 0
transform 1 0 2210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__537_
timestamp 0
transform -1 0 1170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__538_
timestamp 0
transform 1 0 1950 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__539_
timestamp 0
transform 1 0 2450 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__540_
timestamp 0
transform 1 0 890 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__541_
timestamp 0
transform 1 0 1110 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__542_
timestamp 0
transform 1 0 1390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__543_
timestamp 0
transform -1 0 1130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__544_
timestamp 0
transform -1 0 650 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__545_
timestamp 0
transform -1 0 130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__546_
timestamp 0
transform -1 0 130 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__547_
timestamp 0
transform -1 0 130 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__548_
timestamp 0
transform -1 0 390 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__549_
timestamp 0
transform -1 0 370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__550_
timestamp 0
transform -1 0 650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__551_
timestamp 0
transform 1 0 650 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__552_
timestamp 0
transform 1 0 890 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__553_
timestamp 0
transform 1 0 1150 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__554_
timestamp 0
transform 1 0 1430 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__555_
timestamp 0
transform -1 0 370 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__556_
timestamp 0
transform -1 0 130 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__557_
timestamp 0
transform -1 0 130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__558_
timestamp 0
transform 1 0 390 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__559_
timestamp 0
transform -1 0 130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__560_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__561_
timestamp 0
transform 1 0 630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__562_
timestamp 0
transform 1 0 930 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__563_
timestamp 0
transform -1 0 670 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__564_
timestamp 0
transform -1 0 130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__565_
timestamp 0
transform 1 0 110 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__566_
timestamp 0
transform 1 0 110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__567_
timestamp 0
transform 1 0 390 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__568_
timestamp 0
transform -1 0 670 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__569_
timestamp 0
transform -1 0 930 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__570_
timestamp 0
transform 1 0 890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__571_
timestamp 0
transform -1 0 650 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__572_
timestamp 0
transform -1 0 370 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__573_
timestamp 0
transform 1 0 370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__574_
timestamp 0
transform -1 0 390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__575_
timestamp 0
transform 1 0 610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__576_
timestamp 0
transform 1 0 630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__577_
timestamp 0
transform -1 0 130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__578_
timestamp 0
transform -1 0 130 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__579_
timestamp 0
transform 1 0 610 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__580_
timestamp 0
transform -1 0 390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__581_
timestamp 0
transform -1 0 370 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__582_
timestamp 0
transform 1 0 870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__583_
timestamp 0
transform -1 0 650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__584_
timestamp 0
transform 1 0 470 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__585_
timestamp 0
transform -1 0 610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__586_
timestamp 0
transform -1 0 410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__587_
timestamp 0
transform -1 0 130 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__588_
timestamp 0
transform -1 0 130 0 1 250
box -6 -8 26 248
use FILL  FILL_5__589_
timestamp 0
transform -1 0 130 0 1 730
box -6 -8 26 248
use FILL  FILL_5__590_
timestamp 0
transform -1 0 130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__591_
timestamp 0
transform -1 0 390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__592_
timestamp 0
transform -1 0 690 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__593_
timestamp 0
transform 1 0 390 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__594_
timestamp 0
transform -1 0 130 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__595_
timestamp 0
transform -1 0 390 0 1 730
box -6 -8 26 248
use FILL  FILL_5__596_
timestamp 0
transform 1 0 630 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__597_
timestamp 0
transform 1 0 610 0 1 730
box -6 -8 26 248
use FILL  FILL_5__598_
timestamp 0
transform 1 0 670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__599_
timestamp 0
transform 1 0 1230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__600_
timestamp 0
transform -1 0 130 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__601_
timestamp 0
transform -1 0 630 0 1 250
box -6 -8 26 248
use FILL  FILL_5__602_
timestamp 0
transform -1 0 890 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__603_
timestamp 0
transform 1 0 1510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__604_
timestamp 0
transform 1 0 1670 0 1 250
box -6 -8 26 248
use FILL  FILL_5__605_
timestamp 0
transform 1 0 1130 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__606_
timestamp 0
transform -1 0 1670 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__607_
timestamp 0
transform 1 0 1650 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__608_
timestamp 0
transform 1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__609_
timestamp 0
transform -1 0 1150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__610_
timestamp 0
transform 1 0 1370 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__611_
timestamp 0
transform -1 0 1450 0 1 250
box -6 -8 26 248
use FILL  FILL_5__612_
timestamp 0
transform 1 0 1150 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__613_
timestamp 0
transform 1 0 1910 0 1 250
box -6 -8 26 248
use FILL  FILL_5__614_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__615_
timestamp 0
transform 1 0 2190 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__616_
timestamp 0
transform 1 0 2430 0 1 250
box -6 -8 26 248
use FILL  FILL_5__617_
timestamp 0
transform 1 0 2450 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__618_
timestamp 0
transform 1 0 890 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__619_
timestamp 0
transform -1 0 390 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__620_
timestamp 0
transform 1 0 910 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__621_
timestamp 0
transform -1 0 670 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__622_
timestamp 0
transform -1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_5__623_
timestamp 0
transform 1 0 1150 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__624_
timestamp 0
transform 1 0 370 0 1 250
box -6 -8 26 248
use FILL  FILL_5__625_
timestamp 0
transform 1 0 370 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__665_
timestamp 0
transform 1 0 3390 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__666_
timestamp 0
transform 1 0 2750 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__667_
timestamp 0
transform -1 0 4310 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__668_
timestamp 0
transform 1 0 1970 0 1 4570
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert6
timestamp 0
transform -1 0 910 0 1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert7
timestamp 0
transform 1 0 2690 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert8
timestamp 0
transform 1 0 1430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert9
timestamp 0
transform 1 0 1170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert10
timestamp 0
transform -1 0 1930 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert11
timestamp 0
transform 1 0 2450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert12
timestamp 0
transform 1 0 1170 0 1 3130
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert13
timestamp 0
transform 1 0 2170 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert14
timestamp 0
transform -1 0 890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert15
timestamp 0
transform 1 0 2430 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert16
timestamp 0
transform 1 0 3270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert17
timestamp 0
transform 1 0 1910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert18
timestamp 0
transform 1 0 3190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert19
timestamp 0
transform 1 0 2070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert20
timestamp 0
transform 1 0 1790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert0
timestamp 0
transform 1 0 2070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert1
timestamp 0
transform -1 0 1710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert2
timestamp 0
transform 1 0 110 0 1 2170
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert3
timestamp 0
transform 1 0 1850 0 1 3610
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert4
timestamp 0
transform 1 0 1170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert5
timestamp 0
transform 1 0 1190 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__313_
timestamp 0
transform 1 0 1170 0 1 250
box -6 -8 26 248
use FILL  FILL_6__314_
timestamp 0
transform -1 0 1170 0 1 730
box -6 -8 26 248
use FILL  FILL_6__315_
timestamp 0
transform 1 0 890 0 1 730
box -6 -8 26 248
use FILL  FILL_6__316_
timestamp 0
transform -1 0 990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__317_
timestamp 0
transform -1 0 2750 0 1 250
box -6 -8 26 248
use FILL  FILL_6__318_
timestamp 0
transform 1 0 2990 0 1 250
box -6 -8 26 248
use FILL  FILL_6__319_
timestamp 0
transform -1 0 3290 0 1 250
box -6 -8 26 248
use FILL  FILL_6__320_
timestamp 0
transform -1 0 3230 0 1 730
box -6 -8 26 248
use FILL  FILL_6__321_
timestamp 0
transform 1 0 3530 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__322_
timestamp 0
transform 1 0 2950 0 1 730
box -6 -8 26 248
use FILL  FILL_6__323_
timestamp 0
transform -1 0 3030 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__324_
timestamp 0
transform -1 0 2710 0 1 730
box -6 -8 26 248
use FILL  FILL_6__325_
timestamp 0
transform -1 0 3550 0 1 250
box -6 -8 26 248
use FILL  FILL_6__326_
timestamp 0
transform -1 0 3830 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__327_
timestamp 0
transform 1 0 4810 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__328_
timestamp 0
transform 1 0 4330 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__329_
timestamp 0
transform -1 0 4590 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__330_
timestamp 0
transform 1 0 4070 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__331_
timestamp 0
transform -1 0 3030 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__332_
timestamp 0
transform -1 0 2770 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__333_
timestamp 0
transform 1 0 2210 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__334_
timestamp 0
transform 1 0 2190 0 1 250
box -6 -8 26 248
use FILL  FILL_6__335_
timestamp 0
transform -1 0 1950 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__336_
timestamp 0
transform -1 0 3290 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__337_
timestamp 0
transform 1 0 3530 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__338_
timestamp 0
transform -1 0 4110 0 1 250
box -6 -8 26 248
use FILL  FILL_6__339_
timestamp 0
transform 1 0 3810 0 1 250
box -6 -8 26 248
use FILL  FILL_6__340_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 26 248
use FILL  FILL_6__341_
timestamp 0
transform 1 0 4770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__342_
timestamp 0
transform 1 0 4850 0 1 250
box -6 -8 26 248
use FILL  FILL_6__343_
timestamp 0
transform -1 0 4870 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__344_
timestamp 0
transform -1 0 4610 0 1 250
box -6 -8 26 248
use FILL  FILL_6__345_
timestamp 0
transform -1 0 4590 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__346_
timestamp 0
transform 1 0 4270 0 1 730
box -6 -8 26 248
use FILL  FILL_6__347_
timestamp 0
transform -1 0 3490 0 1 730
box -6 -8 26 248
use FILL  FILL_6__348_
timestamp 0
transform -1 0 3770 0 1 730
box -6 -8 26 248
use FILL  FILL_6__349_
timestamp 0
transform 1 0 4790 0 1 730
box -6 -8 26 248
use FILL  FILL_6__350_
timestamp 0
transform 1 0 4530 0 1 730
box -6 -8 26 248
use FILL  FILL_6__351_
timestamp 0
transform 1 0 4570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__352_
timestamp 0
transform 1 0 4550 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__353_
timestamp 0
transform 1 0 4230 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__354_
timestamp 0
transform 1 0 3990 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__355_
timestamp 0
transform 1 0 4490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__356_
timestamp 0
transform -1 0 4230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__357_
timestamp 0
transform -1 0 3690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__358_
timestamp 0
transform -1 0 3950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__359_
timestamp 0
transform -1 0 3550 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__360_
timestamp 0
transform 1 0 4030 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__361_
timestamp 0
transform 1 0 4290 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__362_
timestamp 0
transform -1 0 4030 0 1 730
box -6 -8 26 248
use FILL  FILL_6__363_
timestamp 0
transform -1 0 4990 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__364_
timestamp 0
transform -1 0 4490 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__365_
timestamp 0
transform -1 0 3490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__366_
timestamp 0
transform -1 0 3550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__367_
timestamp 0
transform 1 0 4070 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__368_
timestamp 0
transform 1 0 4590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__369_
timestamp 0
transform 1 0 4070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__370_
timestamp 0
transform 1 0 3770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__371_
timestamp 0
transform 1 0 4050 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__372_
timestamp 0
transform 1 0 4070 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__373_
timestamp 0
transform -1 0 3810 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__374_
timestamp 0
transform -1 0 3830 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__375_
timestamp 0
transform 1 0 3790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__376_
timestamp 0
transform 1 0 3310 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__377_
timestamp 0
transform -1 0 3050 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__378_
timestamp 0
transform 1 0 3530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__379_
timestamp 0
transform -1 0 3270 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__380_
timestamp 0
transform -1 0 3550 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__381_
timestamp 0
transform -1 0 3290 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__382_
timestamp 0
transform 1 0 3250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__383_
timestamp 0
transform -1 0 3010 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__384_
timestamp 0
transform 1 0 3810 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__385_
timestamp 0
transform -1 0 3570 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__386_
timestamp 0
transform -1 0 2730 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__387_
timestamp 0
transform 1 0 2230 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__388_
timestamp 0
transform 1 0 2510 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__389_
timestamp 0
transform -1 0 3010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__390_
timestamp 0
transform -1 0 1930 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__391_
timestamp 0
transform -1 0 2730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__392_
timestamp 0
transform -1 0 2470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__393_
timestamp 0
transform 1 0 1710 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__394_
timestamp 0
transform -1 0 2190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__395_
timestamp 0
transform -1 0 1690 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__396_
timestamp 0
transform 1 0 2250 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__397_
timestamp 0
transform 1 0 2750 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__398_
timestamp 0
transform 1 0 2230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__399_
timestamp 0
transform 1 0 2510 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__400_
timestamp 0
transform -1 0 1910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__401_
timestamp 0
transform -1 0 2190 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__402_
timestamp 0
transform -1 0 2010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__403_
timestamp 0
transform 1 0 2430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__404_
timestamp 0
transform -1 0 2190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__405_
timestamp 0
transform 1 0 1590 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__406_
timestamp 0
transform -1 0 1630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__407_
timestamp 0
transform 1 0 3270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__408_
timestamp 0
transform -1 0 2990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__409_
timestamp 0
transform 1 0 3650 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__410_
timestamp 0
transform -1 0 3770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__411_
timestamp 0
transform -1 0 2470 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__412_
timestamp 0
transform 1 0 2690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__413_
timestamp 0
transform -1 0 3010 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__414_
timestamp 0
transform 1 0 2490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__415_
timestamp 0
transform 1 0 3030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__416_
timestamp 0
transform 1 0 3770 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__417_
timestamp 0
transform -1 0 3930 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__418_
timestamp 0
transform 1 0 4810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__419_
timestamp 0
transform 1 0 4550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__420_
timestamp 0
transform -1 0 4210 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__421_
timestamp 0
transform -1 0 4030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__422_
timestamp 0
transform -1 0 1690 0 1 730
box -6 -8 26 248
use FILL  FILL_6__423_
timestamp 0
transform 1 0 1430 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__424_
timestamp 0
transform 1 0 1390 0 1 730
box -6 -8 26 248
use FILL  FILL_6__425_
timestamp 0
transform 1 0 1430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__426_
timestamp 0
transform -1 0 3410 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__427_
timestamp 0
transform -1 0 2770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__428_
timestamp 0
transform -1 0 3150 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__429_
timestamp 0
transform 1 0 3250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__430_
timestamp 0
transform -1 0 3930 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__431_
timestamp 0
transform 1 0 4010 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__432_
timestamp 0
transform -1 0 3490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__433_
timestamp 0
transform -1 0 3750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__434_
timestamp 0
transform 1 0 4270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__435_
timestamp 0
transform 1 0 4750 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__436_
timestamp 0
transform 1 0 4850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__437_
timestamp 0
transform -1 0 4830 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__438_
timestamp 0
transform -1 0 4310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__439_
timestamp 0
transform -1 0 4290 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__440_
timestamp 0
transform -1 0 3490 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__441_
timestamp 0
transform -1 0 4030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__442_
timestamp 0
transform -1 0 4470 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__443_
timestamp 0
transform 1 0 4690 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__444_
timestamp 0
transform -1 0 4330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__445_
timestamp 0
transform -1 0 4830 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__446_
timestamp 0
transform 1 0 4790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__447_
timestamp 0
transform 1 0 4850 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__448_
timestamp 0
transform -1 0 4630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__449_
timestamp 0
transform 1 0 4190 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__450_
timestamp 0
transform 1 0 4590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__451_
timestamp 0
transform 1 0 4830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__452_
timestamp 0
transform 1 0 4710 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__453_
timestamp 0
transform 1 0 4870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__454_
timestamp 0
transform 1 0 4350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__455_
timestamp 0
transform -1 0 3830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__456_
timestamp 0
transform -1 0 4110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__457_
timestamp 0
transform 1 0 4070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__458_
timestamp 0
transform -1 0 3810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__459_
timestamp 0
transform -1 0 4810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__460_
timestamp 0
transform 1 0 4870 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__461_
timestamp 0
transform 1 0 4570 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__462_
timestamp 0
transform 1 0 4810 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__463_
timestamp 0
transform 1 0 4870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__464_
timestamp 0
transform 1 0 4290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__465_
timestamp 0
transform 1 0 4450 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__466_
timestamp 0
transform 1 0 4550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__467_
timestamp 0
transform 1 0 4590 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__468_
timestamp 0
transform 1 0 4290 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__469_
timestamp 0
transform -1 0 2990 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__470_
timestamp 0
transform -1 0 2450 0 1 730
box -6 -8 26 248
use FILL  FILL_6__471_
timestamp 0
transform -1 0 2650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__472_
timestamp 0
transform 1 0 2170 0 1 730
box -6 -8 26 248
use FILL  FILL_6__473_
timestamp 0
transform 1 0 2470 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__474_
timestamp 0
transform 1 0 2750 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__475_
timestamp 0
transform 1 0 3410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__476_
timestamp 0
transform 1 0 2890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__477_
timestamp 0
transform -1 0 2370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__478_
timestamp 0
transform -1 0 2250 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__479_
timestamp 0
transform -1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__480_
timestamp 0
transform 1 0 3250 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__481_
timestamp 0
transform -1 0 2750 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__482_
timestamp 0
transform 1 0 2850 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__483_
timestamp 0
transform -1 0 1410 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__484_
timestamp 0
transform -1 0 1130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__485_
timestamp 0
transform -1 0 1730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__486_
timestamp 0
transform -1 0 1710 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__487_
timestamp 0
transform -1 0 1450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__488_
timestamp 0
transform -1 0 1170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__489_
timestamp 0
transform -1 0 1990 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__490_
timestamp 0
transform 1 0 1690 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__491_
timestamp 0
transform 1 0 2790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__492_
timestamp 0
transform -1 0 3550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__493_
timestamp 0
transform 1 0 3050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__494_
timestamp 0
transform 1 0 3010 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__495_
timestamp 0
transform 1 0 2190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__496_
timestamp 0
transform 1 0 870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__497_
timestamp 0
transform -1 0 1650 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__498_
timestamp 0
transform 1 0 1010 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__499_
timestamp 0
transform 1 0 1390 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__500_
timestamp 0
transform -1 0 1890 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__501_
timestamp 0
transform 1 0 1230 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__502_
timestamp 0
transform -1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__503_
timestamp 0
transform 1 0 1690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__504_
timestamp 0
transform -1 0 2730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__505_
timestamp 0
transform -1 0 2990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__506_
timestamp 0
transform 1 0 3230 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__507_
timestamp 0
transform 1 0 2970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__508_
timestamp 0
transform -1 0 2870 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__509_
timestamp 0
transform 1 0 3210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__510_
timestamp 0
transform 1 0 3130 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__511_
timestamp 0
transform 1 0 2610 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__512_
timestamp 0
transform 1 0 1710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__513_
timestamp 0
transform -1 0 1530 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__514_
timestamp 0
transform 1 0 1570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__515_
timestamp 0
transform 1 0 1950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__516_
timestamp 0
transform 1 0 1790 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__517_
timestamp 0
transform -1 0 2090 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__518_
timestamp 0
transform -1 0 2790 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__519_
timestamp 0
transform 1 0 2510 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__520_
timestamp 0
transform 1 0 2430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__521_
timestamp 0
transform 1 0 2710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__522_
timestamp 0
transform -1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__523_
timestamp 0
transform 1 0 2310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__524_
timestamp 0
transform 1 0 4350 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__525_
timestamp 0
transform -1 0 4630 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__526_
timestamp 0
transform -1 0 4610 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__527_
timestamp 0
transform -1 0 4550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__528_
timestamp 0
transform -1 0 4290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__529_
timestamp 0
transform -1 0 4350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__530_
timestamp 0
transform 1 0 4310 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__531_
timestamp 0
transform -1 0 1830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__532_
timestamp 0
transform -1 0 950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__533_
timestamp 0
transform -1 0 3830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__534_
timestamp 0
transform -1 0 3270 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__535_
timestamp 0
transform -1 0 2590 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__536_
timestamp 0
transform 1 0 2230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__537_
timestamp 0
transform -1 0 1190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__538_
timestamp 0
transform 1 0 1970 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__539_
timestamp 0
transform 1 0 2470 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__540_
timestamp 0
transform 1 0 910 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__541_
timestamp 0
transform 1 0 1130 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__542_
timestamp 0
transform 1 0 1410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__543_
timestamp 0
transform -1 0 1150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__544_
timestamp 0
transform -1 0 670 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__545_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__546_
timestamp 0
transform -1 0 150 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__547_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__548_
timestamp 0
transform -1 0 410 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__549_
timestamp 0
transform -1 0 390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__550_
timestamp 0
transform -1 0 670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__551_
timestamp 0
transform 1 0 670 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__552_
timestamp 0
transform 1 0 910 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__553_
timestamp 0
transform 1 0 1170 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__554_
timestamp 0
transform 1 0 1450 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__555_
timestamp 0
transform -1 0 390 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__556_
timestamp 0
transform -1 0 150 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__557_
timestamp 0
transform -1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__558_
timestamp 0
transform 1 0 410 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__559_
timestamp 0
transform -1 0 150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__560_
timestamp 0
transform -1 0 950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__561_
timestamp 0
transform 1 0 650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__562_
timestamp 0
transform 1 0 950 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__563_
timestamp 0
transform -1 0 690 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__564_
timestamp 0
transform -1 0 150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__565_
timestamp 0
transform 1 0 130 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__566_
timestamp 0
transform 1 0 130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__567_
timestamp 0
transform 1 0 410 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__568_
timestamp 0
transform -1 0 690 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__569_
timestamp 0
transform -1 0 950 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__570_
timestamp 0
transform 1 0 910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__571_
timestamp 0
transform -1 0 670 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__572_
timestamp 0
transform -1 0 390 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__573_
timestamp 0
transform 1 0 390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__574_
timestamp 0
transform -1 0 410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__575_
timestamp 0
transform 1 0 630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__576_
timestamp 0
transform 1 0 650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__577_
timestamp 0
transform -1 0 150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__578_
timestamp 0
transform -1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__579_
timestamp 0
transform 1 0 630 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__580_
timestamp 0
transform -1 0 410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__581_
timestamp 0
transform -1 0 390 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__582_
timestamp 0
transform 1 0 890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__583_
timestamp 0
transform -1 0 670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__584_
timestamp 0
transform 1 0 490 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__585_
timestamp 0
transform -1 0 630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__586_
timestamp 0
transform -1 0 430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__587_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__588_
timestamp 0
transform -1 0 150 0 1 250
box -6 -8 26 248
use FILL  FILL_6__589_
timestamp 0
transform -1 0 150 0 1 730
box -6 -8 26 248
use FILL  FILL_6__590_
timestamp 0
transform -1 0 150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__591_
timestamp 0
transform -1 0 410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__592_
timestamp 0
transform -1 0 710 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__593_
timestamp 0
transform 1 0 410 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__594_
timestamp 0
transform -1 0 150 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__595_
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_6__596_
timestamp 0
transform 1 0 650 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__597_
timestamp 0
transform 1 0 630 0 1 730
box -6 -8 26 248
use FILL  FILL_6__598_
timestamp 0
transform 1 0 690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__599_
timestamp 0
transform 1 0 1250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__600_
timestamp 0
transform -1 0 150 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__601_
timestamp 0
transform -1 0 650 0 1 250
box -6 -8 26 248
use FILL  FILL_6__602_
timestamp 0
transform -1 0 910 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__603_
timestamp 0
transform 1 0 1530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__604_
timestamp 0
transform 1 0 1690 0 1 250
box -6 -8 26 248
use FILL  FILL_6__605_
timestamp 0
transform 1 0 1150 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__606_
timestamp 0
transform -1 0 1690 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__607_
timestamp 0
transform 1 0 1670 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__608_
timestamp 0
transform 1 0 1170 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__609_
timestamp 0
transform -1 0 1170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__610_
timestamp 0
transform 1 0 1390 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__611_
timestamp 0
transform -1 0 1470 0 1 250
box -6 -8 26 248
use FILL  FILL_6__612_
timestamp 0
transform 1 0 1170 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__613_
timestamp 0
transform 1 0 1930 0 1 250
box -6 -8 26 248
use FILL  FILL_6__614_
timestamp 0
transform 1 0 1930 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__615_
timestamp 0
transform 1 0 2210 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__616_
timestamp 0
transform 1 0 2450 0 1 250
box -6 -8 26 248
use FILL  FILL_6__617_
timestamp 0
transform 1 0 2470 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__618_
timestamp 0
transform 1 0 910 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__619_
timestamp 0
transform -1 0 410 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__620_
timestamp 0
transform 1 0 930 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__621_
timestamp 0
transform -1 0 690 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__622_
timestamp 0
transform -1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_6__623_
timestamp 0
transform 1 0 1170 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__624_
timestamp 0
transform 1 0 390 0 1 250
box -6 -8 26 248
use FILL  FILL_6__625_
timestamp 0
transform 1 0 390 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__665_
timestamp 0
transform 1 0 3410 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__666_
timestamp 0
transform 1 0 2770 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__667_
timestamp 0
transform -1 0 4330 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__668_
timestamp 0
transform 1 0 1990 0 1 4570
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert6
timestamp 0
transform -1 0 930 0 1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert7
timestamp 0
transform 1 0 2710 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert8
timestamp 0
transform 1 0 1450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert9
timestamp 0
transform 1 0 1190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert10
timestamp 0
transform -1 0 1950 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert11
timestamp 0
transform 1 0 2470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert12
timestamp 0
transform 1 0 1190 0 1 3130
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert13
timestamp 0
transform 1 0 2190 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert14
timestamp 0
transform -1 0 910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert15
timestamp 0
transform 1 0 2450 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert16
timestamp 0
transform 1 0 3290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert17
timestamp 0
transform 1 0 1930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert18
timestamp 0
transform 1 0 3210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert19
timestamp 0
transform 1 0 2090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert20
timestamp 0
transform 1 0 1810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert0
timestamp 0
transform 1 0 2090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert1
timestamp 0
transform -1 0 1730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert2
timestamp 0
transform 1 0 130 0 1 2170
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert3
timestamp 0
transform 1 0 1870 0 1 3610
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert4
timestamp 0
transform 1 0 1190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert5
timestamp 0
transform 1 0 1210 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__313_
timestamp 0
transform 1 0 1190 0 1 250
box -6 -8 26 248
use FILL  FILL_7__314_
timestamp 0
transform -1 0 1190 0 1 730
box -6 -8 26 248
use FILL  FILL_7__315_
timestamp 0
transform 1 0 910 0 1 730
box -6 -8 26 248
use FILL  FILL_7__316_
timestamp 0
transform -1 0 1010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__317_
timestamp 0
transform -1 0 2770 0 1 250
box -6 -8 26 248
use FILL  FILL_7__318_
timestamp 0
transform 1 0 3010 0 1 250
box -6 -8 26 248
use FILL  FILL_7__319_
timestamp 0
transform -1 0 3310 0 1 250
box -6 -8 26 248
use FILL  FILL_7__320_
timestamp 0
transform -1 0 3250 0 1 730
box -6 -8 26 248
use FILL  FILL_7__321_
timestamp 0
transform 1 0 3550 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__322_
timestamp 0
transform 1 0 2970 0 1 730
box -6 -8 26 248
use FILL  FILL_7__323_
timestamp 0
transform -1 0 3050 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__324_
timestamp 0
transform -1 0 2730 0 1 730
box -6 -8 26 248
use FILL  FILL_7__325_
timestamp 0
transform -1 0 3570 0 1 250
box -6 -8 26 248
use FILL  FILL_7__326_
timestamp 0
transform -1 0 3850 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__327_
timestamp 0
transform 1 0 4830 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__328_
timestamp 0
transform 1 0 4350 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__329_
timestamp 0
transform -1 0 4610 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__330_
timestamp 0
transform 1 0 4090 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__331_
timestamp 0
transform -1 0 3050 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__332_
timestamp 0
transform -1 0 2790 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__333_
timestamp 0
transform 1 0 2230 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__334_
timestamp 0
transform 1 0 2210 0 1 250
box -6 -8 26 248
use FILL  FILL_7__335_
timestamp 0
transform -1 0 1970 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__336_
timestamp 0
transform -1 0 3310 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__337_
timestamp 0
transform 1 0 3550 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__338_
timestamp 0
transform -1 0 4130 0 1 250
box -6 -8 26 248
use FILL  FILL_7__339_
timestamp 0
transform 1 0 3830 0 1 250
box -6 -8 26 248
use FILL  FILL_7__340_
timestamp 0
transform 1 0 4330 0 1 250
box -6 -8 26 248
use FILL  FILL_7__341_
timestamp 0
transform 1 0 4790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__342_
timestamp 0
transform 1 0 4870 0 1 250
box -6 -8 26 248
use FILL  FILL_7__343_
timestamp 0
transform -1 0 4890 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__344_
timestamp 0
transform -1 0 4630 0 1 250
box -6 -8 26 248
use FILL  FILL_7__345_
timestamp 0
transform -1 0 4610 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__346_
timestamp 0
transform 1 0 4290 0 1 730
box -6 -8 26 248
use FILL  FILL_7__347_
timestamp 0
transform -1 0 3510 0 1 730
box -6 -8 26 248
use FILL  FILL_7__348_
timestamp 0
transform -1 0 3790 0 1 730
box -6 -8 26 248
use FILL  FILL_7__349_
timestamp 0
transform 1 0 4810 0 1 730
box -6 -8 26 248
use FILL  FILL_7__350_
timestamp 0
transform 1 0 4550 0 1 730
box -6 -8 26 248
use FILL  FILL_7__351_
timestamp 0
transform 1 0 4590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__352_
timestamp 0
transform 1 0 4570 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__353_
timestamp 0
transform 1 0 4250 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__354_
timestamp 0
transform 1 0 4010 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__355_
timestamp 0
transform 1 0 4510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__356_
timestamp 0
transform -1 0 4250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__357_
timestamp 0
transform -1 0 3710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__358_
timestamp 0
transform -1 0 3970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__359_
timestamp 0
transform -1 0 3570 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__360_
timestamp 0
transform 1 0 4050 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__361_
timestamp 0
transform 1 0 4310 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__362_
timestamp 0
transform -1 0 4050 0 1 730
box -6 -8 26 248
use FILL  FILL_7__363_
timestamp 0
transform -1 0 5010 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__364_
timestamp 0
transform -1 0 4510 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__365_
timestamp 0
transform -1 0 3510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__366_
timestamp 0
transform -1 0 3570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__367_
timestamp 0
transform 1 0 4090 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__368_
timestamp 0
transform 1 0 4610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__369_
timestamp 0
transform 1 0 4090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__370_
timestamp 0
transform 1 0 3790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__371_
timestamp 0
transform 1 0 4070 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__372_
timestamp 0
transform 1 0 4090 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__373_
timestamp 0
transform -1 0 3830 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__374_
timestamp 0
transform -1 0 3850 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__375_
timestamp 0
transform 1 0 3810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__376_
timestamp 0
transform 1 0 3330 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__377_
timestamp 0
transform -1 0 3070 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__378_
timestamp 0
transform 1 0 3550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__379_
timestamp 0
transform -1 0 3290 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__380_
timestamp 0
transform -1 0 3570 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__381_
timestamp 0
transform -1 0 3310 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__382_
timestamp 0
transform 1 0 3270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__383_
timestamp 0
transform -1 0 3030 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__384_
timestamp 0
transform 1 0 3830 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__385_
timestamp 0
transform -1 0 3590 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__386_
timestamp 0
transform -1 0 2750 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__387_
timestamp 0
transform 1 0 2250 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__388_
timestamp 0
transform 1 0 2530 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__389_
timestamp 0
transform -1 0 3030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__390_
timestamp 0
transform -1 0 1950 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__391_
timestamp 0
transform -1 0 2750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__392_
timestamp 0
transform -1 0 2490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__393_
timestamp 0
transform 1 0 1730 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__394_
timestamp 0
transform -1 0 2210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__395_
timestamp 0
transform -1 0 1710 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__396_
timestamp 0
transform 1 0 2270 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__397_
timestamp 0
transform 1 0 2770 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__398_
timestamp 0
transform 1 0 2250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__399_
timestamp 0
transform 1 0 2530 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__400_
timestamp 0
transform -1 0 1930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__401_
timestamp 0
transform -1 0 2210 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__402_
timestamp 0
transform -1 0 2030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__403_
timestamp 0
transform 1 0 2450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__404_
timestamp 0
transform -1 0 2210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__405_
timestamp 0
transform 1 0 1610 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__406_
timestamp 0
transform -1 0 1650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__407_
timestamp 0
transform 1 0 3290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__408_
timestamp 0
transform -1 0 3010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__409_
timestamp 0
transform 1 0 3670 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__410_
timestamp 0
transform -1 0 3790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__411_
timestamp 0
transform -1 0 2490 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__412_
timestamp 0
transform 1 0 2710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__413_
timestamp 0
transform -1 0 3030 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__414_
timestamp 0
transform 1 0 2510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__415_
timestamp 0
transform 1 0 3050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__416_
timestamp 0
transform 1 0 3790 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__417_
timestamp 0
transform -1 0 3950 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__418_
timestamp 0
transform 1 0 4830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__419_
timestamp 0
transform 1 0 4570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__420_
timestamp 0
transform -1 0 4230 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__421_
timestamp 0
transform -1 0 4050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__422_
timestamp 0
transform -1 0 1710 0 1 730
box -6 -8 26 248
use FILL  FILL_7__423_
timestamp 0
transform 1 0 1450 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__424_
timestamp 0
transform 1 0 1410 0 1 730
box -6 -8 26 248
use FILL  FILL_7__425_
timestamp 0
transform 1 0 1450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__426_
timestamp 0
transform -1 0 3430 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__427_
timestamp 0
transform -1 0 2790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__428_
timestamp 0
transform -1 0 3170 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__429_
timestamp 0
transform 1 0 3270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__430_
timestamp 0
transform -1 0 3950 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__431_
timestamp 0
transform 1 0 4030 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__432_
timestamp 0
transform -1 0 3510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__433_
timestamp 0
transform -1 0 3770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__434_
timestamp 0
transform 1 0 4290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__435_
timestamp 0
transform 1 0 4770 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__436_
timestamp 0
transform 1 0 4870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__437_
timestamp 0
transform -1 0 4850 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__438_
timestamp 0
transform -1 0 4330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__439_
timestamp 0
transform -1 0 4310 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__440_
timestamp 0
transform -1 0 3510 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__441_
timestamp 0
transform -1 0 4050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__442_
timestamp 0
transform -1 0 4490 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__443_
timestamp 0
transform 1 0 4710 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__444_
timestamp 0
transform -1 0 4350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__445_
timestamp 0
transform -1 0 4850 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__446_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__447_
timestamp 0
transform 1 0 4870 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__448_
timestamp 0
transform -1 0 4650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__449_
timestamp 0
transform 1 0 4210 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__450_
timestamp 0
transform 1 0 4610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__451_
timestamp 0
transform 1 0 4850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__452_
timestamp 0
transform 1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__453_
timestamp 0
transform 1 0 4890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__454_
timestamp 0
transform 1 0 4370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__455_
timestamp 0
transform -1 0 3850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__456_
timestamp 0
transform -1 0 4130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__457_
timestamp 0
transform 1 0 4090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__458_
timestamp 0
transform -1 0 3830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__459_
timestamp 0
transform -1 0 4830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__460_
timestamp 0
transform 1 0 4890 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__461_
timestamp 0
transform 1 0 4590 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__462_
timestamp 0
transform 1 0 4830 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__463_
timestamp 0
transform 1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__464_
timestamp 0
transform 1 0 4310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__465_
timestamp 0
transform 1 0 4470 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__466_
timestamp 0
transform 1 0 4570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__467_
timestamp 0
transform 1 0 4610 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__468_
timestamp 0
transform 1 0 4310 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__469_
timestamp 0
transform -1 0 3010 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__470_
timestamp 0
transform -1 0 2470 0 1 730
box -6 -8 26 248
use FILL  FILL_7__471_
timestamp 0
transform -1 0 2670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__472_
timestamp 0
transform 1 0 2190 0 1 730
box -6 -8 26 248
use FILL  FILL_7__473_
timestamp 0
transform 1 0 2490 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__474_
timestamp 0
transform 1 0 2770 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__475_
timestamp 0
transform 1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__476_
timestamp 0
transform 1 0 2910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__477_
timestamp 0
transform -1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__478_
timestamp 0
transform -1 0 2270 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__479_
timestamp 0
transform -1 0 3330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__480_
timestamp 0
transform 1 0 3270 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__481_
timestamp 0
transform -1 0 2770 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__482_
timestamp 0
transform 1 0 2870 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__483_
timestamp 0
transform -1 0 1430 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__484_
timestamp 0
transform -1 0 1150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__485_
timestamp 0
transform -1 0 1750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__486_
timestamp 0
transform -1 0 1730 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__487_
timestamp 0
transform -1 0 1470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__488_
timestamp 0
transform -1 0 1190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__489_
timestamp 0
transform -1 0 2010 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__490_
timestamp 0
transform 1 0 1710 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__491_
timestamp 0
transform 1 0 2810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__492_
timestamp 0
transform -1 0 3570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__493_
timestamp 0
transform 1 0 3070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__494_
timestamp 0
transform 1 0 3030 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__495_
timestamp 0
transform 1 0 2210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__496_
timestamp 0
transform 1 0 890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__497_
timestamp 0
transform -1 0 1670 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__498_
timestamp 0
transform 1 0 1030 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__499_
timestamp 0
transform 1 0 1410 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__500_
timestamp 0
transform -1 0 1910 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__501_
timestamp 0
transform 1 0 1250 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__502_
timestamp 0
transform -1 0 1470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__503_
timestamp 0
transform 1 0 1710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__504_
timestamp 0
transform -1 0 2750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__505_
timestamp 0
transform -1 0 3010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__506_
timestamp 0
transform 1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__507_
timestamp 0
transform 1 0 2990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__508_
timestamp 0
transform -1 0 2890 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__509_
timestamp 0
transform 1 0 3230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__510_
timestamp 0
transform 1 0 3150 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__511_
timestamp 0
transform 1 0 2630 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__512_
timestamp 0
transform 1 0 1730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__513_
timestamp 0
transform -1 0 1550 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__514_
timestamp 0
transform 1 0 1590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__515_
timestamp 0
transform 1 0 1970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__516_
timestamp 0
transform 1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__517_
timestamp 0
transform -1 0 2110 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__518_
timestamp 0
transform -1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__519_
timestamp 0
transform 1 0 2530 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__520_
timestamp 0
transform 1 0 2450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__521_
timestamp 0
transform 1 0 2730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__522_
timestamp 0
transform -1 0 2750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__523_
timestamp 0
transform 1 0 2330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__524_
timestamp 0
transform 1 0 4370 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__525_
timestamp 0
transform -1 0 4650 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__526_
timestamp 0
transform -1 0 4630 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__527_
timestamp 0
transform -1 0 4570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__528_
timestamp 0
transform -1 0 4310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__529_
timestamp 0
transform -1 0 4370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__530_
timestamp 0
transform 1 0 4330 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__531_
timestamp 0
transform -1 0 1850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__532_
timestamp 0
transform -1 0 970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__533_
timestamp 0
transform -1 0 3850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__534_
timestamp 0
transform -1 0 3290 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__535_
timestamp 0
transform -1 0 2610 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__536_
timestamp 0
transform 1 0 2250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__537_
timestamp 0
transform -1 0 1210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__538_
timestamp 0
transform 1 0 1990 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__539_
timestamp 0
transform 1 0 2490 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__540_
timestamp 0
transform 1 0 930 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__541_
timestamp 0
transform 1 0 1150 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__542_
timestamp 0
transform 1 0 1430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__543_
timestamp 0
transform -1 0 1170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__544_
timestamp 0
transform -1 0 690 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__545_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__546_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__547_
timestamp 0
transform -1 0 170 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__548_
timestamp 0
transform -1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__549_
timestamp 0
transform -1 0 410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__550_
timestamp 0
transform -1 0 690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__551_
timestamp 0
transform 1 0 690 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__552_
timestamp 0
transform 1 0 930 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__553_
timestamp 0
transform 1 0 1190 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__554_
timestamp 0
transform 1 0 1470 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__555_
timestamp 0
transform -1 0 410 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__556_
timestamp 0
transform -1 0 170 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__557_
timestamp 0
transform -1 0 170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__558_
timestamp 0
transform 1 0 430 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__559_
timestamp 0
transform -1 0 170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__560_
timestamp 0
transform -1 0 970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__561_
timestamp 0
transform 1 0 670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__562_
timestamp 0
transform 1 0 970 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__563_
timestamp 0
transform -1 0 710 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__564_
timestamp 0
transform -1 0 170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__565_
timestamp 0
transform 1 0 150 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__566_
timestamp 0
transform 1 0 150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__567_
timestamp 0
transform 1 0 430 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__568_
timestamp 0
transform -1 0 710 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__569_
timestamp 0
transform -1 0 970 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__570_
timestamp 0
transform 1 0 930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__571_
timestamp 0
transform -1 0 690 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__572_
timestamp 0
transform -1 0 410 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__573_
timestamp 0
transform 1 0 410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__574_
timestamp 0
transform -1 0 430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__575_
timestamp 0
transform 1 0 650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__576_
timestamp 0
transform 1 0 670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__577_
timestamp 0
transform -1 0 170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__578_
timestamp 0
transform -1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__579_
timestamp 0
transform 1 0 650 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__580_
timestamp 0
transform -1 0 430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__581_
timestamp 0
transform -1 0 410 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__582_
timestamp 0
transform 1 0 910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__583_
timestamp 0
transform -1 0 690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__584_
timestamp 0
transform 1 0 510 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__585_
timestamp 0
transform -1 0 650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__586_
timestamp 0
transform -1 0 450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__587_
timestamp 0
transform -1 0 170 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__588_
timestamp 0
transform -1 0 170 0 1 250
box -6 -8 26 248
use FILL  FILL_7__589_
timestamp 0
transform -1 0 170 0 1 730
box -6 -8 26 248
use FILL  FILL_7__590_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__591_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__592_
timestamp 0
transform -1 0 730 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__593_
timestamp 0
transform 1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__594_
timestamp 0
transform -1 0 170 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__595_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 26 248
use FILL  FILL_7__596_
timestamp 0
transform 1 0 670 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__597_
timestamp 0
transform 1 0 650 0 1 730
box -6 -8 26 248
use FILL  FILL_7__598_
timestamp 0
transform 1 0 710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__599_
timestamp 0
transform 1 0 1270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__600_
timestamp 0
transform -1 0 170 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__601_
timestamp 0
transform -1 0 670 0 1 250
box -6 -8 26 248
use FILL  FILL_7__602_
timestamp 0
transform -1 0 930 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__603_
timestamp 0
transform 1 0 1550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__604_
timestamp 0
transform 1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_7__605_
timestamp 0
transform 1 0 1170 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__606_
timestamp 0
transform -1 0 1710 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__607_
timestamp 0
transform 1 0 1690 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__608_
timestamp 0
transform 1 0 1190 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__609_
timestamp 0
transform -1 0 1190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__610_
timestamp 0
transform 1 0 1410 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__611_
timestamp 0
transform -1 0 1490 0 1 250
box -6 -8 26 248
use FILL  FILL_7__612_
timestamp 0
transform 1 0 1190 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__613_
timestamp 0
transform 1 0 1950 0 1 250
box -6 -8 26 248
use FILL  FILL_7__614_
timestamp 0
transform 1 0 1950 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__615_
timestamp 0
transform 1 0 2230 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__616_
timestamp 0
transform 1 0 2470 0 1 250
box -6 -8 26 248
use FILL  FILL_7__617_
timestamp 0
transform 1 0 2490 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__618_
timestamp 0
transform 1 0 930 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__619_
timestamp 0
transform -1 0 430 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__620_
timestamp 0
transform 1 0 950 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__621_
timestamp 0
transform -1 0 710 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__622_
timestamp 0
transform -1 0 930 0 1 250
box -6 -8 26 248
use FILL  FILL_7__623_
timestamp 0
transform 1 0 1190 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__624_
timestamp 0
transform 1 0 410 0 1 250
box -6 -8 26 248
use FILL  FILL_7__625_
timestamp 0
transform 1 0 410 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__665_
timestamp 0
transform 1 0 3430 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__666_
timestamp 0
transform 1 0 2790 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__667_
timestamp 0
transform -1 0 4350 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__668_
timestamp 0
transform 1 0 2010 0 1 4570
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert6
timestamp 0
transform -1 0 950 0 1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert7
timestamp 0
transform 1 0 2730 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert8
timestamp 0
transform 1 0 1470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert9
timestamp 0
transform 1 0 1210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert10
timestamp 0
transform -1 0 1970 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert11
timestamp 0
transform 1 0 2490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert12
timestamp 0
transform 1 0 1210 0 1 3130
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert13
timestamp 0
transform 1 0 2210 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert14
timestamp 0
transform -1 0 930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert15
timestamp 0
transform 1 0 2470 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert16
timestamp 0
transform 1 0 3310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert17
timestamp 0
transform 1 0 1950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert18
timestamp 0
transform 1 0 3230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert19
timestamp 0
transform 1 0 2110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert20
timestamp 0
transform 1 0 1830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert0
timestamp 0
transform 1 0 2110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert1
timestamp 0
transform -1 0 1750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert2
timestamp 0
transform 1 0 150 0 1 2170
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert3
timestamp 0
transform 1 0 1890 0 1 3610
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert4
timestamp 0
transform 1 0 1210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert5
timestamp 0
transform 1 0 1230 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__313_
timestamp 0
transform 1 0 1210 0 1 250
box -6 -8 26 248
use FILL  FILL_8__314_
timestamp 0
transform -1 0 1210 0 1 730
box -6 -8 26 248
use FILL  FILL_8__316_
timestamp 0
transform -1 0 1030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__317_
timestamp 0
transform -1 0 2790 0 1 250
box -6 -8 26 248
use FILL  FILL_8__318_
timestamp 0
transform 1 0 3030 0 1 250
box -6 -8 26 248
use FILL  FILL_8__319_
timestamp 0
transform -1 0 3330 0 1 250
box -6 -8 26 248
use FILL  FILL_8__321_
timestamp 0
transform 1 0 3570 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__322_
timestamp 0
transform 1 0 2990 0 1 730
box -6 -8 26 248
use FILL  FILL_8__323_
timestamp 0
transform -1 0 3070 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__325_
timestamp 0
transform -1 0 3590 0 1 250
box -6 -8 26 248
use FILL  FILL_8__326_
timestamp 0
transform -1 0 3870 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__327_
timestamp 0
transform 1 0 4850 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__328_
timestamp 0
transform 1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__330_
timestamp 0
transform 1 0 4110 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__331_
timestamp 0
transform -1 0 3070 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__332_
timestamp 0
transform -1 0 2810 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__333_
timestamp 0
transform 1 0 2250 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__335_
timestamp 0
transform -1 0 1990 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__336_
timestamp 0
transform -1 0 3330 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__337_
timestamp 0
transform 1 0 3570 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__339_
timestamp 0
transform 1 0 3850 0 1 250
box -6 -8 26 248
use FILL  FILL_8__340_
timestamp 0
transform 1 0 4350 0 1 250
box -6 -8 26 248
use FILL  FILL_8__341_
timestamp 0
transform 1 0 4810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__342_
timestamp 0
transform 1 0 4890 0 1 250
box -6 -8 26 248
use FILL  FILL_8__344_
timestamp 0
transform -1 0 4650 0 1 250
box -6 -8 26 248
use FILL  FILL_8__345_
timestamp 0
transform -1 0 4630 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__346_
timestamp 0
transform 1 0 4310 0 1 730
box -6 -8 26 248
use FILL  FILL_8__347_
timestamp 0
transform -1 0 3530 0 1 730
box -6 -8 26 248
use FILL  FILL_8__349_
timestamp 0
transform 1 0 4830 0 1 730
box -6 -8 26 248
use FILL  FILL_8__350_
timestamp 0
transform 1 0 4570 0 1 730
box -6 -8 26 248
use FILL  FILL_8__351_
timestamp 0
transform 1 0 4610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__352_
timestamp 0
transform 1 0 4590 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__354_
timestamp 0
transform 1 0 4030 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__355_
timestamp 0
transform 1 0 4530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__356_
timestamp 0
transform -1 0 4270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__358_
timestamp 0
transform -1 0 3990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__359_
timestamp 0
transform -1 0 3590 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__360_
timestamp 0
transform 1 0 4070 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__361_
timestamp 0
transform 1 0 4330 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__363_
timestamp 0
transform -1 0 5030 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__364_
timestamp 0
transform -1 0 4530 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__365_
timestamp 0
transform -1 0 3530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__366_
timestamp 0
transform -1 0 3590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__368_
timestamp 0
transform 1 0 4630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__369_
timestamp 0
transform 1 0 4110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__370_
timestamp 0
transform 1 0 3810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__372_
timestamp 0
transform 1 0 4110 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__373_
timestamp 0
transform -1 0 3850 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__374_
timestamp 0
transform -1 0 3870 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__375_
timestamp 0
transform 1 0 3830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__377_
timestamp 0
transform -1 0 3090 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__378_
timestamp 0
transform 1 0 3570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__379_
timestamp 0
transform -1 0 3310 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__380_
timestamp 0
transform -1 0 3590 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__382_
timestamp 0
transform 1 0 3290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__383_
timestamp 0
transform -1 0 3050 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__384_
timestamp 0
transform 1 0 3850 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__386_
timestamp 0
transform -1 0 2770 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__387_
timestamp 0
transform 1 0 2270 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__388_
timestamp 0
transform 1 0 2550 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__389_
timestamp 0
transform -1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__391_
timestamp 0
transform -1 0 2770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__392_
timestamp 0
transform -1 0 2510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__393_
timestamp 0
transform 1 0 1750 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__394_
timestamp 0
transform -1 0 2230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__396_
timestamp 0
transform 1 0 2290 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__397_
timestamp 0
transform 1 0 2790 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__398_
timestamp 0
transform 1 0 2270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__400_
timestamp 0
transform -1 0 1950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__401_
timestamp 0
transform -1 0 2230 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__402_
timestamp 0
transform -1 0 2050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__403_
timestamp 0
transform 1 0 2470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__405_
timestamp 0
transform 1 0 1630 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__406_
timestamp 0
transform -1 0 1670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__407_
timestamp 0
transform 1 0 3310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__408_
timestamp 0
transform -1 0 3030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__410_
timestamp 0
transform -1 0 3810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__411_
timestamp 0
transform -1 0 2510 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__412_
timestamp 0
transform 1 0 2730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__413_
timestamp 0
transform -1 0 3050 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__415_
timestamp 0
transform 1 0 3070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__416_
timestamp 0
transform 1 0 3810 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__417_
timestamp 0
transform -1 0 3970 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__419_
timestamp 0
transform 1 0 4590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__420_
timestamp 0
transform -1 0 4250 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__421_
timestamp 0
transform -1 0 4070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__422_
timestamp 0
transform -1 0 1730 0 1 730
box -6 -8 26 248
use FILL  FILL_8__424_
timestamp 0
transform 1 0 1430 0 1 730
box -6 -8 26 248
use FILL  FILL_8__425_
timestamp 0
transform 1 0 1470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__426_
timestamp 0
transform -1 0 3450 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__427_
timestamp 0
transform -1 0 2810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__429_
timestamp 0
transform 1 0 3290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__430_
timestamp 0
transform -1 0 3970 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__431_
timestamp 0
transform 1 0 4050 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__433_
timestamp 0
transform -1 0 3790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__434_
timestamp 0
transform 1 0 4310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__435_
timestamp 0
transform 1 0 4790 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__436_
timestamp 0
transform 1 0 4890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__438_
timestamp 0
transform -1 0 4350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__439_
timestamp 0
transform -1 0 4330 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__440_
timestamp 0
transform -1 0 3530 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__441_
timestamp 0
transform -1 0 4070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__443_
timestamp 0
transform 1 0 4730 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__444_
timestamp 0
transform -1 0 4370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__445_
timestamp 0
transform -1 0 4870 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__447_
timestamp 0
transform 1 0 4890 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__448_
timestamp 0
transform -1 0 4670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__449_
timestamp 0
transform 1 0 4230 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__450_
timestamp 0
transform 1 0 4630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__452_
timestamp 0
transform 1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__453_
timestamp 0
transform 1 0 4910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__454_
timestamp 0
transform 1 0 4390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__455_
timestamp 0
transform -1 0 3870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__457_
timestamp 0
transform 1 0 4110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__458_
timestamp 0
transform -1 0 3850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__459_
timestamp 0
transform -1 0 4850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__460_
timestamp 0
transform 1 0 4910 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__462_
timestamp 0
transform 1 0 4850 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__463_
timestamp 0
transform 1 0 4910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__464_
timestamp 0
transform 1 0 4330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__466_
timestamp 0
transform 1 0 4590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__467_
timestamp 0
transform 1 0 4630 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__468_
timestamp 0
transform 1 0 4330 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__469_
timestamp 0
transform -1 0 3030 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__471_
timestamp 0
transform -1 0 2690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__472_
timestamp 0
transform 1 0 2210 0 1 730
box -6 -8 26 248
use FILL  FILL_8__473_
timestamp 0
transform 1 0 2510 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__474_
timestamp 0
transform 1 0 2790 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__476_
timestamp 0
transform 1 0 2930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__477_
timestamp 0
transform -1 0 2410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__478_
timestamp 0
transform -1 0 2290 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__480_
timestamp 0
transform 1 0 3290 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__481_
timestamp 0
transform -1 0 2790 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__482_
timestamp 0
transform 1 0 2890 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__483_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__485_
timestamp 0
transform -1 0 1770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__486_
timestamp 0
transform -1 0 1750 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__487_
timestamp 0
transform -1 0 1490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__488_
timestamp 0
transform -1 0 1210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__490_
timestamp 0
transform 1 0 1730 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__491_
timestamp 0
transform 1 0 2830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__492_
timestamp 0
transform -1 0 3590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__494_
timestamp 0
transform 1 0 3050 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__495_
timestamp 0
transform 1 0 2230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__496_
timestamp 0
transform 1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__497_
timestamp 0
transform -1 0 1690 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__499_
timestamp 0
transform 1 0 1430 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__500_
timestamp 0
transform -1 0 1930 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__501_
timestamp 0
transform 1 0 1270 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__502_
timestamp 0
transform -1 0 1490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__504_
timestamp 0
transform -1 0 2770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__505_
timestamp 0
transform -1 0 3030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__506_
timestamp 0
transform 1 0 3270 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__508_
timestamp 0
transform -1 0 2910 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__509_
timestamp 0
transform 1 0 3250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__510_
timestamp 0
transform 1 0 3170 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__511_
timestamp 0
transform 1 0 2650 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__513_
timestamp 0
transform -1 0 1570 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__514_
timestamp 0
transform 1 0 1610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__515_
timestamp 0
transform 1 0 1990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__516_
timestamp 0
transform 1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__518_
timestamp 0
transform -1 0 2830 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__519_
timestamp 0
transform 1 0 2550 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__520_
timestamp 0
transform 1 0 2470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__521_
timestamp 0
transform 1 0 2750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__523_
timestamp 0
transform 1 0 2350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__524_
timestamp 0
transform 1 0 4390 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__525_
timestamp 0
transform -1 0 4670 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__527_
timestamp 0
transform -1 0 4590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__528_
timestamp 0
transform -1 0 4330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__529_
timestamp 0
transform -1 0 4390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__530_
timestamp 0
transform 1 0 4350 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__532_
timestamp 0
transform -1 0 990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__533_
timestamp 0
transform -1 0 3870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__534_
timestamp 0
transform -1 0 3310 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__535_
timestamp 0
transform -1 0 2630 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__537_
timestamp 0
transform -1 0 1230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__538_
timestamp 0
transform 1 0 2010 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__539_
timestamp 0
transform 1 0 2510 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__541_
timestamp 0
transform 1 0 1170 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__542_
timestamp 0
transform 1 0 1450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__543_
timestamp 0
transform -1 0 1190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__544_
timestamp 0
transform -1 0 710 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__546_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__547_
timestamp 0
transform -1 0 190 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__548_
timestamp 0
transform -1 0 450 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__549_
timestamp 0
transform -1 0 430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__551_
timestamp 0
transform 1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__552_
timestamp 0
transform 1 0 950 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__553_
timestamp 0
transform 1 0 1210 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__555_
timestamp 0
transform -1 0 430 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__556_
timestamp 0
transform -1 0 190 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__557_
timestamp 0
transform -1 0 190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__558_
timestamp 0
transform 1 0 450 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__560_
timestamp 0
transform -1 0 990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__561_
timestamp 0
transform 1 0 690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__562_
timestamp 0
transform 1 0 990 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__563_
timestamp 0
transform -1 0 730 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__565_
timestamp 0
transform 1 0 170 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__566_
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__567_
timestamp 0
transform 1 0 450 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__569_
timestamp 0
transform -1 0 990 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__570_
timestamp 0
transform 1 0 950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__571_
timestamp 0
transform -1 0 710 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__572_
timestamp 0
transform -1 0 430 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__574_
timestamp 0
transform -1 0 450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__575_
timestamp 0
transform 1 0 670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__576_
timestamp 0
transform 1 0 690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__577_
timestamp 0
transform -1 0 190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__579_
timestamp 0
transform 1 0 670 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__580_
timestamp 0
transform -1 0 450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__581_
timestamp 0
transform -1 0 430 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__582_
timestamp 0
transform 1 0 930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__584_
timestamp 0
transform 1 0 530 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__585_
timestamp 0
transform -1 0 670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__586_
timestamp 0
transform -1 0 470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__588_
timestamp 0
transform -1 0 190 0 1 250
box -6 -8 26 248
use FILL  FILL_8__589_
timestamp 0
transform -1 0 190 0 1 730
box -6 -8 26 248
use FILL  FILL_8__590_
timestamp 0
transform -1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__591_
timestamp 0
transform -1 0 450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__593_
timestamp 0
transform 1 0 450 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__594_
timestamp 0
transform -1 0 190 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__595_
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_8__596_
timestamp 0
transform 1 0 690 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__598_
timestamp 0
transform 1 0 730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__599_
timestamp 0
transform 1 0 1290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__600_
timestamp 0
transform -1 0 190 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__602_
timestamp 0
transform -1 0 950 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__603_
timestamp 0
transform 1 0 1570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__604_
timestamp 0
transform 1 0 1730 0 1 250
box -6 -8 26 248
use FILL  FILL_8__605_
timestamp 0
transform 1 0 1190 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__607_
timestamp 0
transform 1 0 1710 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__608_
timestamp 0
transform 1 0 1210 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__609_
timestamp 0
transform -1 0 1210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__610_
timestamp 0
transform 1 0 1430 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__612_
timestamp 0
transform 1 0 1210 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__613_
timestamp 0
transform 1 0 1970 0 1 250
box -6 -8 26 248
use FILL  FILL_8__614_
timestamp 0
transform 1 0 1970 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__616_
timestamp 0
transform 1 0 2490 0 1 250
box -6 -8 26 248
use FILL  FILL_8__617_
timestamp 0
transform 1 0 2510 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__618_
timestamp 0
transform 1 0 950 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__619_
timestamp 0
transform -1 0 450 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__621_
timestamp 0
transform -1 0 730 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__622_
timestamp 0
transform -1 0 950 0 1 250
box -6 -8 26 248
use FILL  FILL_8__623_
timestamp 0
transform 1 0 1210 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__624_
timestamp 0
transform 1 0 430 0 1 250
box -6 -8 26 248
use FILL  FILL_8__665_
timestamp 0
transform 1 0 3450 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__666_
timestamp 0
transform 1 0 2810 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__667_
timestamp 0
transform -1 0 4370 0 1 4570
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert7
timestamp 0
transform 1 0 2750 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert8
timestamp 0
transform 1 0 1490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert9
timestamp 0
transform 1 0 1230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert10
timestamp 0
transform -1 0 1990 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert12
timestamp 0
transform 1 0 1230 0 1 3130
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert13
timestamp 0
transform 1 0 2230 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert14
timestamp 0
transform -1 0 950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert15
timestamp 0
transform 1 0 2490 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert17
timestamp 0
transform 1 0 1970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert18
timestamp 0
transform 1 0 3250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert19
timestamp 0
transform 1 0 2130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert20
timestamp 0
transform 1 0 1850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert0
timestamp 0
transform 1 0 2130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert1
timestamp 0
transform -1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert3
timestamp 0
transform 1 0 1910 0 1 3610
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert4
timestamp 0
transform 1 0 1230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert5
timestamp 0
transform 1 0 1250 0 1 3610
box -6 -8 26 248
<< labels >>
flabel metal1 s 5102 2 5162 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 4397 4857 4403 4863 3 FreeSans 16 90 0 0 Aout[1]
port 2 nsew
flabel metal2 s 4357 4857 4363 4863 3 FreeSans 16 90 0 0 Aout[0]
port 3 nsew
flabel metal3 s -24 2336 -16 2344 7 FreeSans 16 0 0 0 En
port 4 nsew
flabel metal2 s 4637 4857 4643 4863 3 FreeSans 16 90 0 0 FCW[19]
port 5 nsew
flabel metal2 s 4897 4857 4903 4863 3 FreeSans 16 90 0 0 FCW[18]
port 6 nsew
flabel metal3 s 5136 1556 5144 1564 3 FreeSans 16 0 0 0 FCW[17]
port 7 nsew
flabel metal3 s 5136 2036 5144 2044 3 FreeSans 16 0 0 0 FCW[16]
port 8 nsew
flabel metal3 s 5136 3716 5144 3724 3 FreeSans 16 0 0 0 FCW[15]
port 9 nsew
flabel metal3 s 5136 4676 5144 4684 3 FreeSans 16 0 0 0 FCW[14]
port 10 nsew
flabel metal3 s 5136 4716 5144 4724 3 FreeSans 16 0 0 0 FCW[13]
port 11 nsew
flabel metal3 s 5136 4756 5144 4764 3 FreeSans 16 0 0 0 FCW[12]
port 12 nsew
flabel metal3 s 5136 4796 5144 4804 3 FreeSans 16 90 0 0 FCW[11]
port 13 nsew
flabel metal2 s 4877 -23 4883 -17 7 FreeSans 16 270 0 0 FCW[10]
port 14 nsew
flabel metal2 s 3817 -23 3823 -17 7 FreeSans 16 270 0 0 FCW[9]
port 15 nsew
flabel metal2 s 2997 -23 3003 -17 7 FreeSans 16 270 0 0 FCW[8]
port 16 nsew
flabel metal2 s 497 -23 503 -17 7 FreeSans 16 270 0 0 FCW[7]
port 17 nsew
flabel metal2 s 237 -23 243 -17 7 FreeSans 16 270 0 0 FCW[6]
port 18 nsew
flabel metal2 s 197 -23 203 -17 7 FreeSans 16 270 0 0 FCW[5]
port 19 nsew
flabel metal2 s 157 -23 163 -17 7 FreeSans 16 270 0 0 FCW[4]
port 20 nsew
flabel metal3 s -24 4536 -16 4544 7 FreeSans 16 0 0 0 FCW[3]
port 21 nsew
flabel metal3 s -24 4496 -16 4504 7 FreeSans 16 0 0 0 FCW[2]
port 22 nsew
flabel metal3 s -24 4456 -16 4464 7 FreeSans 16 0 0 0 FCW[1]
port 23 nsew
flabel metal3 s -24 4196 -16 4204 7 FreeSans 16 0 0 0 FCW[0]
port 24 nsew
flabel metal2 s 4317 4857 4323 4863 3 FreeSans 16 90 0 0 ISout
port 25 nsew
flabel metal2 s 2057 4857 2063 4863 3 FreeSans 16 90 0 0 Vld
port 26 nsew
flabel metal3 s -24 2296 -16 2304 7 FreeSans 16 0 0 0 clk
port 27 nsew
<< properties >>
string FIXED_BBOX -40 -40 5140 4860
<< end >>
