//      // verilator_coverage annotation
        module cordic_element ( 
        	//timing issue
 003231 	input 			clk,
 000822 	input 	[1:0] 	Xin,
 000836 	output 	[1:0] 	Xout,
 000799 	input 	[1:0] 	Yin,
 000857 	output 	[1:0] 	Yout,
 000815 	input 	[1:0]	Ain,
 000816 	output 	[1:0]	Aout, //13
 000792 	input 			ISin, 
 000107 	output	reg		ISout, //15
%000007 	input	[2:0]	Stg, //20
 000462 	input 			Rdy, 
 000460 	output 			Vld //24
        );
%000001 	reg signed [11:0] oneOverK = 12'd1242;
%000001 	reg signed [11:0] atan0 = 12'd511;//44.96 degree
%000001 	reg signed [11:0] atan1 = 12'd301;//26.50 degree
%000001 	reg signed [11:0] atan2 = 12'd159;//14.02 degree
%000001 	reg signed [11:0] atan3 = 12'd80; // 7.07 degree
%000001 	reg signed [11:0] atan4 = 12'd40; // 3.56 degree
%000001 	reg signed [11:0] atan5 = 12'd19; // 1.71 degree
%000001 	reg signed [11:0] atan6 = 12'd9;  // 0.83 degree
%000001 	reg signed [11:0] atan7 = 12'd4;  // 0.39 degree
        	
        	// Load Control -----------------------------------------------------------
        	integer i;
 000462     reg     [6:0]   LoadCtl;
 001616     always @(posedge clk)
 001616     begin
 001616         LoadCtl[0] <= Rdy;
 009696         for (i=0; i<6; i=i+1)
 009696             LoadCtl[i+1] <= LoadCtl[i];
            end
        	assign Vld = LoadCtl[6];
        	
        	// Invert Sign ------------------------------------------------------------
 001616 	always @(posedge clk) if(LoadCtl[6]) ISout <= ISin;    
        	
        	// Loading Xin, Yin, Ain --------------------------------------------------
 000126 	reg [1:0] Xin5, Xin4, Xin3, Xin2, Xin1, Xin0;
 000119 	reg [1:0] Yin5, Yin4, Yin3, Yin2, Yin1, Yin0;
 000126 	reg [1:0] Ain5, Ain4, Ain3, Ain2, Ain1, Ain0;
        	
 001616 	always @(posedge clk) begin
 000231         if 		(LoadCtl[0]) begin Xin0 <= Xin; Yin0 <= Yin; Ain0 <= Ain; end
 000231         else if (LoadCtl[1]) begin Xin1 <= Xin; Yin1 <= Yin; Ain1 <= Ain; end
 000231 		else if (LoadCtl[2]) begin Xin2 <= Xin; Yin2 <= Yin; Ain2 <= Ain; end
 000231         else if (LoadCtl[3]) begin Xin3 <= Xin; Yin3 <= Yin; Ain3 <= Ain; end
 000230 		else if (LoadCtl[4]) begin Xin4 <= Xin; Yin4 <= Yin; Ain4 <= Ain; end
 000232         else if (LoadCtl[5]) begin Xin5 <= Xin; Yin5 <= Yin; Ain5 <= Ain; end
            end
        	
        	// atan mapping ----------------------------------------------------------
%000006 	reg signed [11:0] atan;
        	
 004839 	always@* begin
 004839 		case(Stg)
 000624 			3'd0:atan = atan0;
 000602 			3'd1:atan = atan1;
 000603 			3'd2:atan = atan2;
 000603 			3'd3:atan = atan3;
 000601 			3'd4:atan = atan4;
 000603 			3'd5:atan = atan5;
 000600 			3'd6:atan = atan6;
 000603 			3'd7:atan = atan7;
        		endcase
        	end
        	
        	// cordic element(shift & add/sub) ---------------------------------------
 000126 	wire signed [11:0] Xin12b = {Xin5, Xin4, Xin3, Xin2, Xin1, Xin0}; 
 000119 	wire signed [11:0] Yin12b = {Yin5, Yin4, Yin3, Yin2, Yin1, Yin0};
 000126 	wire signed [11:0] Ain12b = {Ain5, Ain4, Ain3, Ain2, Ain1, Ain0};
        
 000127 	reg signed [11:0] Xcalc, Ycalc, Acalc;
 001616 	always@(posedge clk) begin
 001386 		if (LoadCtl[6]) begin
 000201 			if(Stg != 3'd0) begin
 000106 				if(Ain12b[11] == 0) begin //postive angle
 000095 					Xcalc <= Xin12b - ( Yin12b >>> Stg );
 000095 					Ycalc <= Yin12b + ( Xin12b >>> Stg );
 000095 					Acalc <= Ain12b - atan;
        				end
 000106 				else begin
 000106 					Xcalc <= Xin12b + ( Yin12b >>> Stg );
 000106 					Ycalc <= Yin12b - ( Xin12b >>> Stg );
 000106 					Acalc <= Ain12b + atan;
        				end
        			end
 000029 			else begin // Stg == 0
 000019 				if(Ain12b[11] == 0) begin //postive angle
 000010 					Xcalc <= oneOverK;
 000010 					Ycalc <= oneOverK;
 000010 					Acalc <= Ain12b - atan;
        				end
 000019 				else begin
 000019 					Xcalc <= oneOverK;
 000019 					Ycalc <= -oneOverK;
 000019 					Acalc <= Ain12b + atan;
        				end
        			end
        		end
        	end
        	
        	// X, Y, A Output -------------------------------------------------------
 000857 	reg [1:0] X_, Y_, A_;
 001617 	always@* begin
 000231 		if 		(LoadCtl[0]) begin X_ = Xcalc[1:0]  ; Y_ = Ycalc[1:0]  ; A_ = Acalc[1:0]  ; end
 000231 		else if (LoadCtl[1]) begin X_ = Xcalc[3:2]  ; Y_ = Ycalc[3:2]  ; A_ = Acalc[3:2]  ; end
 000231 		else if (LoadCtl[2]) begin X_ = Xcalc[5:4]  ; Y_ = Ycalc[5:4]  ; A_ = Acalc[5:4]  ; end
 000231 		else if (LoadCtl[3]) begin X_ = Xcalc[7:6]  ; Y_ = Ycalc[7:6]  ; A_ = Acalc[7:6]  ; end
 000231 		else if (LoadCtl[4]) begin X_ = Xcalc[9:8]  ; Y_ = Ycalc[9:8]  ; A_ = Acalc[9:8]  ; end
 000232 		else if (LoadCtl[5]) begin X_ = Xcalc[11:10]; Y_ = Ycalc[11:10]; A_ = Acalc[11:10]; end
 000232 		else 				 begin X_ = 2'bxx		; Y_ = 2'bxx	   ; A_ = 2'bxx		  ; end			 
        	end
        	
        	assign Xout = X_;
        	assign Yout = Y_;
        	assign Aout = A_;
        	
        endmodule
        
