/* Verilog module written by DEF2Verilog (qflow) */
module output_terminal (
    output [11:0] Dout,
    input ISin,
    input Rdy,
    output Vld,
    input [1:0] Xin,
    input [1:0] Yin,
    input clk,
    input selSign,
    input selXY
);

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire [6:0] LoadCtl ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire ISin ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _256_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _48_ ;
wire _121_ ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire _118_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire _212_ ;
wire _250_ ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire ISreg_bF$buf0 ;
wire ISreg_bF$buf1 ;
wire ISreg_bF$buf2 ;
wire ISreg_bF$buf3 ;
wire ISreg_bF$buf4 ;
wire _80_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _147_ ;
wire _185_ ;
wire selXY ;
wire selSign ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire [11:0] Ycalc ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _96__bF$buf0 ;
wire _96__bF$buf1 ;
wire _96__bF$buf2 ;
wire _96__bF$buf3 ;
wire _96__bF$buf4 ;
wire _138_ ;
wire _30_ ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire ISreg ;
wire _264_ ;
wire [11:0] Dout ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire [11:4] Xin12b ;
wire [1:0] Yin ;
wire _255_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire [11:0] Xcalc ;
wire [1:0] Yin0 ;
wire [1:0] Yin1 ;
wire _214_ ;
wire _252_ ;
wire _117_ ;
wire _155_ ;
wire _193_ ;
wire _249_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire [1:0] Xin0 ;
wire [1:0] Xin1 ;
wire _114_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire _146_ ;
wire _184_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire [11:0] _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire LoadCtl_6_bF$buf0 ;
wire LoadCtl_6_bF$buf1 ;
wire LoadCtl_6_bF$buf2 ;
wire LoadCtl_6_bF$buf3 ;
wire LoadCtl_6_bF$buf4 ;
wire _119_ ;
wire _11_ ;
wire [11:4] Yin12b ;
wire _157_ ;
wire _195_ ;
wire _5_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _116_ ;
wire _154_ ;
wire gnd = 1'b0 ;
wire _192_ ;
wire _248_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire [1:0] Xin ;
wire _245_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire vdd = 1'b1 ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

FILL FILL_2__350_ (
);

FILL FILL_5__494_ (
);

FILL FILL_6__436_ (
);

FILL FILL_1__619_ (
);

DFFPOSX1 _588_ (
    .D(_39_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[4])
);

FILL FILL_1__372_ (
);

FILL FILL_2__406_ (
);

FILL FILL_3__521_ (
);

FILL FILL_7__452_ (
);

FILL FILL_0__394_ (
);

FILL FILL_1__428_ (
);

NOR2X1 _397_ (
    .A(Xin12b[6]),
    .B(Xin12b[7]),
    .Y(_145_)
);

FILL FILL_5__359_ (
);

FILL FILL75150x36150 (
);

FILL FILL_3__330_ (
);

FILL FILL_6__474_ (
);

FILL FILL_7__508_ (
);

FILL FILL_8__623_ (
);

FILL FILL_2__444_ (
);

FILL FILL_9__410_ (
);

FILL FILL_6__283_ (
);

FILL FILL_7__317_ (
);

FILL FILL_7__490_ (
);

FILL FILL_1__466_ (
);

FILL FILL_8__432_ (
);

FILL FILL_5__397_ (
);

FILL FILL_3__615_ (
);

FILL FILL_6__339_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_0_BUFX2_insert21 (
);

FILL FILL_4__402_ (
);

FILL FILL_0_BUFX2_insert22 (
);

FILL FILL_0_BUFX2_insert23 (
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_7__546_ (
);

FILL FILL_0__488_ (
);

FILL FILL_1__275_ (
);

FILL FILL_2__309_ (
);

FILL FILL_2__482_ (
);

FILL FILL_3__424_ (
);

FILL FILL_7__355_ (
);

FILL FILL_0__297_ (
);

FILL FILL_8__470_ (
);

FILL FILL_2__538_ (
);

FILL FILL_9__504_ (
);

FILL FILL_2__291_ (
);

FILL FILL_6__377_ (
);

NAND3X1 _512_ (
    .A(_244_),
    .B(_242_),
    .C(_219_),
    .Y(_245_)
);

FILL FILL_4__440_ (
);

FILL FILL_8__526_ (
);

FILL FILL_2__347_ (
);

FILL FILL_9__313_ (
);

FILL FILL_3__462_ (
);

NAND2X1 _321_ (
    .A(Yin[1]),
    .B(_80_),
    .Y(_83_)
);

FILL FILL_7__393_ (
);

FILL FILL_1__369_ (
);

FILL FILL_8__335_ (
);

FILL FILL_9__542_ (
);

FILL FILL_3__518_ (
);

FILL FILL_4__305_ (
);

FILL FILL_7__449_ (
);

OAI21X1 _550_ (
    .A(_237_),
    .B(_251_),
    .C(_268_),
    .Y(_46_)
);

FILL FILL_5__512_ (
);

FILL FILL_2__385_ (
);

FILL FILL_9__351_ (
);

FILL FILL_3__327_ (
);

DFFPOSX1 _606_ (
    .D(Rdy),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[0])
);

FILL FILL_4__534_ (
);

FILL FILL_5__321_ (
);

FILL FILL_8__373_ (
);

FILL FILL_9__407_ (
);

FILL FILL_0__412_ (
);

FILL FILL_3__556_ (
);

NAND3X1 _415_ (
    .A(ISreg_bF$buf1),
    .B(Xin12b[10]),
    .C(_160_),
    .Y(_161_)
);

FILL FILL_4__343_ (
);

FILL FILL_7__487_ (
);

FILL FILL_8__429_ (
);

FILL FILL_5__550_ (
);

FILL FILL_3__365_ (
);

FILL FILL_7__296_ (
);

FILL FILL_6__301_ (
);

FILL FILL_2__479_ (
);

FILL FILL_9__445_ (
);

FILL FILL74850x57750 (
);

FILL FILL_0__450_ (
);

NOR2X1 _453_ (
    .A(Yin1[0]),
    .B(Yin1[1]),
    .Y(_193_)
);

FILL FILL_4__381_ (
);

FILL FILL_5__415_ (
);

FILL FILL_8__467_ (
);

FILL FILL_6__530_ (
);

FILL FILL_2__288_ (
);

FILL FILL_0__506_ (
);

NAND2X1 _509_ (
    .A(ISreg_bF$buf3),
    .B(Yin12b[10]),
    .Y(_242_)
);

FILL FILL_4__437_ (
);

FILL FILL_2__500_ (
);

FILL FILL_8__276_ (
);

FILL FILL_0__315_ (
);

FILL FILL_3__459_ (
);

NAND2X1 _318_ (
    .A(Yin[0]),
    .B(_80_),
    .Y(_81_)
);

FILL FILL_1__522_ (
);

OR2X2 _491_ (
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

FILL FILL_5__453_ (
);

FILL FILL_0__544_ (
);

NAND2X1 _547_ (
    .A(Yin[0]),
    .B(_251_),
    .Y(_267_)
);

FILL FILL_1__331_ (
);

FILL FILL_4__475_ (
);

FILL FILL_5__509_ (
);

FILL FILL_6__624_ (
);

FILL FILL_7__411_ (
);

FILL FILL_0__353_ (
);

FILL FILL_3__497_ (
);

OAI21X1 _356_ (
    .A(_96__bF$buf2),
    .B(_108_),
    .C(_109_),
    .Y(_11_)
);

FILL FILL_4__284_ (
);

FILL FILL_5__318_ (
);

FILL FILL_5__491_ (
);

FILL FILL_6__433_ (
);

FILL FILL_0__409_ (
);

FILL FILL_1__616_ (
);

DFFPOSX1 _585_ (
    .D(_36_),
    .CLK(clk_bF$buf1),
    .Q(Xin12b[9])
);

FILL FILL_2__403_ (
);

FILL FILL_5__547_ (
);

FILL FILL_9__386_ (
);

FILL FILL_0__391_ (
);

FILL FILL_1__425_ (
);

NAND3X1 _394_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_139_),
    .C(_142_),
    .Y(_143_)
);

FILL FILL_5__356_ (
);

FILL FILL_6__471_ (
);

FILL FILL_7__505_ (
);

FILL FILL_0__447_ (
);

FILL FILL_8__620_ (
);

FILL FILL75150x57750 (
);

FILL FILL_4__378_ (
);

FILL FILL_2__441_ (
);

FILL FILL_6__527_ (
);

FILL FILL_6__280_ (
);

FILL FILL_7__314_ (
);

FILL FILL_1__463_ (
);

FILL FILL_5__394_ (
);

FILL FILL_6__336_ (
);

FILL FILL_7__543_ (
);

FILL FILL_0__485_ (
);

FILL FILL_1__519_ (
);

OAI21X1 _488_ (
    .A(_96__bF$buf0),
    .B(_222_),
    .C(_223_),
    .Y(_29_)
);

FILL FILL_2__306_ (
);

FILL FILL_3__421_ (
);

FILL FILL_9__289_ (
);

FILL FILL_7__352_ (
);

FILL FILL_0__294_ (
);

FILL FILL_1__328_ (
);

INVX1 _297_ (
    .A(Ycalc[8]),
    .Y(_65_)
);

FILL FILL_2__535_ (
);

FILL FILL_9__501_ (
);

FILL FILL75450x10950 (
);

FILL FILL_6__374_ (
);

FILL FILL_7__408_ (
);

FILL FILL_8__523_ (
);

FILL FILL_2__344_ (
);

FILL FILL_5__488_ (
);

FILL FILL_7_CLKBUF1_insert0 (
);

FILL FILL_7_CLKBUF1_insert1 (
);

FILL FILL_7_CLKBUF1_insert2 (
);

FILL FILL_7_CLKBUF1_insert3 (
);

FILL FILL_7_CLKBUF1_insert4 (
);

FILL FILL_7_CLKBUF1_insert5 (
);

FILL FILL_7_CLKBUF1_insert6 (
);

FILL FILL_7__390_ (
);

FILL FILL_1__366_ (
);

FILL FILL_8__332_ (
);

FILL FILL_5__297_ (
);

FILL FILL_3__515_ (
);

FILL FILL_4__302_ (
);

FILL FILL_7__446_ (
);

FILL FILL_0__388_ (
);

FILL FILL_2__382_ (
);

FILL FILL_3__324_ (
);

FILL FILL_6__468_ (
);

DFFPOSX1 _603_ (
    .D(_5_),
    .CLK(clk_bF$buf5),
    .Q(Yin1[1])
);

FILL FILL_4__531_ (
);

FILL FILL_8__617_ (
);

FILL FILL_8__370_ (
);

FILL FILL_2__438_ (
);

FILL FILL_3__553_ (
);

FILL FILL_6__277_ (
);

AND2X2 _412_ (
    .A(_129_),
    .B(_145_),
    .Y(_158_)
);

FILL FILL_4__340_ (
);

FILL FILL_7__484_ (
);

FILL FILL_8__426_ (
);

FILL FILL_3__362_ (
);

FILL FILL_7__293_ (
);

FILL FILL_2__476_ (
);

FILL FILL_3__418_ (
);

FILL FILL_4__625_ (
);

FILL FILL_7__349_ (
);

OR2X2 _450_ (
    .A(_189_),
    .B(Yin1[1]),
    .Y(_191_)
);

FILL FILL_5__412_ (
);

FILL FILL_1__498_ (
);

FILL FILL_8__464_ (
);

FILL FILL_5_BUFX2_insert10 (
);

FILL FILL_5_BUFX2_insert11 (
);

FILL FILL_5_BUFX2_insert12 (
);

FILL FILL_5_BUFX2_insert13 (
);

FILL FILL_5_BUFX2_insert14 (
);

FILL FILL_5_BUFX2_insert15 (
);

FILL FILL_5_BUFX2_insert16 (
);

FILL FILL_5_BUFX2_insert17 (
);

FILL FILL_5_BUFX2_insert18 (
);

FILL FILL_5_BUFX2_insert19 (
);

FILL FILL_2__285_ (
);

FILL FILL_0__503_ (
);

NAND2X1 _506_ (
    .A(Yin12b[11]),
    .B(_169_),
    .Y(_239_)
);

FILL FILL_4__434_ (
);

FILL FILL_8__273_ (
);

FILL FILL_0__312_ (
);

FILL FILL_9__480_ (
);

FILL FILL_3__456_ (
);

INVX1 _315_ (
    .A(Yin12b[4]),
    .Y(_78_)
);

FILL FILL_7__387_ (
);

FILL FILL_8__329_ (
);

FILL FILL_5__450_ (
);

FILL FILL_0__541_ (
);

OAI21X1 _544_ (
    .A(LoadCtl[0]),
    .B(_95_),
    .C(_265_),
    .Y(_43_)
);

FILL FILL_4__472_ (
);

FILL FILL_5__506_ (
);

FILL FILL_6__621_ (
);

FILL FILL_2__379_ (
);

FILL FILL_9__345_ (
);

FILL FILL_0__350_ (
);

FILL FILL_3__494_ (
);

FILL FILL_4__528_ (
);

OAI21X1 _353_ (
    .A(_93_),
    .B(_106_),
    .C(_103_),
    .Y(_107_)
);

FILL FILL_4__281_ (
);

FILL FILL_5__315_ (
);

FILL FILL_8__367_ (
);

FILL FILL_6__430_ (
);

FILL FILL_0__406_ (
);

AOI21X1 _409_ (
    .A(_154_),
    .B(_153_),
    .C(_96__bF$buf3),
    .Y(_156_)
);

FILL FILL_1__613_ (
);

FILL FILL_4__337_ (
);

DFFPOSX1 _582_ (
    .D(_33_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[10])
);

FILL FILL_2__400_ (
);

FILL FILL_5__544_ (
);

FILL FILL_9__383_ (
);

FILL FILL_3__359_ (
);

FILL FILL_1__422_ (
);

INVX1 _391_ (
    .A(Xin12b[7]),
    .Y(_140_)
);

FILL FILL_5__353_ (
);

FILL FILL_9__439_ (
);

FILL FILL_7__502_ (
);

FILL FILL_0__444_ (
);

OAI21X1 _447_ (
    .A(_53_),
    .B(LoadCtl_6_bF$buf4),
    .C(_188_),
    .Y(_23_)
);

FILL FILL_4__375_ (
);

FILL FILL_5__409_ (
);

FILL FILL_6__524_ (
);

FILL FILL_7__311_ (
);

FILL FILL_3__397_ (
);

FILL FILL_1__460_ (
);

FILL FILL_5__391_ (
);

FILL FILL_6__333_ (
);

FILL FILL_0__309_ (
);

FILL FILL_9__477_ (
);

FILL FILL_7__540_ (
);

FILL FILL_0__482_ (
);

FILL FILL_1__516_ (
);

NAND2X1 _485_ (
    .A(_216_),
    .B(_219_),
    .Y(_221_)
);

FILL FILL_2__303_ (
);

FILL FILL_5__447_ (
);

FILL FILL_8__499_ (
);

FILL FILL_0__538_ (
);

FILL FILL_9__286_ (
);

FILL FILL_0__291_ (
);

FILL FILL_1__325_ (
);

FILL FILL_4__469_ (
);

INVX1 _294_ (
    .A(Ycalc[7]),
    .Y(_63_)
);

FILL FILL_2__532_ (
);

FILL FILL_6__618_ (
);

FILL FILL_6__371_ (
);

FILL FILL_7__405_ (
);

FILL FILL_0__347_ (
);

FILL FILL_1__554_ (
);

FILL FILL_8__520_ (
);

FILL FILL_4__278_ (
);

FILL FILL_2__341_ (
);

FILL FILL_5__485_ (
);

FILL FILL_6__427_ (
);

DFFPOSX1 _579_ (
    .D(_30_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[9])
);

FILL FILL_1__363_ (
);

FILL FILL_5__294_ (
);

FILL FILL_3__512_ (
);

FILL FILL_7__443_ (
);

FILL FILL_0__385_ (
);

FILL FILL_1__419_ (
);

INVX1 _388_ (
    .A(Xcalc[7]),
    .Y(_137_)
);

FILL FILL_3__321_ (
);

FILL FILL_6__465_ (
);

DFFPOSX1 _600_ (
    .D(_2_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[4])
);

FILL FILL_8__614_ (
);

FILL FILL_2__435_ (
);

FILL FILL_9__401_ (
);

FILL FILL_3__550_ (
);

FILL FILL_6__274_ (
);

FILL FILL_7__308_ (
);

FILL FILL_7__481_ (
);

FILL FILL_1__457_ (
);

FILL FILL_8__423_ (
);

FILL FILL_5__388_ (
);

FILL FILL_7__537_ (
);

FILL FILL_0__479_ (
);

FILL FILL_7__290_ (
);

FILL FILL_2__473_ (
);

FILL FILL_3__415_ (
);

FILL FILL_4__622_ (
);

FILL FILL_7__346_ (
);

FILL FILL_0__288_ (
);

FILL FILL_1__495_ (
);

FILL FILL_8__461_ (
);

FILL FILL_2__529_ (
);

FILL FILL_2__282_ (
);

FILL FILL_0__500_ (
);

FILL FILL_6__368_ (
);

NAND2X1 _503_ (
    .A(Ycalc[11]),
    .B(_96__bF$buf1),
    .Y(_236_)
);

FILL FILL_4__431_ (
);

FILL FILL_8__517_ (
);

FILL FILL_2__338_ (
);

FILL FILL_9__304_ (
);

FILL FILL_3__453_ (
);

NAND3X1 _312_ (
    .A(_74_),
    .B(LoadCtl[3]),
    .C(_75_),
    .Y(_76_)
);

FILL FILL_7__384_ (
);

FILL FILL_8__326_ (
);

FILL FILL_9__533_ (
);

FILL FILL_3__509_ (
);

OAI21X1 _541_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[1]),
    .Y(_264_)
);

FILL FILL_5__503_ (
);

FILL FILL_8__555_ (
);

FILL FILL_2__376_ (
);

FILL FILL_9__342_ (
);

FILL FILL_3__318_ (
);

FILL FILL73050x10950 (
);

FILL FILL_3__491_ (
);

FILL FILL_4__525_ (
);

OAI21X1 _350_ (
    .A(Xin0[0]),
    .B(Xin0[1]),
    .C(ISreg_bF$buf1),
    .Y(_104_)
);

FILL FILL_5__312_ (
);

FILL FILL_1__398_ (
);

FILL FILL_8__364_ (
);

FILL FILL_0__403_ (
);

FILL FILL_3__547_ (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

INVX1 _406_ (
    .A(Xin12b[9]),
    .Y(_153_)
);

FILL FILL_4__334_ (
);

FILL FILL_7__478_ (
);

FILL FILL_5__541_ (
);

FILL FILL_9__380_ (
);

FILL FILL_3__356_ (
);

FILL FILL_7__287_ (
);

FILL FILL_5__350_ (
);

FILL FILL_9__436_ (
);

FILL FILL_0__441_ (
);

FILL FILL_4__619_ (
);

NOR2X1 _444_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .Y(_186_)
);

FILL FILL_4__372_ (
);

FILL FILL_5__406_ (
);

FILL FILL_8__458_ (
);

FILL FILL_6__521_ (
);

FILL FILL_2__279_ (
);

FILL FILL_3__394_ (
);

FILL FILL_4__428_ (
);

FILL FILL_6__330_ (
);

FILL FILL_0__306_ (
);

FILL FILL_9__474_ (
);

INVX1 _309_ (
    .A(Yin[1]),
    .Y(_73_)
);

FILL FILL_3_BUFX2_insert7 (
);

FILL FILL_3_BUFX2_insert8 (
);

FILL FILL_3_BUFX2_insert9 (
);

FILL FILL_1__513_ (
);

NAND2X1 _482_ (
    .A(_203_),
    .B(_217_),
    .Y(_218_)
);

FILL FILL_2__300_ (
);

FILL FILL_5__444_ (
);

FILL FILL_8__496_ (
);

FILL FILL_0__535_ (
);

FILL FILL_9__283_ (
);

OAI21X1 _538_ (
    .A(_123_),
    .B(_80_),
    .C(_262_),
    .Y(_40_)
);

FILL FILL_1__322_ (
);

FILL FILL_4__466_ (
);

INVX1 _291_ (
    .A(Ycalc[6]),
    .Y(_61_)
);

FILL FILL_6__615_ (
);

FILL FILL_9__339_ (
);

FILL FILL_7__402_ (
);

FILL FILL_0__344_ (
);

FILL FILL_3__488_ (
);

NAND2X1 _347_ (
    .A(Xcalc[1]),
    .B(_96__bF$buf4),
    .Y(_102_)
);

FILL FILL_1__551_ (
);

FILL FILL_4__275_ (
);

FILL FILL_5__309_ (
);

FILL FILL_5__482_ (
);

FILL FILL_6__424_ (
);

FILL FILL_3__297_ (
);

DFFPOSX1 _576_ (
    .D(_27_),
    .CLK(clk_bF$buf4),
    .Q(Ycalc[6])
);

FILL FILL_1__360_ (
);

FILL FILL_5__538_ (
);

FILL FILL_5__291_ (
);

FILL FILL_9__377_ (
);

FILL FILL_7__440_ (
);

FILL FILL_0__382_ (
);

FILL FILL_1__416_ (
);

NAND2X1 _385_ (
    .A(_131_),
    .B(_134_),
    .Y(_135_)
);

FILL FILL_2__623_ (
);

FILL FILL_5__347_ (
);

FILL FILL_8__399_ (
);

FILL FILL_6__462_ (
);

FILL FILL_0__438_ (
);

FILL FILL_4__369_ (
);

FILL FILL_2__432_ (
);

FILL FILL_6__518_ (
);

FILL FILL_7__305_ (
);

FILL FILL73650x28950 (
);

FILL FILL_1__454_ (
);

FILL FILL_8__420_ (
);

FILL FILL_5__385_ (
);

FILL FILL_6__327_ (
);

FILL FILL_5_CLKBUF1_insert0 (
);

FILL FILL_5_CLKBUF1_insert1 (
);

FILL FILL_5_CLKBUF1_insert2 (
);

FILL FILL_5_CLKBUF1_insert3 (
);

FILL FILL_5_CLKBUF1_insert4 (
);

FILL FILL_5_CLKBUF1_insert5 (
);

FILL FILL_5_CLKBUF1_insert6 (
);

FILL FILL_7__534_ (
);

FILL FILL_0__476_ (
);

OAI21X1 _479_ (
    .A(_63_),
    .B(LoadCtl_6_bF$buf2),
    .C(_215_),
    .Y(_28_)
);

FILL FILL_2__470_ (
);

FILL FILL_3__412_ (
);

FILL FILL_6__556_ (
);

FILL FILL_7__343_ (
);

FILL FILL_0__285_ (
);

FILL FILL_1__319_ (
);

INVX1 _288_ (
    .A(Ycalc[5]),
    .Y(_59_)
);

FILL FILL_1__492_ (
);

FILL FILL_2__526_ (
);

FILL FILL_6__365_ (
);

NAND2X1 _500_ (
    .A(_232_),
    .B(_233_),
    .Y(_234_)
);

FILL FILL_1__548_ (
);

FILL FILL_8__514_ (
);

FILL FILL_2__335_ (
);

FILL FILL_9__301_ (
);

FILL FILL_5__479_ (
);

FILL FILL_3__450_ (
);

FILL FILL_7__381_ (
);

FILL FILL_1__357_ (
);

FILL FILL_8__323_ (
);

FILL FILL_9__530_ (
);

FILL FILL_5__288_ (
);

FILL FILL_3__506_ (
);

FILL FILL_7__437_ (
);

FILL FILL_0__379_ (
);

FILL FILL_5__500_ (
);

FILL FILL_8__552_ (
);

FILL FILL_2__373_ (
);

FILL FILL_3__315_ (
);

FILL FILL_6__459_ (
);

FILL FILL_4__522_ (
);

FILL FILL_1__395_ (
);

FILL FILL_8__361_ (
);

FILL FILL_2__429_ (
);

FILL FILL75450x72150 (
);

FILL FILL_0__400_ (
);

FILL FILL_3__544_ (
);

FILL FILL75450x39750 (
);

NAND2X1 _403_ (
    .A(Xcalc[8]),
    .B(_96__bF$buf1),
    .Y(_151_)
);

FILL FILL_4__331_ (
);

FILL FILL_7__475_ (
);

FILL FILL_8__417_ (
);

FILL FILL_9__624_ (
);

FILL FILL_3__353_ (
);

FILL FILL_6__497_ (
);

FILL FILL_7__284_ (
);

FILL FILL_2__467_ (
);

FILL FILL_9__433_ (
);

FILL FILL_3__409_ (
);

FILL FILL_4__616_ (
);

INVX1 _441_ (
    .A(Yin1[0]),
    .Y(_183_)
);

FILL FILL_5__403_ (
);

FILL FILL_1__489_ (
);

FILL FILL_8__455_ (
);

FILL FILL_2__276_ (
);

FILL FILL_3__391_ (
);

FILL FILL_4__425_ (
);

FILL FILL_1__298_ (
);

FILL FILL_0__303_ (
);

FILL FILL_9__471_ (
);

FILL FILL_3__447_ (
);

INVX1 _306_ (
    .A(Ycalc[11]),
    .Y(_71_)
);

FILL FILL_1__510_ (
);

FILL FILL_7__378_ (
);

FILL FILL_5__441_ (
);

FILL FILL_8__493_ (
);

FILL FILL_9__527_ (
);

FILL FILL_0__532_ (
);

NAND2X1 _535_ (
    .A(Xin[0]),
    .B(_80_),
    .Y(_261_)
);

FILL FILL_4__463_ (
);

FILL FILL_8__549_ (
);

FILL FILL_9__336_ (
);

FILL FILL_0__341_ (
);

FILL FILL_3__485_ (
);

FILL FILL_4__519_ (
);

INVX1 _344_ (
    .A(Xin0[1]),
    .Y(_99_)
);

FILL FILL_5__306_ (
);

FILL FILL_8__358_ (
);

FILL FILL_6__421_ (
);

FILL FILL_3__294_ (
);

FILL FILL_4__328_ (
);

DFFPOSX1 _573_ (
    .D(_24_),
    .CLK(clk_bF$buf0),
    .Q(Ycalc[3])
);

FILL FILL_5__535_ (
);

FILL FILL_1__413_ (
);

INVX1 _382_ (
    .A(Xin12b[6]),
    .Y(_132_)
);

FILL FILL_2__620_ (
);

FILL FILL_5__344_ (
);

FILL FILL_8__396_ (
);

FILL FILL_0__435_ (
);

OAI21X1 _438_ (
    .A(_89_),
    .B(_93_),
    .C(_91_),
    .Y(_181_)
);

FILL FILL_4__366_ (
);

FILL FILL_6__515_ (
);

FILL FILL_7__302_ (
);

FILL FILL_3__388_ (
);

FILL FILL_1__451_ (
);

FILL FILL_5__382_ (
);

FILL FILL_6__324_ (
);

FILL FILL_7__531_ (
);

FILL FILL_0__473_ (
);

FILL FILL_1__507_ (
);

NAND2X1 _476_ (
    .A(ISreg_bF$buf4),
    .B(Yin12b[6]),
    .Y(_213_)
);

FILL FILL_5__438_ (
);

FILL FILL_6__553_ (
);

FILL FILL_0__529_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_2_BUFX2_insert21 (
);

FILL FILL_2_BUFX2_insert22 (
);

FILL FILL_2_BUFX2_insert23 (
);

FILL FILL_2_BUFX2_insert24 (
);

FILL FILL_2_BUFX2_insert25 (
);

FILL FILL_7__340_ (
);

FILL FILL_0__282_ (
);

FILL FILL_1__316_ (
);

INVX1 _285_ (
    .A(Ycalc[4]),
    .Y(_57_)
);

FILL FILL_2__523_ (
);

FILL FILL_8__299_ (
);

FILL FILL_6__362_ (
);

FILL FILL_0__338_ (
);

FILL FILL_1__545_ (
);

FILL FILL_8__511_ (
);

FILL FILL_2__332_ (
);

FILL FILL_5__476_ (
);

FILL FILL_6__418_ (
);

FILL FILL_7__625_ (
);

FILL FILL_1__354_ (
);

FILL FILL_8__320_ (
);

FILL FILL_4__498_ (
);

FILL FILL_5__285_ (
);

FILL FILL_3__503_ (
);

FILL FILL_7__434_ (
);

FILL FILL_0__376_ (
);

NOR2X1 _379_ (
    .A(Xin12b[4]),
    .B(Xin12b[5]),
    .Y(_129_)
);

FILL FILL_2__617_ (
);

FILL FILL_2__370_ (
);

FILL FILL_3__312_ (
);

FILL FILL_6__456_ (
);

FILL FILL_1__392_ (
);

FILL FILL_2__426_ (
);

FILL FILL_3__541_ (
);

OR2X2 _400_ (
    .A(_147_),
    .B(_144_),
    .Y(_148_)
);

FILL FILL_7__472_ (
);

FILL FILL_1__448_ (
);

FILL FILL_8__414_ (
);

FILL FILL_9__621_ (
);

FILL FILL_5__379_ (
);

FILL FILL_3__350_ (
);

FILL FILL_6__494_ (
);

FILL FILL_7__528_ (
);

FILL FILL_7__281_ (
);

FILL FILL_2__464_ (
);

FILL FILL_9__430_ (
);

FILL FILL_3__406_ (
);

FILL FILL73950x57750 (
);

FILL FILL_4__613_ (
);

FILL FILL_7__337_ (
);

FILL FILL_0__279_ (
);

FILL FILL_5__400_ (
);

FILL FILL_1__486_ (
);

FILL FILL_8__452_ (
);

FILL FILL_2__273_ (
);

FILL FILL_6__359_ (
);

FILL FILL_4__422_ (
);

FILL FILL_8__508_ (
);

FILL FILL_1__295_ (
);

FILL FILL_2__329_ (
);

FILL FILL_0__300_ (
);

FILL FILL_3__444_ (
);

INVX1 _303_ (
    .A(Ycalc[10]),
    .Y(_69_)
);

FILL FILL_7__375_ (
);

FILL FILL_8__317_ (
);

FILL FILL_8__490_ (
);

FILL FILL_6__397_ (
);

OAI21X1 _532_ (
    .A(_254_),
    .B(_76_),
    .C(_259_),
    .Y(_37_)
);

FILL FILL_4__460_ (
);

FILL FILL_8__546_ (
);

FILL FILL75450x25350 (
);

FILL FILL_2__367_ (
);

FILL FILL_3__309_ (
);

FILL FILL_3__482_ (
);

FILL FILL_4__516_ (
);

NAND2X1 _341_ (
    .A(Xcalc[0]),
    .B(_96__bF$buf4),
    .Y(_97_)
);

FILL FILL_5__303_ (
);

FILL FILL_1__389_ (
);

FILL FILL_8__355_ (
);

FILL FILL_3__538_ (
);

FILL FILL_3__291_ (
);

FILL FILL_4__325_ (
);

FILL FILL_7__469_ (
);

DFFPOSX1 _570_ (
    .D(_21_),
    .CLK(clk_bF$buf3),
    .Q(Ycalc[0])
);

FILL FILL_5__532_ (
);

FILL FILL_0__623_ (
);

FILL FILL_9__371_ (
);

FILL FILL_3__347_ (
);

FILL FILL_1__410_ (
);

FILL FILL_4__554_ (
);

FILL FILL_7__278_ (
);

FILL FILL_5__341_ (
);

FILL FILL_8__393_ (
);

FILL FILL_0__432_ (
);

NAND2X1 _435_ (
    .A(Yin0[0]),
    .B(LoadCtl_6_bF$buf0),
    .Y(_179_)
);

FILL FILL_4__363_ (
);

FILL FILL_8__449_ (
);

FILL FILL_6__512_ (
);

FILL FILL_3__385_ (
);

FILL FILL73050x72150 (
);

FILL FILL_4__419_ (
);

FILL FILL_6__321_ (
);

FILL FILL_2__499_ (
);

FILL FILL_9__465_ (
);

FILL FILL_0__470_ (
);

FILL FILL_1__504_ (
);

NAND3X1 _473_ (
    .A(_206_),
    .B(_203_),
    .C(_197_),
    .Y(_210_)
);

FILL FILL_5__435_ (
);

FILL FILL_8__487_ (
);

FILL FILL_6__550_ (
);

FILL FILL_0__526_ (
);

FILL FILL_9__274_ (
);

NAND2X1 _529_ (
    .A(Xin12b[9]),
    .B(_255_),
    .Y(_258_)
);

FILL FILL_1__313_ (
);

FILL FILL_4__457_ (
);

INVX1 _282_ (
    .A(Ycalc[3]),
    .Y(_55_)
);

FILL FILL_2__520_ (
);

FILL FILL_8__296_ (
);

FILL FILL_0__335_ (
);

FILL FILL_3__479_ (
);

OAI21X1 _338_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_93_),
    .C(_94_),
    .Y(_8_)
);

FILL FILL_1__542_ (
);

FILL FILL_5__473_ (
);

FILL FILL_6__415_ (
);

FILL FILL_7__622_ (
);

FILL FILL_3__288_ (
);

DFFPOSX1 _567_ (
    .D(_18_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[9])
);

FILL FILL_1__351_ (
);

FILL FILL_4__495_ (
);

FILL FILL_5__529_ (
);

FILL FILL_5__282_ (
);

FILL FILL_3__500_ (
);

FILL FILL_9__368_ (
);

FILL FILL_3_CLKBUF1_insert0 (
);

FILL FILL_3_CLKBUF1_insert1 (
);

FILL FILL_3_CLKBUF1_insert2 (
);

FILL FILL_3_CLKBUF1_insert3 (
);

FILL FILL_3_CLKBUF1_insert4 (
);

FILL FILL_3_CLKBUF1_insert5 (
);

FILL FILL_3_CLKBUF1_insert6 (
);

FILL FILL_7__431_ (
);

FILL FILL_0__373_ (
);

FILL FILL_1__407_ (
);

NAND2X1 _376_ (
    .A(_126_),
    .B(_125_),
    .Y(_127_)
);

FILL FILL_2__614_ (
);

FILL FILL_5__338_ (
);

FILL FILL_6__453_ (
);

FILL FILL_0__429_ (
);

FILL FILL_2__423_ (
);

FILL FILL_6__509_ (
);

FILL FILL_1__445_ (
);

FILL FILL_8__411_ (
);

FILL FILL_5__376_ (
);

FILL FILL_6__318_ (
);

FILL FILL_6__491_ (
);

FILL FILL_7__525_ (
);

FILL FILL_0__467_ (
);

FILL FILL_4__398_ (
);

FILL FILL_2__461_ (
);

FILL FILL_3__403_ (
);

FILL FILL_6__547_ (
);

FILL FILL_7__334_ (
);

FILL FILL_0__276_ (
);

INVX1 _279_ (
    .A(Ycalc[2]),
    .Y(_53_)
);

FILL FILL_1__483_ (
);

FILL FILL_2__517_ (
);

FILL FILL_6__356_ (
);

FILL FILL_1__539_ (
);

FILL FILL_8__505_ (
);

FILL FILL_7_BUFX2_insert10 (
);

FILL FILL_7_BUFX2_insert11 (
);

FILL FILL_7_BUFX2_insert12 (
);

FILL FILL_7_BUFX2_insert13 (
);

FILL FILL_7_BUFX2_insert14 (
);

FILL FILL_7_BUFX2_insert15 (
);

FILL FILL_7_BUFX2_insert16 (
);

FILL FILL_1__292_ (
);

FILL FILL_7_BUFX2_insert17 (
);

FILL FILL_7_BUFX2_insert18 (
);

FILL FILL_7_BUFX2_insert19 (
);

FILL FILL_2__326_ (
);

FILL FILL_3__441_ (
);

FILL FILL_7__619_ (
);

INVX1 _300_ (
    .A(Ycalc[9]),
    .Y(_67_)
);

FILL FILL_7__372_ (
);

FILL FILL_1__348_ (
);

FILL FILL_8__314_ (
);

FILL FILL_2__555_ (
);

FILL FILL_5__279_ (
);

FILL FILL_6__394_ (
);

FILL FILL_7__428_ (
);

FILL FILL_8__543_ (
);

FILL FILL_2__364_ (
);

FILL FILL_9__330_ (
);

FILL FILL_3__306_ (
);

FILL FILL_4__513_ (
);

FILL FILL75450x46950 (
);

FILL FILL_5__300_ (
);

FILL FILL_1__386_ (
);

FILL FILL_8__352_ (
);

FILL FILL_3__535_ (
);

FILL FILL74250x28950 (
);

FILL FILL_4__322_ (
);

FILL FILL_7__466_ (
);

FILL FILL_8__408_ (
);

FILL FILL_9__615_ (
);

FILL FILL_0__620_ (
);

FILL FILL_3__344_ (
);

FILL FILL_6__488_ (
);

BUFX2 _623_ (
    .A(_272_[8]),
    .Y(Dout[8])
);

FILL FILL_4__551_ (
);

FILL FILL_7__275_ (
);

FILL FILL_8__390_ (
);

FILL FILL_2__458_ (
);

FILL FILL_9__424_ (
);

FILL FILL_6__297_ (
);

NAND2X1 _432_ (
    .A(_171_),
    .B(_176_),
    .Y(_177_)
);

FILL FILL_4__360_ (
);

FILL FILL_8__446_ (
);

FILL FILL_3__382_ (
);

FILL FILL_4__416_ (
);

FILL FILL_5__623_ (
);

FILL FILL_1__289_ (
);

FILL FILL_2__496_ (
);

FILL FILL_9__462_ (
);

FILL FILL_3__438_ (
);

FILL FILL_1__501_ (
);

FILL FILL_7__369_ (
);

NAND2X1 _470_ (
    .A(_206_),
    .B(_207_),
    .Y(_208_)
);

FILL FILL_5__432_ (
);

FILL FILL_8__484_ (
);

FILL FILL_9__518_ (
);

FILL FILL_0__523_ (
);

NAND2X1 _526_ (
    .A(Xin12b[8]),
    .B(_255_),
    .Y(_256_)
);

FILL FILL_1__310_ (
);

FILL FILL_4__454_ (
);

FILL FILL_8__293_ (
);

FILL FILL_9__327_ (
);

FILL FILL_0__332_ (
);

FILL FILL_3__476_ (
);

OAI21X1 _335_ (
    .A(LoadCtl[0]),
    .B(_91_),
    .C(_92_),
    .Y(_7_)
);

FILL FILL_8__349_ (
);

FILL FILL_5__470_ (
);

FILL FILL_6__412_ (
);

FILL FILL_9__556_ (
);

FILL FILL_3__285_ (
);

FILL FILL_4__319_ (
);

DFFPOSX1 _564_ (
    .D(_15_),
    .CLK(clk_bF$buf5),
    .Q(Xcalc[6])
);

FILL FILL75750x54150 (
);

FILL FILL_4__492_ (
);

FILL FILL_5__526_ (
);

FILL FILL_2__399_ (
);

FILL FILL_0__617_ (
);

FILL FILL_9__365_ (
);

FILL FILL74550x36150 (
);

FILL FILL_0__370_ (
);

FILL FILL_1__404_ (
);

FILL FILL_4__548_ (
);

OAI21X1 _373_ (
    .A(Xin12b[4]),
    .B(_116_),
    .C(ISreg_bF$buf1),
    .Y(_124_)
);

FILL FILL_5__335_ (
);

FILL FILL_8__387_ (
);

FILL FILL_6__450_ (
);

FILL FILL_0__426_ (
);

NAND3X1 _429_ (
    .A(_172_),
    .B(_173_),
    .C(_163_),
    .Y(_174_)
);

FILL FILL_4__357_ (
);

FILL FILL_2__420_ (
);

FILL FILL_6__506_ (
);

FILL FILL_3__379_ (
);

FILL FILL_1__442_ (
);

FILL FILL_5__373_ (
);

FILL FILL_6__315_ (
);

FILL FILL_9__459_ (
);

FILL FILL_7__522_ (
);

FILL FILL_0__464_ (
);

NAND3X1 _467_ (
    .A(ISreg_bF$buf4),
    .B(Yin12b[6]),
    .C(_204_),
    .Y(_205_)
);

FILL FILL_4__395_ (
);

FILL FILL_5__429_ (
);

FILL FILL_3__400_ (
);

FILL FILL_6__544_ (
);

FILL FILL_7__331_ (
);

FILL FILL_0__273_ (
);

FILL FILL_1__307_ (
);

INVX1 _276_ (
    .A(Ycalc[1]),
    .Y(_51_)
);

FILL FILL_1__480_ (
);

FILL FILL_2__514_ (
);

FILL FILL_6__353_ (
);

FILL FILL_0__329_ (
);

FILL FILL_9__497_ (
);

FILL FILL_1__536_ (
);

FILL FILL_8__502_ (
);

FILL FILL_2__323_ (
);

FILL FILL_5__467_ (
);

FILL FILL_6__409_ (
);

FILL FILL_7__616_ (
);

FILL FILL_1__345_ (
);

FILL FILL_8__311_ (
);

FILL FILL_4__489_ (
);

FILL FILL_2__552_ (
);

FILL FILL_5__276_ (
);

FILL FILL_6__391_ (
);

FILL FILL_7__425_ (
);

FILL FILL_0__367_ (
);

FILL FILL_8__540_ (
);

FILL FILL_4__298_ (
);

FILL FILL_2__361_ (
);

FILL FILL_3__303_ (
);

FILL FILL_6__447_ (
);

FILL FILL_4__510_ (
);

DFFPOSX1 _599_ (
    .D(_1_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[7])
);

FILL FILL_1__383_ (
);

FILL FILL_2__417_ (
);

FILL FILL_3__532_ (
);

FILL FILL_7__463_ (
);

FILL FILL_1__439_ (
);

FILL FILL_8__405_ (
);

FILL FILL_3__341_ (
);

FILL FILL_6__485_ (
);

FILL FILL_7__519_ (
);

BUFX2 _620_ (
    .A(_272_[5]),
    .Y(Dout[5])
);

FILL FILL_2__455_ (
);

FILL FILL_9__421_ (
);

FILL FILL_6__294_ (
);

FILL FILL_7__328_ (
);

FILL FILL_1__477_ (
);

FILL FILL_8__443_ (
);

FILL FILL_4__413_ (
);

FILL FILL_0__499_ (
);

FILL FILL_5__620_ (
);

FILL FILL_1__286_ (
);

FILL FILL_2__493_ (
);

FILL FILL_3__435_ (
);

FILL FILL_7__366_ (
);

FILL FILL_8__308_ (
);

FILL FILL_8__481_ (
);

FILL FILL_2__549_ (
);

FILL FILL_9__515_ (
);

FILL FILL_0__520_ (
);

FILL FILL_6__388_ (
);

OAI21X1 _523_ (
    .A(_167_),
    .B(_251_),
    .C(_253_),
    .Y(_34_)
);

FILL FILL_4__451_ (
);

FILL FILL_8__537_ (
);

FILL FILL_8__290_ (
);

FILL FILL_2__358_ (
);

FILL FILL_9__324_ (
);

FILL FILL_3__473_ (
);

FILL FILL_4__507_ (
);

OAI21X1 _332_ (
    .A(LoadCtl[0]),
    .B(_89_),
    .C(_90_),
    .Y(_6_)
);

FILL FILL_8__346_ (
);

FILL FILL_9__553_ (
);

FILL FILL_3__529_ (
);

FILL FILL_3__282_ (
);

FILL FILL_4__316_ (
);

DFFPOSX1 _561_ (
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[3])
);

FILL FILL_5__523_ (
);

FILL FILL_2__396_ (
);

FILL FILL_0__614_ (
);

FILL FILL_9__362_ (
);

FILL FILL_3__338_ (
);

BUFX2 _617_ (
    .A(_272_[2]),
    .Y(Dout[2])
);

FILL FILL_1__401_ (
);

FILL FILL_4__545_ (
);

NAND2X1 _370_ (
    .A(Xcalc[4]),
    .B(_96__bF$buf4),
    .Y(_122_)
);

FILL FILL_5__332_ (
);

FILL FILL_8__384_ (
);

FILL FILL_9__418_ (
);

FILL FILL74550x57750 (
);

FILL FILL_0__423_ (
);

NAND2X1 _426_ (
    .A(_168_),
    .B(_170_),
    .Y(_171_)
);

FILL FILL_4__354_ (
);

FILL FILL_7__498_ (
);

FILL FILL_6__503_ (
);

FILL FILL_3__376_ (
);

FILL FILL_5__617_ (
);

FILL FILL_5__370_ (
);

FILL FILL_6__312_ (
);

FILL FILL_9__456_ (
);

FILL FILL_0__461_ (
);

AOI22X1 _464_ (
    .A(_59_),
    .B(_96__bF$buf1),
    .C(_201_),
    .D(_202_),
    .Y(_26_)
);

FILL FILL_4__392_ (
);

FILL FILL_5__426_ (
);

FILL FILL_8__478_ (
);

FILL FILL_1_CLKBUF1_insert0 (
);

FILL FILL_1_CLKBUF1_insert1 (
);

FILL FILL_1_CLKBUF1_insert2 (
);

FILL FILL_1_CLKBUF1_insert3 (
);

FILL FILL_1_CLKBUF1_insert4 (
);

FILL FILL_1_CLKBUF1_insert5 (
);

FILL FILL_1_CLKBUF1_insert6 (
);

FILL FILL_6__541_ (
);

FILL FILL_2__299_ (
);

FILL FILL_0__517_ (
);

FILL FILL74850x10950 (
);

FILL FILL_1__304_ (
);

FILL FILL_4__448_ (
);

INVX1 _273_ (
    .A(Ycalc[0]),
    .Y(_49_)
);

FILL FILL_2__511_ (
);

FILL FILL_8__287_ (
);

FILL FILL_6__350_ (
);

FILL FILL_0__326_ (
);

OAI21X1 _329_ (
    .A(_73_),
    .B(_86_),
    .C(_88_),
    .Y(_5_)
);

FILL FILL_1__533_ (
);

FILL FILL_2__320_ (
);

FILL FILL_5__464_ (
);

FILL FILL_6__406_ (
);

FILL FILL_7__613_ (
);

FILL FILL_0__555_ (
);

FILL FILL_3__279_ (
);

DFFPOSX1 _558_ (
    .D(_9_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[0])
);

FILL FILL_1__342_ (
);

FILL FILL_4__486_ (
);

FILL FILL_5__273_ (
);

FILL FILL_7__422_ (
);

FILL FILL_0__364_ (
);

AND2X2 _367_ (
    .A(_106_),
    .B(_115_),
    .Y(_119_)
);

FILL FILL_4__295_ (
);

FILL FILL_5__329_ (
);

FILL FILL_3__300_ (
);

FILL FILL_6__444_ (
);

DFFPOSX1 _596_ (
    .D(_47_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[8])
);

FILL FILL_1__380_ (
);

FILL FILL_2__414_ (
);

FILL FILL_7__460_ (
);

FILL FILL_1__436_ (
);

FILL FILL_8__402_ (
);

FILL FILL_5__367_ (
);

FILL FILL_6__309_ (
);

FILL FILL_6__482_ (
);

FILL FILL_7__516_ (
);

FILL FILL_0__458_ (
);

BUFX2 BUFX2_insert7 (
    .A(selXY),
    .Y(selXY_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(selXY),
    .Y(selXY_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(selXY),
    .Y(selXY_bF$buf1)
);

FILL FILL_4__389_ (
);

FILL FILL_2__452_ (
);

FILL FILL_6__538_ (
);

FILL FILL_6__291_ (
);

FILL FILL_7__325_ (
);

FILL FILL_1__474_ (
);

FILL FILL_8__440_ (
);

FILL FILL_2__508_ (
);

FILL FILL75150x10950 (
);

FILL FILL_3__623_ (
);

FILL FILL_6__347_ (
);

FILL FILL_4__410_ (
);

FILL FILL_7__554_ (
);

FILL FILL_0__496_ (
);

NAND2X1 _499_ (
    .A(ISreg_bF$buf3),
    .B(_230_),
    .Y(_233_)
);

FILL FILL_1__283_ (
);

FILL FILL_2__317_ (
);

FILL FILL_2__490_ (
);

FILL FILL_3__432_ (
);

FILL FILL_7__363_ (
);

FILL FILL_1__339_ (
);

FILL FILL_8__305_ (
);

FILL FILL_2__546_ (
);

FILL FILL_9__512_ (
);

FILL FILL_6__385_ (
);

FILL FILL_7__419_ (
);

NAND2X1 _520_ (
    .A(Xin[0]),
    .B(_251_),
    .Y(_252_)
);

FILL FILL_8__534_ (
);

FILL FILL_2__355_ (
);

FILL FILL_9__321_ (
);

FILL FILL_5__499_ (
);

FILL FILL_3__470_ (
);

FILL FILL_4__504_ (
);

FILL FILL_1__377_ (
);

FILL FILL_8__343_ (
);

FILL FILL_9__550_ (
);

FILL FILL_3__526_ (
);

FILL FILL_4__313_ (
);

FILL FILL_7__457_ (
);

FILL FILL_0__399_ (
);

FILL FILL_5__520_ (
);

FILL FILL_2__393_ (
);

FILL FILL_3__335_ (
);

FILL FILL_6__479_ (
);

BUFX2 _614_ (
    .A(_272_[1]),
    .Y(Dout[1])
);

FILL FILL_4__542_ (
);

FILL FILL_8__381_ (
);

FILL FILL_2__449_ (
);

FILL FILL_9__415_ (
);

FILL FILL_0__420_ (
);

FILL FILL_6__288_ (
);

NAND2X1 _423_ (
    .A(selSign),
    .B(_167_),
    .Y(_168_)
);

FILL FILL_4__351_ (
);

FILL FILL_7__495_ (
);

FILL FILL_8__437_ (
);

FILL FILL_6__500_ (
);

FILL FILL_3__373_ (
);

FILL FILL_4__407_ (
);

FILL FILL_5__614_ (
);

FILL FILL_2__487_ (
);

FILL FILL_3__429_ (
);

OAI21X1 _461_ (
    .A(_93_),
    .B(_78_),
    .C(_195_),
    .Y(_200_)
);

FILL FILL_5__423_ (
);

FILL FILL_8__475_ (
);

FILL FILL_2__296_ (
);

FILL FILL_0__514_ (
);

AND2X2 _517_ (
    .A(_75_),
    .B(_248_),
    .Y(_249_)
);

FILL FILL_1__301_ (
);

FILL FILL_4__445_ (
);

FILL FILL_8__284_ (
);

FILL FILL_0__323_ (
);

FILL FILL_3__467_ (
);

FILL FILL_4_BUFX2_insert20 (
);

FILL FILL_4_BUFX2_insert21 (
);

OAI21X1 _326_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[0]),
    .Y(_87_)
);

FILL FILL_4_BUFX2_insert22 (
);

FILL FILL_4_BUFX2_insert23 (
);

FILL FILL_4_BUFX2_insert24 (
);

FILL FILL_4_BUFX2_insert25 (
);

FILL FILL_1__530_ (
);

FILL FILL_7__398_ (
);

FILL FILL_5__461_ (
);

FILL FILL75750x61350 (
);

FILL FILL_6__403_ (
);

FILL FILL75750x28950 (
);

FILL FILL_0__552_ (
);

FILL FILL_3__276_ (
);

NAND2X1 _555_ (
    .A(Yin12b[6]),
    .B(_76_),
    .Y(_271_)
);

FILL FILL_4__483_ (
);

FILL FILL_5__517_ (
);

FILL FILL_9__356_ (
);

FILL FILL_0__361_ (
);

FILL FILL_4__539_ (
);

NAND2X1 _364_ (
    .A(_106_),
    .B(_115_),
    .Y(_116_)
);

FILL FILL_4__292_ (
);

FILL FILL_5__326_ (
);

FILL FILL_8__378_ (
);

FILL FILL_6__441_ (
);

FILL FILL_0__417_ (
);

FILL FILL_1__624_ (
);

FILL FILL_4__348_ (
);

DFFPOSX1 _593_ (
    .D(_44_),
    .CLK(clk_bF$buf2),
    .Q(Xin0[1])
);

FILL FILL_2__411_ (
);

FILL FILL_5__555_ (
);

FILL FILL_9__394_ (
);

FILL FILL_1__433_ (
);

FILL FILL_5__364_ (
);

FILL FILL_6__306_ (
);

FILL FILL_7__513_ (
);

FILL FILL_0__455_ (
);

OAI21X1 _458_ (
    .A(_93_),
    .B(_197_),
    .C(_78_),
    .Y(_198_)
);

FILL FILL_4__386_ (
);

FILL FILL_6__535_ (
);

FILL FILL_7__322_ (
);

FILL FILL_1__471_ (
);

FILL FILL_2__505_ (
);

FILL FILL_3__620_ (
);

FILL FILL_6__344_ (
);

FILL FILL_9__488_ (
);

FILL FILL_7__551_ (
);

FILL FILL_0__493_ (
);

FILL FILL_1__527_ (
);

NAND3X1 _496_ (
    .A(_229_),
    .B(_197_),
    .C(_228_),
    .Y(_230_)
);

FILL FILL_1__280_ (
);

FILL FILL_2__314_ (
);

FILL FILL_5__458_ (
);

FILL FILL_0__549_ (
);

FILL FILL_9__297_ (
);

FILL FILL_7__360_ (
);

FILL FILL_1__336_ (
);

FILL FILL_8__302_ (
);

FILL FILL_2__543_ (
);

FILL FILL_6__382_ (
);

FILL FILL_7__416_ (
);

FILL FILL_0__358_ (
);

FILL FILL75450x7350 (
);

FILL FILL_8__531_ (
);

FILL FILL_4__289_ (
);

FILL FILL_2__352_ (
);

FILL FILL_5__496_ (
);

FILL FILL_6__438_ (
);

FILL FILL_4__501_ (
);

FILL FILL_1__374_ (
);

FILL FILL_8__340_ (
);

FILL FILL_2__408_ (
);

FILL FILL_3__523_ (
);

FILL FILL_4__310_ (
);

FILL FILL_7__454_ (
);

FILL FILL_0__396_ (
);

OAI21X1 _399_ (
    .A(_116_),
    .B(_146_),
    .C(ISreg_bF$buf2),
    .Y(_147_)
);

FILL FILL_2__390_ (
);

FILL FILL_3__332_ (
);

FILL FILL_6__476_ (
);

DFFPOSX1 _611_ (
    .D(LoadCtl[4]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[5])
);

FILL FILL_8__625_ (
);

FILL FILL_2__446_ (
);

FILL FILL_6__285_ (
);

FILL FILL_7__319_ (
);

OAI21X1 _420_ (
    .A(_157_),
    .B(LoadCtl_6_bF$buf4),
    .C(_165_),
    .Y(_19_)
);

FILL FILL_7__492_ (
);

FILL FILL_1__468_ (
);

FILL FILL_8__434_ (
);

FILL FILL_5__399_ (
);

FILL FILL_3__617_ (
);

FILL FILL_3__370_ (
);

FILL FILL_4__404_ (
);

FILL FILL_7__548_ (
);

FILL FILL_1__277_ (
);

FILL FILL_2__484_ (
);

FILL FILL_9__450_ (
);

FILL FILL_3__426_ (
);

FILL FILL_7__357_ (
);

FILL FILL_0__299_ (
);

FILL FILL_5__420_ (
);

FILL FILL_8__472_ (
);

FILL FILL_2__293_ (
);

FILL FILL_0__511_ (
);

FILL FILL_6__379_ (
);

NAND3X1 _514_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_246_),
    .C(_243_),
    .Y(_247_)
);

FILL FILL_4__442_ (
);

FILL FILL_8__528_ (
);

FILL FILL_8__281_ (
);

FILL FILL_2__349_ (
);

FILL FILL_9__315_ (
);

FILL FILL_0__320_ (
);

FILL FILL_3__464_ (
);

INVX1 _323_ (
    .A(Yin[0]),
    .Y(_84_)
);

FILL FILL_7__395_ (
);

FILL FILL_8__337_ (
);

FILL FILL_6__400_ (
);

FILL FILL_9__544_ (
);

FILL FILL_3__273_ (
);

FILL FILL_4__307_ (
);

OAI21X1 _552_ (
    .A(_84_),
    .B(_255_),
    .C(_269_),
    .Y(_47_)
);

FILL FILL_4__480_ (
);

FILL FILL_5__514_ (
);

FILL FILL_2__387_ (
);

FILL FILL_9__353_ (
);

FILL FILL_3__329_ (
);

DFFPOSX1 _608_ (
    .D(LoadCtl[1]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[2])
);

FILL FILL_4__536_ (
);

NAND2X1 _361_ (
    .A(Xcalc[3]),
    .B(_96__bF$buf1),
    .Y(_114_)
);

FILL FILL_5__323_ (
);

FILL FILL_8__375_ (
);

FILL FILL_9__409_ (
);

FILL FILL_0__414_ (
);

NAND2X1 _417_ (
    .A(ISreg_bF$buf2),
    .B(_160_),
    .Y(_163_)
);

FILL FILL_1__621_ (
);

FILL FILL_4__345_ (
);

FILL FILL_7__489_ (
);

DFFPOSX1 _590_ (
    .D(_41_),
    .CLK(clk_bF$buf5),
    .Q(Xin1[0])
);

FILL FILL_5__552_ (
);

FILL FILL_9__391_ (
);

FILL FILL_3__367_ (
);

FILL FILL_1__430_ (
);

FILL FILL_7__298_ (
);

FILL FILL_5__361_ (
);

FILL FILL_6__303_ (
);

FILL FILL_9__447_ (
);

FILL FILL_7__510_ (
);

FILL FILL_0__452_ (
);

NAND2X1 _455_ (
    .A(ISreg_bF$buf3),
    .B(_194_),
    .Y(_195_)
);

FILL FILL_4__383_ (
);

FILL FILL_5__417_ (
);

FILL FILL_8__469_ (
);

FILL FILL_6__532_ (
);

FILL FILL_0__508_ (
);

FILL FILL_4__439_ (
);

FILL FILL_2__502_ (
);

FILL FILL_8__278_ (
);

FILL FILL75750x14550 (
);

FILL FILL_6__341_ (
);

FILL FILL_0__317_ (
);

FILL FILL_9__485_ (
);

FILL FILL_0__490_ (
);

FILL FILL_1__524_ (
);

AOI22X1 _493_ (
    .A(_67_),
    .B(_96__bF$buf0),
    .C(_226_),
    .D(_227_),
    .Y(_30_)
);

FILL FILL_2__311_ (
);

FILL FILL_5__455_ (
);

FILL FILL_0__546_ (
);

FILL FILL_9__294_ (
);

NAND2X1 _549_ (
    .A(Yin[1]),
    .B(_251_),
    .Y(_268_)
);

FILL FILL_1__333_ (
);

FILL FILL_4__477_ (
);

FILL FILL_9_BUFX2_insert11 (
);

FILL FILL_9_BUFX2_insert12 (
);

FILL FILL_9_BUFX2_insert13 (
);

FILL FILL_9_BUFX2_insert15 (
);

FILL FILL_9_BUFX2_insert16 (
);

FILL FILL_9_BUFX2_insert17 (
);

FILL FILL_9_BUFX2_insert19 (
);

FILL FILL_2__540_ (
);

FILL FILL_7__413_ (
);

FILL FILL_0__355_ (
);

FILL FILL_3__499_ (
);

NAND2X1 _358_ (
    .A(Xin1[1]),
    .B(_110_),
    .Y(_111_)
);

FILL FILL_4__286_ (
);

FILL FILL_5__493_ (
);

FILL FILL_6__435_ (
);

FILL FILL74850x72150 (
);

FILL FILL_1__618_ (
);

DFFPOSX1 _587_ (
    .D(_38_),
    .CLK(clk_bF$buf1),
    .Q(Xin12b[7])
);

FILL FILL74850x39750 (
);

FILL FILL_1__371_ (
);

FILL FILL_2__405_ (
);

FILL FILL_5__549_ (
);

FILL FILL_3__520_ (
);

FILL FILL_9__388_ (
);

FILL FILL_7__451_ (
);

FILL FILL_0__393_ (
);

FILL FILL73350x28950 (
);

FILL FILL_1__427_ (
);

INVX1 _396_ (
    .A(Xin12b[8]),
    .Y(_144_)
);

FILL FILL_5__358_ (
);

FILL FILL_6__473_ (
);

FILL FILL_7__507_ (
);

FILL FILL_0__449_ (
);

FILL FILL_8__622_ (
);

FILL FILL_2__443_ (
);

FILL FILL_6__529_ (
);

FILL FILL_6__282_ (
);

FILL FILL_7__316_ (
);

FILL FILL_1__465_ (
);

FILL FILL_8__431_ (
);

FILL FILL_5__396_ (
);

FILL FILL_3__614_ (
);

FILL FILL_6__338_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_4__401_ (
);

FILL FILL_0_BUFX2_insert12 (
);

FILL FILL_0_BUFX2_insert13 (
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

FILL FILL_0_BUFX2_insert16 (
);

FILL FILL_0_BUFX2_insert17 (
);

FILL FILL_0_BUFX2_insert18 (
);

FILL FILL_7__545_ (
);

FILL FILL_0__487_ (
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL_1__274_ (
);

FILL FILL_2__308_ (
);

FILL FILL_2__481_ (
);

FILL FILL_3__423_ (
);

FILL FILL_7__354_ (
);

FILL FILL_0__296_ (
);

OAI21X1 _299_ (
    .A(selXY_bF$buf1),
    .B(_65_),
    .C(_66_),
    .Y(_272_[8])
);

FILL FILL_2__537_ (
);

FILL FILL_9__503_ (
);

FILL FILL_2__290_ (
);

FILL FILL_6__376_ (
);

OAI21X1 _511_ (
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .C(ISreg_bF$buf4),
    .Y(_244_)
);

FILL FILL_8__525_ (
);

FILL FILL_2__346_ (
);

FILL FILL_9__312_ (
);

FILL FILL_8_CLKBUF1_insert0 (
);

FILL FILL_8_CLKBUF1_insert1 (
);

FILL FILL_8_CLKBUF1_insert2 (
);

FILL FILL_8_CLKBUF1_insert3 (
);

FILL FILL_8_CLKBUF1_insert4 (
);

FILL FILL_8_CLKBUF1_insert5 (
);

FILL FILL_8_CLKBUF1_insert6 (
);

FILL FILL_3__461_ (
);

INVX1 _320_ (
    .A(Yin12b[5]),
    .Y(_82_)
);

BUFX2 BUFX2_insert20 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .A(_96_),
    .Y(_96__bF$buf4)
);

BUFX2 BUFX2_insert22 (
    .A(_96_),
    .Y(_96__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .A(_96_),
    .Y(_96__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .A(_96_),
    .Y(_96__bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .A(_96_),
    .Y(_96__bF$buf0)
);

FILL FILL_7__392_ (
);

FILL FILL_1__368_ (
);

FILL FILL_8__334_ (
);

FILL FILL75150x72150 (
);

FILL FILL_9__541_ (
);

FILL FILL_5__299_ (
);

FILL FILL_3__517_ (
);

FILL FILL75150x39750 (
);

FILL FILL_4__304_ (
);

FILL FILL_7__448_ (
);

FILL FILL_5__511_ (
);

FILL FILL_2__384_ (
);

FILL FILL_9__350_ (
);

FILL FILL_3__326_ (
);

DFFPOSX1 _605_ (
    .D(_7_),
    .CLK(clk_bF$buf3),
    .Q(Yin0[1])
);

FILL FILL_4__533_ (
);

FILL FILL_8__619_ (
);

FILL FILL_5__320_ (
);

FILL FILL_8__372_ (
);

FILL FILL_9__406_ (
);

FILL FILL_0__411_ (
);

FILL FILL_3__555_ (
);

FILL FILL_6__279_ (
);

NAND3X1 _414_ (
    .A(_159_),
    .B(_119_),
    .C(_158_),
    .Y(_160_)
);

FILL FILL_4__342_ (
);

FILL FILL_7__486_ (
);

FILL FILL_8__428_ (
);

FILL FILL_3__364_ (
);

FILL FILL_7__295_ (
);

FILL FILL_6__300_ (
);

FILL FILL_2__478_ (
);

FILL FILL_9__444_ (
);

OAI21X1 _452_ (
    .A(_55_),
    .B(LoadCtl_6_bF$buf4),
    .C(_192_),
    .Y(_24_)
);

FILL FILL_4__380_ (
);

FILL FILL_5__414_ (
);

FILL FILL_8__466_ (
);

FILL FILL_2__287_ (
);

FILL FILL_0__505_ (
);

INVX1 _508_ (
    .A(_240_),
    .Y(_241_)
);

FILL FILL_4__436_ (
);

FILL FILL_8__275_ (
);

FILL FILL_9__309_ (
);

FILL FILL_0__314_ (
);

FILL FILL_9__482_ (
);

FILL FILL_3__458_ (
);

NOR2X1 _317_ (
    .A(_74_),
    .B(_79_),
    .Y(_80_)
);

FILL FILL_1__521_ (
);

FILL FILL_7__389_ (
);

OAI21X1 _490_ (
    .A(_93_),
    .B(_216_),
    .C(_219_),
    .Y(_225_)
);

FILL FILL_5__452_ (
);

FILL FILL_9__538_ (
);

FILL FILL_0__543_ (
);

FILL FILL_9__291_ (
);

OAI21X1 _546_ (
    .A(LoadCtl[0]),
    .B(_99_),
    .C(_266_),
    .Y(_44_)
);

FILL FILL_1__330_ (
);

FILL FILL_4__474_ (
);

FILL FILL_5__508_ (
);

FILL FILL_6__623_ (
);

FILL FILL_9__347_ (
);

FILL FILL_7__410_ (
);

FILL FILL_0__352_ (
);

FILL FILL_3__496_ (
);

NAND2X1 _355_ (
    .A(Xcalc[2]),
    .B(_96__bF$buf2),
    .Y(_109_)
);

FILL FILL_4__283_ (
);

FILL FILL_5__317_ (
);

FILL FILL_8__369_ (
);

FILL FILL_5__490_ (
);

FILL FILL_6__432_ (
);

FILL FILL_0__408_ (
);

FILL FILL_1__615_ (
);

FILL FILL_4__339_ (
);

DFFPOSX1 _584_ (
    .D(_35_),
    .CLK(clk_bF$buf5),
    .Q(Xin12b[8])
);

FILL FILL_2__402_ (
);

FILL FILL_5__546_ (
);

FILL FILL_0__390_ (
);

FILL FILL_1__424_ (
);

NAND3X1 _393_ (
    .A(_140_),
    .B(_141_),
    .C(_133_),
    .Y(_142_)
);

FILL FILL_5__355_ (
);

FILL FILL_6__470_ (
);

FILL FILL_7__504_ (
);

FILL FILL_0__446_ (
);

NAND2X1 _449_ (
    .A(Yin1[1]),
    .B(_189_),
    .Y(_190_)
);

FILL FILL_4__377_ (
);

FILL FILL_2__440_ (
);

FILL FILL_6__526_ (
);

FILL FILL_7__313_ (
);

FILL FILL_3__399_ (
);

FILL FILL_1__462_ (
);

FILL FILL_5__393_ (
);

FILL FILL_6__335_ (
);

FILL FILL_7__542_ (
);

FILL FILL_0__484_ (
);

FILL FILL_1__518_ (
);

NAND2X1 _487_ (
    .A(Ycalc[8]),
    .B(_96__bF$buf0),
    .Y(_223_)
);

FILL FILL_2__305_ (
);

FILL FILL_5__449_ (
);

FILL FILL_3__420_ (
);

FILL FILL_7__351_ (
);

FILL FILL_0__293_ (
);

FILL FILL_1__327_ (
);

OAI21X1 _296_ (
    .A(selXY_bF$buf1),
    .B(_63_),
    .C(_64_),
    .Y(_272_[7])
);

FILL FILL_2__534_ (
);

FILL FILL_9__500_ (
);

FILL FILL_6__373_ (
);

FILL FILL74850x25350 (
);

FILL FILL_7__407_ (
);

FILL FILL_0__349_ (
);

FILL FILL_1__556_ (
);

FILL FILL_8__522_ (
);

FILL FILL_2__343_ (
);

FILL FILL_5__487_ (
);

FILL FILL_6__429_ (
);

FILL FILL_1__365_ (
);

FILL FILL_8__331_ (
);

FILL FILL_5__296_ (
);

FILL FILL_3__514_ (
);

FILL FILL_4__301_ (
);

FILL FILL_7__445_ (
);

FILL FILL_0__387_ (
);

FILL FILL_2__381_ (
);

FILL FILL_3__323_ (
);

FILL FILL_6__467_ (
);

DFFPOSX1 _602_ (
    .D(_4_),
    .CLK(clk_bF$buf5),
    .Q(Yin1[0])
);

FILL FILL_4__530_ (
);

FILL FILL_8__616_ (
);

FILL FILL_2__437_ (
);

FILL FILL_9__403_ (
);

FILL FILL73650x57750 (
);

FILL FILL_3__552_ (
);

FILL FILL_6__276_ (
);

INVX1 _411_ (
    .A(Xcalc[10]),
    .Y(_157_)
);

FILL FILL_7__483_ (
);

FILL FILL_1__459_ (
);

FILL FILL_8__425_ (
);

FILL FILL_3__361_ (
);

FILL FILL_7__539_ (
);

FILL FILL_7__292_ (
);

FILL FILL_2__475_ (
);

FILL FILL_9__441_ (
);

FILL FILL_3__417_ (
);

FILL FILL_4__624_ (
);

FILL FILL_7__348_ (
);

FILL FILL_5__411_ (
);

FILL FILL_1__497_ (
);

FILL FILL_8__463_ (
);

FILL FILL_2__284_ (
);

FILL FILL_0__502_ (
);

NAND2X1 _505_ (
    .A(selSign),
    .B(_237_),
    .Y(_238_)
);

FILL FILL_4__433_ (
);

FILL FILL_8__519_ (
);

FILL FILL73950x10950 (
);

FILL FILL75150x25350 (
);

FILL FILL_9__306_ (
);

FILL FILL_0__311_ (
);

FILL FILL_3__455_ (
);

OAI21X1 _314_ (
    .A(_73_),
    .B(_76_),
    .C(_77_),
    .Y(_1_)
);

FILL FILL_7__386_ (
);

FILL FILL_8__328_ (
);

FILL FILL_9__535_ (
);

FILL FILL_0__540_ (
);

NAND2X1 _543_ (
    .A(LoadCtl[0]),
    .B(Xin[0]),
    .Y(_265_)
);

FILL FILL_4__471_ (
);

FILL FILL_5__505_ (
);

FILL FILL_6__620_ (
);

FILL FILL_2__378_ (
);

FILL FILL_3__493_ (
);

FILL FILL_4__527_ (
);

NOR2X1 _352_ (
    .A(Xin0[0]),
    .B(Xin0[1]),
    .Y(_106_)
);

FILL FILL_4__280_ (
);

FILL FILL_5__314_ (
);

FILL FILL_8__366_ (
);

FILL FILL_0__405_ (
);

FILL FILL_3__549_ (
);

OR2X2 _408_ (
    .A(_154_),
    .B(_153_),
    .Y(_155_)
);

FILL FILL_4__336_ (
);

DFFPOSX1 _581_ (
    .D(_32_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[11])
);

FILL FILL_5__543_ (
);

FILL FILL_3__358_ (
);

FILL FILL_1__421_ (
);

FILL FILL_7__289_ (
);

NAND3X1 _390_ (
    .A(ISreg_bF$buf0),
    .B(Xin12b[7]),
    .C(_138_),
    .Y(_139_)
);

FILL FILL_5__352_ (
);

FILL FILL_7__501_ (
);

FILL FILL_0__443_ (
);

NAND3X1 _446_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_187_),
    .C(_185_),
    .Y(_188_)
);

FILL FILL_4__374_ (
);

FILL FILL_5__408_ (
);

FILL FILL_6__523_ (
);

FILL FILL_7__310_ (
);

FILL FILL_3__396_ (
);

FILL FILL_5__390_ (
);

FILL FILL_6__332_ (
);

FILL FILL_0__308_ (
);

FILL FILL_0__481_ (
);

FILL FILL_1__515_ (
);

OR2X2 _484_ (
    .A(_219_),
    .B(_216_),
    .Y(_220_)
);

FILL FILL_2__302_ (
);

FILL FILL_5__446_ (
);

FILL FILL_8__498_ (
);

FILL FILL_0__537_ (
);

FILL FILL_9__285_ (
);

FILL FILL_0__290_ (
);

FILL FILL_1__324_ (
);

FILL FILL_4__468_ (
);

OAI21X1 _293_ (
    .A(selXY_bF$buf2),
    .B(_61_),
    .C(_62_),
    .Y(_272_[6])
);

FILL FILL_2__531_ (
);

FILL FILL_6__617_ (
);

FILL FILL_6__370_ (
);

FILL FILL_7__404_ (
);

FILL FILL_0__346_ (
);

INVX1 _349_ (
    .A(Xin1[0]),
    .Y(_103_)
);

FILL FILL_1__553_ (
);

FILL FILL_4__277_ (
);

FILL FILL_2__340_ (
);

FILL FILL_5__484_ (
);

FILL FILL_6__426_ (
);

FILL FILL_3__299_ (
);

DFFPOSX1 _578_ (
    .D(_29_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[8])
);

FILL FILL_1__362_ (
);

FILL FILL_5__293_ (
);

FILL FILL_3__511_ (
);

FILL FILL_9__379_ (
);

FILL FILL_7__442_ (
);

FILL FILL_0__384_ (
);

FILL FILL_1__418_ (
);

OAI21X1 _387_ (
    .A(_96__bF$buf3),
    .B(_135_),
    .C(_136_),
    .Y(_15_)
);

FILL FILL_2__625_ (
);

FILL FILL_5__349_ (
);

FILL FILL_3__320_ (
);

FILL FILL_6__464_ (
);

FILL FILL_8__613_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_1_BUFX2_insert21 (
);

FILL FILL_1_BUFX2_insert22 (
);

FILL FILL_1_BUFX2_insert23 (
);

FILL FILL_1_BUFX2_insert24 (
);

FILL FILL_1_BUFX2_insert25 (
);

FILL FILL_2__434_ (
);

FILL FILL_6__273_ (
);

FILL FILL_7__307_ (
);

FILL FILL_7__480_ (
);

FILL FILL_1__456_ (
);

FILL FILL_8__422_ (
);

FILL FILL_6_CLKBUF1_insert0 (
);

FILL FILL_6_CLKBUF1_insert1 (
);

FILL FILL_6_CLKBUF1_insert2 (
);

FILL FILL_6_CLKBUF1_insert3 (
);

FILL FILL_6_CLKBUF1_insert4 (
);

FILL FILL_6_CLKBUF1_insert5 (
);

FILL FILL_6_CLKBUF1_insert6 (
);

FILL FILL_5__387_ (
);

FILL FILL_6__329_ (
);

FILL FILL_7__536_ (
);

FILL FILL_0__478_ (
);

FILL FILL_2__472_ (
);

FILL FILL_3__414_ (
);

FILL FILL_4__621_ (
);

FILL FILL_7__345_ (
);

FILL FILL_0__287_ (
);

FILL FILL_1__494_ (
);

FILL FILL_8__460_ (
);

FILL FILL_2__528_ (
);

FILL FILL_2__281_ (
);

FILL FILL_6__367_ (
);

OAI21X1 _502_ (
    .A(_69_),
    .B(LoadCtl_6_bF$buf2),
    .C(_235_),
    .Y(_31_)
);

FILL FILL_4__430_ (
);

FILL FILL_8__516_ (
);

FILL FILL_2__337_ (
);

FILL FILL_3__452_ (
);

NOR2X1 _311_ (
    .A(LoadCtl[0]),
    .B(LoadCtl[1]),
    .Y(_75_)
);

FILL FILL75150x46950 (
);

FILL FILL_7__383_ (
);

FILL FILL_1__359_ (
);

FILL FILL_8__325_ (
);

FILL FILL_3__508_ (
);

FILL FILL_6_BUFX2_insert20 (
);

FILL FILL_6_BUFX2_insert21 (
);

FILL FILL_6_BUFX2_insert22 (
);

FILL FILL_6_BUFX2_insert23 (
);

FILL FILL_6_BUFX2_insert24 (
);

FILL FILL_6_BUFX2_insert25 (
);

FILL FILL_7__439_ (
);

OAI21X1 _540_ (
    .A(_254_),
    .B(_86_),
    .C(_263_),
    .Y(_41_)
);

FILL FILL_5__502_ (
);

FILL FILL_8__554_ (
);

FILL FILL_2__375_ (
);

FILL FILL_9__341_ (
);

FILL FILL_3__317_ (
);

FILL FILL_3__490_ (
);

FILL FILL_4__524_ (
);

FILL FILL_5__311_ (
);

FILL FILL_1__397_ (
);

FILL FILL_8__363_ (
);

FILL FILL_0__402_ (
);

FILL FILL_3__546_ (
);

INVX1 _405_ (
    .A(Xcalc[9]),
    .Y(_152_)
);

FILL FILL_4__333_ (
);

FILL FILL_7__477_ (
);

FILL FILL_8__419_ (
);

FILL FILL_5__540_ (
);

FILL FILL_3__355_ (
);

FILL FILL_6__499_ (
);

FILL FILL_7__286_ (
);

FILL FILL_2__469_ (
);

FILL FILL_9__435_ (
);

FILL FILL_0__440_ (
);

FILL FILL_4__618_ (
);

OR2X2 _443_ (
    .A(_184_),
    .B(_183_),
    .Y(_185_)
);

FILL FILL_4__371_ (
);

FILL FILL_5__405_ (
);

FILL FILL_8__457_ (
);

FILL FILL_6__520_ (
);

FILL FILL_2__278_ (
);

FILL FILL_3__393_ (
);

FILL FILL_4__427_ (
);

FILL FILL_0__305_ (
);

FILL FILL_9__473_ (
);

FILL FILL_3__449_ (
);

OAI21X1 _308_ (
    .A(selXY_bF$buf2),
    .B(_71_),
    .C(_72_),
    .Y(_272_[11])
);

FILL FILL_1__512_ (
);

NOR2X1 _481_ (
    .A(Yin12b[6]),
    .B(Yin12b[7]),
    .Y(_217_)
);

FILL FILL_5__443_ (
);

FILL FILL_8__495_ (
);

FILL FILL_9__529_ (
);

FILL FILL_0__534_ (
);

FILL FILL_9__282_ (
);

NAND2X1 _537_ (
    .A(Xin[1]),
    .B(_80_),
    .Y(_262_)
);

FILL FILL75450x54150 (
);

FILL FILL_1__321_ (
);

FILL FILL_4__465_ (
);

OAI21X1 _290_ (
    .A(selXY_bF$buf2),
    .B(_59_),
    .C(_60_),
    .Y(_272_[5])
);

FILL FILL_6__614_ (
);

FILL FILL_9__338_ (
);

FILL FILL_7__401_ (
);

FILL FILL_0__343_ (
);

FILL FILL_3__487_ (
);

NAND2X1 _346_ (
    .A(_98_),
    .B(_100_),
    .Y(_101_)
);

FILL FILL_1__550_ (
);

FILL FILL_4__274_ (
);

FILL FILL_5__308_ (
);

FILL FILL_5__481_ (
);

FILL FILL_6__423_ (
);

FILL FILL_3__296_ (
);

DFFPOSX1 _575_ (
    .D(_26_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[5])
);

FILL FILL_5__537_ (
);

FILL FILL_5__290_ (
);

FILL FILL_9__376_ (
);

FILL FILL_0__381_ (
);

FILL FILL_1__415_ (
);

NAND2X1 _384_ (
    .A(_132_),
    .B(_133_),
    .Y(_134_)
);

FILL FILL_2__622_ (
);

FILL FILL_5__346_ (
);

FILL FILL_8__398_ (
);

FILL FILL_6__461_ (
);

FILL FILL_0__437_ (
);

FILL FILL_4__368_ (
);

FILL FILL_2__431_ (
);

FILL FILL_6__517_ (
);

FILL FILL_7__304_ (
);

FILL FILL_1__453_ (
);

FILL FILL_5__384_ (
);

FILL FILL_6__326_ (
);

FILL FILL_7__533_ (
);

FILL FILL_0__475_ (
);

FILL FILL_1__509_ (
);

NAND3X1 _478_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_211_),
    .C(_214_),
    .Y(_215_)
);

FILL FILL_3__411_ (
);

FILL FILL_6__555_ (
);

FILL FILL_9__279_ (
);

FILL FILL_7__342_ (
);

FILL FILL_0__284_ (
);

FILL FILL_1__318_ (
);

OAI21X1 _287_ (
    .A(selXY_bF$buf0),
    .B(_57_),
    .C(_58_),
    .Y(_272_[4])
);

FILL FILL_1__491_ (
);

FILL FILL_2__525_ (
);

FILL FILL_6__364_ (
);

FILL FILL_1__547_ (
);

FILL FILL_8__513_ (
);

FILL FILL_2__334_ (
);

FILL FILL_9__300_ (
);

FILL FILL_5__478_ (
);

FILL FILL_7__380_ (
);

FILL FILL_1__356_ (
);

FILL FILL_8__322_ (
);

FILL FILL_5__287_ (
);

FILL FILL_3__505_ (
);

FILL FILL_7__436_ (
);

FILL FILL_0__378_ (
);

FILL FILL_8__551_ (
);

FILL FILL_2__619_ (
);

FILL FILL_2__372_ (
);

FILL FILL_3__314_ (
);

FILL FILL_6__458_ (
);

FILL FILL_4__521_ (
);

FILL FILL_1__394_ (
);

FILL FILL_8__360_ (
);

FILL FILL_2__428_ (
);

FILL FILL_3__543_ (
);

NAND2X1 _402_ (
    .A(_149_),
    .B(_148_),
    .Y(_150_)
);

FILL FILL_4__330_ (
);

FILL FILL_7__474_ (
);

FILL FILL_8__416_ (
);

FILL FILL_9__623_ (
);

FILL FILL_3__352_ (
);

FILL FILL_6__496_ (
);

FILL FILL_7__283_ (
);

FILL FILL_2__466_ (
);

FILL FILL_9__432_ (
);

FILL FILL_3__408_ (
);

FILL FILL_4__615_ (
);

FILL FILL_7__339_ (
);

OAI21X1 _440_ (
    .A(_51_),
    .B(LoadCtl_6_bF$buf4),
    .C(_182_),
    .Y(_22_)
);

FILL FILL_5__402_ (
);

FILL FILL_1__488_ (
);

FILL FILL_8__454_ (
);

FILL FILL_2__275_ (
);

FILL FILL_3__390_ (
);

FILL FILL_4__424_ (
);

FILL FILL_1__297_ (
);

FILL FILL_0__302_ (
);

FILL FILL_9__470_ (
);

FILL FILL_3__446_ (
);

OAI21X1 _305_ (
    .A(selXY_bF$buf1),
    .B(_69_),
    .C(_70_),
    .Y(_272_[10])
);

FILL FILL_7__377_ (
);

FILL FILL_8__319_ (
);

FILL FILL_5__440_ (
);

FILL FILL_8__492_ (
);

FILL FILL_9__526_ (
);

FILL FILL_0__531_ (
);

FILL FILL_6__399_ (
);

OAI21X1 _534_ (
    .A(_257_),
    .B(_76_),
    .C(_260_),
    .Y(_38_)
);

FILL FILL_4__462_ (
);

FILL FILL_8__548_ (
);

FILL FILL_2__369_ (
);

FILL FILL_9__335_ (
);

FILL FILL_0__340_ (
);

FILL FILL_3__484_ (
);

FILL FILL_4__518_ (
);

NAND3X1 _343_ (
    .A(ISreg_bF$buf1),
    .B(Xin0[0]),
    .C(Xin0[1]),
    .Y(_98_)
);

FILL FILL_5__305_ (
);

FILL FILL_8__357_ (
);

FILL FILL74250x57750 (
);

FILL FILL_6__420_ (
);

FILL FILL_3__293_ (
);

FILL FILL_4__327_ (
);

DFFPOSX1 _572_ (
    .D(_23_),
    .CLK(clk_bF$buf0),
    .Q(Ycalc[2])
);

FILL FILL73950x72150 (
);

FILL FILL_5__534_ (
);

FILL FILL_0__625_ (
);

FILL FILL_9__373_ (
);

FILL FILL_3__349_ (
);

FILL FILL_1__412_ (
);

FILL FILL_4__556_ (
);

NAND3X1 _381_ (
    .A(ISreg_bF$buf0),
    .B(Xin12b[6]),
    .C(_130_),
    .Y(_131_)
);

FILL FILL_5__343_ (
);

FILL FILL_8__395_ (
);

FILL FILL_9__429_ (
);

FILL FILL_0__434_ (
);

NAND3X1 _437_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf2),
    .Y(_180_)
);

FILL FILL_4__365_ (
);

FILL FILL_6__514_ (
);

FILL FILL74550x10950 (
);

FILL FILL_7__301_ (
);

FILL FILL_3__387_ (
);

FILL FILL_1__450_ (
);

FILL FILL_5__381_ (
);

FILL FILL_6__323_ (
);

FILL FILL_9__467_ (
);

FILL FILL_7__530_ (
);

FILL FILL_0__472_ (
);

FILL FILL_1__506_ (
);

INVX1 _475_ (
    .A(Yin12b[7]),
    .Y(_212_)
);

FILL FILL_5__437_ (
);

FILL FILL_8__489_ (
);

FILL FILL_6__552_ (
);

FILL FILL_0__528_ (
);

FILL FILL_9__276_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_2_BUFX2_insert12 (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_2_BUFX2_insert17 (
);

FILL FILL_2_BUFX2_insert18 (
);

FILL FILL_2_BUFX2_insert19 (
);

FILL FILL_0__281_ (
);

FILL FILL_1__315_ (
);

FILL FILL_4__459_ (
);

OAI21X1 _284_ (
    .A(selXY_bF$buf0),
    .B(_55_),
    .C(_56_),
    .Y(_272_[3])
);

FILL FILL_2__522_ (
);

FILL FILL_8__298_ (
);

FILL FILL_6__361_ (
);

FILL FILL_0__337_ (
);

FILL FILL_1__544_ (
);

FILL FILL_8__510_ (
);

FILL FILL_2__331_ (
);

FILL FILL_5__475_ (
);

FILL FILL_6__417_ (
);

FILL FILL_7__624_ (
);

DFFPOSX1 _569_ (
    .D(_20_),
    .CLK(clk_bF$buf2),
    .Q(Xcalc[11])
);

FILL FILL_1__353_ (
);

FILL FILL_4__497_ (
);

FILL FILL_4_CLKBUF1_insert0 (
);

FILL FILL_4_CLKBUF1_insert1 (
);

FILL FILL_4_CLKBUF1_insert2 (
);

FILL FILL_4_CLKBUF1_insert3 (
);

FILL FILL_4_CLKBUF1_insert4 (
);

FILL FILL_4_CLKBUF1_insert5 (
);

FILL FILL_4_CLKBUF1_insert6 (
);

FILL FILL_5__284_ (
);

FILL FILL_3__502_ (
);

FILL FILL_7__433_ (
);

FILL FILL_0__375_ (
);

FILL FILL_1__409_ (
);

OAI21X1 _378_ (
    .A(_96__bF$buf2),
    .B(_127_),
    .C(_128_),
    .Y(_14_)
);

FILL FILL_2__616_ (
);

FILL FILL_3__311_ (
);

FILL FILL_6__455_ (
);

FILL FILL_1__391_ (
);

FILL FILL_2__425_ (
);

FILL FILL_3__540_ (
);

FILL FILL_7__471_ (
);

FILL FILL_1__447_ (
);

FILL FILL_8__413_ (
);

FILL FILL_9__620_ (
);

FILL FILL_5__378_ (
);

FILL FILL_6__493_ (
);

FILL FILL_7__527_ (
);

FILL FILL_0__469_ (
);

FILL FILL_7__280_ (
);

FILL FILL_2__463_ (
);

FILL FILL_3__405_ (
);

FILL FILL_6__549_ (
);

FILL FILL_7__336_ (
);

FILL FILL_0__278_ (
);

FILL FILL_1__485_ (
);

FILL FILL_8__451_ (
);

FILL FILL_2__519_ (
);

FILL FILL_6__358_ (
);

FILL FILL_4__421_ (
);

FILL FILL_8__507_ (
);

FILL FILL_1__294_ (
);

FILL FILL_2__328_ (
);

FILL FILL_3__443_ (
);

OAI21X1 _302_ (
    .A(selXY_bF$buf1),
    .B(_67_),
    .C(_68_),
    .Y(_272_[9])
);

FILL FILL_7__374_ (
);

FILL FILL_8__316_ (
);

FILL FILL_9__523_ (
);

FILL FILL_6__396_ (
);

NAND2X1 _531_ (
    .A(Xin12b[6]),
    .B(_76_),
    .Y(_259_)
);

FILL FILL_8__545_ (
);

FILL FILL_2__366_ (
);

FILL FILL_9__332_ (
);

FILL FILL_3__308_ (
);

FILL FILL_3__481_ (
);

FILL FILL_4__515_ (
);

INVX8 _340_ (
    .A(LoadCtl_6_bF$buf4),
    .Y(_96_)
);

FILL FILL_5__302_ (
);

FILL FILL_1__388_ (
);

FILL FILL_8__354_ (
);

FILL FILL_3__537_ (
);

FILL FILL_3__290_ (
);

FILL FILL_4__324_ (
);

FILL FILL_7__468_ (
);

FILL FILL_5__531_ (
);

FILL FILL_9__617_ (
);

FILL FILL_0__622_ (
);

FILL FILL_3__346_ (
);

BUFX2 _625_ (
    .A(LoadCtl_6_bF$buf2),
    .Y(Vld)
);

FILL FILL_4__553_ (
);

FILL FILL_7__277_ (
);

FILL FILL_5__340_ (
);

FILL FILL_8__392_ (
);

FILL FILL_9__426_ (
);

FILL FILL_0__431_ (
);

FILL FILL_6__299_ (
);

NAND2X1 _434_ (
    .A(_166_),
    .B(_178_),
    .Y(_20_)
);

FILL FILL_4__362_ (
);

FILL FILL_8__448_ (
);

FILL FILL_6__511_ (
);

FILL FILL_3__384_ (
);

FILL FILL_4__418_ (
);

FILL FILL_5__625_ (
);

FILL FILL_6__320_ (
);

FILL FILL_2__498_ (
);

FILL FILL_1__503_ (
);

OAI21X1 _472_ (
    .A(_61_),
    .B(LoadCtl_6_bF$buf1),
    .C(_209_),
    .Y(_27_)
);

FILL FILL_5__434_ (
);

FILL FILL_8__486_ (
);

FILL FILL75450x61350 (
);

FILL FILL75450x28950 (
);

FILL FILL_0__525_ (
);

INVX1 _528_ (
    .A(Xin[1]),
    .Y(_257_)
);

FILL FILL_1__312_ (
);

FILL FILL_4__456_ (
);

OAI21X1 _281_ (
    .A(selXY_bF$buf3),
    .B(_53_),
    .C(_54_),
    .Y(_272_[2])
);

FILL FILL_8__295_ (
);

FILL FILL_0__334_ (
);

FILL FILL_3__478_ (
);

NAND2X1 _337_ (
    .A(ISin),
    .B(LoadCtl_6_bF$buf1),
    .Y(_94_)
);

FILL FILL_1__541_ (
);

FILL FILL_5__472_ (
);

FILL FILL_6__414_ (
);

FILL FILL_7__621_ (
);

FILL FILL_3__287_ (
);

DFFPOSX1 _566_ (
    .D(_17_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[8])
);

FILL FILL_1__350_ (
);

FILL FILL_4__494_ (
);

FILL FILL_5__528_ (
);

FILL FILL_5__281_ (
);

FILL FILL_0__619_ (
);

FILL FILL_7__430_ (
);

FILL FILL_0__372_ (
);

FILL FILL_1__406_ (
);

NAND2X1 _375_ (
    .A(_123_),
    .B(_124_),
    .Y(_126_)
);

FILL FILL_2__613_ (
);

FILL FILL_5__337_ (
);

FILL FILL_8__389_ (
);

FILL FILL_6__452_ (
);

FILL FILL_0__428_ (
);

FILL FILL_4__359_ (
);

FILL FILL_2__422_ (
);

FILL FILL_6__508_ (
);

FILL FILL_1__444_ (
);

FILL FILL_8__410_ (
);

FILL FILL_5__375_ (
);

FILL FILL_6__317_ (
);

FILL FILL_6__490_ (
);

FILL FILL_7__524_ (
);

FILL FILL_0__466_ (
);

NAND2X1 _469_ (
    .A(ISreg_bF$buf4),
    .B(_204_),
    .Y(_207_)
);

FILL FILL_4__397_ (
);

FILL FILL_2__460_ (
);

FILL FILL_3__402_ (
);

FILL FILL_6__546_ (
);

FILL FILL_7__333_ (
);

FILL FILL_0__275_ (
);

FILL FILL_1__309_ (
);

OAI21X1 _278_ (
    .A(selXY_bF$buf3),
    .B(_51_),
    .C(_52_),
    .Y(_272_[1])
);

FILL FILL_1__482_ (
);

FILL FILL_2__516_ (
);

FILL FILL75750x36150 (
);

FILL FILL_6__355_ (
);

FILL FILL_9__499_ (
);

FILL FILL_1__538_ (
);

FILL FILL_8__504_ (
);

FILL FILL_1__291_ (
);

FILL FILL_2__325_ (
);

FILL FILL_5__469_ (
);

FILL FILL_3__440_ (
);

FILL FILL_7__618_ (
);

FILL FILL_7__371_ (
);

FILL FILL_1__347_ (
);

FILL FILL_8__313_ (
);

FILL FILL_2__554_ (
);

FILL FILL_9__520_ (
);

FILL FILL_5__278_ (
);

FILL FILL_6__393_ (
);

FILL FILL_7__427_ (
);

FILL FILL_0__369_ (
);

FILL FILL_8__542_ (
);

FILL FILL_2__363_ (
);

FILL FILL_3__305_ (
);

FILL FILL_6__449_ (
);

FILL FILL_4__512_ (
);

FILL FILL_1__385_ (
);

FILL FILL_8__351_ (
);

FILL FILL_2__419_ (
);

FILL FILL_3__534_ (
);

FILL FILL_4__321_ (
);

FILL FILL_7__465_ (
);

FILL FILL_8__407_ (
);

FILL FILL_3__343_ (
);

FILL FILL_6__487_ (
);

BUFX2 _622_ (
    .A(_272_[7]),
    .Y(Dout[7])
);

FILL FILL_4__550_ (
);

FILL FILL_7__274_ (
);

FILL FILL_2__457_ (
);

FILL FILL_6__296_ (
);

NAND3X1 _431_ (
    .A(_175_),
    .B(_173_),
    .C(_147_),
    .Y(_176_)
);

FILL FILL_1__479_ (
);

FILL FILL_8__445_ (
);

FILL FILL_3__381_ (
);

FILL FILL_4__415_ (
);

FILL FILL_5__622_ (
);

FILL FILL_1__288_ (
);

FILL FILL_2__495_ (
);

FILL FILL_3__437_ (
);

FILL FILL_1__500_ (
);

FILL FILL_7__368_ (
);

FILL FILL_5__431_ (
);

FILL FILL_8__483_ (
);

FILL FILL_0__522_ (
);

NAND2X1 _525_ (
    .A(LoadCtl[4]),
    .B(_249_),
    .Y(_255_)
);

FILL FILL_4__453_ (
);

FILL FILL_8__539_ (
);

FILL FILL_8__292_ (
);

FILL FILL_9__326_ (
);

FILL FILL_0__331_ (
);

FILL FILL_3__475_ (
);

FILL FILL_4__509_ (
);

NAND2X1 _334_ (
    .A(LoadCtl[0]),
    .B(Yin[1]),
    .Y(_92_)
);

FILL FILL_8__348_ (
);

FILL FILL_6__411_ (
);

FILL FILL_9__555_ (
);

FILL FILL_3__284_ (
);

FILL FILL_4__318_ (
);

DFFPOSX1 _563_ (
    .D(_14_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[5])
);

FILL FILL_4__491_ (
);

FILL FILL_5__525_ (
);

FILL FILL_2__398_ (
);

FILL FILL_0__616_ (
);

FILL FILL_9__364_ (
);

BUFX2 _619_ (
    .A(_272_[4]),
    .Y(Dout[4])
);

FILL FILL_1__403_ (
);

FILL FILL_4__547_ (
);

INVX1 _372_ (
    .A(Xin12b[5]),
    .Y(_123_)
);

FILL FILL_5__334_ (
);

FILL FILL_8__386_ (
);

FILL FILL_0__425_ (
);

NAND2X1 _428_ (
    .A(ISreg_bF$buf2),
    .B(Xin12b[10]),
    .Y(_173_)
);

FILL FILL_4__356_ (
);

FILL FILL_6__505_ (
);

FILL FILL_3__378_ (
);

FILL FILL_1__441_ (
);

FILL FILL_5__619_ (
);

FILL FILL_3_BUFX2_insert20 (
);

FILL FILL_3_BUFX2_insert21 (
);

FILL FILL_3_BUFX2_insert22 (
);

FILL FILL_3_BUFX2_insert23 (
);

FILL FILL_3_BUFX2_insert24 (
);

FILL FILL_3_BUFX2_insert25 (
);

FILL FILL_5__372_ (
);

FILL FILL_6__314_ (
);

FILL FILL_9__458_ (
);

FILL FILL_7__521_ (
);

FILL FILL_0__463_ (
);

NAND2X1 _466_ (
    .A(_203_),
    .B(_197_),
    .Y(_204_)
);

FILL FILL_2_CLKBUF1_insert0 (
);

FILL FILL_2_CLKBUF1_insert1 (
);

FILL FILL_2_CLKBUF1_insert2 (
);

FILL FILL_2_CLKBUF1_insert3 (
);

FILL FILL_2_CLKBUF1_insert4 (
);

FILL FILL_2_CLKBUF1_insert5 (
);

FILL FILL_2_CLKBUF1_insert6 (
);

FILL FILL_4__394_ (
);

FILL FILL_5__428_ (
);

FILL FILL_6__543_ (
);

FILL FILL_0__519_ (
);

FILL FILL_7__330_ (
);

FILL FILL_1__306_ (
);

OAI21X1 _275_ (
    .A(selXY_bF$buf3),
    .B(_49_),
    .C(_50_),
    .Y(_272_[0])
);

FILL FILL_2__513_ (
);

FILL FILL_8__289_ (
);

FILL FILL_6__352_ (
);

FILL FILL_0__328_ (
);

FILL FILL_9__496_ (
);

FILL FILL_1__535_ (
);

FILL FILL_8__501_ (
);

FILL FILL75750x57750 (
);

FILL FILL_2__322_ (
);

FILL FILL_5__466_ (
);

FILL FILL_6__408_ (
);

FILL FILL_7__615_ (
);

FILL FILL74550x72150 (
);

FILL FILL74550x39750 (
);

FILL FILL_1__344_ (
);

FILL FILL_8__310_ (
);

FILL FILL_4__488_ (
);

FILL FILL_2__551_ (
);

FILL FILL_5__275_ (
);

FILL FILL_6__390_ (
);

FILL FILL_7__424_ (
);

FILL FILL_0__366_ (
);

FILL FILL73050x28950 (
);

NAND2X1 _369_ (
    .A(_117_),
    .B(_120_),
    .Y(_121_)
);

FILL FILL_4__297_ (
);

FILL FILL_2__360_ (
);

FILL FILL_3__302_ (
);

FILL FILL_6__446_ (
);

FILL FILL_8_BUFX2_insert20 (
);

FILL FILL_8_BUFX2_insert21 (
);

FILL FILL_8_BUFX2_insert22 (
);

FILL FILL_8_BUFX2_insert23 (
);

FILL FILL_8_BUFX2_insert24 (
);

FILL FILL_8_BUFX2_insert25 (
);

DFFPOSX1 _598_ (
    .D(_0_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[6])
);

FILL FILL_1__382_ (
);

FILL FILL_2__416_ (
);

FILL FILL_3__531_ (
);

FILL FILL_9__399_ (
);

FILL FILL_7__462_ (
);

FILL FILL_1__438_ (
);

FILL FILL_8__404_ (
);

FILL FILL_5__369_ (
);

FILL FILL_3__340_ (
);

FILL FILL_6__484_ (
);

FILL FILL_7__518_ (
);

FILL FILL_2__454_ (
);

FILL FILL_9__420_ (
);

FILL FILL_6__293_ (
);

FILL FILL_7__327_ (
);

FILL FILL_1__476_ (
);

FILL FILL_8__442_ (
);

FILL FILL_3__625_ (
);

FILL FILL_6__349_ (
);

FILL FILL_4__412_ (
);

FILL FILL_7__556_ (
);

FILL FILL_0__498_ (
);

FILL FILL_1__285_ (
);

FILL FILL_2__319_ (
);

FILL FILL_2__492_ (
);

FILL FILL_3__434_ (
);

FILL FILL_7__365_ (
);

FILL FILL_8__307_ (
);

FILL FILL_8__480_ (
);

FILL FILL_2__548_ (
);

FILL FILL_9__514_ (
);

FILL FILL_6__387_ (
);

NAND2X1 _522_ (
    .A(Xin[1]),
    .B(_251_),
    .Y(_253_)
);

FILL FILL_4__450_ (
);

FILL FILL_8__536_ (
);

FILL FILL_2__357_ (
);

FILL FILL_9__323_ (
);

FILL FILL_3__472_ (
);

FILL FILL_4__506_ (
);

NAND2X1 _331_ (
    .A(LoadCtl[0]),
    .B(Yin[0]),
    .Y(_90_)
);

FILL FILL_1__379_ (
);

FILL FILL_8__345_ (
);

FILL FILL_9__552_ (
);

FILL FILL_3__528_ (
);

FILL FILL_3__281_ (
);

FILL FILL_4__315_ (
);

FILL FILL_7__459_ (
);

DFFPOSX1 _560_ (
    .D(_11_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[2])
);

FILL FILL_5__522_ (
);

FILL FILL_2__395_ (
);

FILL FILL_0__613_ (
);

FILL FILL_9__361_ (
);

FILL FILL_3__337_ (
);

BUFX2 _616_ (
    .A(_272_[11]),
    .Y(Dout[11])
);

FILL FILL_1__400_ (
);

FILL FILL_4__544_ (
);

FILL FILL_5__331_ (
);

FILL FILL_8__383_ (
);

FILL FILL_9__417_ (
);

FILL FILL_0__422_ (
);

NAND2X1 _425_ (
    .A(Xin12b[11]),
    .B(_169_),
    .Y(_170_)
);

FILL FILL_4__353_ (
);

FILL FILL_7__497_ (
);

FILL FILL_8__439_ (
);

FILL FILL_6__502_ (
);

FILL FILL_3__375_ (
);

FILL FILL_4__409_ (
);

FILL FILL_5__616_ (
);

FILL FILL_6__311_ (
);

FILL FILL_2__489_ (
);

FILL FILL_9__455_ (
);

FILL FILL_0__460_ (
);

AOI21X1 _463_ (
    .A(_200_),
    .B(_82_),
    .C(_96__bF$buf1),
    .Y(_202_)
);

FILL FILL_4__391_ (
);

FILL FILL_5__425_ (
);

FILL FILL_8__477_ (
);

FILL FILL_6__540_ (
);

FILL FILL_2__298_ (
);

FILL FILL_0__516_ (
);

NOR2X1 _519_ (
    .A(LoadCtl[4]),
    .B(_250_),
    .Y(_251_)
);

FILL FILL_1__303_ (
);

FILL FILL_4__447_ (
);

FILL FILL_2__510_ (
);

FILL FILL_8__286_ (
);

FILL FILL_0__325_ (
);

FILL FILL_9__493_ (
);

FILL FILL_3__469_ (
);

OAI21X1 _328_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[1]),
    .Y(_88_)
);

FILL FILL_1__532_ (
);

FILL FILL_5__463_ (
);

FILL FILL_6__405_ (
);

FILL FILL_9__549_ (
);

FILL FILL_0__554_ (
);

FILL FILL_3__278_ (
);

DFFPOSX1 _557_ (
    .D(_8_),
    .CLK(clk_bF$buf4),
    .Q(ISreg)
);

FILL FILL_1__341_ (
);

FILL FILL_4__485_ (
);

FILL FILL_5__519_ (
);

FILL FILL_9__358_ (
);

FILL FILL_7__421_ (
);

FILL FILL_0__363_ (
);

INVX1 _366_ (
    .A(Xin12b[4]),
    .Y(_118_)
);

FILL FILL_4__294_ (
);

FILL FILL_5__328_ (
);

FILL FILL75750x7350 (
);

FILL FILL_6__443_ (
);

FILL FILL_0__419_ (
);

DFFPOSX1 _595_ (
    .D(_46_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[11])
);

FILL FILL_2__413_ (
);

FILL FILL_9__396_ (
);

FILL FILL_1__435_ (
);

FILL FILL_8__401_ (
);

FILL FILL_5__366_ (
);

FILL FILL_6__308_ (
);

FILL FILL_6__481_ (
);

FILL FILL_7__515_ (
);

FILL FILL_0__457_ (
);

FILL FILL_4__388_ (
);

FILL FILL_2__451_ (
);

FILL FILL_6__537_ (
);

FILL FILL_6__290_ (
);

FILL FILL_7__324_ (
);

FILL FILL_1__473_ (
);

FILL FILL_2__507_ (
);

FILL FILL_3__622_ (
);

FILL FILL_6__346_ (
);

FILL FILL74550x25350 (
);

FILL FILL_7__553_ (
);

FILL FILL_0__495_ (
);

FILL FILL_1__529_ (
);

INVX1 _498_ (
    .A(Yin12b[10]),
    .Y(_232_)
);

FILL FILL_1__282_ (
);

FILL FILL_2__316_ (
);

FILL FILL_3__431_ (
);

FILL FILL_7__362_ (
);

FILL FILL_1__338_ (
);

FILL FILL_8__304_ (
);

FILL FILL_2__545_ (
);

FILL FILL_9__511_ (
);

FILL FILL_6__384_ (
);

FILL FILL_7__418_ (
);

FILL FILL_8__533_ (
);

FILL FILL_2__354_ (
);

FILL FILL_9__320_ (
);

FILL FILL_5__498_ (
);

FILL FILL_4__503_ (
);

FILL FILL_1__376_ (
);

FILL FILL_8__342_ (
);

FILL FILL_3__525_ (
);

FILL FILL73350x57750 (
);

FILL FILL_4__312_ (
);

FILL FILL_7__456_ (
);

FILL FILL_0__398_ (
);

FILL FILL_2__392_ (
);

FILL FILL_3__334_ (
);

FILL FILL_6__478_ (
);

BUFX2 _613_ (
    .A(_272_[0]),
    .Y(Dout[0])
);

FILL FILL_4__541_ (
);

FILL FILL_8__380_ (
);

FILL FILL_2__448_ (
);

FILL FILL_9__414_ (
);

FILL FILL_6__287_ (
);

INVX1 _422_ (
    .A(Xin12b[11]),
    .Y(_167_)
);

FILL FILL_4__350_ (
);

FILL FILL_7__494_ (
);

FILL FILL_8__436_ (
);

FILL FILL_3__619_ (
);

FILL FILL_3__372_ (
);

FILL FILL_4__406_ (
);

FILL FILL73650x10950 (
);

FILL FILL_5__613_ (
);

FILL FILL_1__279_ (
);

FILL FILL_2__486_ (
);

FILL FILL_9__452_ (
);

FILL FILL_3__428_ (
);

FILL FILL_7__359_ (
);

OAI21X1 _460_ (
    .A(_57_),
    .B(LoadCtl_6_bF$buf0),
    .C(_199_),
    .Y(_25_)
);

FILL FILL_5__422_ (
);

FILL FILL_8__474_ (
);

FILL FILL_9__508_ (
);

FILL FILL_2__295_ (
);

FILL FILL_0__513_ (
);

NOR2X1 _516_ (
    .A(LoadCtl[2]),
    .B(LoadCtl[3]),
    .Y(_248_)
);

FILL FILL_1__300_ (
);

FILL FILL_4__444_ (
);

FILL FILL_8__283_ (
);

FILL FILL_9__317_ (
);

FILL FILL_0__322_ (
);

FILL FILL_9__490_ (
);

FILL FILL_3__466_ (
);

FILL FILL_4_BUFX2_insert10 (
);

FILL FILL_4_BUFX2_insert11 (
);

OR2X2 _325_ (
    .A(_85_),
    .B(LoadCtl[0]),
    .Y(_86_)
);

FILL FILL_4_BUFX2_insert12 (
);

FILL FILL_4_BUFX2_insert13 (
);

FILL FILL_4_BUFX2_insert14 (
);

FILL FILL_4_BUFX2_insert15 (
);

FILL FILL_4_BUFX2_insert16 (
);

FILL FILL_4_BUFX2_insert17 (
);

FILL FILL_4_BUFX2_insert18 (
);

FILL FILL_4_BUFX2_insert19 (
);

FILL FILL_7__397_ (
);

FILL FILL_8__339_ (
);

FILL FILL_5__460_ (
);

FILL FILL_6__402_ (
);

FILL FILL_9__546_ (
);

FILL FILL_0__551_ (
);

FILL FILL_3__275_ (
);

FILL FILL_4__309_ (
);

OAI21X1 _554_ (
    .A(_73_),
    .B(_255_),
    .C(_270_),
    .Y(_48_)
);

FILL FILL_4__482_ (
);

FILL FILL_5__516_ (
);

FILL FILL_2__389_ (
);

FILL FILL_0__360_ (
);

FILL FILL_0_CLKBUF1_insert0 (
);

FILL FILL_0_CLKBUF1_insert1 (
);

FILL FILL_0_CLKBUF1_insert2 (
);

FILL FILL_0_CLKBUF1_insert3 (
);

FILL FILL_0_CLKBUF1_insert4 (
);

FILL FILL_0_CLKBUF1_insert5 (
);

FILL FILL_4__538_ (
);

FILL FILL_0_CLKBUF1_insert6 (
);

NOR2X1 _363_ (
    .A(Xin1[0]),
    .B(Xin1[1]),
    .Y(_115_)
);

FILL FILL_4__291_ (
);

FILL FILL_5__325_ (
);

FILL FILL_8__377_ (
);

FILL FILL_6__440_ (
);

FILL FILL_0__416_ (
);

NAND3X1 _419_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_161_),
    .C(_164_),
    .Y(_165_)
);

FILL FILL_1__623_ (
);

FILL FILL_4__347_ (
);

DFFPOSX1 _592_ (
    .D(_43_),
    .CLK(clk_bF$buf2),
    .Q(Xin0[0])
);

FILL FILL_2__410_ (
);

FILL FILL_5__554_ (
);

FILL FILL_3__369_ (
);

FILL FILL_1__432_ (
);

FILL FILL_5__363_ (
);

FILL FILL_6__305_ (
);

FILL FILL_7__512_ (
);

FILL FILL_0__454_ (
);

AND2X2 _457_ (
    .A(_186_),
    .B(_193_),
    .Y(_197_)
);

FILL FILL_4__385_ (
);

FILL FILL_5__419_ (
);

FILL FILL_6__534_ (
);

FILL FILL_7__321_ (
);

FILL FILL_1__470_ (
);

FILL FILL_2__504_ (
);

FILL FILL_6__343_ (
);

FILL FILL_0__319_ (
);

FILL FILL_7__550_ (
);

FILL FILL_0__492_ (
);

FILL FILL_1__526_ (
);

NOR2X1 _495_ (
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .Y(_229_)
);

FILL FILL_2__313_ (
);

FILL FILL_5__457_ (
);

FILL FILL_0__548_ (
);

FILL FILL_9__296_ (
);

FILL FILL_1__335_ (
);

FILL FILL_8__301_ (
);

FILL FILL_4__479_ (
);

FILL FILL_2__542_ (
);

FILL FILL_6__381_ (
);

FILL FILL_7__415_ (
);

FILL FILL_0__357_ (
);

FILL FILL_8__530_ (
);

FILL FILL_4__288_ (
);

FILL FILL_2__351_ (
);

FILL FILL_5__495_ (
);

FILL FILL_6__437_ (
);

FILL FILL_4__500_ (
);

DFFPOSX1 _589_ (
    .D(_40_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[5])
);

FILL FILL_1__373_ (
);

FILL FILL_2__407_ (
);

FILL FILL_3__522_ (
);

FILL FILL_7__453_ (
);

FILL FILL_0__395_ (
);

FILL FILL_1__429_ (
);

NAND2X1 _398_ (
    .A(_129_),
    .B(_145_),
    .Y(_146_)
);

FILL FILL_3__331_ (
);

FILL FILL_6__475_ (
);

FILL FILL_7__509_ (
);

DFFPOSX1 _610_ (
    .D(LoadCtl[3]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[4])
);

FILL FILL_8__624_ (
);

FILL FILL_2__445_ (
);

FILL FILL_9__411_ (
);

FILL FILL_6__284_ (
);

FILL FILL_7__318_ (
);

FILL FILL_7__491_ (
);

FILL FILL_1__467_ (
);

FILL FILL_8__433_ (
);

FILL FILL_5__398_ (
);

FILL FILL_3__616_ (
);

FILL FILL_8_BUFX2_insert7 (
);

FILL FILL_8_BUFX2_insert8 (
);

FILL FILL_8_BUFX2_insert9 (
);

FILL FILL_4__403_ (
);

FILL FILL_7__547_ (
);

FILL FILL_0__489_ (
);

FILL FILL_1__276_ (
);

FILL FILL_2__483_ (
);

FILL FILL_3__425_ (
);

FILL FILL_7__356_ (
);

FILL FILL_0__298_ (
);

FILL FILL_8__471_ (
);

FILL FILL_2__539_ (
);

FILL FILL_9__505_ (
);

FILL FILL_2__292_ (
);

FILL FILL_0__510_ (
);

FILL FILL_6__378_ (
);

NAND2X1 _513_ (
    .A(_240_),
    .B(_245_),
    .Y(_246_)
);

FILL FILL_4__441_ (
);

FILL FILL_9_CLKBUF1_insert0 (
);

FILL FILL_9_CLKBUF1_insert1 (
);

FILL FILL_9_CLKBUF1_insert2 (
);

FILL FILL_9_CLKBUF1_insert4 (
);

FILL FILL_8__527_ (
);

FILL FILL_9_CLKBUF1_insert5 (
);

FILL FILL_9_CLKBUF1_insert6 (
);

FILL FILL_8__280_ (
);

FILL FILL_2__348_ (
);

FILL FILL_3__463_ (
);

OAI21X1 _322_ (
    .A(_82_),
    .B(_80_),
    .C(_83_),
    .Y(_3_)
);

FILL FILL_7__394_ (
);

FILL FILL_8__336_ (
);

FILL FILL_3__519_ (
);

FILL FILL_4__306_ (
);

NAND2X1 _551_ (
    .A(Yin12b[8]),
    .B(_255_),
    .Y(_269_)
);

FILL FILL_5__513_ (
);

FILL FILL_2__386_ (
);

FILL FILL_3__328_ (
);

DFFPOSX1 _607_ (
    .D(LoadCtl[0]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[1])
);

FILL FILL_4__535_ (
);

NAND2X1 _360_ (
    .A(_111_),
    .B(_112_),
    .Y(_113_)
);

FILL FILL_5__322_ (
);

FILL FILL_8__374_ (
);

FILL FILL_0__413_ (
);

INVX1 _416_ (
    .A(Xin12b[10]),
    .Y(_162_)
);

FILL FILL_1__620_ (
);

FILL FILL_4__344_ (
);

FILL FILL_7__488_ (
);

FILL FILL_5__551_ (
);

FILL FILL_9__390_ (
);

FILL FILL_3__366_ (
);

FILL FILL_7__297_ (
);

FILL FILL_5__360_ (
);

FILL FILL_6__302_ (
);

FILL FILL_0__451_ (
);

NAND2X1 _454_ (
    .A(_186_),
    .B(_193_),
    .Y(_194_)
);

FILL FILL_4__382_ (
);

FILL FILL_5__416_ (
);

FILL FILL_8__468_ (
);

FILL FILL_6__531_ (
);

FILL FILL_2__289_ (
);

FILL FILL_0__507_ (
);

FILL FILL_4__438_ (
);

FILL FILL_2__501_ (
);

FILL FILL_8__277_ (
);

FILL FILL_6__340_ (
);

FILL FILL_0__316_ (
);

FILL FILL_9__484_ (
);

OAI21X1 _319_ (
    .A(_78_),
    .B(_80_),
    .C(_81_),
    .Y(_2_)
);

FILL FILL_1__523_ (
);

AOI21X1 _492_ (
    .A(_225_),
    .B(_224_),
    .C(_96__bF$buf0),
    .Y(_227_)
);

FILL FILL_2__310_ (
);

FILL FILL_5__454_ (
);

FILL FILL_0__545_ (
);

FILL FILL_9__293_ (
);

OAI21X1 _548_ (
    .A(_232_),
    .B(_251_),
    .C(_267_),
    .Y(_45_)
);

FILL FILL_1__332_ (
);

FILL FILL_4__476_ (
);

FILL FILL_6__625_ (
);

FILL FILL_9__349_ (
);

FILL FILL_7__412_ (
);

FILL FILL_0__354_ (
);

FILL FILL_3__498_ (
);

OAI21X1 _357_ (
    .A(_93_),
    .B(_103_),
    .C(_104_),
    .Y(_110_)
);

FILL FILL_4__285_ (
);

FILL FILL_5__319_ (
);

FILL FILL_5__492_ (
);

FILL FILL_6__434_ (
);

FILL FILL_1__617_ (
);

DFFPOSX1 _586_ (
    .D(_37_),
    .CLK(clk_bF$buf5),
    .Q(Xin12b[6])
);

FILL FILL_1__370_ (
);

FILL FILL_2__404_ (
);

FILL FILL_5__548_ (
);

FILL FILL_9__387_ (
);

FILL FILL_7__450_ (
);

FILL FILL_0__392_ (
);

FILL FILL_1__426_ (
);

OAI21X1 _395_ (
    .A(_137_),
    .B(LoadCtl_6_bF$buf3),
    .C(_143_),
    .Y(_16_)
);

FILL FILL_5__357_ (
);

FILL FILL_6__472_ (
);

FILL FILL_7__506_ (
);

FILL FILL_0__448_ (
);

FILL FILL_8__621_ (
);

FILL FILL_4__379_ (
);

FILL FILL75750x50550 (
);

FILL FILL_2__442_ (
);

FILL FILL_6__528_ (
);

FILL FILL_6__281_ (
);

FILL FILL_7__315_ (
);

FILL FILL_1__464_ (
);

FILL FILL_8__430_ (
);

FILL FILL_5__395_ (
);

FILL FILL_3__613_ (
);

FILL FILL_6__337_ (
);

FILL FILL_4__400_ (
);

FILL FILL_7__544_ (
);

FILL FILL_0__486_ (
);

INVX1 _489_ (
    .A(Yin12b[9]),
    .Y(_224_)
);

FILL FILL_1__273_ (
);

FILL FILL_2__307_ (
);

FILL FILL_2__480_ (
);

FILL FILL_3__422_ (
);

FILL FILL_7__353_ (
);

FILL FILL_0__295_ (
);

FILL FILL_1__329_ (
);

NAND2X1 _298_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[8]),
    .Y(_66_)
);

FILL FILL_2__536_ (
);

FILL FILL_6__375_ (
);

FILL FILL_7__409_ (
);

NAND3X1 _510_ (
    .A(_241_),
    .B(_242_),
    .C(_233_),
    .Y(_243_)
);

FILL FILL_8__524_ (
);

FILL FILL_2__345_ (
);

FILL FILL_9__311_ (
);

FILL FILL_5__489_ (
);

FILL FILL_3__460_ (
);

BUFX2 BUFX2_insert10 (
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(ISreg),
    .Y(ISreg_bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .A(ISreg),
    .Y(ISreg_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .A(ISreg),
    .Y(ISreg_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .A(ISreg),
    .Y(ISreg_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .A(ISreg),
    .Y(ISreg_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf4)
);

FILL FILL_7__391_ (
);

BUFX2 BUFX2_insert17 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf1)
);

FILL FILL_1__367_ (
);

FILL FILL_8__333_ (
);

FILL FILL_9__540_ (
);

FILL FILL_5__298_ (
);

FILL FILL_3__516_ (
);

FILL FILL_4__303_ (
);

FILL FILL_7__447_ (
);

FILL FILL_0__389_ (
);

FILL FILL_5__510_ (
);

FILL FILL75150x7350 (
);

FILL FILL_2__383_ (
);

FILL FILL_3__325_ (
);

FILL FILL_6__469_ (
);

DFFPOSX1 _604_ (
    .D(_6_),
    .CLK(clk_bF$buf3),
    .Q(Yin0[0])
);

FILL FILL_4__532_ (
);

FILL FILL_8__618_ (
);

FILL FILL_8__371_ (
);

FILL FILL_2__439_ (
);

FILL FILL_9__405_ (
);

FILL FILL_0__410_ (
);

FILL FILL_3__554_ (
);

FILL FILL_6__278_ (
);

NOR2X1 _413_ (
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .Y(_159_)
);

FILL FILL_4__341_ (
);

FILL FILL_7__485_ (
);

FILL FILL_8__427_ (
);

FILL FILL_3__363_ (
);

FILL FILL_7__294_ (
);

FILL FILL_2__477_ (
);

FILL FILL_9__443_ (
);

FILL FILL_3__419_ (
);

NAND3X1 _451_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_190_),
    .C(_191_),
    .Y(_192_)
);

FILL FILL_5__413_ (
);

FILL FILL_1__499_ (
);

FILL FILL_8__465_ (
);

FILL FILL_5_BUFX2_insert20 (
);

FILL FILL_5_BUFX2_insert21 (
);

FILL FILL_5_BUFX2_insert22 (
);

FILL FILL_5_BUFX2_insert23 (
);

FILL FILL_5_BUFX2_insert24 (
);

FILL FILL_5_BUFX2_insert25 (
);

FILL FILL_2__286_ (
);

FILL FILL_0__504_ (
);

NAND2X1 _507_ (
    .A(_238_),
    .B(_239_),
    .Y(_240_)
);

FILL FILL_4__435_ (
);

FILL FILL_8__274_ (
);

FILL FILL_9__308_ (
);

FILL FILL_0__313_ (
);

FILL FILL_9__481_ (
);

FILL FILL_3__457_ (
);

INVX1 _316_ (
    .A(_75_),
    .Y(_79_)
);

FILL FILL_1__520_ (
);

FILL FILL_7__388_ (
);

FILL FILL_5__451_ (
);

FILL FILL_9__537_ (
);

FILL FILL_0__542_ (
);

FILL FILL_9__290_ (
);

NAND2X1 _545_ (
    .A(LoadCtl[0]),
    .B(Xin[1]),
    .Y(_266_)
);

FILL FILL73650x72150 (
);

FILL FILL_4__473_ (
);

FILL FILL_5__507_ (
);

FILL FILL_6__622_ (
);

FILL FILL_9__346_ (
);

FILL FILL_0__351_ (
);

FILL FILL_3__495_ (
);

FILL FILL_4__529_ (
);

NAND2X1 _354_ (
    .A(_107_),
    .B(_105_),
    .Y(_108_)
);

FILL FILL_4__282_ (
);

FILL FILL_5__316_ (
);

FILL FILL_8__368_ (
);

FILL FILL_6__431_ (
);

FILL FILL_0__407_ (
);

FILL FILL_1__614_ (
);

FILL FILL_4__338_ (
);

DFFPOSX1 _583_ (
    .D(_34_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[11])
);

FILL FILL_2__401_ (
);

FILL FILL_5__545_ (
);

FILL FILL_9__384_ (
);

FILL FILL74250x10950 (
);

FILL FILL_1__423_ (
);

NAND2X1 _392_ (
    .A(ISreg_bF$buf0),
    .B(Xin12b[6]),
    .Y(_141_)
);

FILL FILL_5__354_ (
);

FILL FILL_7__503_ (
);

FILL FILL_0__445_ (
);

OAI21X1 _448_ (
    .A(_93_),
    .B(_183_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_4__376_ (
);

FILL FILL_6__525_ (
);

FILL FILL_7__312_ (
);

FILL FILL_3__398_ (
);

FILL FILL_1__461_ (
);

FILL FILL_5__392_ (
);

FILL FILL_6__334_ (
);

FILL FILL_9__478_ (
);

FILL FILL_7__541_ (
);

FILL FILL_0__483_ (
);

FILL FILL_1__517_ (
);

NAND2X1 _486_ (
    .A(_221_),
    .B(_220_),
    .Y(_222_)
);

FILL FILL_2__304_ (
);

FILL FILL_5__448_ (
);

FILL FILL_0__539_ (
);

FILL FILL_9__287_ (
);

FILL FILL_7__350_ (
);

FILL FILL_0__292_ (
);

FILL FILL_1__326_ (
);

NAND2X1 _295_ (
    .A(selXY_bF$buf2),
    .B(Xcalc[7]),
    .Y(_64_)
);

FILL FILL_2__533_ (
);

FILL FILL_6__619_ (
);

FILL FILL_6__372_ (
);

FILL FILL_7__406_ (
);

FILL FILL_0__348_ (
);

FILL FILL_1__555_ (
);

FILL FILL_8__521_ (
);

FILL FILL_4__279_ (
);

FILL FILL_2__342_ (
);

FILL FILL_5__486_ (
);

FILL FILL_6__428_ (
);

FILL FILL_1__364_ (
);

FILL FILL_8__330_ (
);

FILL FILL_5__295_ (
);

FILL FILL_3__513_ (
);

FILL FILL_4__300_ (
);

FILL FILL_7__444_ (
);

FILL FILL_0__386_ (
);

NAND3X1 _389_ (
    .A(_132_),
    .B(_129_),
    .C(_119_),
    .Y(_138_)
);

FILL FILL_2__380_ (
);

FILL FILL_3__322_ (
);

FILL FILL_6__466_ (
);

DFFPOSX1 _601_ (
    .D(_3_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[5])
);

FILL FILL_8__615_ (
);

FILL FILL_2__436_ (
);

FILL FILL_9__402_ (
);

FILL FILL_3__551_ (
);

FILL FILL_6__275_ (
);

FILL FILL_7__309_ (
);

AOI22X1 _410_ (
    .A(_152_),
    .B(_96__bF$buf3),
    .C(_155_),
    .D(_156_),
    .Y(_18_)
);

FILL FILL_7__482_ (
);

FILL FILL_1__458_ (
);

FILL FILL_8__424_ (
);

FILL FILL_5__389_ (
);

FILL FILL_3__360_ (
);

FILL FILL_7__538_ (
);

FILL FILL_7__291_ (
);

FILL FILL_2__474_ (
);

FILL FILL_9__440_ (
);

FILL FILL_3__416_ (
);

FILL FILL_4__623_ (
);

FILL FILL74850x28950 (
);

FILL FILL_7__347_ (
);

FILL FILL_0__289_ (
);

FILL FILL_5__410_ (
);

FILL FILL_1__496_ (
);

FILL FILL_8__462_ (
);

FILL FILL_2__283_ (
);

FILL FILL_0__501_ (
);

FILL FILL_6__369_ (
);

INVX1 _504_ (
    .A(Yin12b[11]),
    .Y(_237_)
);

FILL FILL_4__432_ (
);

FILL FILL_8__518_ (
);

FILL FILL_2__339_ (
);

FILL FILL_9__305_ (
);

FILL FILL_0__310_ (
);

FILL FILL_3__454_ (
);

NAND2X1 _313_ (
    .A(Yin12b[7]),
    .B(_76_),
    .Y(_77_)
);

FILL FILL_7__385_ (
);

FILL FILL_8__327_ (
);

FILL FILL_9__534_ (
);

OAI21X1 _542_ (
    .A(_257_),
    .B(_86_),
    .C(_264_),
    .Y(_42_)
);

FILL FILL_4__470_ (
);

FILL FILL_5__504_ (
);

FILL FILL_8__556_ (
);

FILL FILL_2__377_ (
);

FILL FILL_9__343_ (
);

FILL FILL_3__319_ (
);

FILL FILL_3__492_ (
);

FILL FILL_4__526_ (
);

OR2X2 _351_ (
    .A(_104_),
    .B(_103_),
    .Y(_105_)
);

FILL FILL_5__313_ (
);

FILL FILL_1__399_ (
);

FILL FILL_8__365_ (
);

FILL FILL_0__404_ (
);

FILL FILL_3__548_ (
);

OAI21X1 _407_ (
    .A(_93_),
    .B(_144_),
    .C(_147_),
    .Y(_154_)
);

FILL FILL_4__335_ (
);

FILL FILL_7__479_ (
);

DFFPOSX1 _580_ (
    .D(_31_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[10])
);

FILL FILL_5__542_ (
);

FILL FILL_9__381_ (
);

FILL FILL_3__357_ (
);

FILL FILL_1__420_ (
);

FILL FILL_7__288_ (
);

FILL FILL_5__351_ (
);

FILL FILL_9__437_ (
);

FILL FILL_7__500_ (
);

FILL FILL_0__442_ (
);

OAI21X1 _445_ (
    .A(_93_),
    .B(_186_),
    .C(_183_),
    .Y(_187_)
);

FILL FILL_4__373_ (
);

FILL FILL_5__407_ (
);

FILL FILL_8__459_ (
);

FILL FILL75150x28950 (
);

FILL FILL_6__522_ (
);

FILL FILL_3__395_ (
);

FILL FILL_4__429_ (
);

FILL FILL_6__331_ (
);

FILL FILL_0__307_ (
);

FILL FILL_9__475_ (
);

FILL FILL_0__480_ (
);

FILL FILL_1__514_ (
);

OAI21X1 _483_ (
    .A(_194_),
    .B(_218_),
    .C(ISreg_bF$buf3),
    .Y(_219_)
);

FILL FILL_2__301_ (
);

FILL FILL_5__445_ (
);

FILL FILL_8__497_ (
);

FILL FILL_0__536_ (
);

OAI21X1 _539_ (
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[0]),
    .Y(_263_)
);

FILL FILL_1__323_ (
);

FILL FILL_4__467_ (
);

NAND2X1 _292_ (
    .A(selXY_bF$buf1),
    .B(Xcalc[6]),
    .Y(_62_)
);

FILL FILL_2__530_ (
);

FILL FILL_6__616_ (
);

FILL FILL_7__403_ (
);

FILL FILL_0__345_ (
);

FILL FILL_3__489_ (
);

OAI21X1 _348_ (
    .A(_96__bF$buf4),
    .B(_101_),
    .C(_102_),
    .Y(_10_)
);

FILL FILL_1__552_ (
);

FILL FILL_4__276_ (
);

FILL FILL_5__483_ (
);

FILL FILL_6__425_ (
);

FILL FILL_3__298_ (
);

DFFPOSX1 _577_ (
    .D(_28_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[7])
);

FILL FILL_1__361_ (
);

FILL FILL_5__539_ (
);

FILL FILL_5__292_ (
);

FILL FILL_3__510_ (
);

FILL FILL_7__441_ (
);

FILL FILL_0__383_ (
);

FILL FILL_1__417_ (
);

NAND2X1 _386_ (
    .A(Xcalc[6]),
    .B(_96__bF$buf3),
    .Y(_136_)
);

FILL FILL_2__624_ (
);

FILL FILL_5__348_ (
);

FILL FILL_6__463_ (
);

FILL FILL_0__439_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_2__433_ (
);

FILL FILL_1_BUFX2_insert18 (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_6__519_ (
);

FILL FILL_7__306_ (
);

FILL FILL_1__455_ (
);

FILL FILL_8__421_ (
);

FILL FILL_5__386_ (
);

FILL FILL75450x36150 (
);

FILL FILL_6__328_ (
);

FILL FILL_7__535_ (
);

FILL FILL_0__477_ (
);

FILL FILL72750x10950 (
);

FILL FILL_2__471_ (
);

FILL FILL_3__413_ (
);

FILL FILL_4__620_ (
);

FILL FILL_7__344_ (
);

FILL FILL_0__286_ (
);

NAND2X1 _289_ (
    .A(selXY_bF$buf0),
    .B(Xcalc[5]),
    .Y(_60_)
);

FILL FILL_1__493_ (
);

FILL FILL_2__527_ (
);

FILL FILL_2__280_ (
);

FILL FILL_6__366_ (
);

NAND3X1 _501_ (
    .A(LoadCtl_6_bF$buf2),
    .B(_231_),
    .C(_234_),
    .Y(_235_)
);

FILL FILL_1__549_ (
);

FILL FILL_8__515_ (
);

FILL FILL_2__336_ (
);

FILL FILL_9__302_ (
);

FILL FILL_3__451_ (
);

INVX1 _310_ (
    .A(LoadCtl[2]),
    .Y(_74_)
);

FILL FILL_7__382_ (
);

FILL FILL_1__358_ (
);

FILL FILL_8__324_ (
);

FILL FILL_9__531_ (
);

FILL FILL_5__289_ (
);

FILL FILL_3__507_ (
);

FILL FILL_6_BUFX2_insert10 (
);

FILL FILL_6_BUFX2_insert11 (
);

FILL FILL_6_BUFX2_insert12 (
);

FILL FILL_6_BUFX2_insert13 (
);

FILL FILL_6_BUFX2_insert14 (
);

FILL FILL_6_BUFX2_insert15 (
);

FILL FILL_6_BUFX2_insert16 (
);

FILL FILL_6_BUFX2_insert17 (
);

FILL FILL_6_BUFX2_insert18 (
);

FILL FILL_6_BUFX2_insert19 (
);

FILL FILL_7__438_ (
);

FILL FILL_5__501_ (
);

FILL FILL_8__553_ (
);

FILL FILL_2__374_ (
);

FILL FILL_3__316_ (
);

FILL FILL_4__523_ (
);

FILL FILL_5__310_ (
);

FILL FILL_1__396_ (
);

FILL FILL_8__362_ (
);

FILL FILL_0__401_ (
);

FILL FILL_3__545_ (
);

OAI21X1 _404_ (
    .A(_96__bF$buf0),
    .B(_150_),
    .C(_151_),
    .Y(_17_)
);

FILL FILL_4__332_ (
);

FILL FILL_7__476_ (
);

FILL FILL_8__418_ (
);

FILL FILL_9__625_ (
);

FILL FILL_3__354_ (
);

FILL FILL_6__498_ (
);

FILL FILL_7__285_ (
);

FILL FILL_2__468_ (
);

FILL FILL_4__617_ (
);

OAI21X1 _442_ (
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf2),
    .Y(_184_)
);

FILL FILL_4__370_ (
);

FILL FILL_5__404_ (
);

FILL FILL_8__456_ (
);

FILL FILL_2__277_ (
);

FILL FILL_3__392_ (
);

FILL FILL_4__426_ (
);

FILL FILL_1__299_ (
);

FILL FILL_0__304_ (
);

FILL FILL_3__448_ (
);

NAND2X1 _307_ (
    .A(selXY_bF$buf2),
    .B(Xcalc[11]),
    .Y(_72_)
);

FILL FILL_1__511_ (
);

FILL FILL_7__379_ (
);

INVX1 _480_ (
    .A(Yin12b[8]),
    .Y(_216_)
);

FILL FILL_5__442_ (
);

FILL FILL_8__494_ (
);

FILL FILL_0__533_ (
);

FILL FILL_9__281_ (
);

OAI21X1 _536_ (
    .A(_118_),
    .B(_80_),
    .C(_261_),
    .Y(_39_)
);

FILL FILL_1__320_ (
);

FILL FILL_4__464_ (
);

FILL FILL_6__613_ (
);

FILL FILL_7__400_ (
);

FILL FILL_0__342_ (
);

FILL FILL_3__486_ (
);

OAI21X1 _345_ (
    .A(_93_),
    .B(_95_),
    .C(_99_),
    .Y(_100_)
);

FILL FILL_4__273_ (
);

FILL FILL_5__307_ (
);

FILL FILL_8__359_ (
);

FILL FILL_5__480_ (
);

FILL FILL_6__422_ (
);

FILL FILL_3__295_ (
);

FILL FILL_4__329_ (
);

DFFPOSX1 _574_ (
    .D(_25_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[4])
);

FILL FILL_5__536_ (
);

FILL FILL_9__375_ (
);

FILL FILL_0__380_ (
);

FILL FILL_1__414_ (
);

NAND2X1 _383_ (
    .A(ISreg_bF$buf0),
    .B(_130_),
    .Y(_133_)
);

FILL FILL_2__621_ (
);

FILL FILL_5__345_ (
);

FILL FILL_8__397_ (
);

FILL FILL_6__460_ (
);

FILL FILL_0__436_ (
);

NAND3X1 _439_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_180_),
    .C(_181_),
    .Y(_182_)
);

FILL FILL_4__367_ (
);

FILL FILL_2__430_ (
);

FILL FILL_6__516_ (
);

FILL FILL_7__303_ (
);

FILL FILL_3__389_ (
);

FILL FILL_1__452_ (
);

FILL FILL_5__383_ (
);

FILL FILL_6__325_ (
);

FILL FILL_9__469_ (
);

FILL FILL_7__532_ (
);

FILL FILL_0__474_ (
);

FILL FILL_5_BUFX2_insert7 (
);

FILL FILL_1__508_ (
);

FILL FILL_5_BUFX2_insert8 (
);

FILL FILL_5_BUFX2_insert9 (
);

NAND3X1 _477_ (
    .A(_212_),
    .B(_213_),
    .C(_207_),
    .Y(_214_)
);

FILL FILL75450x57750 (
);

FILL FILL_5__439_ (
);

FILL FILL_3__410_ (
);

FILL FILL_6__554_ (
);

FILL FILL_9__278_ (
);

FILL FILL74250x72150 (
);

FILL FILL74250x39750 (
);

FILL FILL_7__341_ (
);

FILL FILL_0__283_ (
);

FILL FILL_1__317_ (
);

NAND2X1 _286_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[4]),
    .Y(_58_)
);

FILL FILL_1__490_ (
);

FILL FILL_2__524_ (
);

FILL FILL_6__363_ (
);

FILL FILL_0__339_ (
);

FILL FILL_1__546_ (
);

FILL FILL_8__512_ (
);

FILL FILL_2__333_ (
);

FILL FILL_5__477_ (
);

FILL FILL_6__419_ (
);

FILL FILL_1__355_ (
);

FILL FILL_8__321_ (
);

FILL FILL_4__499_ (
);

FILL FILL_5__286_ (
);

FILL FILL_3__504_ (
);

FILL FILL75750x10950 (
);

FILL FILL_7__435_ (
);

FILL FILL_0__377_ (
);

FILL FILL_7_BUFX2_insert7 (
);

FILL FILL_7_BUFX2_insert8 (
);

FILL FILL_7_BUFX2_insert9 (
);

FILL FILL_8__550_ (
);

FILL FILL_2__618_ (
);

FILL FILL_2__371_ (
);

FILL FILL_3__313_ (
);

FILL FILL_6__457_ (
);

FILL FILL_4__520_ (
);

FILL FILL_1__393_ (
);

FILL FILL_2__427_ (
);

FILL FILL_3__542_ (
);

NAND2X1 _401_ (
    .A(_144_),
    .B(_147_),
    .Y(_149_)
);

FILL FILL_7__473_ (
);

FILL FILL_1__449_ (
);

FILL FILL_8__415_ (
);

FILL FILL_3__351_ (
);

FILL FILL_6__495_ (
);

FILL FILL_7__529_ (
);

FILL FILL_7__282_ (
);

FILL FILL_2__465_ (
);

FILL FILL_3__407_ (
);

FILL FILL_4__614_ (
);

FILL FILL_7__338_ (
);

FILL FILL_9_BUFX2_insert8 (
);

FILL FILL_9_BUFX2_insert9 (
);

FILL FILL_5__401_ (
);

FILL FILL_1__487_ (
);

FILL FILL_8__453_ (
);

FILL FILL_2__274_ (
);

FILL FILL_4__423_ (
);

FILL FILL_8__509_ (
);

FILL FILL_1__296_ (
);

FILL FILL_0__301_ (
);

FILL FILL_3__445_ (
);

NAND2X1 _304_ (
    .A(selXY_bF$buf2),
    .B(Xcalc[10]),
    .Y(_70_)
);

FILL FILL_7__376_ (
);

FILL FILL_8__318_ (
);

FILL FILL_8__491_ (
);

FILL FILL_9__525_ (
);

FILL FILL_0__530_ (
);

FILL FILL_6__398_ (
);

NAND2X1 _533_ (
    .A(Xin12b[7]),
    .B(_76_),
    .Y(_260_)
);

FILL FILL_4__461_ (
);

FILL FILL_8__547_ (
);

FILL FILL_2__368_ (
);

FILL FILL_9__334_ (
);

FILL FILL_3__483_ (
);

FILL FILL_4__517_ (
);

OAI21X1 _342_ (
    .A(_95_),
    .B(_96__bF$buf2),
    .C(_97_),
    .Y(_9_)
);

FILL FILL_5__304_ (
);

FILL FILL_8__356_ (
);

FILL FILL_3__539_ (
);

FILL FILL_3__292_ (
);

FILL FILL_4__326_ (
);

DFFPOSX1 _571_ (
    .D(_22_),
    .CLK(clk_bF$buf3),
    .Q(Ycalc[1])
);

FILL FILL_5__533_ (
);

FILL FILL_9__619_ (
);

FILL FILL_0__624_ (
);

FILL FILL_9__372_ (
);

FILL FILL_3__348_ (
);

FILL FILL_1__411_ (
);

FILL FILL_4__555_ (
);

FILL FILL_7__279_ (
);

NAND2X1 _380_ (
    .A(_129_),
    .B(_119_),
    .Y(_130_)
);

FILL FILL_5__342_ (
);

FILL FILL_8__394_ (
);

FILL FILL_9__428_ (
);

FILL FILL_0__433_ (
);

OAI21X1 _436_ (
    .A(LoadCtl_6_bF$buf4),
    .B(_49_),
    .C(_179_),
    .Y(_21_)
);

FILL FILL_4__364_ (
);

FILL FILL_6__513_ (
);

FILL FILL_7__300_ (
);

FILL FILL_3__386_ (
);

FILL FILL_5__380_ (
);

FILL FILL_6__322_ (
);

FILL FILL_9__466_ (
);

FILL FILL_0__471_ (
);

FILL FILL_1__505_ (
);

NAND3X1 _474_ (
    .A(ISreg_bF$buf4),
    .B(Yin12b[7]),
    .C(_210_),
    .Y(_211_)
);

FILL FILL_5__436_ (
);

FILL FILL_8__488_ (
);

FILL FILL_6__551_ (
);

FILL FILL_0__527_ (
);

FILL FILL_9__275_ (
);

FILL FILL_0__280_ (
);

FILL FILL_1__314_ (
);

FILL FILL_4__458_ (
);

NAND2X1 _283_ (
    .A(selXY_bF$buf0),
    .B(Xcalc[3]),
    .Y(_56_)
);

FILL FILL_2__521_ (
);

FILL FILL_8__297_ (
);

FILL FILL_6__360_ (
);

FILL FILL_0__336_ (
);

INVX1 _339_ (
    .A(Xin0[0]),
    .Y(_95_)
);

FILL FILL_1__543_ (
);

FILL FILL_2__330_ (
);

FILL FILL_5__474_ (
);

FILL FILL_6__416_ (
);

FILL FILL_7__623_ (
);

FILL FILL_3__289_ (
);

DFFPOSX1 _568_ (
    .D(_19_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[10])
);

FILL FILL_1__352_ (
);

FILL FILL_4__496_ (
);

FILL FILL_5__283_ (
);

FILL FILL_3__501_ (
);

FILL FILL_9__369_ (
);

FILL FILL_7__432_ (
);

FILL FILL_0__374_ (
);

FILL FILL_1__408_ (
);

NAND2X1 _377_ (
    .A(Xcalc[5]),
    .B(_96__bF$buf2),
    .Y(_128_)
);

FILL FILL_2__615_ (
);

FILL FILL_5__339_ (
);

FILL FILL_3__310_ (
);

FILL FILL_6__454_ (
);

FILL FILL_1__390_ (
);

FILL FILL_2__424_ (
);

FILL FILL_7__470_ (
);

FILL FILL_1__446_ (
);

FILL FILL_8__412_ (
);

FILL FILL_5__377_ (
);

FILL FILL_6__319_ (
);

FILL FILL74250x25350 (
);

FILL FILL_6__492_ (
);

FILL FILL_7__526_ (
);

FILL FILL_0__468_ (
);

FILL FILL_4__399_ (
);

FILL FILL_2__462_ (
);

FILL FILL_3__404_ (
);

FILL FILL_6__548_ (
);

FILL FILL_7__335_ (
);

FILL FILL_0__277_ (
);

FILL FILL_1__484_ (
);

FILL FILL_8__450_ (
);

FILL FILL_2__518_ (
);

FILL FILL_6__357_ (
);

FILL FILL_4__420_ (
);

FILL FILL_8__506_ (
);

FILL FILL_7_BUFX2_insert20 (
);

FILL FILL_7_BUFX2_insert21 (
);

FILL FILL_7_BUFX2_insert22 (
);

FILL FILL_7_BUFX2_insert23 (
);

FILL FILL_7_BUFX2_insert24 (
);

FILL FILL_7_BUFX2_insert25 (
);

FILL FILL_1__293_ (
);

FILL FILL_2__327_ (
);

FILL FILL_3__442_ (
);

NAND2X1 _301_ (
    .A(selXY_bF$buf0),
    .B(Xcalc[9]),
    .Y(_68_)
);

FILL FILL_7__373_ (
);

FILL FILL_1__349_ (
);

FILL FILL_8__315_ (
);

FILL FILL_2__556_ (
);

FILL FILL_9__522_ (
);

FILL FILL_6__395_ (
);

FILL FILL_7__429_ (
);

OAI21X1 _530_ (
    .A(_257_),
    .B(_255_),
    .C(_258_),
    .Y(_36_)
);

FILL FILL_8__544_ (
);

FILL FILL72750x72150 (
);

FILL FILL_2__365_ (
);

FILL FILL_9__331_ (
);

FILL FILL_3__307_ (
);

FILL FILL_3__480_ (
);

FILL FILL_4__514_ (
);

FILL FILL_5__301_ (
);

FILL FILL_1__387_ (
);

FILL FILL_8__353_ (
);

FILL FILL_3__536_ (
);

FILL FILL_4__323_ (
);

FILL FILL_7__467_ (
);

FILL FILL_8__409_ (
);

FILL FILL_5__530_ (
);

FILL FILL_9__616_ (
);

FILL FILL_0__621_ (
);

FILL FILL_3__345_ (
);

FILL FILL_6__489_ (
);

BUFX2 _624_ (
    .A(_272_[9]),
    .Y(Dout[9])
);

FILL FILL73350x10950 (
);

FILL FILL_4__552_ (
);

FILL FILL_7__276_ (
);

FILL FILL75750x18150 (
);

FILL FILL_8__391_ (
);

FILL FILL_2__459_ (
);

FILL FILL_9__425_ (
);

FILL FILL_0__430_ (
);

FILL FILL_6__298_ (
);

NAND3X1 _433_ (
    .A(LoadCtl_6_bF$buf3),
    .B(_177_),
    .C(_174_),
    .Y(_178_)
);

FILL FILL_4__361_ (
);

FILL FILL_8__447_ (
);

FILL FILL_6__510_ (
);

FILL FILL_3__383_ (
);

FILL FILL_4__417_ (
);

FILL FILL_5__624_ (
);

FILL FILL_2__497_ (
);

FILL FILL_9__463_ (
);

FILL FILL_3__439_ (
);

FILL FILL_1__502_ (
);

NAND3X1 _471_ (
    .A(LoadCtl_6_bF$buf1),
    .B(_205_),
    .C(_208_),
    .Y(_209_)
);

FILL FILL_5__433_ (
);

FILL FILL_8__485_ (
);

FILL FILL_9__519_ (
);

FILL FILL_0__524_ (
);

OAI21X1 _527_ (
    .A(_254_),
    .B(_255_),
    .C(_256_),
    .Y(_35_)
);

FILL FILL_1__311_ (
);

FILL FILL_4__455_ (
);

NAND2X1 _280_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[2]),
    .Y(_54_)
);

FILL FILL_8__294_ (
);

FILL FILL_9__328_ (
);

FILL FILL_0__333_ (
);

FILL FILL_3__477_ (
);

INVX4 _336_ (
    .A(ISreg_bF$buf4),
    .Y(_93_)
);

FILL FILL_1__540_ (
);

FILL FILL_5__471_ (
);

FILL FILL_6__413_ (
);

FILL FILL_7__620_ (
);

FILL FILL_3__286_ (
);

DFFPOSX1 _565_ (
    .D(_16_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[7])
);

FILL FILL_4__493_ (
);

FILL FILL_5__527_ (
);

FILL FILL_5__280_ (
);

FILL FILL_0__618_ (
);

FILL FILL_9__366_ (
);

FILL FILL_0__371_ (
);

FILL FILL_1__405_ (
);

FILL FILL_4__549_ (
);

OR2X2 _374_ (
    .A(_124_),
    .B(_123_),
    .Y(_125_)
);

FILL FILL_5__336_ (
);

FILL FILL_8__388_ (
);

FILL FILL_6__451_ (
);

FILL FILL_0__427_ (
);

FILL FILL_4__358_ (
);

FILL FILL_2__421_ (
);

FILL FILL_6__507_ (
);

FILL FILL_1__443_ (
);

FILL FILL_5__374_ (
);

FILL FILL_6__316_ (
);

FILL FILL_7__523_ (
);

FILL FILL_0__465_ (
);

INVX1 _468_ (
    .A(Yin12b[6]),
    .Y(_206_)
);

FILL FILL_4__396_ (
);

FILL FILL_3__401_ (
);

FILL FILL_6__545_ (
);

FILL FILL_7__332_ (
);

FILL FILL_0__274_ (
);

FILL FILL_1__308_ (
);

NAND2X1 _277_ (
    .A(selXY_bF$buf3),
    .B(Xcalc[1]),
    .Y(_52_)
);

FILL FILL73950x28950 (
);

FILL FILL_1__481_ (
);

FILL FILL_2__515_ (
);

FILL FILL_6__354_ (
);

FILL FILL_1__537_ (
);

FILL FILL_8__503_ (
);

FILL FILL_1__290_ (
);

FILL FILL_2__324_ (
);

FILL FILL_5__468_ (
);

FILL FILL_7__617_ (
);

FILL FILL_7__370_ (
);

FILL FILL_1__346_ (
);

FILL FILL_8__312_ (
);

FILL FILL_2__553_ (
);

FILL FILL_5__277_ (
);

FILL FILL_6__392_ (
);

FILL FILL_7__426_ (
);

FILL FILL_0__368_ (
);

FILL FILL_8__541_ (
);

FILL FILL_4__299_ (
);

FILL FILL_2__362_ (
);

FILL FILL_3__304_ (
);

FILL FILL_6__448_ (
);

FILL FILL_4__511_ (
);

FILL FILL_1__384_ (
);

FILL FILL_8__350_ (
);

FILL FILL_2__418_ (
);

FILL FILL_3__533_ (
);

FILL FILL_4__320_ (
);

FILL FILL_7__464_ (
);

FILL FILL_8__406_ (
);

FILL FILL_9__613_ (
);

FILL FILL_3__342_ (
);

FILL FILL_6__486_ (
);

BUFX2 _621_ (
    .A(_272_[6]),
    .Y(Dout[6])
);

FILL FILL_7__273_ (
);

FILL FILL_2__456_ (
);

FILL FILL_9__422_ (
);

FILL FILL75750x72150 (
);

FILL FILL75750x39750 (
);

FILL FILL_6__295_ (
);

FILL FILL_7__329_ (
);

OAI21X1 _430_ (
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .C(ISreg_bF$buf0),
    .Y(_175_)
);

FILL FILL_1__478_ (
);

FILL FILL_8__444_ (
);

FILL FILL_3__380_ (
);

FILL FILL_4__414_ (
);

FILL FILL_5__621_ (
);

FILL FILL_1__287_ (
);

FILL FILL_2__494_ (
);

FILL FILL_9__460_ (
);

FILL FILL_3__436_ (
);

FILL FILL_7__367_ (
);

FILL FILL_8__309_ (
);

FILL FILL_5__430_ (
);

FILL FILL_8__482_ (
);

FILL FILL_9__516_ (
);

FILL FILL_0__521_ (
);

FILL FILL_6__389_ (
);

INVX1 _524_ (
    .A(Xin[0]),
    .Y(_254_)
);

FILL FILL_4__452_ (
);

FILL FILL_8__538_ (
);

FILL FILL_8__291_ (
);

FILL FILL_2__359_ (
);

FILL FILL_0__330_ (
);

FILL FILL_3__474_ (
);

FILL FILL_4__508_ (
);

INVX1 _333_ (
    .A(Yin0[1]),
    .Y(_91_)
);

FILL FILL_8__347_ (
);

FILL FILL_6__410_ (
);

FILL FILL_3__283_ (
);

FILL FILL_4__317_ (
);

DFFPOSX1 _562_ (
    .D(_13_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[4])
);

FILL FILL_4__490_ (
);

FILL FILL_5__524_ (
);

FILL FILL_2__397_ (
);

FILL FILL_0__615_ (
);

FILL FILL_3__339_ (
);

BUFX2 _618_ (
    .A(_272_[3]),
    .Y(Dout[3])
);

FILL FILL_1__402_ (
);

FILL FILL_4__546_ (
);

OAI21X1 _371_ (
    .A(_96__bF$buf4),
    .B(_121_),
    .C(_122_),
    .Y(_13_)
);

FILL FILL_5__333_ (
);

FILL FILL_8__385_ (
);

FILL FILL_0__424_ (
);

INVX1 _427_ (
    .A(_171_),
    .Y(_172_)
);

FILL FILL_4__355_ (
);

FILL FILL_7__499_ (
);

FILL FILL_6__504_ (
);

FILL FILL_3__377_ (
);

FILL FILL_1__440_ (
);

FILL FILL_5__618_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_3_BUFX2_insert11 (
);

FILL FILL_3_BUFX2_insert12 (
);

FILL FILL_3_BUFX2_insert13 (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert15 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_3_BUFX2_insert18 (
);

FILL FILL_3_BUFX2_insert19 (
);

FILL FILL_5__371_ (
);

FILL FILL_6__313_ (
);

FILL FILL_7__520_ (
);

FILL FILL_0__462_ (
);

NOR2X1 _465_ (
    .A(Yin12b[4]),
    .B(Yin12b[5]),
    .Y(_203_)
);

FILL FILL_4__393_ (
);

FILL FILL_5__427_ (
);

FILL FILL_8__479_ (
);

FILL FILL_6__542_ (
);

FILL FILL_0__518_ (
);

FILL FILL_1__305_ (
);

FILL FILL_4__449_ (
);

NAND2X1 _274_ (
    .A(Xcalc[0]),
    .B(selXY_bF$buf0),
    .Y(_50_)
);

FILL FILL_2__512_ (
);

FILL FILL_8__288_ (
);

FILL FILL_6__351_ (
);

FILL FILL_0__327_ (
);

FILL FILL_9__495_ (
);

FILL FILL_1__534_ (
);

FILL FILL_8__500_ (
);

FILL FILL_2__321_ (
);

FILL FILL_5__465_ (
);

FILL FILL_6__407_ (
);

FILL FILL_7__614_ (
);

FILL FILL_0__556_ (
);

DFFPOSX1 _559_ (
    .D(_10_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[1])
);

FILL FILL_1__343_ (
);

FILL FILL_4__487_ (
);

FILL FILL_2__550_ (
);

FILL FILL_5__274_ (
);

FILL FILL_7__423_ (
);

FILL FILL_0__365_ (
);

OAI21X1 _368_ (
    .A(_93_),
    .B(_119_),
    .C(_118_),
    .Y(_120_)
);

FILL FILL_4__296_ (
);

FILL FILL_3__301_ (
);

FILL FILL_6__445_ (
);

FILL FILL_8_BUFX2_insert10 (
);

FILL FILL_8_BUFX2_insert11 (
);

FILL FILL_8_BUFX2_insert12 (
);

FILL FILL_8_BUFX2_insert13 (
);

FILL FILL_8_BUFX2_insert14 (
);

FILL FILL_8_BUFX2_insert15 (
);

FILL FILL_8_BUFX2_insert16 (
);

FILL FILL_8_BUFX2_insert17 (
);

FILL FILL_8_BUFX2_insert18 (
);

FILL FILL_8_BUFX2_insert19 (
);

DFFPOSX1 _597_ (
    .D(_48_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[9])
);

FILL FILL75450x50550 (
);

FILL FILL_1__381_ (
);

FILL FILL_2__415_ (
);

FILL FILL_3__530_ (
);

FILL FILL_9__398_ (
);

FILL FILL_7__461_ (
);

FILL FILL_1__437_ (
);

FILL FILL_8__403_ (
);

FILL FILL_5__368_ (
);

FILL FILL_6__483_ (
);

FILL FILL_7__517_ (
);

FILL FILL_0__459_ (
);

FILL FILL_2__453_ (
);

FILL FILL_6__539_ (
);

FILL FILL_6__292_ (
);

FILL FILL_7__326_ (
);

FILL FILL_1__475_ (
);

FILL FILL_8__441_ (
);

FILL FILL_2__509_ (
);

FILL FILL_3__624_ (
);

FILL FILL_6__348_ (
);

FILL FILL_4__411_ (
);

FILL FILL_7__555_ (
);

FILL FILL_0__497_ (
);

FILL FILL_1__284_ (
);

FILL FILL_2__318_ (
);

FILL FILL_2__491_ (
);

FILL FILL_3__433_ (
);

FILL FILL_7__364_ (
);

FILL FILL_8__306_ (
);

FILL FILL_2__547_ (
);

FILL FILL_6__386_ (
);

OAI21X1 _521_ (
    .A(_162_),
    .B(_251_),
    .C(_252_),
    .Y(_33_)
);

FILL FILL_8__535_ (
);

FILL FILL_2__356_ (
);

FILL FILL_3__471_ (
);

FILL FILL_4__505_ (
);

INVX1 _330_ (
    .A(Yin0[0]),
    .Y(_89_)
);

FILL FILL_1__378_ (
);

FILL FILL_8__344_ (
);

FILL FILL_3__527_ (
);

FILL FILL_3__280_ (
);

FILL FILL_4__314_ (
);

FILL FILL_7__458_ (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_5__521_ (
);

FILL FILL75750x25350 (
);

FILL FILL_2__394_ (
);

FILL FILL_9__360_ (
);

FILL FILL_3__336_ (
);

BUFX2 _615_ (
    .A(_272_[10]),
    .Y(Dout[10])
);

FILL FILL_4__543_ (
);

FILL FILL_5__330_ (
);

FILL FILL_8__382_ (
);

FILL FILL_0__421_ (
);

FILL FILL_6__289_ (
);

INVX1 _424_ (
    .A(selSign),
    .Y(_169_)
);

FILL FILL_4__352_ (
);

FILL FILL_7__496_ (
);

FILL FILL_8__438_ (
);

FILL FILL_6__501_ (
);

FILL FILL_3__374_ (
);

FILL FILL_4__408_ (
);

FILL FILL_5__615_ (
);

FILL FILL_6__310_ (
);

FILL FILL_2__488_ (
);

FILL FILL_9__454_ (
);

OR2X2 _462_ (
    .A(_200_),
    .B(_82_),
    .Y(_201_)
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_4__390_ (
);

FILL FILL_2_BUFX2_insert9 (
);

FILL FILL_5__424_ (
);

FILL FILL_8__476_ (
);

FILL FILL_2__297_ (
);

FILL FILL_0__515_ (
);

NAND2X1 _518_ (
    .A(LoadCtl[5]),
    .B(_249_),
    .Y(_250_)
);

FILL FILL73350x72150 (
);

FILL FILL_1__302_ (
);

FILL FILL_4__446_ (
);

FILL FILL_8__285_ (
);

FILL FILL_9__319_ (
);

FILL FILL_0__324_ (
);

FILL FILL_9__492_ (
);

FILL FILL_3__468_ (
);

OAI21X1 _327_ (
    .A(_84_),
    .B(_86_),
    .C(_87_),
    .Y(_4_)
);

FILL FILL_1__531_ (
);

FILL FILL_7__399_ (
);

FILL FILL_5__462_ (
);

FILL FILL_6__404_ (
);

FILL FILL_9__548_ (
);

FILL FILL_0__553_ (
);

FILL FILL_3__277_ (
);

OAI21X1 _556_ (
    .A(_84_),
    .B(_76_),
    .C(_271_),
    .Y(_0_)
);

FILL FILL_1__340_ (
);

FILL FILL_4__484_ (
);

FILL FILL_5__518_ (
);

FILL FILL_9__357_ (
);

FILL FILL_7__420_ (
);

FILL FILL_0__362_ (
);

NAND3X1 _365_ (
    .A(ISreg_bF$buf1),
    .B(Xin12b[4]),
    .C(_116_),
    .Y(_117_)
);

FILL FILL_4__293_ (
);

FILL FILL_5__327_ (
);

FILL FILL_8__379_ (
);

FILL FILL_4_BUFX2_insert7 (
);

FILL FILL_4_BUFX2_insert8 (
);

FILL FILL_4_BUFX2_insert9 (
);

FILL FILL_6__442_ (
);

FILL FILL_0__418_ (
);

FILL FILL_1__625_ (
);

FILL FILL_4__349_ (
);

DFFPOSX1 _594_ (
    .D(_45_),
    .CLK(clk_bF$buf3),
    .Q(Yin12b[10])
);

FILL FILL_2__412_ (
);

FILL FILL_5__556_ (
);

FILL FILL_9__395_ (
);

FILL FILL_1__434_ (
);

FILL FILL_8__400_ (
);

FILL FILL_5__365_ (
);

FILL FILL_6__307_ (
);

FILL FILL_6__480_ (
);

FILL FILL_7__514_ (
);

FILL FILL_0__456_ (
);

NAND3X1 _459_ (
    .A(LoadCtl_6_bF$buf0),
    .B(_198_),
    .C(_196_),
    .Y(_199_)
);

FILL FILL_4__387_ (
);

FILL FILL_2__450_ (
);

FILL FILL_6__536_ (
);

FILL FILL_7__323_ (
);

FILL FILL_1__472_ (
);

FILL FILL_2__506_ (
);

FILL FILL_6_BUFX2_insert7 (
);

FILL FILL_6_BUFX2_insert8 (
);

FILL FILL_6_BUFX2_insert9 (
);

FILL FILL_3__621_ (
);

FILL FILL_6__345_ (
);

FILL FILL_9__489_ (
);

FILL FILL_7__552_ (
);

FILL FILL_0__494_ (
);

FILL FILL_1__528_ (
);

NAND3X1 _497_ (
    .A(ISreg_bF$buf3),
    .B(Yin12b[10]),
    .C(_230_),
    .Y(_231_)
);

FILL FILL_1__281_ (
);

FILL FILL_2__315_ (
);

FILL FILL_5__459_ (
);

FILL FILL_3__430_ (
);

FILL FILL_9__298_ (
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert6 (
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_7__361_ (
);

FILL FILL_1__337_ (
);

FILL FILL_8__303_ (
);

FILL FILL_2__544_ (
);

FILL FILL_9__510_ (
);

FILL FILL_6__383_ (
);

FILL FILL_7__417_ (
);

FILL FILL_0__359_ (
);

FILL FILL_8__532_ (
);

FILL FILL_2__353_ (
);

FILL FILL_5__497_ (
);

FILL FILL_6__439_ (
);

FILL FILL_4__502_ (
);

FILL FILL_1__375_ (
);

FILL FILL_8__341_ (
);

FILL FILL_2__409_ (
);

FILL FILL_3__524_ (
);

FILL FILL_4__311_ (
);

FILL FILL_7__455_ (
);

FILL FILL_0__397_ (
);

FILL FILL_2__391_ (
);

FILL FILL_3__333_ (
);

FILL FILL_6__477_ (
);

DFFPOSX1 _612_ (
    .D(LoadCtl[5]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[6])
);

FILL FILL_4__540_ (
);

FILL FILL75750x46950 (
);

FILL FILL_2__447_ (
);

FILL FILL_9__413_ (
);

FILL FILL_6__286_ (
);

NAND2X1 _421_ (
    .A(Xcalc[11]),
    .B(_96__bF$buf4),
    .Y(_166_)
);

FILL FILL74550x28950 (
);

FILL FILL_7__493_ (
);

FILL FILL_1__469_ (
);

FILL FILL_8__435_ (
);

FILL FILL_3__618_ (
);

FILL FILL_3__371_ (
);

FILL FILL_4__405_ (
);

FILL FILL_7__549_ (
);

FILL FILL_1__278_ (
);

FILL FILL_2__485_ (
);

FILL FILL_9__451_ (
);

FILL FILL_3__427_ (
);

FILL FILL_7__358_ (
);

FILL FILL_5__421_ (
);

FILL FILL_8__473_ (
);

FILL FILL_9__507_ (
);

FILL FILL_2__294_ (
);

FILL FILL_0__512_ (
);

NAND2X1 _515_ (
    .A(_236_),
    .B(_247_),
    .Y(_32_)
);

FILL FILL_4__443_ (
);

FILL FILL_8__529_ (
);

FILL FILL_8__282_ (
);

FILL FILL_9__316_ (
);

FILL FILL_0__321_ (
);

FILL FILL_3__465_ (
);

INVX2 _324_ (
    .A(LoadCtl[1]),
    .Y(_85_)
);

FILL FILL_7__396_ (
);

FILL FILL_8__338_ (
);

FILL FILL_6__401_ (
);

FILL FILL_9__545_ (
);

FILL FILL_0__550_ (
);

FILL FILL_3__274_ (
);

FILL FILL_4__308_ (
);

NAND2X1 _553_ (
    .A(Yin12b[9]),
    .B(_255_),
    .Y(_270_)
);

FILL FILL_4__481_ (
);

FILL FILL_5__515_ (
);

FILL FILL_2__388_ (
);

FILL FILL_9__354_ (
);

DFFPOSX1 _609_ (
    .D(LoadCtl[2]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[3])
);

FILL FILL_4__537_ (
);

OAI21X1 _362_ (
    .A(_96__bF$buf3),
    .B(_113_),
    .C(_114_),
    .Y(_12_)
);

FILL FILL_4__290_ (
);

FILL FILL_5__324_ (
);

FILL FILL_8__376_ (
);

FILL FILL_0__415_ (
);

NAND2X1 _418_ (
    .A(_162_),
    .B(_163_),
    .Y(_164_)
);

FILL FILL_1__622_ (
);

FILL FILL_4__346_ (
);

DFFPOSX1 _591_ (
    .D(_42_),
    .CLK(clk_bF$buf5),
    .Q(Xin1[1])
);

FILL FILL_5__553_ (
);

FILL FILL_9__392_ (
);

FILL FILL_3__368_ (
);

FILL FILL74850x36150 (
);

FILL FILL_1__431_ (
);

FILL FILL_7__299_ (
);

FILL FILL_5__362_ (
);

FILL FILL_6__304_ (
);

FILL FILL_9__448_ (
);

FILL FILL_7__511_ (
);

FILL FILL_0__453_ (
);

OR2X2 _456_ (
    .A(_195_),
    .B(_78_),
    .Y(_196_)
);

FILL FILL_4__384_ (
);

FILL FILL_5__418_ (
);

FILL FILL_6__533_ (
);

FILL FILL_0__509_ (
);

FILL FILL_7__320_ (
);

FILL FILL_2__503_ (
);

FILL FILL_8__279_ (
);

FILL FILL_6__342_ (
);

FILL FILL_0__318_ (
);

FILL FILL_9__486_ (
);

FILL FILL_0__491_ (
);

FILL FILL_1__525_ (
);

AND2X2 _494_ (
    .A(_203_),
    .B(_217_),
    .Y(_228_)
);

FILL FILL_2__312_ (
);

FILL FILL_5__456_ (
);

FILL FILL_0__547_ (
);

FILL FILL_1__334_ (
);

FILL FILL_8__300_ (
);

FILL FILL_4__478_ (
);

FILL FILL_9_BUFX2_insert20 (
);

FILL FILL_9_BUFX2_insert21 (
);

FILL FILL_9_BUFX2_insert23 (
);

FILL FILL_9_BUFX2_insert24 (
);

FILL FILL_9_BUFX2_insert25 (
);

FILL FILL_2__541_ (
);

FILL FILL_6__380_ (
);

FILL FILL_7__414_ (
);

FILL FILL_0__356_ (
);

OR2X2 _359_ (
    .A(_110_),
    .B(Xin1[1]),
    .Y(_112_)
);

FILL FILL_4__287_ (
);

endmodule
