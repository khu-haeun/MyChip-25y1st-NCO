/* Verilog module written by vlog2Verilog (qflow) */

module phase_accumulator(
    output [1:0] Aout,
    input En,
    input [19:0] FCW,
    output ISout,
    output Vld,
    input clk
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _73__bF$buf0 ;
wire _73__bF$buf1 ;
wire _73__bF$buf2 ;
wire _73__bF$buf3 ;
wire _73__bF$buf4 ;
wire _218_ ;
wire _256_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _197_ ;
wire _7_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire ISout ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire [11:0] Atmp ;
wire _309_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _288_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire [19:0] acc_reg ;
wire _212_ ;
wire _250_ ;
wire _306_ ;
wire En_bF$buf0 ;
wire En_bF$buf1 ;
wire En_bF$buf2 ;
wire En_bF$buf3 ;
wire En_bF$buf4 ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire _282_ ;
wire _147_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _273_ ;
wire _138_ ;
wire _30_ ;
wire En ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _264_ ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _299_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _255_ ;
wire _293_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire [1:0] _311_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire _214_ ;
wire _252_ ;
wire _308_ ;
wire _117_ ;
wire _290_ ;
wire _155_ ;
wire [1:0] Aout ;
wire _193_ ;
wire _249_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire _305_ ;
wire _114_ ;
wire [19:0] FCW ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _284_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire RdyCtl_6_bF$buf0 ;
wire RdyCtl_6_bF$buf1 ;
wire RdyCtl_6_bF$buf2 ;
wire RdyCtl_6_bF$buf3 ;
wire RdyCtl_6_bF$buf4 ;
wire _281_ ;
wire _146_ ;
wire _184_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _275_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire [6:0] RdyCtl ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _298_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _157_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _310_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _307_ ;
wire _116_ ;
wire _154_ ;
wire _192_ ;
wire _248_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _245_ ;
wire _283_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _301_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _280_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

FILL FILL_2__350_ (
);

FILL FILL_5__494_ (
);

FILL FILL_6__436_ (
);

FILL FILL_0__585_ (
);

FILL FILL_1__619_ (
);

NOR2X1 _588_ (
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_118_)
);

FILL FILL_1__372_ (
);

FILL FILL_2__406_ (
);

FILL FILL_3__521_ (
);

FILL FILL_6__665_ (
);

FILL FILL_7__452_ (
);

FILL FILL_0__394_ (
);

FILL FILL_1__428_ (
);

INVX1 _397_ (
    .A(_229_),
    .Y(_230_)
);

FILL FILL_5__359_ (
);

FILL FILL75150x36150 (
);

FILL FILL_3__330_ (
);

FILL FILL_6__474_ (
);

FILL FILL_7__508_ (
);

FILL FILL_8__623_ (
);

FILL FILL_2__444_ (
);

FILL FILL_5__588_ (
);

FILL FILL_7__317_ (
);

FILL FILL_7__490_ (
);

FILL FILL_1__466_ (
);

FILL FILL_5__397_ (
);

FILL FILL_3__615_ (
);

FILL FILL_6__339_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_4__402_ (
);

FILL FILL_7__546_ (
);

FILL FILL_0__488_ (
);

FILL FILL_2__482_ (
);

FILL FILL_3__424_ (
);

FILL FILL_6__568_ (
);

FILL FILL_7__355_ (
);

FILL FILL_2__538_ (
);

FILL FILL_6__377_ (
);

INVX1 _512_ (
    .A(Atmp[9]),
    .Y(_56_)
);

FILL FILL_4__440_ (
);

FILL FILL_7__584_ (
);

FILL FILL_2__347_ (
);

FILL FILL_3__462_ (
);

NAND2X1 _321_ (
    .A(_159_),
    .B(_156_),
    .Y(_161_)
);

FILL FILL76050x50550 (
);

FILL FILL_7__393_ (
);

FILL FILL_1__369_ (
);

FILL FILL_8__335_ (
);

FILL FILL_2__576_ (
);

FILL FILL_3__518_ (
);

FILL FILL_7__449_ (
);

NOR2X1 _550_ (
    .A(_78_),
    .B(_83_),
    .Y(_84_)
);

FILL FILL_5__512_ (
);

FILL FILL_1__598_ (
);

FILL FILL74550x14550 (
);

FILL FILL_2__385_ (
);

FILL FILL_0__603_ (
);

FILL FILL_3__327_ (
);

OAI21X1 _606_ (
    .A(_133_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

FILL FILL_4__534_ (
);

FILL FILL_5__321_ (
);

FILL FILL_8__373_ (
);

FILL FILL_0__412_ (
);

FILL FILL_3__556_ (
);

NAND2X1 _415_ (
    .A(_246_),
    .B(_245_),
    .Y(_247_)
);

FILL FILL_4__343_ (
);

FILL FILL_7__487_ (
);

FILL FILL_8__429_ (
);

FILL FILL_5__550_ (
);

FILL FILL_3__365_ (
);

DFFPOSX1 _644_ (
    .D(_18_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[11])
);

FILL FILL_4__572_ (
);

FILL FILL_5__606_ (
);

FILL FILL_2__479_ (
);

FILL FILL74850x57750 (
);

FILL FILL_0__450_ (
);

FILL FILL_3__594_ (
);

OAI21X1 _453_ (
    .A(_276_),
    .B(_277_),
    .C(_282_),
    .Y(_283_)
);

FILL FILL_4__381_ (
);

FILL FILL_5__415_ (
);

FILL FILL_8__467_ (
);

FILL FILL_6__530_ (
);

FILL FILL_0__506_ (
);

NAND2X1 _509_ (
    .A(Atmp[0]),
    .B(RdyCtl[0]),
    .Y(_54_)
);

FILL FILL_4__437_ (
);

FILL FILL_2__500_ (
);

FILL FILL_0__315_ (
);

FILL FILL_3__459_ (
);

OR2X2 _318_ (
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_158_)
);

FILL FILL_1__522_ (
);

FILL FILL_4__666_ (
);

NOR2X1 _491_ (
    .A(Atmp[11]),
    .B(RdyCtl_6_bF$buf2),
    .Y(_309_)
);

FILL FILL_5__453_ (
);

FILL FILL_7__602_ (
);

FILL FILL_0__544_ (
);

NOR2X1 _547_ (
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_81_)
);

FILL FILL_1__331_ (
);

FILL FILL_4__475_ (
);

FILL FILL_5__509_ (
);

FILL FILL_6__624_ (
);

FILL FILL_7__411_ (
);

FILL FILL_0__353_ (
);

FILL FILL_3__497_ (
);

AOI21X1 _356_ (
    .A(_187_),
    .B(_191_),
    .C(_73__bF$buf2),
    .Y(_193_)
);

FILL FILL_1__560_ (
);

FILL FILL_5__318_ (
);

FILL FILL_5__491_ (
);

FILL FILL_6__433_ (
);

FILL FILL_0__409_ (
);

FILL FILL_0__582_ (
);

FILL FILL_1__616_ (
);

AOI21X1 _585_ (
    .A(_114_),
    .B(RdyCtl_6_bF$buf4),
    .C(_115_),
    .Y(_11_)
);

FILL FILL_2__403_ (
);

FILL FILL_5__547_ (
);

FILL FILL_8__599_ (
);

FILL FILL_0__391_ (
);

FILL FILL_1__425_ (
);

FILL FILL_4__569_ (
);

AOI21X1 _394_ (
    .A(_226_),
    .B(RdyCtl_6_bF$buf1),
    .C(_227_),
    .Y(_21_)
);

FILL FILL_5__356_ (
);

FILL FILL_6__471_ (
);

FILL FILL_7__505_ (
);

FILL FILL_0__447_ (
);

FILL FILL75150x57750 (
);

FILL FILL_4__378_ (
);

FILL FILL_2__441_ (
);

FILL FILL_5__585_ (
);

FILL FILL_6__527_ (
);

FILL FILL_7__314_ (
);

FILL FILL_1__463_ (
);

FILL FILL_5__394_ (
);

FILL FILL_3__612_ (
);

FILL FILL_6__336_ (
);

FILL FILL_7__543_ (
);

FILL FILL_0__485_ (
);

FILL FILL_1__519_ (
);

AOI21X1 _488_ (
    .A(_43_),
    .B(_73__bF$buf3),
    .C(_307_),
    .Y(_35_)
);

FILL FILL_3__421_ (
);

FILL FILL_6__565_ (
);

FILL FILL_7__352_ (
);

FILL FILL_1__328_ (
);

FILL FILL_2__535_ (
);

FILL FILL75450x10950 (
);

FILL FILL_6__374_ (
);

FILL FILL_7__408_ (
);

FILL FILL_7__581_ (
);

FILL FILL_1__557_ (
);

FILL FILL_8__523_ (
);

FILL FILL_2__344_ (
);

FILL FILL_5__488_ (
);

FILL FILL_0__579_ (
);

FILL FILL_7_CLKBUF1_insert0 (
);

FILL FILL_7_CLKBUF1_insert1 (
);

FILL FILL_7_CLKBUF1_insert2 (
);

FILL FILL_7_CLKBUF1_insert3 (
);

FILL FILL_7_CLKBUF1_insert4 (
);

FILL FILL_7_CLKBUF1_insert5 (
);

FILL FILL_7__390_ (
);

FILL FILL_1__366_ (
);

FILL FILL_8__332_ (
);

FILL FILL_2__573_ (
);

FILL FILL_3__515_ (
);

FILL FILL_7__446_ (
);

FILL FILL_0__388_ (
);

FILL FILL_1__595_ (
);

FILL FILL_8__561_ (
);

FILL FILL_2__382_ (
);

FILL FILL_0__600_ (
);

FILL FILL_3__324_ (
);

FILL FILL_6__468_ (
);

OR2X2 _603_ (
    .A(_128_),
    .B(_131_),
    .Y(_132_)
);

FILL FILL_4__531_ (
);

FILL FILL_8__617_ (
);

FILL FILL_8__370_ (
);

FILL FILL_2__438_ (
);

FILL FILL_3__553_ (
);

AND2X2 _412_ (
    .A(_243_),
    .B(_217_),
    .Y(_244_)
);

FILL FILL_4__340_ (
);

FILL FILL_7__484_ (
);

FILL FILL_8__426_ (
);

FILL FILL_2__667_ (
);

FILL FILL_3__609_ (
);

FILL FILL_3__362_ (
);

DFFPOSX1 _641_ (
    .D(_15_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[8])
);

FILL FILL_5__603_ (
);

FILL FILL_2__476_ (
);

FILL FILL_3__418_ (
);

FILL FILL_3__591_ (
);

FILL FILL_4__625_ (
);

FILL FILL_7__349_ (
);

INVX1 _450_ (
    .A(_272_),
    .Y(_280_)
);

FILL FILL_5__412_ (
);

FILL FILL_1__498_ (
);

FILL FILL_8__464_ (
);

FILL FILL_5_BUFX2_insert10 (
);

FILL FILL_5_BUFX2_insert11 (
);

FILL FILL_5_BUFX2_insert12 (
);

FILL FILL_5_BUFX2_insert13 (
);

FILL FILL_5_BUFX2_insert14 (
);

FILL FILL_5_BUFX2_insert15 (
);

FILL FILL_5_BUFX2_insert16 (
);

FILL FILL_5_BUFX2_insert17 (
);

FILL FILL_5_BUFX2_insert18 (
);

FILL FILL_5_BUFX2_insert19 (
);

FILL FILL_0__503_ (
);

INVX1 _506_ (
    .A(Atmp[2]),
    .Y(_51_)
);

FILL FILL_4__434_ (
);

FILL FILL_7__578_ (
);

FILL FILL_3__456_ (
);

OAI21X1 _315_ (
    .A(_152_),
    .B(_149_),
    .C(_154_),
    .Y(_155_)
);

FILL FILL_7__387_ (
);

FILL FILL_5__450_ (
);

FILL FILL_0__541_ (
);

NAND2X1 _544_ (
    .A(acc_reg[0]),
    .B(FCW[0]),
    .Y(_78_)
);

FILL FILL_4__472_ (
);

FILL FILL_5__506_ (
);

FILL FILL_8__558_ (
);

FILL FILL_6__621_ (
);

FILL FILL_2__379_ (
);

FILL FILL_0__350_ (
);

FILL FILL_3__494_ (
);

FILL FILL_4__528_ (
);

NOR2X1 _353_ (
    .A(_189_),
    .B(_188_),
    .Y(_190_)
);

FILL FILL_5__315_ (
);

FILL FILL_6__430_ (
);

FILL FILL_0__406_ (
);

OR2X2 _409_ (
    .A(_197_),
    .B(_240_),
    .Y(_241_)
);

FILL FILL_1__613_ (
);

FILL FILL_4__337_ (
);

NAND2X1 _582_ (
    .A(_112_),
    .B(_111_),
    .Y(_113_)
);

FILL FILL_2__400_ (
);

FILL FILL_5__544_ (
);

FILL FILL_8__596_ (
);

FILL FILL_3__359_ (
);

DFFPOSX1 _638_ (
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[5])
);

FILL FILL_1__422_ (
);

FILL FILL_4__566_ (
);

OAI21X1 _391_ (
    .A(_221_),
    .B(_222_),
    .C(_220_),
    .Y(_225_)
);

FILL FILL_5__353_ (
);

FILL FILL_7__502_ (
);

FILL FILL_0__444_ (
);

FILL FILL_3__588_ (
);

NOR2X1 _447_ (
    .A(acc_reg[18]),
    .B(FCW[18]),
    .Y(_277_)
);

FILL FILL_4__375_ (
);

FILL FILL_5__409_ (
);

FILL FILL_5__582_ (
);

FILL FILL_6__524_ (
);

FILL FILL_3__397_ (
);

FILL FILL_1__460_ (
);

FILL FILL_5__391_ (
);

FILL FILL_6__333_ (
);

FILL FILL_7__540_ (
);

FILL FILL_0__482_ (
);

FILL FILL_1__516_ (
);

OAI21X1 _485_ (
    .A(acc_reg[15]),
    .B(_73__bF$buf0),
    .C(En_bF$buf3),
    .Y(_306_)
);

FILL FILL_5__447_ (
);

FILL FILL_8__499_ (
);

FILL FILL_6__562_ (
);

FILL FILL_0__538_ (
);

FILL FILL_1__325_ (
);

FILL FILL_4__469_ (
);

FILL FILL_2__532_ (
);

FILL FILL_6__618_ (
);

FILL FILL_6__371_ (
);

FILL FILL_7__405_ (
);

FILL FILL_0__347_ (
);

FILL FILL_1__554_ (
);

FILL FILL_8__520_ (
);

FILL FILL_2__341_ (
);

FILL FILL_5__485_ (
);

FILL FILL_6__427_ (
);

FILL FILL_0__576_ (
);

OAI21X1 _579_ (
    .A(_108_),
    .B(_109_),
    .C(_107_),
    .Y(_110_)
);

FILL FILL_1__363_ (
);

FILL FILL_2__570_ (
);

FILL FILL_3__512_ (
);

FILL FILL_7__443_ (
);

FILL FILL_0__385_ (
);

FILL FILL_1__419_ (
);

NOR2X1 _388_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_222_)
);

FILL FILL_1__592_ (
);

FILL FILL_3__321_ (
);

FILL FILL_6__465_ (
);

NAND2X1 _600_ (
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_129_)
);

FILL FILL_8__614_ (
);

FILL FILL_2__435_ (
);

FILL FILL_5__579_ (
);

FILL FILL_3__550_ (
);

FILL FILL_7__481_ (
);

FILL FILL_1__457_ (
);

FILL FILL75750x150 (
);

FILL FILL_5__388_ (
);

FILL FILL_3__606_ (
);

FILL FILL75750x3750 (
);

FILL FILL_7__537_ (
);

FILL FILL_0__479_ (
);

FILL FILL_5__600_ (
);

FILL FILL_2__473_ (
);

FILL FILL_3__415_ (
);

FILL FILL_6__559_ (
);

FILL FILL_4__622_ (
);

FILL FILL_7__346_ (
);

FILL FILL_1__495_ (
);

FILL FILL_2__529_ (
);

FILL FILL_0__500_ (
);

FILL FILL_6__368_ (
);

OAI21X1 _503_ (
    .A(_41_),
    .B(_42_),
    .C(_47_),
    .Y(_48_)
);

FILL FILL_4__431_ (
);

FILL FILL_7__575_ (
);

FILL FILL_2__338_ (
);

FILL FILL_3__453_ (
);

FILL FILL_6__597_ (
);

FILL FILL_7__384_ (
);

FILL FILL_8__326_ (
);

FILL FILL_2__567_ (
);

FILL FILL_3__509_ (
);

NAND2X1 _541_ (
    .A(FCW[0]),
    .B(RdyCtl_6_bF$buf1),
    .Y(_76_)
);

FILL FILL_5__503_ (
);

FILL FILL_1__589_ (
);

FILL FILL_8__555_ (
);

FILL FILL_2__376_ (
);

FILL FILL_3__318_ (
);

FILL FILL_3__491_ (
);

FILL FILL_4__525_ (
);

NAND2X1 _350_ (
    .A(_186_),
    .B(_182_),
    .Y(_187_)
);

FILL FILL75450x18150 (
);

FILL FILL_1__398_ (
);

FILL FILL_8__364_ (
);

FILL FILL_0__403_ (
);

FILL FILL_3__547_ (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

AOI21X1 _406_ (
    .A(_233_),
    .B(_237_),
    .C(_238_),
    .Y(_22_)
);

FILL FILL_1__610_ (
);

FILL FILL_4__334_ (
);

FILL FILL_7__478_ (
);

FILL FILL_5__541_ (
);

FILL FILL_8__593_ (
);

FILL FILL_3__356_ (
);

DFFPOSX1 _635_ (
    .D(_9_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[2])
);

FILL FILL_4__563_ (
);

FILL FILL_5__350_ (
);

FILL FILL_0__441_ (
);

FILL FILL_3__585_ (
);

FILL FILL_4__619_ (
);

OAI21X1 _444_ (
    .A(_272_),
    .B(_261_),
    .C(_273_),
    .Y(_274_)
);

FILL FILL_4__372_ (
);

FILL FILL_5__406_ (
);

FILL FILL_8__458_ (
);

FILL FILL_6__521_ (
);

FILL FILL_3__394_ (
);

FILL FILL_4__428_ (
);

FILL FILL_6__330_ (
);

FILL FILL_3_BUFX2_insert6 (
);

FILL FILL_3_BUFX2_insert7 (
);

FILL FILL_3_BUFX2_insert8 (
);

FILL FILL_3_BUFX2_insert9 (
);

FILL FILL_1__513_ (
);

AOI21X1 _482_ (
    .A(_55_),
    .B(_73__bF$buf4),
    .C(_304_),
    .Y(_32_)
);

FILL FILL_5__444_ (
);

FILL FILL_8__496_ (
);

FILL FILL_0__535_ (
);

NAND2X1 _538_ (
    .A(En_bF$buf3),
    .B(_44_),
    .Y(_5_)
);

FILL FILL_1__322_ (
);

FILL FILL_4__466_ (
);

FILL FILL_6__615_ (
);

FILL FILL_7__402_ (
);

FILL FILL_0__344_ (
);

FILL FILL_3__488_ (
);

OAI21X1 _347_ (
    .A(acc_reg[10]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_185_)
);

FILL FILL_1__551_ (
);

FILL FILL_5__482_ (
);

FILL FILL_6__424_ (
);

FILL FILL_0__573_ (
);

FILL FILL_1__607_ (
);

AND2X2 _576_ (
    .A(_104_),
    .B(_106_),
    .Y(_107_)
);

FILL FILL_1__360_ (
);

FILL FILL_5__538_ (
);

FILL FILL_7__440_ (
);

FILL FILL_0__382_ (
);

FILL FILL_1__416_ (
);

OAI21X1 _385_ (
    .A(_203_),
    .B(_218_),
    .C(_211_),
    .Y(_219_)
);

FILL FILL_2__623_ (
);

FILL FILL_5__347_ (
);

FILL FILL75150x64950 (
);

FILL FILL_6__462_ (
);

FILL FILL_0__438_ (
);

FILL FILL_4__369_ (
);

FILL FILL_2__432_ (
);

FILL FILL_5__576_ (
);

FILL FILL_6__518_ (
);

FILL FILL_0__667_ (
);

FILL FILL_1__454_ (
);

FILL FILL_8__420_ (
);

FILL FILL_4__598_ (
);

FILL FILL_5__385_ (
);

FILL FILL_3__603_ (
);

FILL FILL_6__327_ (
);

FILL FILL_5_CLKBUF1_insert0 (
);

FILL FILL_5_CLKBUF1_insert1 (
);

FILL FILL_5_CLKBUF1_insert2 (
);

FILL FILL_5_CLKBUF1_insert3 (
);

FILL FILL_5_CLKBUF1_insert4 (
);

FILL FILL_5_CLKBUF1_insert5 (
);

FILL FILL_7__534_ (
);

FILL FILL_0__476_ (
);

OAI21X1 _479_ (
    .A(acc_reg[12]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_303_)
);

FILL FILL_2__470_ (
);

FILL FILL_3__412_ (
);

FILL FILL_6__556_ (
);

FILL FILL_7__343_ (
);

FILL FILL_1__319_ (
);

FILL FILL_1__492_ (
);

FILL FILL_2__526_ (
);

FILL FILL_6__365_ (
);

NAND2X1 _500_ (
    .A(Atmp[11]),
    .B(_44_),
    .Y(_45_)
);

FILL FILL_7__572_ (
);

FILL FILL_1__548_ (
);

FILL FILL_8__514_ (
);

FILL FILL_2__335_ (
);

FILL FILL_5__479_ (
);

FILL FILL_3__450_ (
);

FILL FILL_6__594_ (
);

FILL FILL_7__381_ (
);

FILL FILL_1__357_ (
);

FILL FILL_8__323_ (
);

FILL FILL_2__564_ (
);

FILL FILL_3__506_ (
);

FILL FILL_7__437_ (
);

FILL FILL_0__379_ (
);

FILL FILL_5__500_ (
);

FILL FILL_1__586_ (
);

FILL FILL_8__552_ (
);

FILL FILL_2__373_ (
);

FILL FILL_3__315_ (
);

FILL FILL_6__459_ (
);

FILL FILL_4__522_ (
);

FILL FILL_7__666_ (
);

FILL FILL_8__608_ (
);

FILL FILL_1__395_ (
);

FILL FILL_8__361_ (
);

FILL FILL_2__429_ (
);

FILL FILL_0__400_ (
);

FILL FILL_3__544_ (
);

FILL FILL75450x39750 (
);

NAND2X1 _403_ (
    .A(_229_),
    .B(_235_),
    .Y(_236_)
);

FILL FILL_4__331_ (
);

FILL FILL_7__475_ (
);

FILL FILL_8__417_ (
);

FILL FILL_8__590_ (
);

FILL FILL_3__353_ (
);

FILL FILL_6__497_ (
);

DFFPOSX1 _632_ (
    .D(_6_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[6])
);

FILL FILL_4__560_ (
);

FILL FILL73950x36150 (
);

FILL FILL_2__467_ (
);

FILL FILL_3__409_ (
);

FILL FILL_3__582_ (
);

FILL FILL_4__616_ (
);

AOI21X1 _441_ (
    .A(_269_),
    .B(_270_),
    .C(_271_),
    .Y(_24_)
);

FILL FILL_5__403_ (
);

FILL FILL76050x10950 (
);

FILL FILL_1__489_ (
);

FILL FILL_8__455_ (
);

FILL FILL_3__391_ (
);

FILL FILL_4__425_ (
);

FILL FILL_7__569_ (
);

FILL FILL_3__447_ (
);

FILL FILL_1__510_ (
);

FILL FILL_7__378_ (
);

FILL FILL_5__441_ (
);

FILL FILL_0__532_ (
);

AND2X2 _535_ (
    .A(RdyCtl[1]),
    .B(En_bF$buf4),
    .Y(_2_)
);

FILL FILL_4__463_ (
);

FILL FILL_8__549_ (
);

FILL FILL_6__612_ (
);

FILL FILL_0__341_ (
);

FILL FILL_3__485_ (
);

FILL FILL_4__519_ (
);

NAND2X1 _344_ (
    .A(_181_),
    .B(_178_),
    .Y(_182_)
);

FILL FILL_8__358_ (
);

FILL FILL_6__421_ (
);

FILL FILL_2__599_ (
);

FILL FILL74850x50550 (
);

FILL FILL_0__570_ (
);

FILL FILL_1__604_ (
);

FILL FILL_4__328_ (
);

NAND3X1 _573_ (
    .A(_88_),
    .B(_91_),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_5__535_ (
);

DFFPOSX1 _629_ (
    .D(_3_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[3])
);

FILL FILL_1__413_ (
);

FILL FILL_4__557_ (
);

AOI21X1 _382_ (
    .A(_214_),
    .B(_215_),
    .C(_216_),
    .Y(_20_)
);

FILL FILL_2__620_ (
);

FILL FILL_5__344_ (
);

FILL FILL_8__396_ (
);

FILL FILL_0__435_ (
);

FILL FILL_3__579_ (
);

OR2X2 _438_ (
    .A(_265_),
    .B(_268_),
    .Y(_269_)
);

FILL FILL_4__366_ (
);

FILL FILL_5__573_ (
);

FILL FILL_6__515_ (
);

FILL FILL_3__388_ (
);

BUFX2 _667_ (
    .A(_312_),
    .Y(ISout)
);

FILL FILL_1__451_ (
);

FILL FILL_4__595_ (
);

FILL FILL_5__382_ (
);

FILL FILL_3__600_ (
);

FILL FILL_6__324_ (
);

FILL FILL_7__531_ (
);

FILL FILL_0__473_ (
);

FILL FILL_1__507_ (
);

AOI21X1 _476_ (
    .A(_51_),
    .B(_73__bF$buf1),
    .C(_301_),
    .Y(_29_)
);

FILL FILL_5__438_ (
);

FILL FILL_6__553_ (
);

FILL FILL_0__529_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_7__340_ (
);

FILL FILL_1__316_ (
);

FILL FILL_2__523_ (
);

FILL FILL_5__667_ (
);

FILL FILL_6__609_ (
);

FILL FILL_6__362_ (
);

FILL FILL_0__338_ (
);

FILL FILL_1__545_ (
);

FILL FILL_8__511_ (
);

FILL FILL_2__332_ (
);

FILL FILL_5__476_ (
);

FILL FILL_6__418_ (
);

FILL FILL_6__591_ (
);

FILL FILL74550x7350 (
);

FILL FILL_7__625_ (
);

FILL FILL_0__567_ (
);

FILL FILL_1__354_ (
);

FILL FILL75150x50550 (
);

FILL FILL_4__498_ (
);

FILL FILL_2__561_ (
);

FILL FILL_3__503_ (
);

FILL FILL76050x150 (
);

FILL FILL_7__434_ (
);

FILL FILL_0__376_ (
);

OR2X2 _379_ (
    .A(_210_),
    .B(_213_),
    .Y(_214_)
);

FILL FILL_1__583_ (
);

FILL FILL_2__617_ (
);

FILL FILL_2__370_ (
);

FILL FILL_6__456_ (
);

FILL FILL_8__605_ (
);

FILL FILL_1__392_ (
);

FILL FILL_2__426_ (
);

FILL FILL_3__541_ (
);

NAND3X1 _400_ (
    .A(_228_),
    .B(_232_),
    .C(_224_),
    .Y(_233_)
);

FILL FILL_7__472_ (
);

FILL FILL_1__448_ (
);

FILL FILL_5__379_ (
);

FILL FILL_3__350_ (
);

FILL FILL_6__494_ (
);

FILL FILL_7__528_ (
);

FILL FILL_2__464_ (
);

FILL FILL_3__406_ (
);

FILL FILL73950x57750 (
);

FILL FILL_4__613_ (
);

FILL FILL_7__337_ (
);

FILL FILL_5__400_ (
);

FILL FILL_1__486_ (
);

FILL FILL_8__452_ (
);

FILL FILL_6__359_ (
);

FILL FILL_4__422_ (
);

FILL FILL_7__566_ (
);

FILL FILL_8__508_ (
);

FILL FILL_2__329_ (
);

FILL FILL_3__444_ (
);

FILL FILL_6__588_ (
);

FILL FILL_7__375_ (
);

FILL FILL_8__317_ (
);

FILL FILL_8__490_ (
);

FILL FILL_2__558_ (
);

FILL FILL_6__397_ (
);

INVX2 _532_ (
    .A(En_bF$buf1),
    .Y(_74_)
);

FILL FILL_4__460_ (
);

FILL FILL_8__546_ (
);

FILL FILL75450x25350 (
);

FILL FILL_2__367_ (
);

FILL FILL_3__482_ (
);

FILL FILL_4__516_ (
);

AND2X2 _341_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_179_)
);

FILL FILL_1__389_ (
);

FILL FILL_8__355_ (
);

FILL FILL_2__596_ (
);

FILL FILL_3__538_ (
);

FILL FILL_1__601_ (
);

FILL FILL_4__325_ (
);

FILL FILL_7__469_ (
);

OAI21X1 _570_ (
    .A(_97_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_5__532_ (
);

FILL FILL_8__584_ (
);

FILL FILL_0__623_ (
);

FILL FILL_3__347_ (
);

DFFPOSX1 _626_ (
    .D(_0_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[0])
);

FILL FILL_1__410_ (
);

FILL FILL_4__554_ (
);

FILL FILL_5__341_ (
);

FILL FILL75750x68550 (
);

FILL FILL_8__393_ (
);

FILL FILL_0__432_ (
);

FILL FILL_3__576_ (
);

AND2X2 _435_ (
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_266_)
);

FILL FILL_4__363_ (
);

FILL FILL_8__449_ (
);

FILL FILL_5__570_ (
);

FILL FILL_6__512_ (
);

FILL FILL75150x3750 (
);

FILL FILL_3__385_ (
);

FILL FILL_4__419_ (
);

DFFPOSX1 _664_ (
    .D(_38_),
    .CLK(clk_bF$buf2),
    .Q(_312_)
);

FILL FILL73050x39750 (
);

FILL FILL_4__592_ (
);

FILL FILL_6__321_ (
);

FILL FILL_2__499_ (
);

FILL FILL_0__470_ (
);

FILL FILL_1__504_ (
);

OAI21X1 _473_ (
    .A(acc_reg[9]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_300_)
);

FILL FILL_5__435_ (
);

FILL FILL_8__487_ (
);

FILL FILL_6__550_ (
);

FILL FILL_0__526_ (
);

NAND2X1 _529_ (
    .A(_312_),
    .B(_66_),
    .Y(_72_)
);

FILL FILL_1__313_ (
);

FILL FILL_4__457_ (
);

FILL FILL_2__520_ (
);

FILL FILL_6__606_ (
);

FILL FILL76050x18150 (
);

FILL FILL_0__335_ (
);

FILL FILL_3__479_ (
);

INVX1 _338_ (
    .A(_175_),
    .Y(_176_)
);

FILL FILL_1__542_ (
);

FILL FILL_5__473_ (
);

FILL FILL_6__415_ (
);

FILL FILL_7__622_ (
);

FILL FILL_0__564_ (
);

NOR2X1 _567_ (
    .A(_98_),
    .B(_97_),
    .Y(_99_)
);

FILL FILL_1__351_ (
);

FILL FILL_4__495_ (
);

FILL FILL_5__529_ (
);

FILL FILL_3__500_ (
);

FILL FILL_3_CLKBUF1_insert0 (
);

FILL FILL_3_CLKBUF1_insert1 (
);

FILL FILL_3_CLKBUF1_insert2 (
);

FILL FILL_3_CLKBUF1_insert3 (
);

FILL FILL_3_CLKBUF1_insert4 (
);

FILL FILL_3_CLKBUF1_insert5 (
);

FILL FILL_7__431_ (
);

FILL FILL_0__373_ (
);

FILL FILL_1__407_ (
);

NAND2X1 _376_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_211_)
);

FILL FILL_1__580_ (
);

FILL FILL_2__614_ (
);

FILL FILL_5__338_ (
);

FILL FILL_6__453_ (
);

FILL FILL_0__429_ (
);

FILL FILL_8__602_ (
);

FILL FILL_2__423_ (
);

FILL FILL_5__567_ (
);

FILL FILL_6__509_ (
);

FILL FILL_1__445_ (
);

FILL FILL_8__411_ (
);

FILL FILL_4__589_ (
);

FILL FILL_5__376_ (
);

FILL FILL_6__318_ (
);

FILL FILL_6__491_ (
);

FILL FILL_7__525_ (
);

FILL FILL_0__467_ (
);

FILL FILL_4__398_ (
);

FILL FILL_2__461_ (
);

FILL FILL_3__403_ (
);

FILL FILL_6__547_ (
);

FILL FILL_4__610_ (
);

FILL FILL_7__334_ (
);

FILL FILL_1__483_ (
);

FILL FILL_2__517_ (
);

FILL FILL_6__356_ (
);

FILL FILL_7__563_ (
);

FILL FILL_1__539_ (
);

FILL FILL_8__505_ (
);

FILL FILL_7_BUFX2_insert10 (
);

FILL FILL_7_BUFX2_insert11 (
);

FILL FILL_7_BUFX2_insert12 (
);

FILL FILL_7_BUFX2_insert13 (
);

FILL FILL_7_BUFX2_insert14 (
);

FILL FILL_7_BUFX2_insert15 (
);

FILL FILL_7_BUFX2_insert16 (
);

FILL FILL_7_BUFX2_insert17 (
);

FILL FILL_7_BUFX2_insert18 (
);

FILL FILL_7_BUFX2_insert19 (
);

FILL FILL_2__326_ (
);

FILL FILL_3__441_ (
);

FILL FILL_6__585_ (
);

FILL FILL_7__619_ (
);

FILL FILL_7__372_ (
);

FILL FILL_1__348_ (
);

FILL FILL_8__314_ (
);

FILL FILL_2__555_ (
);

FILL FILL_6__394_ (
);

FILL FILL_7__428_ (
);

FILL FILL_1__577_ (
);

FILL FILL_8__543_ (
);

FILL FILL_2__364_ (
);

FILL FILL_4__513_ (
);

FILL FILL_0__599_ (
);

FILL FILL75450x46950 (
);

FILL FILL_1__386_ (
);

FILL FILL_8__352_ (
);

FILL FILL_2__593_ (
);

FILL FILL74250x61350 (
);

FILL FILL_3__535_ (
);

FILL FILL74250x28950 (
);

FILL FILL_4__322_ (
);

FILL FILL_7__466_ (
);

FILL FILL_8__408_ (
);

FILL FILL_8__581_ (
);

FILL FILL_0__620_ (
);

FILL FILL_3__344_ (
);

FILL FILL_6__488_ (
);

NOR2X1 _623_ (
    .A(_145_),
    .B(_149_),
    .Y(_150_)
);

FILL FILL_4__551_ (
);

FILL FILL_2__458_ (
);

FILL FILL_3__573_ (
);

FILL FILL_4__607_ (
);

OAI21X1 _432_ (
    .A(acc_reg[16]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_264_)
);

FILL FILL_4__360_ (
);

FILL FILL_3__382_ (
);

FILL FILL_4__416_ (
);

DFFPOSX1 _661_ (
    .D(_35_),
    .CLK(clk_bF$buf3),
    .Q(Atmp[8])
);

FILL FILL_5__623_ (
);

FILL FILL_2__496_ (
);

FILL FILL_3__438_ (
);

FILL FILL_1__501_ (
);

FILL FILL_7__369_ (
);

OAI21X1 _470_ (
    .A(acc_reg[8]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_298_)
);

FILL FILL_5__432_ (
);

FILL FILL_0__523_ (
);

FILL FILL_3__667_ (
);

INVX1 _526_ (
    .A(acc_reg[19]),
    .Y(_69_)
);

FILL FILL_4__454_ (
);

FILL FILL_7__598_ (
);

FILL FILL_6__603_ (
);

FILL FILL_0__332_ (
);

FILL FILL_3__476_ (
);

AOI21X1 _335_ (
    .A(_172_),
    .B(_170_),
    .C(_173_),
    .Y(_16_)
);

FILL FILL_8__349_ (
);

FILL FILL76050x39750 (
);

FILL FILL_5__470_ (
);

FILL FILL_6__412_ (
);

FILL FILL_0__561_ (
);

FILL FILL_4__319_ (
);

OAI21X1 _564_ (
    .A(acc_reg[3]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_96_)
);

FILL FILL75750x54150 (
);

FILL FILL_4__492_ (
);

FILL FILL_5__526_ (
);

FILL FILL_2__399_ (
);

FILL FILL_0__617_ (
);

FILL FILL74550x36150 (
);

FILL FILL_0__370_ (
);

FILL FILL_1__404_ (
);

FILL FILL_4__548_ (
);

AOI21X1 _373_ (
    .A(_208_),
    .B(_195_),
    .C(_74_),
    .Y(_19_)
);

FILL FILL_2__611_ (
);

FILL FILL_5__335_ (
);

FILL FILL_8__387_ (
);

FILL FILL_6__450_ (
);

FILL FILL_0__426_ (
);

AOI21X1 _429_ (
    .A(_257_),
    .B(_258_),
    .C(_260_),
    .Y(_261_)
);

FILL FILL_4__357_ (
);

FILL FILL_2__420_ (
);

FILL FILL_5__564_ (
);

FILL FILL_6__506_ (
);

FILL FILL_3__379_ (
);

DFFPOSX1 _658_ (
    .D(_32_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[5])
);

FILL FILL_1__442_ (
);

FILL FILL_4__586_ (
);

FILL FILL_5__373_ (
);

FILL FILL_6__315_ (
);

FILL FILL_7__522_ (
);

FILL FILL_0__464_ (
);

AOI21X1 _467_ (
    .A(_294_),
    .B(_295_),
    .C(_73__bF$buf2),
    .Y(_296_)
);

FILL FILL_4__395_ (
);

FILL FILL_5__429_ (
);

FILL FILL_3__400_ (
);

FILL FILL_6__544_ (
);

FILL FILL_7__331_ (
);

FILL FILL_1__480_ (
);

FILL FILL_2__514_ (
);

FILL FILL_6__353_ (
);

FILL FILL_0__329_ (
);

FILL FILL_7__560_ (
);

FILL FILL_1__536_ (
);

FILL FILL_8__502_ (
);

FILL FILL_2__323_ (
);

FILL FILL_5__467_ (
);

FILL FILL_6__409_ (
);

FILL FILL_6__582_ (
);

FILL FILL_7__616_ (
);

FILL FILL_0__558_ (
);

FILL FILL_1__345_ (
);

FILL FILL_4__489_ (
);

FILL FILL_2__552_ (
);

FILL FILL_6__391_ (
);

FILL FILL_7__425_ (
);

FILL FILL_0__367_ (
);

FILL FILL_1__574_ (
);

FILL FILL_2__608_ (
);

FILL FILL74850x3750 (
);

FILL FILL_2__361_ (
);

FILL FILL_6__447_ (
);

FILL FILL_4__510_ (
);

FILL FILL_0__596_ (
);

AOI21X1 _599_ (
    .A(_111_),
    .B(_127_),
    .C(_126_),
    .Y(_128_)
);

FILL FILL_1__383_ (
);

FILL FILL_2__417_ (
);

FILL FILL_2__590_ (
);

FILL FILL_3__532_ (
);

FILL FILL_7__463_ (
);

FILL FILL_1__439_ (
);

FILL FILL_8__405_ (
);

FILL FILL_3__341_ (
);

FILL FILL_6__485_ (
);

FILL FILL_7__519_ (
);

NOR2X1 _620_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_147_)
);

FILL FILL_1__668_ (
);

FILL FILL_2__455_ (
);

FILL FILL_5__599_ (
);

FILL FILL_3__570_ (
);

FILL FILL_4__604_ (
);

FILL FILL_7__328_ (
);

FILL FILL_1__477_ (
);

FILL FILL_8__443_ (
);

FILL FILL_4__413_ (
);

FILL FILL_7__557_ (
);

FILL FILL_0__499_ (
);

FILL FILL_5__620_ (
);

FILL FILL_2__493_ (
);

FILL FILL_3__435_ (
);

FILL FILL_6__579_ (
);

FILL FILL_7__366_ (
);

FILL FILL_8__481_ (
);

FILL FILL_2__549_ (
);

FILL FILL_0__520_ (
);

FILL FILL_6__388_ (
);

INVX1 _523_ (
    .A(RdyCtl[5]),
    .Y(_66_)
);

FILL FILL_4__451_ (
);

FILL FILL_7__595_ (
);

FILL FILL_8__537_ (
);

FILL FILL_6__600_ (
);

FILL FILL_2__358_ (
);

FILL FILL74250x14550 (
);

FILL FILL_3__473_ (
);

FILL FILL_4__507_ (
);

NOR2X1 _332_ (
    .A(_169_),
    .B(_164_),
    .Y(_171_)
);

FILL FILL_8__346_ (
);

FILL FILL_2__587_ (
);

FILL FILL_3__529_ (
);

FILL FILL_4__316_ (
);

OAI21X1 _561_ (
    .A(_88_),
    .B(_91_),
    .C(_93_),
    .Y(_94_)
);

FILL FILL_5__523_ (
);

FILL FILL_8__575_ (
);

FILL FILL_2__396_ (
);

FILL FILL_0__614_ (
);

FILL FILL_3__338_ (
);

AOI21X1 _617_ (
    .A(_142_),
    .B(_143_),
    .C(_144_),
    .Y(_14_)
);

FILL FILL_1__401_ (
);

FILL FILL_4__545_ (
);

NOR2X1 _370_ (
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

FILL FILL_5__332_ (
);

FILL FILL_8__384_ (
);

FILL FILL74550x57750 (
);

FILL FILL_0__423_ (
);

FILL FILL_3__567_ (
);

NOR2X1 _426_ (
    .A(_197_),
    .B(_240_),
    .Y(_258_)
);

FILL FILL_4__354_ (
);

FILL FILL_7__498_ (
);

FILL FILL_5__561_ (
);

FILL FILL_6__503_ (
);

FILL FILL_3__376_ (
);

DFFPOSX1 _655_ (
    .D(_29_),
    .CLK(clk_bF$buf4),
    .Q(Atmp[2])
);

FILL FILL_4__583_ (
);

FILL FILL_5__617_ (
);

FILL FILL_5__370_ (
);

FILL FILL_0__461_ (
);

NAND2X1 _464_ (
    .A(_292_),
    .B(_289_),
    .Y(_293_)
);

FILL FILL_4__392_ (
);

FILL FILL_5__426_ (
);

FILL FILL_8__478_ (
);

FILL FILL_1_CLKBUF1_insert0 (
);

FILL FILL_1_CLKBUF1_insert1 (
);

FILL FILL_1_CLKBUF1_insert2 (
);

FILL FILL_1_CLKBUF1_insert3 (
);

FILL FILL_1_CLKBUF1_insert4 (
);

FILL FILL_1_CLKBUF1_insert5 (
);

FILL FILL_6__541_ (
);

FILL FILL_0__517_ (
);

FILL FILL74850x10950 (
);

FILL FILL_4__448_ (
);

FILL FILL76050x25350 (
);

FILL FILL_2__511_ (
);

FILL FILL_6__350_ (
);

FILL FILL_0__326_ (
);

NAND2X1 _329_ (
    .A(_166_),
    .B(_167_),
    .Y(_168_)
);

FILL FILL_1__533_ (
);

FILL FILL_2__320_ (
);

FILL FILL_5__464_ (
);

FILL FILL_6__406_ (
);

FILL FILL_7__613_ (
);

FILL FILL_0__555_ (
);

NOR2X1 _558_ (
    .A(_90_),
    .B(_89_),
    .Y(_91_)
);

FILL FILL_1__342_ (
);

FILL FILL_4__486_ (
);

FILL FILL_7__422_ (
);

FILL FILL_0__364_ (
);

NAND2X1 _367_ (
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_203_)
);

FILL FILL_1__571_ (
);

FILL FILL_2__605_ (
);

FILL FILL_5__329_ (
);

FILL FILL_6__444_ (
);

FILL FILL_0__593_ (
);

INVX1 _596_ (
    .A(_117_),
    .Y(_125_)
);

FILL FILL_1__380_ (
);

FILL FILL_2__414_ (
);

FILL FILL_5__558_ (
);

FILL FILL_7__460_ (
);

FILL FILL_1__436_ (
);

FILL FILL_8__402_ (
);

FILL FILL_5__367_ (
);

FILL FILL_6__482_ (
);

FILL FILL_7__516_ (
);

FILL FILL_0__458_ (
);

BUFX2 BUFX2_insert6 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf1)
);

FILL FILL_1__665_ (
);

FILL FILL_4__389_ (
);

FILL FILL_2__452_ (
);

FILL FILL_5__596_ (
);

FILL FILL_6__538_ (
);

FILL FILL_4__601_ (
);

FILL FILL_7__325_ (
);

FILL FILL_1__474_ (
);

FILL FILL_8__440_ (
);

FILL FILL_2__508_ (
);

FILL FILL75150x10950 (
);

FILL FILL_3__623_ (
);

FILL FILL_6__347_ (
);

FILL FILL_4__410_ (
);

FILL FILL_7__554_ (
);

FILL FILL_0__496_ (
);

INVX1 _499_ (
    .A(RdyCtl[4]),
    .Y(_44_)
);

FILL FILL_2__317_ (
);

FILL FILL_2__490_ (
);

FILL FILL_3__432_ (
);

FILL FILL_6__576_ (
);

FILL FILL_7__363_ (
);

FILL FILL_1__339_ (
);

FILL FILL_2__546_ (
);

FILL FILL_6__385_ (
);

FILL FILL_7__419_ (
);

OAI21X1 _520_ (
    .A(RdyCtl[1]),
    .B(_61_),
    .C(_63_),
    .Y(_64_)
);

FILL FILL_7__592_ (
);

FILL FILL_1__568_ (
);

FILL FILL_8__534_ (
);

FILL FILL_2__355_ (
);

FILL FILL_5__499_ (
);

FILL FILL_3__470_ (
);

FILL FILL_4__504_ (
);

FILL FILL_1__377_ (
);

FILL FILL_2__584_ (
);

FILL FILL_3__526_ (
);

FILL FILL73950x50550 (
);

FILL FILL_4__313_ (
);

FILL FILL_7__457_ (
);

FILL FILL_0__399_ (
);

FILL FILL_5__520_ (
);

FILL FILL_8__572_ (
);

FILL FILL_2__393_ (
);

FILL FILL_0__611_ (
);

FILL FILL_3__335_ (
);

FILL FILL_6__479_ (
);

OR2X2 _614_ (
    .A(_138_),
    .B(_141_),
    .Y(_142_)
);

FILL FILL_4__542_ (
);

FILL FILL_2__449_ (
);

FILL FILL_0__420_ (
);

FILL FILL_3__564_ (
);

NAND2X1 _423_ (
    .A(_254_),
    .B(_127_),
    .Y(_255_)
);

FILL FILL_4__351_ (
);

FILL FILL_7__495_ (
);

FILL FILL_6__500_ (
);

FILL FILL_3__373_ (
);

FILL FILL_4__407_ (
);

DFFPOSX1 _652_ (
    .D(_26_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[19])
);

FILL FILL_4__580_ (
);

FILL FILL_5__614_ (
);

FILL FILL_8__666_ (
);

FILL FILL_2__487_ (
);

FILL FILL_3__429_ (
);

NAND2X1 _461_ (
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_290_)
);

FILL FILL_5__423_ (
);

FILL FILL_0__514_ (
);

OAI21X1 _517_ (
    .A(_40_),
    .B(_55_),
    .C(_60_),
    .Y(_61_)
);

FILL FILL_4__445_ (
);

FILL FILL_7__589_ (
);

FILL FILL_0__323_ (
);

FILL FILL76050x46950 (
);

FILL FILL_3__467_ (
);

FILL FILL_4_BUFX2_insert20 (
);

NAND2X1 _326_ (
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_165_)
);

FILL FILL_1__530_ (
);

FILL FILL_7__398_ (
);

FILL FILL_5__461_ (
);

FILL FILL75750x61350 (
);

FILL FILL_6__403_ (
);

FILL FILL75750x28950 (
);

FILL FILL_7__610_ (
);

FILL FILL_0__552_ (
);

OAI21X1 _555_ (
    .A(_78_),
    .B(_81_),
    .C(_79_),
    .Y(_88_)
);

FILL FILL_4__483_ (
);

FILL FILL_5__517_ (
);

FILL FILL_8__569_ (
);

FILL FILL_0__608_ (
);

FILL FILL_0__361_ (
);

FILL FILL_4__539_ (
);

AOI21X1 _364_ (
    .A(_199_),
    .B(_179_),
    .C(_188_),
    .Y(_200_)
);

FILL FILL_2__602_ (
);

FILL FILL_5__326_ (
);

FILL FILL_8__378_ (
);

FILL FILL_6__441_ (
);

FILL FILL_0__417_ (
);

FILL FILL_0__590_ (
);

FILL FILL_1__624_ (
);

FILL FILL_4__348_ (
);

OAI21X1 _593_ (
    .A(acc_reg[5]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_123_)
);

FILL FILL_2__411_ (
);

FILL FILL_5__555_ (
);

DFFPOSX1 _649_ (
    .D(_23_),
    .CLK(clk_bF$buf5),
    .Q(acc_reg[16])
);

FILL FILL_1__433_ (
);

FILL FILL_4__577_ (
);

FILL FILL_5__364_ (
);

FILL FILL_7__513_ (
);

FILL FILL_0__455_ (
);

FILL FILL_3__599_ (
);

NAND2X1 _458_ (
    .A(acc_reg[19]),
    .B(En_bF$buf4),
    .Y(_287_)
);

FILL FILL_4__386_ (
);

FILL FILL_5__593_ (
);

FILL FILL_6__535_ (
);

FILL FILL_7__322_ (
);

FILL FILL_1__471_ (
);

FILL FILL_2__505_ (
);

FILL FILL_3__620_ (
);

FILL FILL_6__344_ (
);

FILL FILL_7__551_ (
);

FILL FILL_0__493_ (
);

FILL FILL_1__527_ (
);

INVX1 _496_ (
    .A(Atmp[6]),
    .Y(_41_)
);

FILL FILL_2__314_ (
);

FILL FILL_5__458_ (
);

FILL FILL_6__573_ (
);

FILL FILL_7__607_ (
);

FILL FILL_0__549_ (
);

FILL FILL_7__360_ (
);

FILL FILL_1__336_ (
);

FILL FILL_2__543_ (
);

FILL FILL_6__382_ (
);

FILL FILL_7__416_ (
);

FILL FILL_0__358_ (
);

FILL FILL75450x7350 (
);

FILL FILL_1__565_ (
);

FILL FILL74850x18150 (
);

FILL FILL_2__352_ (
);

FILL FILL_5__496_ (
);

FILL FILL_6__438_ (
);

FILL FILL_4__501_ (
);

FILL FILL_0__587_ (
);

FILL FILL_1__374_ (
);

FILL FILL_8__340_ (
);

FILL FILL_2__408_ (
);

FILL FILL_2__581_ (
);

FILL FILL_3__523_ (
);

FILL FILL_6__667_ (
);

FILL FILL_7__454_ (
);

FILL FILL_0__396_ (
);

NOR2X1 _399_ (
    .A(_231_),
    .B(_230_),
    .Y(_232_)
);

FILL FILL_2__390_ (
);

FILL FILL_3__332_ (
);

FILL FILL_6__476_ (
);

NAND2X1 _611_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_139_)
);

FILL FILL_2__446_ (
);

FILL FILL_3__561_ (
);

FILL FILL_7__319_ (
);

NOR2X1 _420_ (
    .A(_251_),
    .B(_250_),
    .Y(_252_)
);

FILL FILL_7__492_ (
);

FILL FILL_1__468_ (
);

FILL FILL_8__434_ (
);

FILL FILL_5__399_ (
);

FILL FILL_3__617_ (
);

FILL FILL_3__370_ (
);

FILL FILL_4__404_ (
);

FILL FILL_7__548_ (
);

FILL FILL_5__611_ (
);

FILL FILL_2__484_ (
);

FILL FILL_3__426_ (
);

FILL FILL_7__357_ (
);

FILL FILL_5__420_ (
);

FILL FILL_8__472_ (
);

FILL FILL_0__511_ (
);

FILL FILL_6__379_ (
);

INVX1 _514_ (
    .A(Atmp[7]),
    .Y(_58_)
);

FILL FILL_4__442_ (
);

FILL FILL_7__586_ (
);

FILL FILL_8__528_ (
);

FILL FILL_2__349_ (
);

FILL FILL_0__320_ (
);

FILL FILL_3__464_ (
);

OAI21X1 _323_ (
    .A(acc_reg[8]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_163_)
);

FILL FILL75150x18150 (
);

FILL FILL_7__395_ (
);

FILL FILL_8__337_ (
);

FILL FILL_6__400_ (
);

FILL FILL_2__578_ (
);

NAND2X1 _552_ (
    .A(_82_),
    .B(_85_),
    .Y(_86_)
);

FILL FILL_4__480_ (
);

FILL FILL_5__514_ (
);

FILL FILL_8__566_ (
);

FILL FILL_2__387_ (
);

FILL FILL_0__605_ (
);

FILL FILL_3__329_ (
);

OAI21X1 _608_ (
    .A(acc_reg[6]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_137_)
);

FILL FILL_4__536_ (
);

NAND3X1 _361_ (
    .A(_181_),
    .B(_190_),
    .C(_196_),
    .Y(_197_)
);

FILL FILL_5__323_ (
);

FILL FILL_8__375_ (
);

FILL FILL_0__414_ (
);

FILL FILL_3__558_ (
);

OAI21X1 _417_ (
    .A(_156_),
    .B(_241_),
    .C(_248_),
    .Y(_249_)
);

FILL FILL_1__621_ (
);

FILL FILL_4__345_ (
);

FILL FILL_7__489_ (
);

NAND2X1 _590_ (
    .A(_119_),
    .B(_116_),
    .Y(_120_)
);

FILL FILL_5__552_ (
);

FILL FILL_3__367_ (
);

DFFPOSX1 _646_ (
    .D(_20_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[13])
);

FILL FILL_1__430_ (
);

FILL FILL_4__574_ (
);

FILL FILL_5__608_ (
);

FILL FILL_5__361_ (
);

FILL FILL_7__510_ (
);

FILL FILL_0__452_ (
);

FILL FILL_3__596_ (
);

OAI21X1 _455_ (
    .A(acc_reg[18]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf4),
    .Y(_285_)
);

FILL FILL76050x3750 (
);

FILL FILL_4__383_ (
);

FILL FILL_5__417_ (
);

FILL FILL_8__469_ (
);

FILL FILL_5__590_ (
);

FILL FILL_6__532_ (
);

FILL FILL_0__508_ (
);

FILL FILL_4__439_ (
);

FILL FILL_2__502_ (
);

FILL FILL75750x14550 (
);

FILL FILL_6__341_ (
);

FILL FILL_0__317_ (
);

FILL FILL_0__490_ (
);

FILL FILL_1__524_ (
);

FILL FILL_4__668_ (
);

NOR2X1 _493_ (
    .A(_309_),
    .B(_310_),
    .Y(_37_)
);

FILL FILL_5__455_ (
);

FILL FILL_6__570_ (
);

FILL FILL_7__604_ (
);

FILL FILL_0__546_ (
);

OR2X2 _549_ (
    .A(_80_),
    .B(_81_),
    .Y(_83_)
);

FILL FILL_1__333_ (
);

FILL FILL_4__477_ (
);

FILL FILL_2__540_ (
);

FILL FILL_7__413_ (
);

FILL FILL_0__355_ (
);

FILL FILL_3__499_ (
);

AOI21X1 _358_ (
    .A(_192_),
    .B(_193_),
    .C(_194_),
    .Y(_18_)
);

FILL FILL_1__562_ (
);

FILL FILL_5__493_ (
);

FILL FILL_6__435_ (
);

FILL FILL_0__584_ (
);

FILL FILL_1__618_ (
);

AND2X2 _587_ (
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_117_)
);

FILL FILL74850x39750 (
);

FILL FILL_1__371_ (
);

FILL FILL_2__405_ (
);

FILL FILL_5__549_ (
);

FILL FILL_3__520_ (
);

FILL FILL_7__451_ (
);

FILL FILL_0__393_ (
);

FILL FILL_1__427_ (
);

NAND2X1 _396_ (
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_229_)
);

FILL FILL_5__358_ (
);

FILL FILL_6__473_ (
);

FILL FILL_7__507_ (
);

FILL FILL_0__449_ (
);

FILL FILL_8__622_ (
);

FILL FILL_2__443_ (
);

FILL FILL_5__587_ (
);

FILL FILL_6__529_ (
);

FILL FILL_7__316_ (
);

FILL FILL_1__465_ (
);

FILL FILL_8__431_ (
);

FILL FILL_5__396_ (
);

FILL FILL_3__614_ (
);

FILL FILL_6__338_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_4__401_ (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_0_BUFX2_insert12 (
);

FILL FILL_0_BUFX2_insert13 (
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

FILL FILL_0_BUFX2_insert16 (
);

FILL FILL_0_BUFX2_insert17 (
);

FILL FILL_7__545_ (
);

FILL FILL_0_BUFX2_insert18 (
);

FILL FILL_0__487_ (
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL_2__481_ (
);

FILL FILL_3__423_ (
);

FILL FILL_6__567_ (
);

FILL FILL_7__354_ (
);

FILL FILL_2__537_ (
);

FILL FILL_6__376_ (
);

INVX1 _511_ (
    .A(Atmp[5]),
    .Y(_55_)
);

FILL FILL_7__583_ (
);

FILL FILL_1__559_ (
);

FILL FILL_8__525_ (
);

FILL FILL_2__346_ (
);

FILL FILL_8_CLKBUF1_insert0 (
);

FILL FILL_8_CLKBUF1_insert1 (
);

FILL FILL_8_CLKBUF1_insert3 (
);

FILL FILL_8_CLKBUF1_insert4 (
);

FILL FILL_8_CLKBUF1_insert5 (
);

FILL FILL_3__461_ (
);

OR2X2 _320_ (
    .A(_156_),
    .B(_159_),
    .Y(_160_)
);

BUFX2 BUFX2_insert20 (
    .A(_73_),
    .Y(_73__bF$buf0)
);

FILL FILL_7__392_ (
);

FILL FILL_1__368_ (
);

FILL FILL_2__575_ (
);

FILL FILL_3__517_ (
);

FILL FILL75150x39750 (
);

FILL FILL_7__448_ (
);

FILL FILL_5__511_ (
);

FILL FILL_1__597_ (
);

FILL FILL_8__563_ (
);

FILL FILL_2__384_ (
);

FILL FILL_0__602_ (
);

FILL FILL_3__326_ (
);

INVX1 _605_ (
    .A(_130_),
    .Y(_134_)
);

FILL FILL_4__533_ (
);

FILL FILL_8__619_ (
);

FILL FILL_5__320_ (
);

FILL FILL_8__372_ (
);

FILL FILL_0__411_ (
);

FILL FILL_3__555_ (
);

AOI21X1 _414_ (
    .A(_235_),
    .B(_221_),
    .C(_230_),
    .Y(_246_)
);

FILL FILL_4__342_ (
);

FILL FILL_7__486_ (
);

FILL FILL_3__364_ (
);

DFFPOSX1 _643_ (
    .D(_17_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[10])
);

FILL FILL_4__571_ (
);

FILL FILL_5__605_ (
);

FILL FILL_2__478_ (
);

FILL FILL_3__593_ (
);

AOI21X1 _452_ (
    .A(_249_),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

FILL FILL_4__380_ (
);

FILL FILL_5__414_ (
);

FILL FILL_8__466_ (
);

FILL FILL_0__505_ (
);

OAI21X1 _508_ (
    .A(RdyCtl[1]),
    .B(_50_),
    .C(_52_),
    .Y(_53_)
);

FILL FILL_4__436_ (
);

FILL FILL_0__314_ (
);

FILL FILL_3__458_ (
);

NAND2X1 _317_ (
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_157_)
);

FILL FILL_1__521_ (
);

FILL FILL_4__665_ (
);

FILL FILL_7__389_ (
);

AOI21X1 _490_ (
    .A(_56_),
    .B(_73__bF$buf3),
    .C(_308_),
    .Y(_36_)
);

FILL FILL_5__452_ (
);

FILL FILL74550x50550 (
);

FILL FILL_7__601_ (
);

FILL FILL_0__543_ (
);

INVX1 _546_ (
    .A(_79_),
    .Y(_80_)
);

FILL FILL_1__330_ (
);

FILL FILL_4__474_ (
);

FILL FILL_5__508_ (
);

FILL FILL_6__623_ (
);

FILL FILL_7__410_ (
);

FILL FILL_0__352_ (
);

FILL FILL_3__496_ (
);

OR2X2 _355_ (
    .A(_187_),
    .B(_191_),
    .Y(_192_)
);

FILL FILL_5__317_ (
);

FILL FILL_8__369_ (
);

FILL FILL_5__490_ (
);

FILL FILL_6__432_ (
);

FILL FILL_0__408_ (
);

FILL FILL_0__581_ (
);

FILL FILL_1__615_ (
);

FILL FILL_4__339_ (
);

OAI21X1 _584_ (
    .A(acc_reg[4]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_115_)
);

FILL FILL_2__402_ (
);

FILL FILL_5__546_ (
);

FILL FILL_8__598_ (
);

FILL FILL_0__390_ (
);

FILL FILL_1__424_ (
);

FILL FILL_4__568_ (
);

OAI21X1 _393_ (
    .A(acc_reg[14]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf3),
    .Y(_227_)
);

FILL FILL_5__355_ (
);

FILL FILL_6__470_ (
);

FILL FILL_7__504_ (
);

FILL FILL_0__446_ (
);

NAND2X1 _449_ (
    .A(_278_),
    .B(_274_),
    .Y(_279_)
);

FILL FILL_4__377_ (
);

FILL FILL_2__440_ (
);

FILL FILL_5__584_ (
);

FILL FILL_6__526_ (
);

FILL FILL_7__313_ (
);

FILL FILL_3__399_ (
);

FILL FILL_1__462_ (
);

FILL FILL_5__393_ (
);

FILL FILL_3__611_ (
);

FILL FILL_6__335_ (
);

FILL FILL_7__542_ (
);

FILL FILL_0__484_ (
);

FILL FILL_1__518_ (
);

OAI21X1 _487_ (
    .A(acc_reg[16]),
    .B(_73__bF$buf3),
    .C(En_bF$buf1),
    .Y(_307_)
);

FILL FILL_5__449_ (
);

FILL FILL_3__420_ (
);

FILL FILL_6__564_ (
);

FILL FILL_7__351_ (
);

FILL FILL_1__327_ (
);

FILL FILL_2__534_ (
);

FILL FILL_6__373_ (
);

FILL FILL74850x25350 (
);

FILL FILL_7__407_ (
);

FILL FILL_0__349_ (
);

FILL FILL_7__580_ (
);

FILL FILL_1__556_ (
);

FILL FILL_2__343_ (
);

FILL FILL_5__487_ (
);

FILL FILL_6__429_ (
);

FILL FILL_0__578_ (
);

FILL FILL_1__365_ (
);

FILL FILL_8__331_ (
);

FILL FILL_2__572_ (
);

FILL FILL_3__514_ (
);

FILL FILL_7__445_ (
);

FILL FILL_0__387_ (
);

FILL FILL_1__594_ (
);

FILL FILL_8__560_ (
);

FILL FILL_2__381_ (
);

FILL FILL_3__323_ (
);

FILL FILL_6__467_ (
);

NAND2X1 _602_ (
    .A(_129_),
    .B(_130_),
    .Y(_131_)
);

FILL FILL_4__530_ (
);

FILL FILL_8__616_ (
);

FILL FILL_2__437_ (
);

FILL FILL73650x57750 (
);

FILL FILL_3__552_ (
);

NOR2X1 _411_ (
    .A(_223_),
    .B(_236_),
    .Y(_243_)
);

FILL FILL_7__483_ (
);

FILL FILL_1__459_ (
);

FILL FILL_8__425_ (
);

FILL FILL_2__666_ (
);

FILL FILL_3__608_ (
);

FILL FILL_3__361_ (
);

FILL FILL_7__539_ (
);

DFFPOSX1 _640_ (
    .D(_14_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[7])
);

FILL FILL_5__602_ (
);

FILL FILL_2__475_ (
);

FILL FILL_3__417_ (
);

FILL FILL_3__590_ (
);

FILL FILL_4__624_ (
);

FILL FILL_7__348_ (
);

FILL FILL_5__411_ (
);

FILL FILL_1__497_ (
);

FILL FILL_8__463_ (
);

FILL FILL_0__502_ (
);

OAI21X1 _505_ (
    .A(_39_),
    .B(_40_),
    .C(_49_),
    .Y(_50_)
);

FILL FILL_4__433_ (
);

FILL FILL_7__577_ (
);

FILL FILL_8__519_ (
);

FILL FILL73950x10950 (
);

FILL FILL75150x25350 (
);

FILL FILL_3__455_ (
);

FILL FILL_6__599_ (
);

INVX1 _314_ (
    .A(_153_),
    .Y(_154_)
);

FILL FILL_7__386_ (
);

FILL FILL_8__328_ (
);

FILL FILL_2__569_ (
);

FILL FILL_0__540_ (
);

AOI21X1 _543_ (
    .A(_75_),
    .B(_76_),
    .C(_77_),
    .Y(_7_)
);

FILL FILL_4__471_ (
);

FILL FILL_5__505_ (
);

FILL FILL_8__557_ (
);

FILL FILL_6__620_ (
);

FILL FILL_2__378_ (
);

FILL FILL_3__493_ (
);

FILL FILL_4__527_ (
);

NOR2X1 _352_ (
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_189_)
);

FILL FILL_5__314_ (
);

FILL FILL_8__366_ (
);

FILL FILL75450x68550 (
);

FILL FILL_0__405_ (
);

FILL FILL_3__549_ (
);

NAND3X1 _408_ (
    .A(_239_),
    .B(_232_),
    .C(_217_),
    .Y(_240_)
);

FILL FILL_1__612_ (
);

FILL FILL_4__336_ (
);

NOR2X1 _581_ (
    .A(_109_),
    .B(_108_),
    .Y(_112_)
);

FILL FILL_5__543_ (
);

FILL FILL_8__595_ (
);

FILL FILL_3__358_ (
);

DFFPOSX1 _637_ (
    .D(_11_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[4])
);

FILL FILL_1__421_ (
);

FILL FILL_4__565_ (
);

OR2X2 _390_ (
    .A(_220_),
    .B(_223_),
    .Y(_224_)
);

FILL FILL_5__352_ (
);

FILL FILL_7__501_ (
);

FILL FILL_0__443_ (
);

FILL FILL_3__587_ (
);

NOR2X1 _446_ (
    .A(_68_),
    .B(_275_),
    .Y(_276_)
);

FILL FILL_4__374_ (
);

FILL FILL_5__408_ (
);

FILL FILL_5__581_ (
);

FILL FILL_6__523_ (
);

FILL FILL75750x21750 (
);

FILL FILL_3__396_ (
);

FILL FILL_5__390_ (
);

FILL FILL_6__332_ (
);

FILL FILL_0__481_ (
);

FILL FILL_1__515_ (
);

AOI21X1 _484_ (
    .A(_41_),
    .B(_73__bF$buf0),
    .C(_305_),
    .Y(_33_)
);

FILL FILL_5__446_ (
);

FILL FILL_6__561_ (
);

FILL FILL_0__537_ (
);

FILL FILL_1__324_ (
);

FILL FILL_4__468_ (
);

FILL FILL_2__531_ (
);

FILL FILL_6__617_ (
);

FILL FILL_6__370_ (
);

FILL FILL_7__404_ (
);

FILL FILL_0__346_ (
);

NAND2X1 _349_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_186_)
);

FILL FILL_1__553_ (
);

FILL FILL_2__340_ (
);

FILL FILL_5__484_ (
);

FILL FILL_6__426_ (
);

FILL FILL_0__575_ (
);

FILL FILL_1__609_ (
);

NOR2X1 _578_ (
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_109_)
);

FILL FILL_1__362_ (
);

FILL FILL_3__511_ (
);

FILL FILL_7__442_ (
);

FILL FILL_0__384_ (
);

FILL FILL_1__418_ (
);

AND2X2 _387_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_221_)
);

FILL FILL_1__591_ (
);

FILL FILL_2__625_ (
);

FILL FILL_5__349_ (
);

FILL FILL_3__320_ (
);

FILL FILL_6__464_ (
);

FILL FILL_8__613_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_2__434_ (
);

FILL FILL_5__578_ (
);

FILL FILL_7__480_ (
);

FILL FILL_1__456_ (
);

FILL FILL_8__422_ (
);

FILL FILL_6_CLKBUF1_insert0 (
);

FILL FILL_6_CLKBUF1_insert1 (
);

FILL FILL_6_CLKBUF1_insert2 (
);

FILL FILL_6_CLKBUF1_insert3 (
);

FILL FILL_6_CLKBUF1_insert4 (
);

FILL FILL_6_CLKBUF1_insert5 (
);

FILL FILL_5__387_ (
);

FILL FILL_3__605_ (
);

FILL FILL_6__329_ (
);

FILL FILL_7__536_ (
);

FILL FILL_0__478_ (
);

FILL FILL_2__472_ (
);

FILL FILL_3__414_ (
);

FILL FILL_6__558_ (
);

FILL FILL_4__621_ (
);

FILL FILL_7__345_ (
);

FILL FILL_1__494_ (
);

FILL FILL_8__460_ (
);

FILL FILL_2__528_ (
);

FILL FILL_6__367_ (
);

NAND2X1 _502_ (
    .A(_42_),
    .B(_46_),
    .Y(_47_)
);

FILL FILL_4__430_ (
);

FILL FILL_7__574_ (
);

FILL FILL_8__516_ (
);

FILL FILL_2__337_ (
);

FILL FILL_3__452_ (
);

FILL FILL_6__596_ (
);

FILL FILL_7__383_ (
);

FILL FILL_1__359_ (
);

FILL FILL_8__325_ (
);

FILL FILL_2__566_ (
);

FILL FILL_3__508_ (
);

FILL FILL_6_BUFX2_insert20 (
);

FILL FILL_7__439_ (
);

INVX1 _540_ (
    .A(acc_reg[0]),
    .Y(_75_)
);

FILL FILL_5__502_ (
);

FILL FILL_1__588_ (
);

FILL FILL_2__375_ (
);

FILL FILL_3__317_ (
);

FILL FILL_3__490_ (
);

FILL FILL_4__524_ (
);

FILL FILL_7__668_ (
);

FILL FILL_1__397_ (
);

FILL FILL_8__363_ (
);

FILL FILL_0__402_ (
);

FILL FILL_3__546_ (
);

OAI21X1 _405_ (
    .A(acc_reg[15]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf3),
    .Y(_238_)
);

FILL FILL_4__333_ (
);

FILL FILL_7__477_ (
);

FILL FILL_8__419_ (
);

FILL FILL_5__540_ (
);

FILL FILL_3__355_ (
);

FILL FILL_6__499_ (
);

DFFPOSX1 _634_ (
    .D(_8_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[1])
);

FILL FILL_4__562_ (
);

FILL FILL_2__469_ (
);

FILL FILL_0__440_ (
);

FILL FILL_3__584_ (
);

FILL FILL_4__618_ (
);

AOI21X1 _443_ (
    .A(_268_),
    .B(_250_),
    .C(_266_),
    .Y(_273_)
);

FILL FILL_4__371_ (
);

FILL FILL_5__405_ (
);

FILL FILL_8__457_ (
);

FILL FILL_6__520_ (
);

FILL FILL_3__393_ (
);

FILL FILL_4__427_ (
);

FILL FILL_3__449_ (
);

FILL FILL_1__512_ (
);

OAI21X1 _481_ (
    .A(acc_reg[13]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_304_)
);

FILL FILL_5__443_ (
);

FILL FILL_8__495_ (
);

FILL FILL_0__534_ (
);

NOR2X1 _537_ (
    .A(_42_),
    .B(_74_),
    .Y(_4_)
);

FILL FILL75450x54150 (
);

FILL FILL_1__321_ (
);

FILL FILL_4__465_ (
);

FILL FILL_6__614_ (
);

FILL FILL74250x36150 (
);

FILL FILL_7__401_ (
);

FILL FILL_0__343_ (
);

FILL FILL_3__487_ (
);

NAND2X1 _346_ (
    .A(_182_),
    .B(_183_),
    .Y(_184_)
);

FILL FILL_1__550_ (
);

FILL FILL_5__481_ (
);

FILL FILL_6__423_ (
);

FILL FILL73950x18150 (
);

FILL FILL_0__572_ (
);

FILL FILL_1__606_ (
);

AOI21X1 _575_ (
    .A(_105_),
    .B(_89_),
    .C(_97_),
    .Y(_106_)
);

FILL FILL_5__537_ (
);

FILL FILL_8__589_ (
);

FILL FILL_0__381_ (
);

FILL FILL_1__415_ (
);

FILL FILL_4__559_ (
);

NOR2X1 _384_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_218_)
);

FILL FILL_2__622_ (
);

FILL FILL_5__346_ (
);

FILL FILL_8__398_ (
);

FILL FILL_6__461_ (
);

FILL FILL_0__437_ (
);

FILL FILL_8__610_ (
);

FILL FILL_4__368_ (
);

FILL FILL_2__431_ (
);

FILL FILL_5__575_ (
);

FILL FILL_6__517_ (
);

FILL FILL_0__666_ (
);

FILL FILL_1__453_ (
);

FILL FILL_4__597_ (
);

FILL FILL_5__384_ (
);

FILL FILL_3__602_ (
);

FILL FILL_6__326_ (
);

FILL FILL_7__533_ (
);

FILL FILL_0__475_ (
);

FILL FILL_1__509_ (
);

AOI21X1 _478_ (
    .A(_62_),
    .B(_73__bF$buf3),
    .C(_302_),
    .Y(_30_)
);

FILL FILL_3__411_ (
);

FILL FILL_6__555_ (
);

FILL FILL_7__342_ (
);

FILL FILL_1__318_ (
);

FILL FILL_1__491_ (
);

FILL FILL_2__525_ (
);

FILL FILL_6__364_ (
);

FILL FILL_7__571_ (
);

FILL FILL_1__547_ (
);

FILL FILL_8__513_ (
);

FILL FILL_2__334_ (
);

FILL FILL_5__478_ (
);

FILL FILL_6__593_ (
);

FILL FILL_0__569_ (
);

FILL FILL_7__380_ (
);

FILL FILL_1__356_ (
);

FILL FILL_8__322_ (
);

FILL FILL_2__563_ (
);

FILL FILL_3__505_ (
);

FILL FILL_7__436_ (
);

FILL FILL_0__378_ (
);

FILL FILL_1__585_ (
);

FILL FILL_8__551_ (
);

FILL FILL_2__619_ (
);

FILL FILL_2__372_ (
);

FILL FILL_3__314_ (
);

FILL FILL_6__458_ (
);

FILL FILL_4__521_ (
);

FILL FILL_7__665_ (
);

FILL FILL_8__607_ (
);

FILL FILL_1__394_ (
);

FILL FILL_8__360_ (
);

FILL FILL_2__428_ (
);

FILL FILL_3__543_ (
);

INVX1 _402_ (
    .A(_231_),
    .Y(_235_)
);

FILL FILL_4__330_ (
);

FILL FILL_7__474_ (
);

FILL FILL_8__416_ (
);

FILL FILL_3__352_ (
);

FILL FILL_6__496_ (
);

DFFPOSX1 _631_ (
    .D(_5_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[5])
);

FILL FILL_2__466_ (
);

FILL FILL_3__408_ (
);

FILL FILL_3__581_ (
);

FILL FILL_4__615_ (
);

FILL FILL_7__339_ (
);

OAI21X1 _440_ (
    .A(acc_reg[17]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_271_)
);

FILL FILL_5__402_ (
);

FILL FILL_1__488_ (
);

FILL FILL_8__454_ (
);

FILL FILL_3__390_ (
);

FILL FILL_4__424_ (
);

FILL FILL_7__568_ (
);

FILL FILL_3__446_ (
);

FILL FILL_7__377_ (
);

FILL FILL_8__319_ (
);

FILL FILL_5__440_ (
);

FILL FILL_8__492_ (
);

FILL FILL_0__531_ (
);

FILL FILL_6__399_ (
);

AND2X2 _534_ (
    .A(RdyCtl[0]),
    .B(En_bF$buf2),
    .Y(_1_)
);

FILL FILL_4__462_ (
);

FILL FILL_8__548_ (
);

FILL FILL_6__611_ (
);

FILL FILL_2__369_ (
);

FILL FILL_0__340_ (
);

FILL FILL_3__484_ (
);

FILL FILL_4__518_ (
);

NOR2X1 _343_ (
    .A(_180_),
    .B(_179_),
    .Y(_181_)
);

FILL FILL74250x57750 (
);

FILL FILL_6__420_ (
);

FILL FILL_2__598_ (
);

FILL FILL_1__603_ (
);

FILL FILL_4__327_ (
);

AOI21X1 _572_ (
    .A(_103_),
    .B(RdyCtl_6_bF$buf4),
    .C(_96_),
    .Y(_10_)
);

FILL FILL_5__534_ (
);

FILL FILL73950x39750 (
);

FILL FILL_8__586_ (
);

FILL FILL_0__625_ (
);

FILL FILL_3__349_ (
);

DFFPOSX1 _628_ (
    .D(_2_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[2])
);

FILL FILL_1__412_ (
);

FILL FILL_4__556_ (
);

OAI21X1 _381_ (
    .A(acc_reg[13]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf4),
    .Y(_216_)
);

FILL FILL_5__343_ (
);

FILL FILL_0__434_ (
);

FILL FILL_3__578_ (
);

NOR2X1 _437_ (
    .A(_267_),
    .B(_266_),
    .Y(_268_)
);

FILL FILL_4__365_ (
);

FILL FILL_5__572_ (
);

FILL FILL_6__514_ (
);

FILL FILL74550x10950 (
);

FILL FILL_3__387_ (
);

BUFX2 _666_ (
    .A(_311_[1]),
    .Y(Aout[1])
);

FILL FILL_1__450_ (
);

FILL FILL_4__594_ (
);

FILL FILL_5__381_ (
);

FILL FILL_6__323_ (
);

FILL FILL_7__530_ (
);

FILL FILL_0__472_ (
);

FILL FILL_1__506_ (
);

OAI21X1 _475_ (
    .A(acc_reg[10]),
    .B(_73__bF$buf2),
    .C(En_bF$buf2),
    .Y(_301_)
);

FILL FILL_5__437_ (
);

FILL FILL_6__552_ (
);

FILL FILL_0__528_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_2_BUFX2_insert12 (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_2_BUFX2_insert17 (
);

FILL FILL_2_BUFX2_insert18 (
);

FILL FILL_2_BUFX2_insert19 (
);

FILL FILL_1__315_ (
);

FILL FILL_4__459_ (
);

FILL FILL_2__522_ (
);

FILL FILL_5__666_ (
);

FILL FILL_6__608_ (
);

FILL FILL_6__361_ (
);

FILL FILL_0__337_ (
);

FILL FILL76050x68550 (
);

FILL FILL_1__544_ (
);

FILL FILL_8__510_ (
);

FILL FILL_2__331_ (
);

FILL FILL_5__475_ (
);

FILL FILL_6__417_ (
);

FILL FILL_6__590_ (
);

FILL FILL_7__624_ (
);

FILL FILL_0__566_ (
);

NOR2X1 _569_ (
    .A(_89_),
    .B(_92_),
    .Y(_101_)
);

FILL FILL_1__353_ (
);

FILL FILL_4__497_ (
);

FILL FILL_4_CLKBUF1_insert0 (
);

FILL FILL_4_CLKBUF1_insert1 (
);

FILL FILL_4_CLKBUF1_insert2 (
);

FILL FILL_4_CLKBUF1_insert3 (
);

FILL FILL_4_CLKBUF1_insert4 (
);

FILL FILL_4_CLKBUF1_insert5 (
);

FILL FILL_2__560_ (
);

FILL FILL_3__502_ (
);

FILL FILL_7__433_ (
);

FILL FILL_0__375_ (
);

FILL FILL_1__409_ (
);

NAND2X1 _378_ (
    .A(_211_),
    .B(_212_),
    .Y(_213_)
);

FILL FILL_1__582_ (
);

FILL FILL_2__616_ (
);

FILL FILL_6__455_ (
);

FILL FILL_8__604_ (
);

FILL FILL_1__391_ (
);

FILL FILL_2__425_ (
);

FILL FILL_5__569_ (
);

FILL FILL_3__540_ (
);

FILL FILL_7__471_ (
);

FILL FILL_1__447_ (
);

FILL FILL_8__413_ (
);

FILL FILL_5__378_ (
);

FILL FILL_6__493_ (
);

FILL FILL_7__527_ (
);

FILL FILL_0__469_ (
);

FILL FILL_2__463_ (
);

FILL FILL_3__405_ (
);

FILL FILL_6__549_ (
);

FILL FILL_4__612_ (
);

FILL FILL_7__336_ (
);

FILL FILL_1__485_ (
);

FILL FILL_2__519_ (
);

FILL FILL_6__358_ (
);

FILL FILL_4__421_ (
);

FILL FILL_7__565_ (
);

FILL FILL_2__328_ (
);

FILL FILL_3__443_ (
);

FILL FILL_6__587_ (
);

FILL FILL_7__374_ (
);

FILL FILL_8__316_ (
);

FILL FILL_2__557_ (
);

FILL FILL73650x50550 (
);

FILL FILL_6__396_ (
);

INVX8 _531_ (
    .A(RdyCtl_6_bF$buf0),
    .Y(_73_)
);

FILL FILL_1__579_ (
);

FILL FILL_2__366_ (
);

FILL FILL_3__481_ (
);

FILL FILL_4__515_ (
);

OAI21X1 _340_ (
    .A(_177_),
    .B(_156_),
    .C(_176_),
    .Y(_178_)
);

FILL FILL_1__388_ (
);

FILL FILL_8__354_ (
);

FILL FILL_2__595_ (
);

FILL FILL_3__537_ (
);

FILL FILL_1__600_ (
);

FILL FILL_4__324_ (
);

FILL FILL_7__468_ (
);

FILL FILL_5__531_ (
);

FILL FILL_0__622_ (
);

FILL FILL_3__346_ (
);

AOI21X1 _625_ (
    .A(_151_),
    .B(_108_),
    .C(_117_),
    .Y(_152_)
);

FILL FILL_4__553_ (
);

FILL FILL_5__340_ (
);

FILL FILL_8__392_ (
);

FILL FILL_0__431_ (
);

FILL FILL_3__575_ (
);

FILL FILL_4__609_ (
);

AOI21X1 _434_ (
    .A(_249_),
    .B(_252_),
    .C(_250_),
    .Y(_265_)
);

FILL FILL_4__362_ (
);

FILL FILL_8__448_ (
);

FILL FILL_6__511_ (
);

FILL FILL_3__384_ (
);

FILL FILL_4__418_ (
);

DFFPOSX1 _663_ (
    .D(_37_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[11])
);

FILL FILL_4__591_ (
);

FILL FILL_5__625_ (
);

FILL FILL_6__320_ (
);

FILL FILL_2__498_ (
);

FILL FILL_1__503_ (
);

NOR2X1 _472_ (
    .A(Atmp[1]),
    .B(RdyCtl_6_bF$buf0),
    .Y(_299_)
);

FILL FILL_5__434_ (
);

FILL FILL_8__486_ (
);

FILL FILL75450x61350 (
);

FILL FILL75450x28950 (
);

FILL FILL_0__525_ (
);

NAND2X1 _528_ (
    .A(_67_),
    .B(_70_),
    .Y(_71_)
);

FILL FILL_4__456_ (
);

FILL FILL_6__605_ (
);

FILL FILL_0__334_ (
);

FILL FILL_3__478_ (
);

OAI21X1 _337_ (
    .A(_157_),
    .B(_174_),
    .C(_165_),
    .Y(_175_)
);

FILL FILL73950x25350 (
);

FILL FILL_1__541_ (
);

FILL FILL_5__472_ (
);

FILL FILL_6__414_ (
);

FILL FILL_7__621_ (
);

FILL FILL_0__563_ (
);

NOR2X1 _566_ (
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_98_)
);

FILL FILL_1__350_ (
);

FILL FILL_4__494_ (
);

FILL FILL_5__528_ (
);

FILL FILL_0__619_ (
);

FILL FILL_7__430_ (
);

FILL FILL_0__372_ (
);

FILL FILL_1__406_ (
);

OAI21X1 _375_ (
    .A(_205_),
    .B(_209_),
    .C(_203_),
    .Y(_210_)
);

FILL FILL_2__613_ (
);

FILL FILL_5__337_ (
);

FILL FILL_8__389_ (
);

FILL FILL_6__452_ (
);

FILL FILL_0__428_ (
);

FILL FILL_4__359_ (
);

FILL FILL_2__422_ (
);

FILL FILL_5__566_ (
);

FILL FILL_6__508_ (
);

FILL FILL_1__444_ (
);

FILL FILL_8__410_ (
);

FILL FILL_4__588_ (
);

FILL FILL_5__375_ (
);

FILL FILL_6__317_ (
);

FILL FILL_6__490_ (
);

FILL FILL_7__524_ (
);

FILL FILL_0__466_ (
);

NOR2X1 _469_ (
    .A(Atmp[0]),
    .B(RdyCtl_6_bF$buf0),
    .Y(_297_)
);

FILL FILL_4__397_ (
);

FILL FILL_2__460_ (
);

FILL FILL_3__402_ (
);

FILL FILL_6__546_ (
);

FILL FILL76050x54150 (
);

FILL FILL_7__333_ (
);

FILL FILL_1__482_ (
);

FILL FILL_2__516_ (
);

FILL FILL75750x36150 (
);

FILL FILL_6__355_ (
);

FILL FILL_7__562_ (
);

FILL FILL_1__538_ (
);

FILL FILL_8__504_ (
);

FILL FILL74550x18150 (
);

FILL FILL_2__325_ (
);

FILL FILL_5__469_ (
);

FILL FILL_3__440_ (
);

FILL FILL_6__584_ (
);

FILL FILL_7__618_ (
);

FILL FILL_7__371_ (
);

FILL FILL_1__347_ (
);

FILL FILL_8__313_ (
);

FILL FILL_2__554_ (
);

FILL FILL_6__393_ (
);

FILL FILL_7__427_ (
);

FILL FILL_0__369_ (
);

FILL FILL_1__576_ (
);

FILL FILL_8__542_ (
);

FILL FILL_2__363_ (
);

FILL FILL_6__449_ (
);

FILL FILL_4__512_ (
);

FILL FILL_0__598_ (
);

FILL FILL_1__385_ (
);

FILL FILL_8__351_ (
);

FILL FILL_2__419_ (
);

FILL FILL_2__592_ (
);

FILL FILL_3__534_ (
);

FILL FILL_4__321_ (
);

FILL FILL_7__465_ (
);

FILL FILL_8__407_ (
);

FILL FILL_8__580_ (
);

FILL FILL_3__343_ (
);

FILL FILL_6__487_ (
);

NAND3X1 _622_ (
    .A(_129_),
    .B(_130_),
    .C(_148_),
    .Y(_149_)
);

FILL FILL_4__550_ (
);

FILL FILL_2__457_ (
);

FILL FILL_3__572_ (
);

FILL FILL_4__606_ (
);

NAND2X1 _431_ (
    .A(_262_),
    .B(_253_),
    .Y(_263_)
);

FILL FILL_1__479_ (
);

FILL FILL_8__445_ (
);

FILL FILL_3__381_ (
);

FILL FILL_4__415_ (
);

FILL FILL_7__559_ (
);

DFFPOSX1 _660_ (
    .D(_34_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[7])
);

FILL FILL_5__622_ (
);

FILL FILL_2__495_ (
);

FILL FILL_3__437_ (
);

FILL FILL_1__500_ (
);

FILL FILL_7__368_ (
);

FILL FILL_5__431_ (
);

FILL FILL_8__483_ (
);

FILL FILL_0__522_ (
);

FILL FILL_3__666_ (
);

INVX1 _525_ (
    .A(acc_reg[18]),
    .Y(_68_)
);

FILL FILL_4__453_ (
);

FILL FILL_7__597_ (
);

FILL FILL_8__539_ (
);

FILL FILL_6__602_ (
);

FILL FILL_0__331_ (
);

FILL FILL_3__475_ (
);

FILL FILL_4__509_ (
);

OAI21X1 _334_ (
    .A(acc_reg[9]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_173_)
);

FILL FILL_6__411_ (
);

FILL FILL_2__589_ (
);

FILL FILL_0__560_ (
);

FILL FILL_4__318_ (
);

AOI21X1 _563_ (
    .A(_94_),
    .B(_95_),
    .C(_74_),
    .Y(_9_)
);

FILL FILL_4__491_ (
);

FILL FILL_5__525_ (
);

FILL FILL_8__577_ (
);

FILL FILL_2__398_ (
);

FILL FILL_0__616_ (
);

AND2X2 _619_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_146_)
);

FILL FILL_1__403_ (
);

FILL FILL_4__547_ (
);

OAI21X1 _372_ (
    .A(_206_),
    .B(_207_),
    .C(RdyCtl_6_bF$buf2),
    .Y(_208_)
);

FILL FILL_2__610_ (
);

FILL FILL_5__334_ (
);

FILL FILL_8__386_ (
);

FILL FILL_0__425_ (
);

FILL FILL_3__569_ (
);

OAI21X1 _428_ (
    .A(_240_),
    .B(_201_),
    .C(_259_),
    .Y(_260_)
);

FILL FILL_4__356_ (
);

FILL FILL_5__563_ (
);

FILL FILL_6__505_ (
);

FILL FILL_3__378_ (
);

DFFPOSX1 _657_ (
    .D(_31_),
    .CLK(clk_bF$buf2),
    .Q(Atmp[4])
);

FILL FILL_1__441_ (
);

FILL FILL_4__585_ (
);

FILL FILL_5__619_ (
);

FILL FILL75450x14550 (
);

FILL FILL_3_BUFX2_insert20 (
);

FILL FILL_5__372_ (
);

FILL FILL_6__314_ (
);

FILL FILL_7__521_ (
);

FILL FILL_0__463_ (
);

INVX1 _466_ (
    .A(_292_),
    .Y(_295_)
);

FILL FILL_2_CLKBUF1_insert0 (
);

FILL FILL_2_CLKBUF1_insert1 (
);

FILL FILL_2_CLKBUF1_insert2 (
);

FILL FILL_2_CLKBUF1_insert3 (
);

FILL FILL_2_CLKBUF1_insert4 (
);

FILL FILL_2_CLKBUF1_insert5 (
);

FILL FILL_4__394_ (
);

FILL FILL_5__428_ (
);

FILL FILL_6__543_ (
);

FILL FILL_0__519_ (
);

FILL FILL_7__330_ (
);

FILL FILL_2__513_ (
);

FILL FILL_6__352_ (
);

FILL FILL_0__328_ (
);

FILL FILL_1__535_ (
);

FILL FILL_8__501_ (
);

FILL FILL75750x57750 (
);

FILL FILL_2__322_ (
);

FILL FILL_5__466_ (
);

FILL FILL_6__408_ (
);

FILL FILL_6__581_ (
);

FILL FILL_7__615_ (
);

FILL FILL_0__557_ (
);

FILL FILL74550x39750 (
);

FILL FILL_1__344_ (
);

FILL FILL_4__488_ (
);

FILL FILL_2__551_ (
);

FILL FILL_6__390_ (
);

FILL FILL_7__424_ (
);

FILL FILL_0__366_ (
);

NAND2X1 _369_ (
    .A(_203_),
    .B(_204_),
    .Y(_205_)
);

FILL FILL_1__573_ (
);

FILL FILL_2__607_ (
);

FILL FILL_2__360_ (
);

FILL FILL_6__446_ (
);

FILL FILL_8_BUFX2_insert20 (
);

FILL FILL_0__595_ (
);

AND2X2 _598_ (
    .A(_112_),
    .B(_119_),
    .Y(_127_)
);

FILL FILL_1__382_ (
);

FILL FILL_2__416_ (
);

FILL FILL_3__531_ (
);

FILL FILL_7__462_ (
);

FILL FILL_1__438_ (
);

FILL FILL_5__369_ (
);

FILL FILL_3__340_ (
);

FILL FILL_6__484_ (
);

FILL FILL_7__518_ (
);

FILL FILL_1__667_ (
);

FILL FILL_2__454_ (
);

FILL FILL_5__598_ (
);

FILL FILL_4__603_ (
);

FILL FILL_7__327_ (
);

FILL FILL_1__476_ (
);

FILL FILL_3__625_ (
);

FILL FILL_6__349_ (
);

FILL FILL_4__412_ (
);

FILL FILL_7__556_ (
);

FILL FILL_0__498_ (
);

FILL FILL_2__319_ (
);

FILL FILL_2__492_ (
);

FILL FILL_3__434_ (
);

FILL FILL_6__578_ (
);

FILL FILL_7__365_ (
);

FILL FILL_8__480_ (
);

FILL FILL_2__548_ (
);

FILL FILL_6__387_ (
);

OAI21X1 _522_ (
    .A(RdyCtl[0]),
    .B(_64_),
    .C(_65_),
    .Y(_311_[1])
);

FILL FILL_4__450_ (
);

FILL FILL_7__594_ (
);

FILL FILL_2__357_ (
);

FILL FILL_3__472_ (
);

FILL FILL_4__506_ (
);

NAND2X1 _331_ (
    .A(_169_),
    .B(_164_),
    .Y(_170_)
);

FILL FILL_1__379_ (
);

FILL FILL_8__345_ (
);

FILL FILL_2__586_ (
);

FILL FILL_3__528_ (
);

FILL FILL_4__315_ (
);

FILL FILL_7__459_ (
);

NOR2X1 _560_ (
    .A(_73__bF$buf0),
    .B(_92_),
    .Y(_93_)
);

FILL FILL_5__522_ (
);

FILL FILL_8__574_ (
);

FILL FILL_2__395_ (
);

FILL FILL_0__613_ (
);

FILL FILL_3__337_ (
);

OAI21X1 _616_ (
    .A(acc_reg[7]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_144_)
);

FILL FILL_1__400_ (
);

FILL FILL_4__544_ (
);

FILL FILL_5__331_ (
);

FILL FILL_8__383_ (
);

FILL FILL_0__422_ (
);

FILL FILL_3__566_ (
);

OAI21X1 _425_ (
    .A(_255_),
    .B(_107_),
    .C(_256_),
    .Y(_257_)
);

FILL FILL_4__353_ (
);

FILL FILL_7__497_ (
);

FILL FILL_8__439_ (
);

FILL FILL_5__560_ (
);

FILL FILL_6__502_ (
);

FILL FILL_3__375_ (
);

FILL FILL_4__409_ (
);

DFFPOSX1 _654_ (
    .D(_28_),
    .CLK(clk_bF$buf4),
    .Q(Atmp[1])
);

FILL FILL_4__582_ (
);

FILL FILL_5__616_ (
);

FILL FILL_2__489_ (
);

FILL FILL_0__460_ (
);

NAND2X1 _463_ (
    .A(_290_),
    .B(_291_),
    .Y(_292_)
);

FILL FILL_4__391_ (
);

FILL FILL_5__425_ (
);

FILL FILL_8__477_ (
);

FILL FILL74250x50550 (
);

FILL FILL_6__540_ (
);

FILL FILL_0__516_ (
);

NAND2X1 _519_ (
    .A(RdyCtl[1]),
    .B(_62_),
    .Y(_63_)
);

FILL FILL_4__447_ (
);

FILL FILL_2__510_ (
);

FILL FILL_0__325_ (
);

FILL FILL_3__469_ (
);

INVX1 _328_ (
    .A(FCW[9]),
    .Y(_167_)
);

FILL FILL_1__532_ (
);

FILL FILL_5__463_ (
);

FILL FILL_6__405_ (
);

FILL FILL_7__612_ (
);

FILL FILL_0__554_ (
);

NOR2X1 _557_ (
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_90_)
);

FILL FILL_1__341_ (
);

FILL FILL_4__485_ (
);

FILL FILL_5__519_ (
);

FILL FILL_7__421_ (
);

FILL FILL_0__363_ (
);

OAI21X1 _366_ (
    .A(_197_),
    .B(_156_),
    .C(_201_),
    .Y(_202_)
);

FILL FILL_1__570_ (
);

FILL FILL_2__604_ (
);

FILL FILL_5__328_ (
);

FILL FILL75750x7350 (
);

FILL FILL_6__443_ (
);

FILL FILL_0__419_ (
);

FILL FILL_0__592_ (
);

INVX1 _595_ (
    .A(_108_),
    .Y(_124_)
);

FILL FILL_2__413_ (
);

FILL FILL_5__557_ (
);

FILL FILL_1__435_ (
);

FILL FILL_8__401_ (
);

FILL FILL_4__579_ (
);

FILL FILL_5__366_ (
);

FILL FILL_6__481_ (
);

FILL FILL_7__515_ (
);

FILL FILL_0__457_ (
);

FILL FILL76050x61350 (
);

FILL FILL_4__388_ (
);

FILL FILL76050x28950 (
);

FILL FILL_2__451_ (
);

FILL FILL_5__595_ (
);

FILL FILL_6__537_ (
);

FILL FILL_4__600_ (
);

FILL FILL_7__324_ (
);

FILL FILL75750x43350 (
);

FILL FILL_1__473_ (
);

FILL FILL_2__507_ (
);

FILL FILL_3__622_ (
);

FILL FILL_6__346_ (
);

FILL FILL74550x25350 (
);

FILL FILL_7__553_ (
);

FILL FILL_0__495_ (
);

FILL FILL_1__529_ (
);

INVX1 _498_ (
    .A(Atmp[8]),
    .Y(_43_)
);

FILL FILL_2__316_ (
);

FILL FILL_3__431_ (
);

FILL FILL_6__575_ (
);

FILL FILL_7__609_ (
);

FILL FILL_7__362_ (
);

FILL FILL_1__338_ (
);

FILL FILL_2__545_ (
);

FILL FILL_6__384_ (
);

FILL FILL_7__418_ (
);

FILL FILL_7__591_ (
);

FILL FILL_1__567_ (
);

FILL FILL_8__533_ (
);

FILL FILL_2__354_ (
);

FILL FILL_5__498_ (
);

FILL FILL74850x68550 (
);

FILL FILL_4__503_ (
);

FILL FILL_0__589_ (
);

FILL FILL_1__376_ (
);

FILL FILL_8__342_ (
);

FILL FILL_2__583_ (
);

FILL FILL_3__525_ (
);

FILL FILL_7__456_ (
);

FILL FILL_0__398_ (
);

FILL FILL_8__571_ (
);

FILL FILL_2__392_ (
);

FILL FILL_0__610_ (
);

FILL FILL_3__334_ (
);

FILL FILL_6__478_ (
);

NAND2X1 _613_ (
    .A(_139_),
    .B(_140_),
    .Y(_141_)
);

FILL FILL_4__541_ (
);

FILL FILL_8__380_ (
);

FILL FILL_2__448_ (
);

FILL FILL_3__563_ (
);

NOR2X1 _422_ (
    .A(_141_),
    .B(_131_),
    .Y(_254_)
);

FILL FILL_4__350_ (
);

FILL FILL_7__494_ (
);

FILL FILL_8__436_ (
);

FILL FILL_3__619_ (
);

FILL FILL_3__372_ (
);

FILL FILL_4__406_ (
);

DFFPOSX1 _651_ (
    .D(_25_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[18])
);

FILL FILL_5__613_ (
);

FILL FILL_8__665_ (
);

FILL FILL_2__486_ (
);

FILL FILL_3__428_ (
);

FILL FILL_7__359_ (
);

OAI21X1 _460_ (
    .A(_277_),
    .B(_282_),
    .C(_288_),
    .Y(_289_)
);

FILL FILL_5__422_ (
);

FILL FILL_8__474_ (
);

FILL FILL_0__513_ (
);

OAI21X1 _516_ (
    .A(RdyCtl[3]),
    .B(_57_),
    .C(_59_),
    .Y(_60_)
);

FILL FILL_4__444_ (
);

FILL FILL_7__588_ (
);

FILL FILL_0__322_ (
);

FILL FILL_3__466_ (
);

FILL FILL_4_BUFX2_insert10 (
);

FILL FILL_4_BUFX2_insert11 (
);

OAI21X1 _325_ (
    .A(_159_),
    .B(_156_),
    .C(_157_),
    .Y(_164_)
);

FILL FILL_4_BUFX2_insert12 (
);

FILL FILL_4_BUFX2_insert13 (
);

FILL FILL_4_BUFX2_insert14 (
);

FILL FILL_4_BUFX2_insert15 (
);

FILL FILL_4_BUFX2_insert16 (
);

FILL FILL_4_BUFX2_insert17 (
);

FILL FILL_4_BUFX2_insert18 (
);

FILL FILL_4_BUFX2_insert19 (
);

FILL FILL_7__397_ (
);

FILL FILL_8__339_ (
);

FILL FILL75150x68550 (
);

FILL FILL_5__460_ (
);

FILL FILL_6__402_ (
);

FILL FILL_0__551_ (
);

AOI21X1 _554_ (
    .A(_86_),
    .B(RdyCtl_6_bF$buf1),
    .C(_87_),
    .Y(_8_)
);

FILL FILL_4__482_ (
);

FILL FILL_5__516_ (
);

FILL FILL_2__389_ (
);

FILL FILL_0__607_ (
);

FILL FILL_0__360_ (
);

FILL FILL_0_CLKBUF1_insert0 (
);

FILL FILL_0_CLKBUF1_insert1 (
);

FILL FILL_0_CLKBUF1_insert2 (
);

FILL FILL_0_CLKBUF1_insert3 (
);

FILL FILL_0_CLKBUF1_insert4 (
);

FILL FILL_0_CLKBUF1_insert5 (
);

FILL FILL_4__538_ (
);

INVX1 _363_ (
    .A(_189_),
    .Y(_199_)
);

FILL FILL_2__601_ (
);

FILL FILL_5__325_ (
);

FILL FILL_8__377_ (
);

FILL FILL_6__440_ (
);

FILL FILL_0__416_ (
);

NOR2X1 _419_ (
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_251_)
);

FILL FILL_1__623_ (
);

FILL FILL_4__347_ (
);

NOR2X1 _592_ (
    .A(_73__bF$buf3),
    .B(_121_),
    .Y(_122_)
);

FILL FILL_2__410_ (
);

FILL FILL_5__554_ (
);

FILL FILL75450x21750 (
);

FILL FILL_3__369_ (
);

DFFPOSX1 _648_ (
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[15])
);

FILL FILL_1__432_ (
);

FILL FILL_4__576_ (
);

FILL FILL_5__363_ (
);

FILL FILL_7__512_ (
);

FILL FILL_0__454_ (
);

FILL FILL_3__598_ (
);

INVX1 _457_ (
    .A(_0_),
    .Y(_286_)
);

FILL FILL_4__385_ (
);

FILL FILL_5__419_ (
);

FILL FILL_5__592_ (
);

FILL FILL_6__534_ (
);

FILL FILL_7__321_ (
);

FILL FILL_1__470_ (
);

FILL FILL_2__504_ (
);

FILL FILL75750x64950 (
);

FILL FILL_6__343_ (
);

FILL FILL_0__319_ (
);

FILL FILL_7__550_ (
);

FILL FILL_0__492_ (
);

FILL FILL_1__526_ (
);

INVX1 _495_ (
    .A(RdyCtl[2]),
    .Y(_40_)
);

FILL FILL_2__313_ (
);

FILL FILL_5__457_ (
);

FILL FILL_6__572_ (
);

FILL FILL_7__606_ (
);

FILL FILL_0__548_ (
);

FILL FILL_1__335_ (
);

FILL FILL_4__479_ (
);

FILL FILL_2__542_ (
);

FILL FILL_6__381_ (
);

FILL FILL_7__415_ (
);

FILL FILL_0__357_ (
);

FILL FILL_1__564_ (
);

FILL FILL_8__530_ (
);

FILL FILL_2__351_ (
);

FILL FILL_5__495_ (
);

FILL FILL_6__437_ (
);

FILL FILL_4__500_ (
);

FILL FILL_0__586_ (
);

NOR2X1 _589_ (
    .A(_118_),
    .B(_117_),
    .Y(_119_)
);

FILL FILL_1__373_ (
);

FILL FILL_2__407_ (
);

FILL FILL_2__580_ (
);

FILL FILL_3__522_ (
);

FILL FILL_6__666_ (
);

FILL FILL76050x14550 (
);

FILL FILL_7__453_ (
);

FILL FILL_0__395_ (
);

FILL FILL_1__429_ (
);

NOR2X1 _398_ (
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_231_)
);

FILL FILL_3__331_ (
);

FILL FILL_6__475_ (
);

FILL FILL_7__509_ (
);

OAI21X1 _610_ (
    .A(_134_),
    .B(_128_),
    .C(_129_),
    .Y(_138_)
);

FILL FILL_8__624_ (
);

FILL FILL_2__445_ (
);

FILL FILL_5__589_ (
);

FILL FILL_3__560_ (
);

FILL FILL_7__318_ (
);

FILL FILL_7__491_ (
);

FILL FILL_1__467_ (
);

FILL FILL_8__433_ (
);

FILL FILL_5__398_ (
);

FILL FILL_3__616_ (
);

FILL FILL_8_BUFX2_insert7 (
);

FILL FILL_8_BUFX2_insert8 (
);

FILL FILL_8_BUFX2_insert9 (
);

FILL FILL_4__403_ (
);

FILL FILL_7__547_ (
);

FILL FILL_0__489_ (
);

FILL FILL_5__610_ (
);

FILL FILL_2__483_ (
);

FILL FILL_3__425_ (
);

FILL FILL_6__569_ (
);

FILL FILL_7__356_ (
);

FILL FILL_8__471_ (
);

FILL FILL_2__539_ (
);

FILL FILL74850x54150 (
);

FILL FILL_0__510_ (
);

FILL FILL_6__378_ (
);

OAI21X1 _513_ (
    .A(_44_),
    .B(_56_),
    .C(_45_),
    .Y(_57_)
);

FILL FILL_4__441_ (
);

FILL FILL_7__585_ (
);

FILL FILL_8__527_ (
);

FILL FILL_2__348_ (
);

FILL FILL_3__463_ (
);

NAND2X1 _322_ (
    .A(_161_),
    .B(_160_),
    .Y(_162_)
);

FILL FILL_7__394_ (
);

FILL FILL_8__336_ (
);

FILL FILL_2__577_ (
);

FILL FILL_3__519_ (
);

INVX1 _551_ (
    .A(_84_),
    .Y(_85_)
);

FILL FILL_5__513_ (
);

FILL FILL_1__599_ (
);

FILL FILL_8__565_ (
);

FILL FILL_2__386_ (
);

FILL FILL_0__604_ (
);

FILL FILL_3__328_ (
);

NAND2X1 _607_ (
    .A(_135_),
    .B(_132_),
    .Y(_136_)
);

FILL FILL_4__535_ (
);

NOR2X1 _360_ (
    .A(_159_),
    .B(_169_),
    .Y(_196_)
);

FILL FILL_5__322_ (
);

FILL FILL_8__374_ (
);

FILL FILL_0__413_ (
);

FILL FILL_3__557_ (
);

AOI21X1 _416_ (
    .A(_244_),
    .B(_242_),
    .C(_247_),
    .Y(_248_)
);

FILL FILL_1__620_ (
);

FILL FILL_4__344_ (
);

FILL FILL_7__488_ (
);

FILL FILL_5__551_ (
);

FILL FILL_3__366_ (
);

DFFPOSX1 _645_ (
    .D(_19_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[12])
);

FILL FILL_4__573_ (
);

FILL FILL_5__607_ (
);

FILL FILL_5__360_ (
);

FILL FILL_0__451_ (
);

FILL FILL_3__595_ (
);

NAND2X1 _454_ (
    .A(_279_),
    .B(_283_),
    .Y(_284_)
);

FILL FILL_4__382_ (
);

FILL FILL_5__416_ (
);

FILL FILL_8__468_ (
);

FILL FILL_6__531_ (
);

FILL FILL_0__507_ (
);

FILL FILL75150x54150 (
);

FILL FILL_4__438_ (
);

FILL FILL_2__501_ (
);

FILL FILL_6__340_ (
);

FILL FILL_0__316_ (
);

NAND2X1 _319_ (
    .A(_157_),
    .B(_158_),
    .Y(_159_)
);

FILL FILL_1__523_ (
);

FILL FILL_4__667_ (
);

OAI21X1 _492_ (
    .A(acc_reg[18]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_310_)
);

FILL FILL_5__454_ (
);

FILL FILL73650x18150 (
);

FILL FILL_7__603_ (
);

FILL FILL_0__545_ (
);

OAI21X1 _548_ (
    .A(_81_),
    .B(_80_),
    .C(_78_),
    .Y(_82_)
);

FILL FILL_1__332_ (
);

FILL FILL_4__476_ (
);

FILL FILL_6__625_ (
);

FILL FILL_7__412_ (
);

FILL FILL_0__354_ (
);

FILL FILL_3__498_ (
);

OAI21X1 _357_ (
    .A(acc_reg[11]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_194_)
);

FILL FILL_1__561_ (
);

FILL FILL_5__319_ (
);

FILL FILL_5__492_ (
);

FILL FILL_6__434_ (
);

FILL FILL_0__583_ (
);

FILL FILL_1__617_ (
);

AOI21X1 _586_ (
    .A(_111_),
    .B(_112_),
    .C(_108_),
    .Y(_116_)
);

FILL FILL_1__370_ (
);

FILL FILL_2__404_ (
);

FILL FILL_5__548_ (
);

FILL FILL_7__450_ (
);

FILL FILL_0__392_ (
);

FILL FILL_1__426_ (
);

NAND2X1 _395_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_228_)
);

FILL FILL_5__357_ (
);

FILL FILL_6__472_ (
);

FILL FILL_7__506_ (
);

FILL FILL_0__448_ (
);

FILL FILL_8__621_ (
);

FILL FILL_4__379_ (
);

FILL FILL75750x50550 (
);

FILL FILL_2__442_ (
);

FILL FILL_5__586_ (
);

FILL FILL_6__528_ (
);

FILL FILL_7__315_ (
);

FILL FILL_1__464_ (
);

FILL FILL_8__430_ (
);

FILL FILL_5__395_ (
);

FILL FILL_3__613_ (
);

FILL FILL_6__337_ (
);

FILL FILL_4__400_ (
);

FILL FILL_7__544_ (
);

FILL FILL_0__486_ (
);

OAI21X1 _489_ (
    .A(acc_reg[17]),
    .B(_73__bF$buf3),
    .C(En_bF$buf2),
    .Y(_308_)
);

FILL FILL_2__480_ (
);

FILL FILL_3__422_ (
);

FILL FILL_6__566_ (
);

FILL FILL_7__353_ (
);

FILL FILL_1__329_ (
);

FILL FILL_2__536_ (
);

FILL FILL_6__375_ (
);

FILL FILL_7__409_ (
);

OAI21X1 _510_ (
    .A(RdyCtl[0]),
    .B(_53_),
    .C(_54_),
    .Y(_311_[0])
);

FILL FILL_7__582_ (
);

FILL FILL_1__558_ (
);

FILL FILL_8__524_ (
);

FILL FILL_2__345_ (
);

FILL FILL_5__489_ (
);

FILL FILL_3__460_ (
);

BUFX2 BUFX2_insert10 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(En),
    .Y(En_bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .A(En),
    .Y(En_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .A(En),
    .Y(En_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .A(En),
    .Y(En_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .A(En),
    .Y(En_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .A(_73_),
    .Y(_73__bF$buf4)
);

FILL FILL_7__391_ (
);

BUFX2 BUFX2_insert17 (
    .A(_73_),
    .Y(_73__bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .A(_73_),
    .Y(_73__bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .A(_73_),
    .Y(_73__bF$buf1)
);

FILL FILL_1__367_ (
);

FILL FILL_8__333_ (
);

FILL FILL_2__574_ (
);

FILL FILL_3__516_ (
);

FILL FILL_7__447_ (
);

FILL FILL_0__389_ (
);

FILL FILL_5__510_ (
);

FILL FILL_1__596_ (
);

FILL FILL_8__562_ (
);

FILL FILL75150x7350 (
);

FILL FILL_2__383_ (
);

FILL FILL_0__601_ (
);

FILL FILL_3__325_ (
);

FILL FILL_6__469_ (
);

INVX1 _604_ (
    .A(_129_),
    .Y(_133_)
);

FILL FILL_4__532_ (
);

FILL FILL_8__618_ (
);

FILL FILL_2__439_ (
);

FILL FILL_0__410_ (
);

FILL FILL_3__554_ (
);

NAND3X1 _413_ (
    .A(_219_),
    .B(_239_),
    .C(_232_),
    .Y(_245_)
);

FILL FILL_4__341_ (
);

FILL FILL_7__485_ (
);

FILL FILL_8__427_ (
);

FILL FILL_2__668_ (
);

FILL FILL_3__363_ (
);

DFFPOSX1 _642_ (
    .D(_16_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[9])
);

FILL FILL_4__570_ (
);

FILL FILL_5__604_ (
);

FILL FILL_2__477_ (
);

FILL FILL_3__419_ (
);

FILL FILL_3__592_ (
);

INVX1 _451_ (
    .A(_273_),
    .Y(_281_)
);

FILL FILL_5__413_ (
);

FILL FILL_1__499_ (
);

FILL FILL_5_BUFX2_insert20 (
);

FILL FILL_0__504_ (
);

NAND2X1 _507_ (
    .A(RdyCtl[1]),
    .B(_51_),
    .Y(_52_)
);

FILL FILL_4__435_ (
);

FILL FILL_7__579_ (
);

FILL FILL74550x150 (
);

FILL FILL_0__313_ (
);

FILL FILL_3__457_ (
);

AOI21X1 _316_ (
    .A(_150_),
    .B(_111_),
    .C(_155_),
    .Y(_156_)
);

FILL FILL_1__520_ (
);

FILL FILL_7__388_ (
);

FILL FILL_5__451_ (
);

FILL FILL_7__600_ (
);

FILL FILL_0__542_ (
);

NAND2X1 _545_ (
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_79_)
);

FILL FILL_4__473_ (
);

FILL FILL_5__507_ (
);

FILL FILL73650x39750 (
);

FILL FILL_6__622_ (
);

FILL FILL_0__351_ (
);

FILL FILL_3__495_ (
);

FILL FILL_4__529_ (
);

INVX1 _354_ (
    .A(_190_),
    .Y(_191_)
);

FILL FILL_5__316_ (
);

FILL FILL_8__368_ (
);

FILL FILL_6__431_ (
);

FILL FILL_0__407_ (
);

FILL FILL_0__580_ (
);

FILL FILL_1__614_ (
);

FILL FILL_4__338_ (
);

NAND2X1 _583_ (
    .A(_113_),
    .B(_110_),
    .Y(_114_)
);

FILL FILL_2__401_ (
);

FILL FILL_5__545_ (
);

FILL FILL74250x10950 (
);

DFFPOSX1 _639_ (
    .D(_13_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[6])
);

FILL FILL_1__423_ (
);

FILL FILL_4__567_ (
);

NAND2X1 _392_ (
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

FILL FILL_5__354_ (
);

FILL FILL_7__503_ (
);

FILL FILL_0__445_ (
);

FILL FILL_3__589_ (
);

NOR2X1 _448_ (
    .A(_277_),
    .B(_276_),
    .Y(_278_)
);

FILL FILL_4__376_ (
);

FILL FILL_5__583_ (
);

FILL FILL_6__525_ (
);

FILL FILL_3__398_ (
);

FILL FILL_1__461_ (
);

FILL FILL_5__392_ (
);

FILL FILL_3__610_ (
);

FILL FILL_6__334_ (
);

FILL FILL_7__541_ (
);

FILL FILL_0__483_ (
);

FILL FILL_1__517_ (
);

AOI21X1 _486_ (
    .A(_58_),
    .B(_73__bF$buf0),
    .C(_306_),
    .Y(_34_)
);

FILL FILL_5__448_ (
);

FILL FILL_6__563_ (
);

FILL FILL_0__539_ (
);

FILL FILL_7__350_ (
);

FILL FILL_1__326_ (
);

FILL FILL_2__533_ (
);

FILL FILL_6__619_ (
);

FILL FILL_6__372_ (
);

FILL FILL_7__406_ (
);

FILL FILL_0__348_ (
);

FILL FILL_1__555_ (
);

FILL FILL_8__521_ (
);

FILL FILL_2__342_ (
);

FILL FILL_5__486_ (
);

FILL FILL_6__428_ (
);

FILL FILL_0__577_ (
);

FILL FILL_1__364_ (
);

FILL FILL_8__330_ (
);

FILL FILL76050x21750 (
);

FILL FILL_2__571_ (
);

FILL FILL_3__513_ (
);

FILL FILL_7__444_ (
);

FILL FILL_0__386_ (
);

OR2X2 _389_ (
    .A(_221_),
    .B(_222_),
    .Y(_223_)
);

FILL FILL_1__593_ (
);

FILL FILL_2__380_ (
);

FILL FILL_3__322_ (
);

FILL FILL_6__466_ (
);

OR2X2 _601_ (
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_130_)
);

FILL FILL_2__436_ (
);

FILL FILL_3__551_ (
);

NAND2X1 _410_ (
    .A(_200_),
    .B(_198_),
    .Y(_242_)
);

FILL FILL_7__482_ (
);

FILL FILL_1__458_ (
);

FILL FILL_8__424_ (
);

FILL FILL_2__665_ (
);

FILL FILL_5__389_ (
);

FILL FILL_3__607_ (
);

FILL FILL_3__360_ (
);

FILL FILL_7__538_ (
);

FILL FILL_5__601_ (
);

FILL FILL_2__474_ (
);

FILL FILL_3__416_ (
);

FILL FILL74850x61350 (
);

FILL FILL_4__623_ (
);

FILL FILL74850x28950 (
);

FILL FILL_7__347_ (
);

FILL FILL_5__410_ (
);

FILL FILL_1__496_ (
);

FILL FILL_8__462_ (
);

FILL FILL_0__501_ (
);

FILL FILL_6__369_ (
);

NAND2X1 _504_ (
    .A(_40_),
    .B(_48_),
    .Y(_49_)
);

FILL FILL_4__432_ (
);

FILL FILL_7__576_ (
);

FILL FILL_8__518_ (
);

FILL FILL_2__339_ (
);

FILL FILL_3__454_ (
);

FILL FILL_6__598_ (
);

OAI21X1 _313_ (
    .A(_129_),
    .B(_147_),
    .C(_139_),
    .Y(_153_)
);

FILL FILL_7__385_ (
);

FILL FILL_8__327_ (
);

FILL FILL_2__568_ (
);

OAI21X1 _542_ (
    .A(_75_),
    .B(_76_),
    .C(En_bF$buf3),
    .Y(_77_)
);

FILL FILL_4__470_ (
);

FILL FILL_5__504_ (
);

FILL FILL_8__556_ (
);

FILL FILL_2__377_ (
);

FILL FILL_3__319_ (
);

FILL FILL_3__492_ (
);

FILL FILL_4__526_ (
);

AND2X2 _351_ (
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_188_)
);

FILL FILL_5__313_ (
);

FILL FILL_1__399_ (
);

FILL FILL_8__365_ (
);

FILL FILL_0__404_ (
);

FILL FILL_3__548_ (
);

NOR2X1 _407_ (
    .A(_222_),
    .B(_221_),
    .Y(_239_)
);

FILL FILL_1__611_ (
);

FILL FILL_4__335_ (
);

FILL FILL_7__479_ (
);

NAND2X1 _580_ (
    .A(_106_),
    .B(_104_),
    .Y(_111_)
);

FILL FILL_5__542_ (
);

FILL FILL_8__594_ (
);

FILL FILL_3__357_ (
);

DFFPOSX1 _636_ (
    .D(_10_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[3])
);

FILL FILL_1__420_ (
);

FILL FILL_4__564_ (
);

FILL FILL_5__351_ (
);

FILL FILL_7__500_ (
);

FILL FILL_0__442_ (
);

FILL FILL_3__586_ (
);

INVX1 _445_ (
    .A(FCW[18]),
    .Y(_275_)
);

FILL FILL_4__373_ (
);

FILL FILL_5__407_ (
);

FILL FILL_8__459_ (
);

FILL FILL75150x61350 (
);

FILL FILL_5__580_ (
);

FILL FILL75150x28950 (
);

FILL FILL_6__522_ (
);

FILL FILL_3__395_ (
);

FILL FILL_4__429_ (
);

FILL FILL_6__331_ (
);

FILL FILL_0__480_ (
);

FILL FILL_1__514_ (
);

OAI21X1 _483_ (
    .A(acc_reg[14]),
    .B(_73__bF$buf0),
    .C(En_bF$buf3),
    .Y(_305_)
);

FILL FILL74850x7350 (
);

FILL FILL_5__445_ (
);

FILL FILL_8__497_ (
);

FILL FILL_6__560_ (
);

FILL FILL_0__536_ (
);

NOR2X1 _539_ (
    .A(_66_),
    .B(_74_),
    .Y(_6_)
);

FILL FILL_1__323_ (
);

FILL FILL_4__467_ (
);

FILL FILL_2__530_ (
);

FILL FILL_6__616_ (
);

FILL FILL_7__403_ (
);

FILL FILL_0__345_ (
);

FILL FILL_3__489_ (
);

AOI21X1 _348_ (
    .A(_184_),
    .B(RdyCtl_6_bF$buf3),
    .C(_185_),
    .Y(_17_)
);

FILL FILL_1__552_ (
);

FILL FILL_5__483_ (
);

FILL FILL_6__425_ (
);

FILL FILL_0__574_ (
);

FILL FILL_1__608_ (
);

AND2X2 _577_ (
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_108_)
);

FILL FILL_1__361_ (
);

FILL FILL_5__539_ (
);

FILL FILL_3__510_ (
);

FILL FILL_7__441_ (
);

FILL FILL_0__383_ (
);

FILL FILL_1__417_ (
);

AOI21X1 _386_ (
    .A(_202_),
    .B(_217_),
    .C(_219_),
    .Y(_220_)
);

FILL FILL_1__590_ (
);

FILL FILL_2__624_ (
);

FILL FILL_5__348_ (
);

FILL FILL_6__463_ (
);

FILL FILL_0__439_ (
);

FILL FILL_8__612_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_2__433_ (
);

FILL FILL_1_BUFX2_insert18 (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_5__577_ (
);

FILL FILL_6__519_ (
);

FILL FILL_0__668_ (
);

FILL FILL_1__455_ (
);

FILL FILL_8__421_ (
);

FILL FILL_4__599_ (
);

FILL FILL_5__386_ (
);

FILL FILL_3__604_ (
);

FILL FILL75450x36150 (
);

FILL FILL_6__328_ (
);

FILL FILL_7__535_ (
);

FILL FILL_0__477_ (
);

FILL FILL74250x18150 (
);

FILL FILL_2__471_ (
);

FILL FILL_3__413_ (
);

FILL FILL_6__557_ (
);

FILL FILL_4__620_ (
);

FILL FILL_7__344_ (
);

FILL FILL_1__493_ (
);

FILL FILL_2__527_ (
);

FILL FILL_6__366_ (
);

OAI21X1 _501_ (
    .A(_43_),
    .B(_44_),
    .C(_45_),
    .Y(_46_)
);

FILL FILL_7__573_ (
);

FILL FILL_1__549_ (
);

FILL FILL_8__515_ (
);

FILL FILL_2__336_ (
);

FILL FILL_3__451_ (
);

FILL FILL_6__595_ (
);

FILL FILL_7__382_ (
);

FILL FILL_1__358_ (
);

FILL FILL_2__565_ (
);

FILL FILL_3__507_ (
);

FILL FILL_6_BUFX2_insert10 (
);

FILL FILL_6_BUFX2_insert11 (
);

FILL FILL_6_BUFX2_insert12 (
);

FILL FILL_6_BUFX2_insert13 (
);

FILL FILL_6_BUFX2_insert14 (
);

FILL FILL_6_BUFX2_insert15 (
);

FILL FILL_6_BUFX2_insert16 (
);

FILL FILL_6_BUFX2_insert17 (
);

FILL FILL_6_BUFX2_insert18 (
);

FILL FILL_6_BUFX2_insert19 (
);

FILL FILL_7__438_ (
);

FILL FILL_5__501_ (
);

FILL FILL_1__587_ (
);

FILL FILL_8__553_ (
);

FILL FILL_2__374_ (
);

FILL FILL_3__316_ (
);

FILL FILL_4__523_ (
);

FILL FILL_7__667_ (
);

FILL FILL_8__609_ (
);

FILL FILL_1__396_ (
);

FILL FILL_0__401_ (
);

FILL FILL_3__545_ (
);

AOI21X1 _404_ (
    .A(_234_),
    .B(_236_),
    .C(_73__bF$buf4),
    .Y(_237_)
);

FILL FILL_4__332_ (
);

FILL FILL_7__476_ (
);

FILL FILL75450x3750 (
);

FILL FILL_8__591_ (
);

FILL FILL74850x14550 (
);

FILL FILL_3__354_ (
);

FILL FILL_6__498_ (
);

DFFPOSX1 _633_ (
    .D(_7_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[0])
);

FILL FILL_4__561_ (
);

FILL FILL_2__468_ (
);

FILL FILL_3__583_ (
);

FILL FILL_4__617_ (
);

NAND2X1 _442_ (
    .A(_252_),
    .B(_268_),
    .Y(_272_)
);

FILL FILL_4__370_ (
);

FILL FILL_5__404_ (
);

FILL FILL_3__392_ (
);

FILL FILL_4__426_ (
);

FILL FILL_3__448_ (
);

FILL FILL_1__511_ (
);

FILL FILL_7__379_ (
);

AOI21X1 _480_ (
    .A(_39_),
    .B(_73__bF$buf2),
    .C(_303_),
    .Y(_31_)
);

FILL FILL_5__442_ (
);

FILL FILL_8__494_ (
);

FILL FILL_0__533_ (
);

NOR2X1 _536_ (
    .A(_40_),
    .B(_74_),
    .Y(_3_)
);

FILL FILL_1__320_ (
);

FILL FILL_4__464_ (
);

FILL FILL_6__613_ (
);

FILL FILL_7__400_ (
);

FILL FILL_0__342_ (
);

FILL FILL_3__486_ (
);

OR2X2 _345_ (
    .A(_178_),
    .B(_181_),
    .Y(_183_)
);

FILL FILL_8__359_ (
);

FILL FILL_5__480_ (
);

FILL FILL_6__422_ (
);

FILL FILL_0__571_ (
);

FILL FILL_1__605_ (
);

FILL FILL_4__329_ (
);

INVX1 _574_ (
    .A(_98_),
    .Y(_105_)
);

FILL FILL_5__536_ (
);

FILL FILL_8__588_ (
);

FILL FILL_0__380_ (
);

FILL FILL_1__414_ (
);

FILL FILL_4__558_ (
);

NOR2X1 _383_ (
    .A(_205_),
    .B(_213_),
    .Y(_217_)
);

FILL FILL75150x14550 (
);

FILL FILL_2__621_ (
);

FILL FILL_5__345_ (
);

FILL FILL_8__397_ (
);

FILL FILL_6__460_ (
);

FILL FILL_0__436_ (
);

AOI21X1 _439_ (
    .A(_265_),
    .B(_268_),
    .C(_73__bF$buf2),
    .Y(_270_)
);

FILL FILL_4__367_ (
);

FILL FILL_2__430_ (
);

FILL FILL_5__574_ (
);

FILL FILL_6__516_ (
);

FILL FILL_0__665_ (
);

FILL FILL_3__389_ (
);

BUFX2 _668_ (
    .A(RdyCtl_6_bF$buf1),
    .Y(Vld)
);

FILL FILL_1__452_ (
);

FILL FILL_4__596_ (
);

FILL FILL_5__383_ (
);

FILL FILL_3__601_ (
);

FILL FILL_6__325_ (
);

FILL FILL_7__532_ (
);

FILL FILL_0__474_ (
);

FILL FILL_5_BUFX2_insert6 (
);

FILL FILL_5_BUFX2_insert7 (
);

FILL FILL_5_BUFX2_insert8 (
);

FILL FILL_1__508_ (
);

FILL FILL_5_BUFX2_insert9 (
);

OAI21X1 _477_ (
    .A(acc_reg[11]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_302_)
);

FILL FILL75450x57750 (
);

FILL FILL_5__439_ (
);

FILL FILL_3__410_ (
);

FILL FILL_6__554_ (
);

FILL FILL74250x39750 (
);

FILL FILL_7__341_ (
);

FILL FILL_1__317_ (
);

FILL FILL_1__490_ (
);

FILL FILL_2__524_ (
);

FILL FILL_5__668_ (
);

FILL FILL_6__363_ (
);

FILL FILL_0__339_ (
);

FILL FILL_7__570_ (
);

FILL FILL_1__546_ (
);

FILL FILL_2__333_ (
);

FILL FILL_5__477_ (
);

FILL FILL_6__419_ (
);

FILL FILL_6__592_ (
);

FILL FILL_0__568_ (
);

FILL FILL_1__355_ (
);

FILL FILL_8__321_ (
);

FILL FILL_4__499_ (
);

FILL FILL_2__562_ (
);

FILL FILL_3__504_ (
);

FILL FILL75750x10950 (
);

FILL FILL_7__435_ (
);

FILL FILL_0__377_ (
);

FILL FILL_7_BUFX2_insert6 (
);

FILL FILL_7_BUFX2_insert7 (
);

FILL FILL_7_BUFX2_insert8 (
);

FILL FILL_7_BUFX2_insert9 (
);

FILL FILL74850x150 (
);

FILL FILL_1__584_ (
);

FILL FILL_2__618_ (
);

FILL FILL_2__371_ (
);

FILL FILL_3__313_ (
);

FILL FILL_6__457_ (
);

FILL FILL_4__520_ (
);

FILL FILL_1__393_ (
);

FILL FILL_2__427_ (
);

FILL FILL_3__542_ (
);

OAI21X1 _401_ (
    .A(_223_),
    .B(_220_),
    .C(_228_),
    .Y(_234_)
);

FILL FILL_7__473_ (
);

FILL FILL_1__449_ (
);

FILL FILL_8__415_ (
);

FILL FILL_3__351_ (
);

FILL FILL_6__495_ (
);

FILL FILL_7__529_ (
);

DFFPOSX1 _630_ (
    .D(_4_),
    .CLK(clk_bF$buf3),
    .Q(RdyCtl[4])
);

FILL FILL_2__465_ (
);

FILL FILL_3__407_ (
);

FILL FILL_3__580_ (
);

FILL FILL_4__614_ (
);

FILL FILL_7__338_ (
);

FILL FILL_5__401_ (
);

FILL FILL_1__487_ (
);

FILL FILL_8__453_ (
);

FILL FILL_4__423_ (
);

FILL FILL_7__567_ (
);

FILL FILL_8__509_ (
);

FILL FILL_3__445_ (
);

FILL FILL_6__589_ (
);

FILL FILL_7__376_ (
);

FILL FILL_8__318_ (
);

FILL FILL_8__491_ (
);

FILL FILL_2__559_ (
);

FILL FILL_0__530_ (
);

FILL FILL_6__398_ (
);

NOR2X1 _533_ (
    .A(_73__bF$buf2),
    .B(_74_),
    .Y(_0_)
);

FILL FILL_4__461_ (
);

FILL FILL_8__547_ (
);

FILL FILL_6__610_ (
);

FILL FILL_2__368_ (
);

FILL FILL_3__483_ (
);

FILL FILL_4__517_ (
);

NOR2X1 _342_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_180_)
);

FILL FILL_8__356_ (
);

FILL FILL_2__597_ (
);

FILL FILL_3__539_ (
);

FILL FILL_1__602_ (
);

FILL FILL_4__326_ (
);

NAND2X1 _571_ (
    .A(_100_),
    .B(_102_),
    .Y(_103_)
);

FILL FILL_5__533_ (
);

FILL FILL_8__585_ (
);

FILL FILL_0__624_ (
);

FILL FILL_3__348_ (
);

DFFPOSX1 _627_ (
    .D(_1_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[1])
);

FILL FILL_1__411_ (
);

FILL FILL_4__555_ (
);

AOI21X1 _380_ (
    .A(_210_),
    .B(_213_),
    .C(_73__bF$buf4),
    .Y(_215_)
);

FILL FILL_5__342_ (
);

FILL FILL_8__394_ (
);

FILL FILL_0__433_ (
);

FILL FILL_3__577_ (
);

NOR2X1 _436_ (
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_267_)
);

FILL FILL_4__364_ (
);

FILL FILL_5__571_ (
);

FILL FILL_6__513_ (
);

FILL FILL_3__386_ (
);

BUFX2 _665_ (
    .A(_311_[0]),
    .Y(Aout[0])
);

FILL FILL_4__593_ (
);

FILL FILL_5__380_ (
);

FILL FILL_6__322_ (
);

FILL FILL_0__471_ (
);

FILL FILL_1__505_ (
);

NOR2X1 _474_ (
    .A(_299_),
    .B(_300_),
    .Y(_28_)
);

FILL FILL_5__436_ (
);

FILL FILL_8__488_ (
);

FILL FILL_6__551_ (
);

FILL FILL_0__527_ (
);

FILL FILL_1__314_ (
);

FILL FILL_4__458_ (
);

FILL FILL_2__521_ (
);

FILL FILL_5__665_ (
);

FILL FILL_6__607_ (
);

FILL FILL_6__360_ (
);

FILL FILL_0__336_ (
);

OR2X2 _339_ (
    .A(_169_),
    .B(_159_),
    .Y(_177_)
);

FILL FILL_1__543_ (
);

FILL FILL_2__330_ (
);

FILL FILL_5__474_ (
);

FILL FILL_6__416_ (
);

FILL FILL_7__623_ (
);

FILL FILL_0__565_ (
);

OAI21X1 _568_ (
    .A(_89_),
    .B(_92_),
    .C(_99_),
    .Y(_100_)
);

FILL FILL_1__352_ (
);

FILL FILL_4__496_ (
);

FILL FILL_3__501_ (
);

FILL FILL_7__432_ (
);

FILL FILL_0__374_ (
);

FILL FILL_1__408_ (
);

OR2X2 _377_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_212_)
);

FILL FILL_1__581_ (
);

FILL FILL_2__615_ (
);

FILL FILL_5__339_ (
);

FILL FILL_6__454_ (
);

FILL FILL_8__603_ (
);

FILL FILL_1__390_ (
);

FILL FILL_2__424_ (
);

FILL FILL_5__568_ (
);

FILL FILL75450x43350 (
);

FILL FILL73950x150 (
);

FILL FILL_7__470_ (
);

FILL FILL_1__446_ (
);

FILL FILL_8__412_ (
);

FILL FILL_5__377_ (
);

FILL FILL_6__319_ (
);

FILL FILL74250x25350 (
);

FILL FILL_6__492_ (
);

FILL FILL_7__526_ (
);

FILL FILL_0__468_ (
);

FILL FILL_4__399_ (
);

FILL FILL_2__462_ (
);

FILL FILL_3__404_ (
);

FILL FILL_6__548_ (
);

FILL FILL_4__611_ (
);

FILL FILL_7__335_ (
);

FILL FILL_1__484_ (
);

FILL FILL_8__450_ (
);

FILL FILL_2__518_ (
);

FILL FILL_6__357_ (
);

FILL FILL_4__420_ (
);

FILL FILL_7__564_ (
);

FILL FILL_8__506_ (
);

FILL FILL_7_BUFX2_insert20 (
);

FILL FILL_2__327_ (
);

FILL FILL74550x68550 (
);

FILL FILL_3__442_ (
);

FILL FILL_6__586_ (
);

FILL FILL_7__373_ (
);

FILL FILL_1__349_ (
);

FILL FILL_2__556_ (
);

FILL FILL_6__395_ (
);

FILL FILL_7__429_ (
);

OAI21X1 _530_ (
    .A(_66_),
    .B(_71_),
    .C(_72_),
    .Y(_38_)
);

FILL FILL_1__578_ (
);

FILL FILL_8__544_ (
);

FILL FILL_2__365_ (
);

FILL FILL_3__480_ (
);

FILL FILL_4__514_ (
);

FILL FILL_1__387_ (
);

FILL FILL_2__594_ (
);

FILL FILL_3__536_ (
);

FILL FILL76050x7350 (
);

FILL FILL_4__323_ (
);

FILL FILL74850x21750 (
);

FILL FILL_7__467_ (
);

FILL FILL76050x36150 (
);

FILL FILL_5__530_ (
);

FILL FILL_8__582_ (
);

FILL FILL_0__621_ (
);

FILL FILL_3__345_ (
);

FILL FILL_6__489_ (
);

INVX1 _624_ (
    .A(_118_),
    .Y(_151_)
);

FILL FILL_4__552_ (
);

FILL FILL75750x18150 (
);

FILL FILL_8__391_ (
);

FILL FILL_2__459_ (
);

FILL FILL_0__430_ (
);

FILL FILL_3__574_ (
);

FILL FILL_4__608_ (
);

AOI21X1 _433_ (
    .A(_263_),
    .B(RdyCtl_6_bF$buf3),
    .C(_264_),
    .Y(_23_)
);

FILL FILL_4__361_ (
);

FILL FILL_8__447_ (
);

FILL FILL_6__510_ (
);

FILL FILL_3__383_ (
);

FILL FILL_4__417_ (
);

DFFPOSX1 _662_ (
    .D(_36_),
    .CLK(clk_bF$buf3),
    .Q(Atmp[9])
);

FILL FILL_4__590_ (
);

FILL FILL_5__624_ (
);

FILL FILL_2__497_ (
);

FILL FILL_3__439_ (
);

FILL FILL_1__502_ (
);

NOR2X1 _471_ (
    .A(_297_),
    .B(_298_),
    .Y(_27_)
);

FILL FILL_5__433_ (
);

FILL FILL_8__485_ (
);

FILL FILL_0__524_ (
);

FILL FILL_3__668_ (
);

NAND2X1 _527_ (
    .A(_68_),
    .B(_69_),
    .Y(_70_)
);

FILL FILL_4__455_ (
);

FILL FILL_7__599_ (
);

FILL FILL_6__604_ (
);

FILL FILL_0__333_ (
);

FILL FILL_3__477_ (
);

NOR2X1 _336_ (
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_174_)
);

FILL FILL_1__540_ (
);

FILL FILL_5__471_ (
);

FILL FILL_6__413_ (
);

FILL FILL_7__620_ (
);

FILL FILL_0__562_ (
);

AND2X2 _565_ (
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_97_)
);

FILL FILL_4__493_ (
);

FILL FILL_5__527_ (
);

FILL FILL_8__579_ (
);

FILL FILL75150x21750 (
);

FILL FILL_0__618_ (
);

FILL FILL_0__371_ (
);

FILL FILL_1__405_ (
);

FILL FILL_4__549_ (
);

INVX1 _374_ (
    .A(_202_),
    .Y(_209_)
);

FILL FILL_2__612_ (
);

FILL FILL_5__336_ (
);

FILL FILL_8__388_ (
);

FILL FILL_6__451_ (
);

FILL FILL_0__427_ (
);

FILL FILL_8__600_ (
);

FILL FILL_4__358_ (
);

FILL FILL_2__421_ (
);

FILL FILL_5__565_ (
);

FILL FILL_6__507_ (
);

DFFPOSX1 _659_ (
    .D(_33_),
    .CLK(clk_bF$buf0),
    .Q(Atmp[6])
);

FILL FILL_1__443_ (
);

FILL FILL_4__587_ (
);

FILL FILL_5__374_ (
);

FILL FILL_6__316_ (
);

FILL FILL75450x64950 (
);

FILL FILL_7__523_ (
);

FILL FILL_0__465_ (
);

AOI22X1 _468_ (
    .A(_286_),
    .B(_287_),
    .C(_296_),
    .D(_293_),
    .Y(_26_)
);

FILL FILL_4__396_ (
);

FILL FILL_3__401_ (
);

FILL FILL_6__545_ (
);

FILL FILL_7__332_ (
);

FILL FILL73950x61350 (
);

FILL FILL_1__481_ (
);

FILL FILL_2__515_ (
);

FILL FILL75150x150 (
);

FILL FILL_6__354_ (
);

FILL FILL_7__561_ (
);

FILL FILL_1__537_ (
);

FILL FILL_2__324_ (
);

FILL FILL_5__468_ (
);

FILL FILL_6__583_ (
);

FILL FILL_7__617_ (
);

FILL FILL_0__559_ (
);

FILL FILL_7__370_ (
);

FILL FILL_1__346_ (
);

FILL FILL_2__553_ (
);

FILL FILL_6__392_ (
);

FILL FILL_7__426_ (
);

FILL FILL_0__368_ (
);

FILL FILL_1__575_ (
);

FILL FILL_8__541_ (
);

FILL FILL_2__609_ (
);

FILL FILL_2__362_ (
);

FILL FILL_6__448_ (
);

FILL FILL_4__511_ (
);

FILL FILL_0__597_ (
);

FILL FILL_1__384_ (
);

FILL FILL_8__350_ (
);

FILL FILL_2__418_ (
);

FILL FILL_2__591_ (
);

FILL FILL_3__533_ (
);

FILL FILL_4__320_ (
);

FILL FILL_7__464_ (
);

FILL FILL_8__406_ (
);

FILL FILL_3__342_ (
);

FILL FILL_6__486_ (
);

NOR2X1 _621_ (
    .A(_147_),
    .B(_146_),
    .Y(_148_)
);

FILL FILL76050x57750 (
);

FILL FILL_2__456_ (
);

FILL FILL75750x39750 (
);

FILL FILL_3__571_ (
);

FILL FILL_4__605_ (
);

FILL FILL_7__329_ (
);

OAI21X1 _430_ (
    .A(_250_),
    .B(_251_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__478_ (
);

FILL FILL_8__444_ (
);

FILL FILL_3__380_ (
);

FILL FILL_4__414_ (
);

FILL FILL_7__558_ (
);

FILL FILL_5__621_ (
);

FILL FILL_2__494_ (
);

FILL FILL_3__436_ (
);

FILL FILL_7__367_ (
);

FILL FILL_5__430_ (
);

FILL FILL_8__482_ (
);

FILL FILL_0__521_ (
);

FILL FILL_3__665_ (
);

FILL FILL_6__389_ (
);

NAND2X1 _524_ (
    .A(acc_reg[18]),
    .B(acc_reg[19]),
    .Y(_67_)
);

FILL FILL_4__452_ (
);

FILL FILL_7__596_ (
);

FILL FILL_8__538_ (
);

FILL FILL_6__601_ (
);

FILL FILL_2__359_ (
);

FILL FILL_0__330_ (
);

FILL FILL_3__474_ (
);

FILL FILL_4__508_ (
);

NOR2X1 _333_ (
    .A(_73__bF$buf1),
    .B(_171_),
    .Y(_172_)
);

FILL FILL_8__347_ (
);

FILL FILL_6__410_ (
);

FILL FILL_2__588_ (
);

FILL FILL_4__317_ (
);

NAND2X1 _562_ (
    .A(acc_reg[2]),
    .B(_73__bF$buf0),
    .Y(_95_)
);

FILL FILL_4__490_ (
);

FILL FILL_5__524_ (
);

FILL FILL_8__576_ (
);

FILL FILL_2__397_ (
);

FILL FILL_0__615_ (
);

FILL FILL_3__339_ (
);

NAND2X1 _618_ (
    .A(_112_),
    .B(_119_),
    .Y(_145_)
);

FILL FILL_1__402_ (
);

FILL FILL_4__546_ (
);

AND2X2 _371_ (
    .A(_202_),
    .B(_205_),
    .Y(_207_)
);

FILL FILL_5__333_ (
);

FILL FILL_0__424_ (
);

FILL FILL_3__568_ (
);

AND2X2 _427_ (
    .A(_245_),
    .B(_246_),
    .Y(_259_)
);

FILL FILL_4__355_ (
);

FILL FILL_7__499_ (
);

FILL FILL_5__562_ (
);

FILL FILL_6__504_ (
);

FILL FILL_3__377_ (
);

DFFPOSX1 _656_ (
    .D(_30_),
    .CLK(clk_bF$buf5),
    .Q(Atmp[3])
);

FILL FILL_1__440_ (
);

FILL FILL_4__584_ (
);

FILL FILL_5__618_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_3_BUFX2_insert11 (
);

FILL FILL_3_BUFX2_insert12 (
);

FILL FILL_3_BUFX2_insert13 (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert15 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_3_BUFX2_insert18 (
);

FILL FILL_3_BUFX2_insert19 (
);

FILL FILL_5__371_ (
);

FILL FILL_6__313_ (
);

FILL FILL_7__520_ (
);

FILL FILL_0__462_ (
);

AOI21X1 _465_ (
    .A(_274_),
    .B(_278_),
    .C(_276_),
    .Y(_294_)
);

FILL FILL_4__393_ (
);

FILL FILL_5__427_ (
);

FILL FILL_6__542_ (
);

FILL FILL_0__518_ (
);

FILL FILL_4__449_ (
);

FILL FILL_2__512_ (
);

FILL FILL_6__351_ (
);

FILL FILL_0__327_ (
);

FILL FILL_1__534_ (
);

FILL FILL_8__500_ (
);

FILL FILL_2__321_ (
);

FILL FILL_5__465_ (
);

FILL FILL_6__407_ (
);

FILL FILL_6__580_ (
);

FILL FILL_7__614_ (
);

FILL FILL_0__556_ (
);

AND2X2 _559_ (
    .A(_91_),
    .B(_88_),
    .Y(_92_)
);

FILL FILL_1__343_ (
);

FILL FILL_4__487_ (
);

FILL FILL74250x150 (
);

FILL FILL_2__550_ (
);

FILL FILL_7__423_ (
);

FILL FILL_0__365_ (
);

OR2X2 _368_ (
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_204_)
);

FILL FILL_1__572_ (
);

FILL FILL_2__606_ (
);

FILL FILL_6__445_ (
);

FILL FILL_8_BUFX2_insert10 (
);

FILL FILL_8_BUFX2_insert12 (
);

FILL FILL_8_BUFX2_insert13 (
);

FILL FILL_8_BUFX2_insert14 (
);

FILL FILL_8_BUFX2_insert15 (
);

FILL FILL_8_BUFX2_insert17 (
);

FILL FILL_8_BUFX2_insert18 (
);

FILL FILL_8_BUFX2_insert19 (
);

FILL FILL_0__594_ (
);

OAI21X1 _597_ (
    .A(_118_),
    .B(_124_),
    .C(_125_),
    .Y(_126_)
);

FILL FILL75450x50550 (
);

FILL FILL_1__381_ (
);

FILL FILL_2__415_ (
);

FILL FILL_5__559_ (
);

FILL FILL_3__530_ (
);

FILL FILL_7__461_ (
);

FILL FILL_1__437_ (
);

FILL FILL_8__403_ (
);

FILL FILL_5__368_ (
);

FILL FILL_6__483_ (
);

FILL FILL_7__517_ (
);

FILL FILL_0__459_ (
);

FILL FILL73950x14550 (
);

FILL FILL_1__666_ (
);

FILL FILL_2__453_ (
);

FILL FILL_5__597_ (
);

FILL FILL_6__539_ (
);

FILL FILL_4__602_ (
);

FILL FILL_7__326_ (
);

FILL FILL_1__475_ (
);

FILL FILL_8__441_ (
);

FILL FILL_2__509_ (
);

FILL FILL_3__624_ (
);

FILL FILL_6__348_ (
);

FILL FILL_4__411_ (
);

FILL FILL_7__555_ (
);

FILL FILL_0__497_ (
);

FILL FILL_2__318_ (
);

FILL FILL_2__491_ (
);

FILL FILL_3__433_ (
);

FILL FILL_6__577_ (
);

FILL FILL_7__364_ (
);

FILL FILL_2__547_ (
);

FILL FILL_6__386_ (
);

NAND2X1 _521_ (
    .A(RdyCtl[0]),
    .B(Atmp[1]),
    .Y(_65_)
);

FILL FILL_7__593_ (
);

FILL FILL_1__569_ (
);

FILL FILL_8__535_ (
);

FILL FILL_2__356_ (
);

FILL FILL_3__471_ (
);

FILL FILL_4__505_ (
);

NAND2X1 _330_ (
    .A(_165_),
    .B(_168_),
    .Y(_169_)
);

FILL FILL_1__378_ (
);

FILL FILL_8__344_ (
);

FILL FILL_2__585_ (
);

FILL FILL76050x43350 (
);

FILL FILL_3__527_ (
);

FILL FILL_4__314_ (
);

FILL FILL_7__458_ (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_5__521_ (
);

FILL FILL75750x25350 (
);

FILL FILL_2__394_ (
);

FILL FILL_0__612_ (
);

FILL FILL_3__336_ (
);

AOI21X1 _615_ (
    .A(_138_),
    .B(_141_),
    .C(_73__bF$buf1),
    .Y(_143_)
);

FILL FILL_4__543_ (
);

FILL FILL_5__330_ (
);

FILL FILL_8__382_ (
);

FILL FILL_0__421_ (
);

FILL FILL_3__565_ (
);

AOI21X1 _424_ (
    .A(_254_),
    .B(_126_),
    .C(_153_),
    .Y(_256_)
);

FILL FILL_4__352_ (
);

FILL FILL_7__496_ (
);

FILL FILL_8__438_ (
);

FILL FILL_6__501_ (
);

FILL FILL_3__374_ (
);

FILL FILL_4__408_ (
);

DFFPOSX1 _653_ (
    .D(_27_),
    .CLK(clk_bF$buf5),
    .Q(Atmp[0])
);

FILL FILL_4__581_ (
);

FILL FILL_5__615_ (
);

FILL FILL_8__667_ (
);

FILL FILL_2__488_ (
);

OR2X2 _462_ (
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_291_)
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_4__390_ (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_2_BUFX2_insert9 (
);

FILL FILL_5__424_ (
);

FILL FILL_8__476_ (
);

FILL FILL_0__515_ (
);

INVX1 _518_ (
    .A(Atmp[3]),
    .Y(_62_)
);

FILL FILL_4__446_ (
);

FILL FILL73350x39750 (
);

FILL FILL_0__324_ (
);

FILL FILL_3__468_ (
);

INVX1 _327_ (
    .A(acc_reg[9]),
    .Y(_166_)
);

FILL FILL_1__531_ (
);

FILL FILL_7__399_ (
);

FILL FILL_5__462_ (
);

FILL FILL_6__404_ (
);

FILL FILL_7__611_ (
);

FILL FILL_0__553_ (
);

AND2X2 _556_ (
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_89_)
);

FILL FILL_1__340_ (
);

FILL FILL_4__484_ (
);

FILL FILL_5__518_ (
);

FILL FILL_0__609_ (
);

FILL FILL_7__420_ (
);

FILL FILL_0__362_ (
);

AND2X2 _365_ (
    .A(_198_),
    .B(_200_),
    .Y(_201_)
);

FILL FILL_2__603_ (
);

FILL FILL_5__327_ (
);

FILL FILL_8__379_ (
);

FILL FILL_4_BUFX2_insert6 (
);

FILL FILL_4_BUFX2_insert7 (
);

FILL FILL_4_BUFX2_insert8 (
);

FILL FILL_4_BUFX2_insert9 (
);

FILL FILL_6__442_ (
);

FILL FILL_0__418_ (
);

FILL FILL_0__591_ (
);

FILL FILL_1__625_ (
);

FILL FILL_4__349_ (
);

AOI21X1 _594_ (
    .A(_122_),
    .B(_120_),
    .C(_123_),
    .Y(_12_)
);

FILL FILL_2__412_ (
);

FILL FILL_5__556_ (
);

FILL FILL_1__434_ (
);

FILL FILL_8__400_ (
);

FILL FILL_4__578_ (
);

FILL FILL_5__365_ (
);

FILL FILL_6__480_ (
);

FILL FILL_7__514_ (
);

FILL FILL_0__456_ (
);

INVX1 _459_ (
    .A(_276_),
    .Y(_288_)
);

FILL FILL_4__387_ (
);

FILL FILL_2__450_ (
);

FILL FILL_5__594_ (
);

FILL FILL_6__536_ (
);

FILL FILL_7__323_ (
);

FILL FILL_1__472_ (
);

FILL FILL_2__506_ (
);

FILL FILL_6_BUFX2_insert6 (
);

FILL FILL_6_BUFX2_insert7 (
);

FILL FILL_6_BUFX2_insert8 (
);

FILL FILL_6_BUFX2_insert9 (
);

FILL FILL_3__621_ (
);

FILL FILL_6__345_ (
);

FILL FILL_7__552_ (
);

FILL FILL_0__494_ (
);

FILL FILL_1__528_ (
);

INVX1 _497_ (
    .A(RdyCtl[3]),
    .Y(_42_)
);

FILL FILL_2__315_ (
);

FILL FILL_5__459_ (
);

FILL FILL_3__430_ (
);

FILL FILL_6__574_ (
);

FILL FILL_7__608_ (
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_7__361_ (
);

FILL FILL_1__337_ (
);

FILL FILL_2__544_ (
);

FILL FILL_6__383_ (
);

FILL FILL_7__417_ (
);

FILL FILL_0__359_ (
);

FILL FILL_7__590_ (
);

FILL FILL_1__566_ (
);

FILL FILL_8__532_ (
);

FILL FILL_2__353_ (
);

FILL FILL_5__497_ (
);

FILL FILL_6__439_ (
);

FILL FILL_4__502_ (
);

FILL FILL_0__588_ (
);

FILL FILL_1__375_ (
);

FILL FILL_8__341_ (
);

FILL FILL_2__409_ (
);

FILL FILL_2__582_ (
);

FILL FILL_3__524_ (
);

FILL FILL_6__668_ (
);

FILL FILL_7__455_ (
);

FILL FILL_0__397_ (
);

FILL FILL76050x64950 (
);

FILL FILL_8__570_ (
);

FILL FILL_2__391_ (
);

FILL FILL_3__333_ (
);

FILL FILL_6__477_ (
);

OR2X2 _612_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_140_)
);

FILL FILL_4__540_ (
);

FILL FILL75750x46950 (
);

FILL FILL_2__447_ (
);

FILL FILL74550x61350 (
);

FILL FILL_3__562_ (
);

NAND2X1 _421_ (
    .A(_252_),
    .B(_249_),
    .Y(_253_)
);

FILL FILL74550x28950 (
);

FILL FILL_7__493_ (
);

FILL FILL_1__469_ (
);

FILL FILL_8__435_ (
);

FILL FILL_3__618_ (
);

FILL FILL_3__371_ (
);

FILL FILL_4__405_ (
);

FILL FILL_7__549_ (
);

DFFPOSX1 _650_ (
    .D(_24_),
    .CLK(clk_bF$buf5),
    .Q(acc_reg[17])
);

FILL FILL_5__612_ (
);

FILL FILL_2__485_ (
);

FILL FILL_3__427_ (
);

FILL FILL_7__358_ (
);

FILL FILL_5__421_ (
);

FILL FILL_8__473_ (
);

FILL FILL_0__512_ (
);

AOI21X1 _515_ (
    .A(_58_),
    .B(RdyCtl[3]),
    .C(RdyCtl[2]),
    .Y(_59_)
);

FILL FILL_4__443_ (
);

FILL FILL_7__587_ (
);

FILL FILL_8__529_ (
);

FILL FILL_0__321_ (
);

FILL FILL_3__465_ (
);

AOI21X1 _324_ (
    .A(_162_),
    .B(RdyCtl_6_bF$buf3),
    .C(_163_),
    .Y(_15_)
);

FILL FILL_7__396_ (
);

FILL FILL_6__401_ (
);

FILL FILL_2__579_ (
);

FILL FILL_0__550_ (
);

OAI21X1 _553_ (
    .A(acc_reg[1]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf3),
    .Y(_87_)
);

FILL FILL_4__481_ (
);

FILL FILL_5__515_ (
);

FILL FILL_8__567_ (
);

FILL FILL75450x150 (
);

FILL FILL_2__388_ (
);

FILL FILL_0__606_ (
);

AOI21X1 _609_ (
    .A(_136_),
    .B(RdyCtl_6_bF$buf4),
    .C(_137_),
    .Y(_13_)
);

FILL FILL_4__537_ (
);

NAND3X1 _362_ (
    .A(_175_),
    .B(_181_),
    .C(_190_),
    .Y(_198_)
);

FILL FILL_2__600_ (
);

FILL FILL_5__324_ (
);

FILL FILL_0__415_ (
);

FILL FILL_3__559_ (
);

AND2X2 _418_ (
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_250_)
);

FILL FILL_1__622_ (
);

FILL FILL_4__346_ (
);

NOR2X1 _591_ (
    .A(_119_),
    .B(_116_),
    .Y(_121_)
);

FILL FILL_5__553_ (
);

FILL FILL_3__368_ (
);

DFFPOSX1 _647_ (
    .D(_21_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[14])
);

FILL FILL74850x36150 (
);

FILL FILL_1__431_ (
);

FILL FILL_4__575_ (
);

FILL FILL_5__609_ (
);

FILL FILL_5__362_ (
);

FILL FILL_7__511_ (
);

FILL FILL_0__453_ (
);

FILL FILL_3__597_ (
);

AOI21X1 _456_ (
    .A(_284_),
    .B(RdyCtl_6_bF$buf2),
    .C(_285_),
    .Y(_25_)
);

FILL FILL_4__384_ (
);

FILL FILL_5__418_ (
);

FILL FILL_5__591_ (
);

FILL FILL_6__533_ (
);

FILL FILL_0__509_ (
);

FILL FILL_7__320_ (
);

FILL FILL_2__503_ (
);

FILL FILL_6__342_ (
);

FILL FILL_0__318_ (
);

FILL FILL_0__491_ (
);

FILL FILL_1__525_ (
);

INVX1 _494_ (
    .A(Atmp[4]),
    .Y(_39_)
);

FILL FILL_5__456_ (
);

FILL FILL_6__571_ (
);

FILL FILL_7__605_ (
);

FILL FILL_0__547_ (
);

FILL FILL_1__334_ (
);

FILL FILL_4__478_ (
);

FILL FILL_2__541_ (
);

FILL FILL_6__380_ (
);

FILL FILL_7__414_ (
);

FILL FILL_0__356_ (
);

NAND2X1 _359_ (
    .A(acc_reg[12]),
    .B(_73__bF$buf4),
    .Y(_195_)
);

FILL FILL_1__563_ (
);

endmodule
