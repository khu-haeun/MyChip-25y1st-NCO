magic
tech scmos
magscale 1 3
timestamp 1569543463
<< checkpaint >>
rect -485 -485 485 550
<< metal2 >>
rect -425 425 425 490
use pad80_CDNS_704676826050$3  pad80_CDNS_704676826050$3_0
timestamp 1569543463
transform 1 0 -425 0 1 -425
box 0 0 850 850
<< end >>
