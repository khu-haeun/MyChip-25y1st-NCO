magic
tech scmos
magscale 1 3
timestamp 1569533753
<< checkpaint >>
rect -52 -52 332 108
<< pseudo_rpoly2 >>
rect 8 8 272 48
use poly2cont_CDNS_704676826057$1  poly2cont_CDNS_704676826057$1_0
timestamp 1569533753
transform 1 0 254 0 1 8
box 0 0 18 40
use poly2cont_CDNS_704676826057$1  poly2cont_CDNS_704676826057$1_1
timestamp 1569533753
transform 1 0 8 0 1 8
box 0 0 18 40
<< end >>
