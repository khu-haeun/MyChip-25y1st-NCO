/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module nco(
    output [11:0] Dout,
    input En,
    input [19:0] FCW,
    output Vld,
    input clk,
    input selSign,
    input selXY
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire \genblk1[0].u_ce.Vld_bF$buf4  ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire [1:0] \a[5]  ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire \genblk1[2].u_ce.Vld_bF$buf0  ;
wire [1:0] \genblk1[2].u_ce.Y_  ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _7004_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire \u_ot.ISreg_bF$buf3  ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire [1:0] \genblk1[5].u_ce.Yin0  ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _7042_ ;
wire _6833__bF$buf0 ;
wire _6833__bF$buf1 ;
wire _6833__bF$buf2 ;
wire _6833__bF$buf3 ;
wire _6833__bF$buf4 ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6771_ ;
wire _6351_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf1  ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf2  ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire [1:0] \genblk1[2].u_ce.Xin1  ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire \genblk1[0].u_ce.Vld_bF$buf1  ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7001_ ;
wire [11:0] \u_pa.Atmp  ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire \u_ot.ISreg_bF$buf0  ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire \genblk1[2].u_ce.ISout  ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire [11:0] \genblk1[5].u_ce.Xcalc  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6956_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _1834__bF$buf0 ;
wire _1834__bF$buf1 ;
wire _1834__bF$buf2 ;
wire _1834__bF$buf3 ;
wire _1834__bF$buf4 ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf2  ;
wire _4925_ ;
wire _4505_ ;
wire \genblk1[5].u_ce.Vld_bF$buf2  ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _3524__bF$buf0 ;
wire _3524__bF$buf1 ;
wire _3524__bF$buf2 ;
wire _3524__bF$buf3 ;
wire _3524__bF$buf4 ;
wire _3524__bF$buf5 ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5151__bF$buf0 ;
wire _5151__bF$buf1 ;
wire _5151__bF$buf2 ;
wire _5151__bF$buf3 ;
wire _5151__bF$buf4 ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _197_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf1  ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire \u_ot.ISreg  ;
wire _6821_ ;
wire _6401_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire [11:0] \u_ot.Xcalc  ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire [1:0] \genblk1[0].u_ce.Ain1  ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire [1:0] \genblk1[3].u_ce.Y_  ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf2  ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _7033_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf3  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire [11:0] \genblk1[0].u_ce.Yin12b  ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire [1:0] \genblk1[1].u_ce.Xin0  ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire [11:0] _7071_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _158__bF$buf0 ;
wire _158__bF$buf1 ;
wire _158__bF$buf2 ;
wire _158__bF$buf3 ;
wire _158__bF$buf4 ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire [11:0] \genblk1[2].u_ce.Yin12b  ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire \genblk1[2].u_ce.Vld  ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _7068_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire [11:0] \genblk1[4].u_ce.Yin12b  ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire [1:0] \a[0]  ;
wire _2679_ ;
wire _2259_ ;
wire [1:0] \genblk1[3].u_ce.Yin1  ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire [1:0] \genblk1[6].u_ce.Ain0  ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire [11:0] \u_ot.Yin12b  ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire [11:0] \genblk1[6].u_ce.Yin12b  ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _4348__bF$buf0 ;
wire _4348__bF$buf1 ;
wire _4348__bF$buf2 ;
wire _4348__bF$buf3 ;
wire _4348__bF$buf4 ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _6912_ ;
wire _2832_ ;
wire _2412_ ;
wire [11:0] \genblk1[7].u_ce.Ycalc  ;
wire _3617_ ;
wire _6089_ ;
wire _7030_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf0  ;
wire _6721_ ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire En_bF$buf0 ;
wire En_bF$buf1 ;
wire En_bF$buf2 ;
wire En_bF$buf3 ;
wire En_bF$buf4 ;
wire _5704_ ;
wire \genblk1[3].u_ce.Vld_bF$buf2  ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _973__bF$buf0 ;
wire _973__bF$buf1 ;
wire _973__bF$buf2 ;
wire _973__bF$buf3 ;
wire _973__bF$buf4 ;
wire _6718_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf1  ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _7065_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire [11:0] \genblk1[2].u_ce.Xcalc  ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire \genblk1[7].u_ce.Vld  ;
wire _896_ ;
wire [6:0] \genblk1[1].u_ce.LoadCtl  ;
wire _476_ ;
wire _3711_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf2  ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire [1:0] \genblk1[6].u_ce.Xin1  ;
wire _5683_ ;
wire _5263_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf3  ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _6812_ ;
wire _2732_ ;
wire _2312_ ;
wire \genblk1[1].u_ce.Vld_bF$buf3  ;
wire _3937_ ;
wire _3517_ ;
wire [1:0] \a[7]  ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire [1:0] \genblk1[4].u_ce.Y_  ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _39_ ;
wire _6906_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _7024_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _2649__bF$buf0 ;
wire _2649__bF$buf1 ;
wire _2649__bF$buf2 ;
wire _2649__bF$buf3 ;
wire _2649__bF$buf4 ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire \genblk1[6].u_ce.ISout  ;
wire _3649_ ;
wire _3229_ ;
wire _7062_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire [1:0] \genblk1[2].u_ce.Yin0  ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _172__bF$buf0 ;
wire _244_ ;
wire _172__bF$buf1 ;
wire _172__bF$buf2 ;
wire _172__bF$buf3 ;
wire _172__bF$buf4 ;
wire _172__bF$buf5 ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire [6:0] \u_pa.RdyCtl  ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf0  ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _7059_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _2672__bF$buf0 ;
wire _2672__bF$buf1 ;
wire _2672__bF$buf2 ;
wire _2672__bF$buf3 ;
wire _2672__bF$buf4 ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire selXY ;
wire _4625_ ;
wire _4205_ ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire \genblk1[1].u_ce.Vld_bF$buf0  ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire selSign ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf3  ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _6903_ ;
wire _4090_ ;
wire _4362__bF$buf0 ;
wire _4362__bF$buf1 ;
wire _2823_ ;
wire _4362__bF$buf2 ;
wire _2403_ ;
wire _4362__bF$buf3 ;
wire _4362__bF$buf4 ;
wire _4362__bF$buf5 ;
wire _5295_ ;
wire _3608_ ;
wire _7021_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf2  ;
wire _5601_ ;
wire [1:0] \genblk1[4].u_ce.Ain1  ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire [11:0] \genblk1[4].u_ce.Ycalc  ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf3  ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire [1:0] \genblk1[5].u_ce.Xin0  ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire [11:0] \genblk1[5].u_ce.Acalc  ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7056_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire \genblk1[0].u_ce.Vld  ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf0  ;
wire \genblk1[6].u_ce.Vld_bF$buf1  ;
wire [1:0] \genblk1[7].u_ce.Yin1  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _6900_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire [1:0] \u_ot.Yin1  ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _6803_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf0  ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire [1:0] \genblk1[5].u_ce.Y_  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _7053_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire [11:0] \genblk1[1].u_ce.Yin12b  ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \u_ot.LoadCtl_6_bF$buf4  ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf3  ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire \genblk1[4].u_ce.Vld_bF$buf2  ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire \genblk1[3].u_ce.ISout  ;
wire _4713_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire [11:0] \genblk1[6].u_ce.Xcalc  ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire En ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf2  ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire [1:0] \a[2]  ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire \genblk1[5].u_ce.Vld  ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire _2088_ ;
wire _5174__bF$buf0 ;
wire _5174__bF$buf1 ;
wire _5174__bF$buf2 ;
wire _5174__bF$buf3 ;
wire _5174__bF$buf4 ;
wire [1:0] \genblk1[0].u_ce.Yin1  ;
wire \genblk1[0].u_ce.Rdy_bF$buf2  ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire [1:0] \genblk1[3].u_ce.Ain0  ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire [1:0] \genblk1[0].u_ce.X_  ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf3  ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _7012_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf4  ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _7050_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire \u_ot.LoadCtl_6_bF$buf1  ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf0  ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire [6:0] \genblk1[3].u_ce.LoadCtl  ;
wire _690_ ;
wire _270_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _6929_ ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire [1:0] \genblk1[6].u_ce.Yin0  ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _7047_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire [11:0] \genblk1[1].u_ce.Ycalc  ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _3487__bF$buf0 ;
wire _3487__bF$buf1 ;
wire _3487__bF$buf2 ;
wire _3487__bF$buf3 ;
wire _3487__bF$buf4 ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf0  ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf1  ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _1679_ ;
wire _1259_ ;
wire [1:0] \genblk1[3].u_ce.Xin1  ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _6603_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire \genblk1[2].u_ce.Vld_bF$buf2  ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire [11:0] \genblk1[6].u_ce.Ain12b  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire [1:0] \genblk1[6].u_ce.Y_  ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _7044_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _6773_ ;
wire _6353_ ;
wire _2693_ ;
wire _2273_ ;
wire _996__bF$buf0 ;
wire _996__bF$buf1 ;
wire _996__bF$buf2 ;
wire _996__bF$buf3 ;
wire _996__bF$buf4 ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf3  ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire [11:0] Dout ;
wire _5909_ ;
wire _3096_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf4  ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire \genblk1[0].u_ce.ISout  ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire \genblk1[0].u_ce.Vld_bF$buf3  ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire [11:0] \genblk1[3].u_ce.Xcalc  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire [1:0] \genblk1[1].u_ce.X_  ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7003_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire \u_ot.ISreg_bF$buf2  ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _7041_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf0  ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire [1:0] \genblk1[1].u_ce.Ain1  ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf1  ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire \genblk1[7].u_ce.ISout  ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire [1:0] \genblk1[2].u_ce.Xin0  ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire \genblk1[0].u_ce.Vld_bF$buf0  ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf4  ;
wire _4927_ ;
wire _4507_ ;
wire \genblk1[5].u_ce.Vld_bF$buf4  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7000_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire [1:0] \genblk1[4].u_ce.Yin1  ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire \genblk1[3].u_ce.Vld  ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _199_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf3  ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _6823_ ;
wire _6403_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire [1:0] \genblk1[7].u_ce.Y_  ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire [11:0] \genblk1[5].u_ce.Ycalc  ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf1  ;
wire _4924_ ;
wire _4504_ ;
wire \genblk1[5].u_ce.Vld_bF$buf1  ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire [11:0] \genblk1[6].u_ce.Acalc  ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _1810__bF$buf0 ;
wire _1810__bF$buf1 ;
wire _1810__bF$buf2 ;
wire _1810__bF$buf3 ;
wire _1810__bF$buf4 ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire [6:0] \genblk1[0].u_ce.LoadCtl  ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _196_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf0  ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire [1:0] \a[4]  ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire [19:0] \u_pa.acc_reg  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire [1:0] \genblk1[2].u_ce.X_  ;
wire [1:0] \genblk1[7].u_ce.Xin1  ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire [1:0] \genblk1[0].u_ce.Ain0  ;
wire _1188_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf1  ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire [6:0] \genblk1[5].u_ce.LoadCtl  ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _6914_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire [11:0] \genblk1[0].u_ce.Xcalc  ;
wire _7032_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf2  ;
wire _6723_ ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire [1:0] \u_ot.Xin1  ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _7070_ ;
wire _5803_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _2686__bF$buf0 ;
wire _2686__bF$buf1 ;
wire _2686__bF$buf2 ;
wire _2686__bF$buf3 ;
wire _2686__bF$buf4 ;
wire _2686__bF$buf5 ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire \genblk1[3].u_ce.Vld_bF$buf4  ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf3  ;
wire _5744_ ;
wire _5324_ ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _7067_ ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire [1:0] \genblk1[3].u_ce.Yin0  ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire _134__bF$buf0 ;
wire clk_bF$buf76 ;
wire _134__bF$buf1 ;
wire clk_bF$buf77 ;
wire _134__bF$buf2 ;
wire clk_bF$buf78 ;
wire _134__bF$buf3 ;
wire _134__bF$buf4 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire [11:0] \genblk1[1].u_ce.Ain12b  ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire \genblk1[4].u_ce.ISout  ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [11:0] \genblk1[3].u_ce.Ain12b  ;
wire _1185_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire [11:0] \genblk1[7].u_ce.Xcalc  ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _6911_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire [1:0] \genblk1[0].u_ce.Xin1  ;
wire [11:0] \genblk1[5].u_ce.Ain12b  ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire \genblk1[0].u_ce.ISin  ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _4324__bF$buf0 ;
wire _4324__bF$buf1 ;
wire _4324__bF$buf2 ;
wire _4324__bF$buf3 ;
wire _4324__bF$buf4 ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire [11:0] \genblk1[7].u_ce.Ain12b  ;
wire _5703_ ;
wire \genblk1[3].u_ce.Vld_bF$buf1  ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _5949__bF$buf0 ;
wire _5949__bF$buf1 ;
wire _5949__bF$buf2 ;
wire _5949__bF$buf3 ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire [19:0] FCW ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf0  ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _7064_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire [1:0] \genblk1[5].u_ce.Ain1  ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf1  ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire [1:0] \genblk1[6].u_ce.Xin0  ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf2  ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire [11:0] \genblk1[2].u_ce.Ycalc  ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire [11:0] \genblk1[7].u_ce.Xin12b  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire [11:0] \genblk1[3].u_ce.Acalc  ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _2731_ ;
wire _2311_ ;
wire \genblk1[1].u_ce.Vld_bF$buf2  ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire [1:0] \genblk1[3].u_ce.X_  ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _3510__bF$buf0 ;
wire _3510__bF$buf1 ;
wire _3510__bF$buf2 ;
wire _3510__bF$buf3 ;
wire _3510__bF$buf4 ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7023_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire \genblk1[1].u_ce.Vld  ;
wire _6714_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _7061_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _7058_ ;
wire _2193_ ;
wire \genblk1[0].u_ce.Rdy  ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _5829_ ;
wire _5409_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf2  ;
wire \genblk1[6].u_ce.Vld_bF$buf3  ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _6902_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7020_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire \genblk1[1].u_ce.ISout  ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire [1:0] \genblk1[1].u_ce.Yin1  ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf1  ;
wire _4239_ ;
wire _5600_ ;
wire [1:0] \genblk1[4].u_ce.Ain0  ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire [11:0] \genblk1[4].u_ce.Xcalc  ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf2  ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _7055_ ;
wire _2190_ ;
wire _3395_ ;
wire _5963__bF$buf0 ;
wire _5963__bF$buf1 ;
wire _5963__bF$buf2 ;
wire _5963__bF$buf3 ;
wire _5963__bF$buf4 ;
wire _5963__bF$buf5 ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _4621_ ;
wire _4201_ ;
wire [6:0] \genblk1[2].u_ce.LoadCtl  ;
wire _5826_ ;
wire _5406_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire \genblk1[4].u_ce.Vld_bF$buf4  ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire \genblk1[6].u_ce.Vld_bF$buf0  ;
wire _1649_ ;
wire _1229_ ;
wire [1:0] \genblk1[7].u_ce.Yin0  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire [6:0] \genblk1[7].u_ce.LoadCtl  ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire [1:0] \u_ot.Yin0  ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf4  ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire [1:0] \a[6]  ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire [1:0] \genblk1[4].u_ce.X_  ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7014_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire [1:0] \genblk1[4].u_ce.Xin1  ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire [11:0] \genblk1[0].u_ce.Acalc  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _7052_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \u_ot.LoadCtl_6_bF$buf3  ;
wire _3677_ ;
wire _3257_ ;
wire _5823_ ;
wire _5403_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf2  ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire \genblk1[4].u_ce.Vld_bF$buf1  ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire [11:0] \genblk1[0].u_ce.Ain12b  ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _7049_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf1  ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire [11:0] \genblk1[2].u_ce.Ain12b  ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire [11:0] \genblk1[6].u_ce.Ycalc  ;
wire [1:0] \genblk1[0].u_ce.Yin0  ;
wire \genblk1[0].u_ce.Rdy_bF$buf1  ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf2  ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire [11:0] \genblk1[4].u_ce.Ain12b  ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _7011_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf3  ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _5150__bF$buf0 ;
wire _5150__bF$buf1 ;
wire _5150__bF$buf2 ;
wire _5150__bF$buf3 ;
wire _5150__bF$buf4 ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1848__bF$buf0 ;
wire _1848__bF$buf1 ;
wire _1848__bF$buf2 ;
wire _1848__bF$buf3 ;
wire _1848__bF$buf4 ;
wire _1848__bF$buf5 ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire \u_ot.LoadCtl_6_bF$buf0  ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire \genblk1[2].u_ce.Vld_bF$buf4  ;
wire [11:0] \genblk1[2].u_ce.Xin12b  ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _5723_ ;
wire _5303_ ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _6562__bF$buf0 ;
wire _6562__bF$buf1 ;
wire _6562__bF$buf2 ;
wire _6562__bF$buf3 ;
wire _6562__bF$buf4 ;
wire [11:0] \genblk1[1].u_ce.Xcalc  ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7046_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire [11:0] \genblk1[4].u_ce.Xin12b  ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire Vld ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire [1:0] \genblk1[2].u_ce.Ain1  ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire _3098_ ;
wire [11:0] \genblk1[6].u_ce.Xin12b  ;
wire _5664_ ;
wire _5244_ ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf0  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _1678_ ;
wire _1258_ ;
wire [1:0] \genblk1[3].u_ce.Xin0  ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire \genblk1[2].u_ce.Vld_bF$buf1  ;
wire [1:0] \genblk1[5].u_ce.X_  ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire \u_ot.ISreg_bF$buf4  ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire [1:0] \genblk1[5].u_ce.Yin1  ;
wire _2425_ ;
wire _2005_ ;
wire _7043_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf2  ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf3  ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire [1:0] \a[1]  ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _972__bF$buf0 ;
wire _972__bF$buf1 ;
wire _972__bF$buf2 ;
wire _972__bF$buf3 ;
wire _972__bF$buf4 ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6998_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire \genblk1[0].u_ce.Vld_bF$buf2  ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7002_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [11:0] \genblk1[3].u_ce.Ycalc  ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire \u_ot.ISreg_bF$buf1  ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7040_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire [11:0] \genblk1[4].u_ce.Acalc  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire [6:0] \genblk1[4].u_ce.LoadCtl  ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire [1:0] \genblk1[1].u_ce.Ain0  ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf0  ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _2648__bF$buf0 ;
wire _2648__bF$buf1 ;
wire _4641_ ;
wire _2648__bF$buf2 ;
wire _4221_ ;
wire _2648__bF$buf3 ;
wire _2648__bF$buf4 ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf3  ;
wire _4926_ ;
wire _4506_ ;
wire \genblk1[5].u_ce.Vld_bF$buf3  ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire [1:0] \genblk1[4].u_ce.Yin0  ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _198_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf2  ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire [1:0] \genblk1[6].u_ce.X_  ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire [11:0] \u_ot.Ycalc  ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf3  ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _7034_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf4  ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire [1:0] \genblk1[1].u_ce.Xin1  ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf0  ;
wire _4923_ ;
wire _4503_ ;
wire \genblk1[5].u_ce.Vld_bF$buf0  ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _7069_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire [1:0] \genblk1[6].u_ce.Ain1  ;
wire _5784_ ;
wire _5364_ ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire [1:0] \genblk1[7].u_ce.Xin0  ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire \genblk1[7].u_ce.Ain12b_11_bF$buf0  ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _6913_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _7031_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf1  ;
wire _6722_ ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire [1:0] \u_ot.Xin0  ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire [11:0] \genblk1[1].u_ce.Xin12b  ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire [11:0] \genblk1[0].u_ce.Ycalc  ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire [11:0] \genblk1[3].u_ce.Xin12b  ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire \genblk1[3].u_ce.Vld_bF$buf3  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire [11:0] \genblk1[1].u_ce.Acalc  ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf2  ;
wire _5743_ ;
wire _5323_ ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _7066_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire [11:0] \genblk1[5].u_ce.Xin12b  ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf3  ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf4  ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _6910_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire [1:0] \genblk1[0].u_ce.Xin0  ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire \genblk1[1].u_ce.Vld_bF$buf4  ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire [1:0] \genblk1[7].u_ce.X_  ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire \genblk1[3].u_ce.Vld_bF$buf0  ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _7063_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire [1:0] \genblk1[2].u_ce.Yin1  ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _5605_ ;
wire [1:0] \genblk1[5].u_ce.Ain0  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _5188__bF$buf0 ;
wire _5188__bF$buf1 ;
wire _5188__bF$buf2 ;
wire _5188__bF$buf3 ;
wire _5188__bF$buf4 ;
wire _5188__bF$buf5 ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf0  ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _5925__bF$buf0 ;
wire _5925__bF$buf1 ;
wire _5925__bF$buf2 ;
wire _5925__bF$buf3 ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf1  ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire [1:0] \a[3]  ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _3486__bF$buf0 ;
wire _3486__bF$buf1 ;
wire _3486__bF$buf2 ;
wire _6598_ ;
wire _3486__bF$buf3 ;
wire _6178_ ;
wire _3486__bF$buf4 ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire \genblk1[1].u_ce.Vld_bF$buf1  ;
wire _3935_ ;
wire _3515_ ;
wire [6:0] \genblk1[6].u_ce.LoadCtl  ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _1598_ ;
wire _1178_ ;
wire [1:0] \genblk1[0].u_ce.Y_  ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _6904_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7022_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _7060_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire \genblk1[6].u_ce.Vld  ;
wire _6751_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf3  ;
wire _5602_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf4  ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1811__bF$buf0 ;
wire _1811__bF$buf1 ;
wire _1811__bF$buf2 ;
wire _1811__bF$buf3 ;
wire _1811__bF$buf4 ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire _1845_ ;
wire [1:0] \genblk1[5].u_ce.Xin1  ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _7057_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire \genblk1[7].u_ce.LoadCtl_0_bF$buf1  ;
wire \genblk1[6].u_ce.Vld_bF$buf2  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _6901_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [1:0] \genblk1[1].u_ce.Yin0  ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf0  ;
wire _4238_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _6613_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf1  ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _135__bF$buf0 ;
wire _135__bF$buf1 ;
wire _135__bF$buf2 ;
wire _135__bF$buf3 ;
wire _135__bF$buf4 ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _7054_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _1010__bF$buf0 ;
wire _1010__bF$buf1 ;
wire _1010__bF$buf2 ;
wire _1010__bF$buf3 ;
wire _1010__bF$buf4 ;
wire _847_ ;
wire _1010__bF$buf5 ;
wire _427_ ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _2283_ ;
wire [6:0] \u_ot.LoadCtl  ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf4  ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire \genblk1[4].u_ce.Vld_bF$buf3  ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf3  ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _4325__bF$buf0 ;
wire _4325__bF$buf1 ;
wire _4325__bF$buf2 ;
wire _4325__bF$buf3 ;
wire _4325__bF$buf4 ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf3  ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire [1:0] \genblk1[3].u_ce.Ain1  ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire [1:0] \genblk1[1].u_ce.Y_  ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire [11:0] \genblk1[0].u_ce.Xin12b  ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _7013_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire [1:0] \genblk1[4].u_ce.Xin0  ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _7051_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \u_ot.LoadCtl_6_bF$buf2  ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf1  ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire \genblk1[4].u_ce.Vld_bF$buf0  ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _1645_ ;
wire _1225_ ;
wire [1:0] \genblk1[6].u_ce.Yin1  ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _7048_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire [11:0] \genblk1[3].u_ce.Yin12b  ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf0  ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire [11:0] \u_ot.Xin12b  ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire \genblk1[0].u_ce.Rdy_bF$buf0  ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire [11:0] \genblk1[5].u_ce.Yin12b  ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf1  ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7010_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf2  ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire [11:0] \genblk1[7].u_ce.Yin12b  ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire \genblk1[5].u_ce.ISout  ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire \genblk1[2].u_ce.Vld_bF$buf3  ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire _5926__bF$buf0 ;
wire _5926__bF$buf1 ;
wire _5926__bF$buf2 ;
wire _5926__bF$buf3 ;
wire _5926__bF$buf4 ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7045_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire \genblk1[4].u_ce.Vld  ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire [1:0] \genblk1[2].u_ce.Ain0  ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire [11:0] \genblk1[2].u_ce.Acalc  ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;

CLKBUF1 CLKBUF1_insert391 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert390 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert389 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert388 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert387 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert386 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert385 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert384 (
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

BUFX2 BUFX2_insert383 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert382 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert381 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert380 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert379 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert378 (
    .A(_973_),
    .Y(_973__bF$buf0)
);

BUFX2 BUFX2_insert377 (
    .A(_973_),
    .Y(_973__bF$buf1)
);

BUFX2 BUFX2_insert376 (
    .A(_973_),
    .Y(_973__bF$buf2)
);

BUFX2 BUFX2_insert375 (
    .A(_973_),
    .Y(_973__bF$buf3)
);

BUFX2 BUFX2_insert374 (
    .A(_973_),
    .Y(_973__bF$buf4)
);

BUFX2 BUFX2_insert373 (
    .A(_6833_),
    .Y(_6833__bF$buf0)
);

BUFX2 BUFX2_insert372 (
    .A(_6833_),
    .Y(_6833__bF$buf1)
);

BUFX2 BUFX2_insert371 (
    .A(_6833_),
    .Y(_6833__bF$buf2)
);

BUFX2 BUFX2_insert370 (
    .A(_6833_),
    .Y(_6833__bF$buf3)
);

BUFX2 BUFX2_insert369 (
    .A(_6833_),
    .Y(_6833__bF$buf4)
);

BUFX2 BUFX2_insert368 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert367 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert366 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert365 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert364 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert363 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert362 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert361 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert360 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert359 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert358 (
    .A(_5963_),
    .Y(_5963__bF$buf0)
);

BUFX2 BUFX2_insert357 (
    .A(_5963_),
    .Y(_5963__bF$buf1)
);

BUFX2 BUFX2_insert356 (
    .A(_5963_),
    .Y(_5963__bF$buf2)
);

BUFX2 BUFX2_insert355 (
    .A(_5963_),
    .Y(_5963__bF$buf3)
);

BUFX2 BUFX2_insert354 (
    .A(_5963_),
    .Y(_5963__bF$buf4)
);

BUFX2 BUFX2_insert353 (
    .A(_5963_),
    .Y(_5963__bF$buf5)
);

BUFX2 BUFX2_insert352 (
    .A(_5925_),
    .Y(_5925__bF$buf0)
);

BUFX2 BUFX2_insert351 (
    .A(_5925_),
    .Y(_5925__bF$buf1)
);

BUFX2 BUFX2_insert350 (
    .A(_5925_),
    .Y(_5925__bF$buf2)
);

BUFX2 BUFX2_insert349 (
    .A(_5925_),
    .Y(_5925__bF$buf3)
);

BUFX2 BUFX2_insert348 (
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert347 (
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert346 (
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert345 (
    .A(\genblk1[6].u_ce.Vld ),
    .Y(\genblk1[6].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert344 (
    .A(_1810_),
    .Y(_1810__bF$buf0)
);

BUFX2 BUFX2_insert343 (
    .A(_1810_),
    .Y(_1810__bF$buf1)
);

BUFX2 BUFX2_insert342 (
    .A(_1810_),
    .Y(_1810__bF$buf2)
);

BUFX2 BUFX2_insert341 (
    .A(_1810_),
    .Y(_1810__bF$buf3)
);

BUFX2 BUFX2_insert340 (
    .A(_1810_),
    .Y(_1810__bF$buf4)
);

BUFX2 BUFX2_insert339 (
    .A(_1848_),
    .Y(_1848__bF$buf0)
);

BUFX2 BUFX2_insert338 (
    .A(_1848_),
    .Y(_1848__bF$buf1)
);

BUFX2 BUFX2_insert337 (
    .A(_1848_),
    .Y(_1848__bF$buf2)
);

BUFX2 BUFX2_insert336 (
    .A(_1848_),
    .Y(_1848__bF$buf3)
);

BUFX2 BUFX2_insert335 (
    .A(_1848_),
    .Y(_1848__bF$buf4)
);

BUFX2 BUFX2_insert334 (
    .A(_1848_),
    .Y(_1848__bF$buf5)
);

BUFX2 BUFX2_insert333 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert332 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert331 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert330 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert329 (
    .A(_3524_),
    .Y(_3524__bF$buf0)
);

BUFX2 BUFX2_insert328 (
    .A(_3524_),
    .Y(_3524__bF$buf1)
);

BUFX2 BUFX2_insert327 (
    .A(_3524_),
    .Y(_3524__bF$buf2)
);

BUFX2 BUFX2_insert326 (
    .A(_3524_),
    .Y(_3524__bF$buf3)
);

BUFX2 BUFX2_insert325 (
    .A(_3524_),
    .Y(_3524__bF$buf4)
);

BUFX2 BUFX2_insert324 (
    .A(_3524_),
    .Y(_3524__bF$buf5)
);

BUFX2 BUFX2_insert323 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert322 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert321 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert320 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert319 (
    .A(_2686_),
    .Y(_2686__bF$buf0)
);

BUFX2 BUFX2_insert318 (
    .A(_2686_),
    .Y(_2686__bF$buf1)
);

BUFX2 BUFX2_insert317 (
    .A(_2686_),
    .Y(_2686__bF$buf2)
);

BUFX2 BUFX2_insert316 (
    .A(_2686_),
    .Y(_2686__bF$buf3)
);

BUFX2 BUFX2_insert315 (
    .A(_2686_),
    .Y(_2686__bF$buf4)
);

BUFX2 BUFX2_insert314 (
    .A(_2686_),
    .Y(_2686__bF$buf5)
);

BUFX2 BUFX2_insert313 (
    .A(_2648_),
    .Y(_2648__bF$buf0)
);

BUFX2 BUFX2_insert312 (
    .A(_2648_),
    .Y(_2648__bF$buf1)
);

BUFX2 BUFX2_insert311 (
    .A(_2648_),
    .Y(_2648__bF$buf2)
);

BUFX2 BUFX2_insert310 (
    .A(_2648_),
    .Y(_2648__bF$buf3)
);

BUFX2 BUFX2_insert309 (
    .A(_2648_),
    .Y(_2648__bF$buf4)
);

BUFX2 BUFX2_insert308 (
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf0 )
);

BUFX2 BUFX2_insert307 (
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf1 )
);

BUFX2 BUFX2_insert306 (
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf2 )
);

BUFX2 BUFX2_insert305 (
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf3 )
);

BUFX2 BUFX2_insert304 (
    .A(\u_ot.LoadCtl [6]),
    .Y(\u_ot.LoadCtl_6_bF$buf4 )
);

BUFX2 BUFX2_insert303 (
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert302 (
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert301 (
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert300 (
    .A(\genblk1[7].u_ce.LoadCtl [0]),
    .Y(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert299 (
    .A(_4362_),
    .Y(_4362__bF$buf0)
);

BUFX2 BUFX2_insert298 (
    .A(_4362_),
    .Y(_4362__bF$buf1)
);

BUFX2 BUFX2_insert297 (
    .A(_4362_),
    .Y(_4362__bF$buf2)
);

BUFX2 BUFX2_insert296 (
    .A(_4362_),
    .Y(_4362__bF$buf3)
);

BUFX2 BUFX2_insert295 (
    .A(_4362_),
    .Y(_4362__bF$buf4)
);

BUFX2 BUFX2_insert294 (
    .A(_4362_),
    .Y(_4362__bF$buf5)
);

BUFX2 BUFX2_insert293 (
    .A(_5949_),
    .Y(_5949__bF$buf0)
);

BUFX2 BUFX2_insert292 (
    .A(_5949_),
    .Y(_5949__bF$buf1)
);

BUFX2 BUFX2_insert291 (
    .A(_5949_),
    .Y(_5949__bF$buf2)
);

BUFX2 BUFX2_insert290 (
    .A(_5949_),
    .Y(_5949__bF$buf3)
);

BUFX2 BUFX2_insert289 (
    .A(_4324_),
    .Y(_4324__bF$buf0)
);

BUFX2 BUFX2_insert288 (
    .A(_4324_),
    .Y(_4324__bF$buf1)
);

BUFX2 BUFX2_insert287 (
    .A(_4324_),
    .Y(_4324__bF$buf2)
);

BUFX2 BUFX2_insert286 (
    .A(_4324_),
    .Y(_4324__bF$buf3)
);

BUFX2 BUFX2_insert285 (
    .A(_4324_),
    .Y(_4324__bF$buf4)
);

BUFX2 BUFX2_insert284 (
    .A(_5150_),
    .Y(_5150__bF$buf0)
);

BUFX2 BUFX2_insert283 (
    .A(_5150_),
    .Y(_5150__bF$buf1)
);

BUFX2 BUFX2_insert282 (
    .A(_5150_),
    .Y(_5150__bF$buf2)
);

BUFX2 BUFX2_insert281 (
    .A(_5150_),
    .Y(_5150__bF$buf3)
);

BUFX2 BUFX2_insert280 (
    .A(_5150_),
    .Y(_5150__bF$buf4)
);

BUFX2 BUFX2_insert279 (
    .A(_172_),
    .Y(_172__bF$buf0)
);

BUFX2 BUFX2_insert278 (
    .A(_172_),
    .Y(_172__bF$buf1)
);

BUFX2 BUFX2_insert277 (
    .A(_172_),
    .Y(_172__bF$buf2)
);

BUFX2 BUFX2_insert276 (
    .A(_172_),
    .Y(_172__bF$buf3)
);

BUFX2 BUFX2_insert275 (
    .A(_172_),
    .Y(_172__bF$buf4)
);

BUFX2 BUFX2_insert274 (
    .A(_172_),
    .Y(_172__bF$buf5)
);

BUFX2 BUFX2_insert273 (
    .A(_134_),
    .Y(_134__bF$buf0)
);

BUFX2 BUFX2_insert272 (
    .A(_134_),
    .Y(_134__bF$buf1)
);

BUFX2 BUFX2_insert271 (
    .A(_134_),
    .Y(_134__bF$buf2)
);

BUFX2 BUFX2_insert270 (
    .A(_134_),
    .Y(_134__bF$buf3)
);

BUFX2 BUFX2_insert269 (
    .A(_134_),
    .Y(_134__bF$buf4)
);

BUFX2 BUFX2_insert268 (
    .A(_1834_),
    .Y(_1834__bF$buf0)
);

BUFX2 BUFX2_insert267 (
    .A(_1834_),
    .Y(_1834__bF$buf1)
);

BUFX2 BUFX2_insert266 (
    .A(_1834_),
    .Y(_1834__bF$buf2)
);

BUFX2 BUFX2_insert265 (
    .A(_1834_),
    .Y(_1834__bF$buf3)
);

BUFX2 BUFX2_insert264 (
    .A(_1834_),
    .Y(_1834__bF$buf4)
);

BUFX2 BUFX2_insert263 (
    .A(_5188_),
    .Y(_5188__bF$buf0)
);

BUFX2 BUFX2_insert262 (
    .A(_5188_),
    .Y(_5188__bF$buf1)
);

BUFX2 BUFX2_insert261 (
    .A(_5188_),
    .Y(_5188__bF$buf2)
);

BUFX2 BUFX2_insert260 (
    .A(_5188_),
    .Y(_5188__bF$buf3)
);

BUFX2 BUFX2_insert259 (
    .A(_5188_),
    .Y(_5188__bF$buf4)
);

BUFX2 BUFX2_insert258 (
    .A(_5188_),
    .Y(_5188__bF$buf5)
);

BUFX2 BUFX2_insert257 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert256 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert255 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert254 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert253 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert252 (
    .A(_3486_),
    .Y(_3486__bF$buf0)
);

BUFX2 BUFX2_insert251 (
    .A(_3486_),
    .Y(_3486__bF$buf1)
);

BUFX2 BUFX2_insert250 (
    .A(_3486_),
    .Y(_3486__bF$buf2)
);

BUFX2 BUFX2_insert249 (
    .A(_3486_),
    .Y(_3486__bF$buf3)
);

BUFX2 BUFX2_insert248 (
    .A(_3486_),
    .Y(_3486__bF$buf4)
);

BUFX2 BUFX2_insert247 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert246 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert245 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert244 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert243 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert242 (
    .A(_3510_),
    .Y(_3510__bF$buf0)
);

BUFX2 BUFX2_insert241 (
    .A(_3510_),
    .Y(_3510__bF$buf1)
);

BUFX2 BUFX2_insert240 (
    .A(_3510_),
    .Y(_3510__bF$buf2)
);

BUFX2 BUFX2_insert239 (
    .A(_3510_),
    .Y(_3510__bF$buf3)
);

BUFX2 BUFX2_insert238 (
    .A(_3510_),
    .Y(_3510__bF$buf4)
);

BUFX2 BUFX2_insert237 (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf0 )
);

BUFX2 BUFX2_insert236 (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf1 )
);

BUFX2 BUFX2_insert235 (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf2 )
);

BUFX2 BUFX2_insert234 (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf3 )
);

BUFX2 BUFX2_insert233 (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(\genblk1[0].u_ce.Rdy_bF$buf4 )
);

BUFX2 BUFX2_insert232 (
    .A(_5926_),
    .Y(_5926__bF$buf0)
);

BUFX2 BUFX2_insert231 (
    .A(_5926_),
    .Y(_5926__bF$buf1)
);

BUFX2 BUFX2_insert230 (
    .A(_5926_),
    .Y(_5926__bF$buf2)
);

BUFX2 BUFX2_insert229 (
    .A(_5926_),
    .Y(_5926__bF$buf3)
);

BUFX2 BUFX2_insert228 (
    .A(_5926_),
    .Y(_5926__bF$buf4)
);

BUFX2 BUFX2_insert227 (
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert226 (
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert225 (
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert224 (
    .A(\genblk1[7].u_ce.Ain12b [11]),
    .Y(\genblk1[7].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert223 (
    .A(_2672_),
    .Y(_2672__bF$buf0)
);

BUFX2 BUFX2_insert222 (
    .A(_2672_),
    .Y(_2672__bF$buf1)
);

BUFX2 BUFX2_insert221 (
    .A(_2672_),
    .Y(_2672__bF$buf2)
);

BUFX2 BUFX2_insert220 (
    .A(_2672_),
    .Y(_2672__bF$buf3)
);

BUFX2 BUFX2_insert219 (
    .A(_2672_),
    .Y(_2672__bF$buf4)
);

BUFX2 BUFX2_insert218 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert217 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert216 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert215 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert214 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert213 (
    .A(_1811_),
    .Y(_1811__bF$buf0)
);

BUFX2 BUFX2_insert212 (
    .A(_1811_),
    .Y(_1811__bF$buf1)
);

BUFX2 BUFX2_insert211 (
    .A(_1811_),
    .Y(_1811__bF$buf2)
);

BUFX2 BUFX2_insert210 (
    .A(_1811_),
    .Y(_1811__bF$buf3)
);

BUFX2 BUFX2_insert209 (
    .A(_1811_),
    .Y(_1811__bF$buf4)
);

BUFX2 BUFX2_insert208 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert207 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert206 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert205 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert204 (
    .A(_4348_),
    .Y(_4348__bF$buf0)
);

BUFX2 BUFX2_insert203 (
    .A(_4348_),
    .Y(_4348__bF$buf1)
);

BUFX2 BUFX2_insert202 (
    .A(_4348_),
    .Y(_4348__bF$buf2)
);

BUFX2 BUFX2_insert201 (
    .A(_4348_),
    .Y(_4348__bF$buf3)
);

BUFX2 BUFX2_insert200 (
    .A(_4348_),
    .Y(_4348__bF$buf4)
);

BUFX2 BUFX2_insert199 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert198 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert197 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert196 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert195 (
    .A(_5174_),
    .Y(_5174__bF$buf0)
);

BUFX2 BUFX2_insert194 (
    .A(_5174_),
    .Y(_5174__bF$buf1)
);

BUFX2 BUFX2_insert193 (
    .A(_5174_),
    .Y(_5174__bF$buf2)
);

BUFX2 BUFX2_insert192 (
    .A(_5174_),
    .Y(_5174__bF$buf3)
);

BUFX2 BUFX2_insert191 (
    .A(_5174_),
    .Y(_5174__bF$buf4)
);

BUFX2 BUFX2_insert190 (
    .A(_158_),
    .Y(_158__bF$buf0)
);

BUFX2 BUFX2_insert189 (
    .A(_158_),
    .Y(_158__bF$buf1)
);

BUFX2 BUFX2_insert188 (
    .A(_158_),
    .Y(_158__bF$buf2)
);

BUFX2 BUFX2_insert187 (
    .A(_158_),
    .Y(_158__bF$buf3)
);

BUFX2 BUFX2_insert186 (
    .A(_158_),
    .Y(_158__bF$buf4)
);

BUFX2 BUFX2_insert185 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert184 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert183 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert182 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert181 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert180 (
    .A(_2649_),
    .Y(_2649__bF$buf0)
);

BUFX2 BUFX2_insert179 (
    .A(_2649_),
    .Y(_2649__bF$buf1)
);

BUFX2 BUFX2_insert178 (
    .A(_2649_),
    .Y(_2649__bF$buf2)
);

BUFX2 BUFX2_insert177 (
    .A(_2649_),
    .Y(_2649__bF$buf3)
);

BUFX2 BUFX2_insert176 (
    .A(_2649_),
    .Y(_2649__bF$buf4)
);

BUFX2 BUFX2_insert175 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert174 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert173 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert172 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert171 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert170 (
    .A(_972_),
    .Y(_972__bF$buf0)
);

BUFX2 BUFX2_insert169 (
    .A(_972_),
    .Y(_972__bF$buf1)
);

BUFX2 BUFX2_insert168 (
    .A(_972_),
    .Y(_972__bF$buf2)
);

BUFX2 BUFX2_insert167 (
    .A(_972_),
    .Y(_972__bF$buf3)
);

BUFX2 BUFX2_insert166 (
    .A(_972_),
    .Y(_972__bF$buf4)
);

BUFX2 BUFX2_insert165 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert164 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert163 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert162 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert161 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert160 (
    .A(_4325_),
    .Y(_4325__bF$buf0)
);

BUFX2 BUFX2_insert159 (
    .A(_4325_),
    .Y(_4325__bF$buf1)
);

BUFX2 BUFX2_insert158 (
    .A(_4325_),
    .Y(_4325__bF$buf2)
);

BUFX2 BUFX2_insert157 (
    .A(_4325_),
    .Y(_4325__bF$buf3)
);

BUFX2 BUFX2_insert156 (
    .A(_4325_),
    .Y(_4325__bF$buf4)
);

BUFX2 BUFX2_insert155 (
    .A(_5151_),
    .Y(_5151__bF$buf0)
);

BUFX2 BUFX2_insert154 (
    .A(_5151_),
    .Y(_5151__bF$buf1)
);

BUFX2 BUFX2_insert153 (
    .A(_5151_),
    .Y(_5151__bF$buf2)
);

BUFX2 BUFX2_insert152 (
    .A(_5151_),
    .Y(_5151__bF$buf3)
);

BUFX2 BUFX2_insert151 (
    .A(_5151_),
    .Y(_5151__bF$buf4)
);

BUFX2 BUFX2_insert150 (
    .A(_135_),
    .Y(_135__bF$buf0)
);

BUFX2 BUFX2_insert149 (
    .A(_135_),
    .Y(_135__bF$buf1)
);

BUFX2 BUFX2_insert148 (
    .A(_135_),
    .Y(_135__bF$buf2)
);

BUFX2 BUFX2_insert147 (
    .A(_135_),
    .Y(_135__bF$buf3)
);

BUFX2 BUFX2_insert146 (
    .A(_135_),
    .Y(_135__bF$buf4)
);

BUFX2 BUFX2_insert145 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert144 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert143 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert142 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert141 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert140 (
    .A(En),
    .Y(En_bF$buf0)
);

BUFX2 BUFX2_insert139 (
    .A(En),
    .Y(En_bF$buf1)
);

BUFX2 BUFX2_insert138 (
    .A(En),
    .Y(En_bF$buf2)
);

BUFX2 BUFX2_insert137 (
    .A(En),
    .Y(En_bF$buf3)
);

BUFX2 BUFX2_insert136 (
    .A(En),
    .Y(En_bF$buf4)
);

BUFX2 BUFX2_insert135 (
    .A(_3487_),
    .Y(_3487__bF$buf0)
);

BUFX2 BUFX2_insert134 (
    .A(_3487_),
    .Y(_3487__bF$buf1)
);

BUFX2 BUFX2_insert133 (
    .A(_3487_),
    .Y(_3487__bF$buf2)
);

BUFX2 BUFX2_insert132 (
    .A(_3487_),
    .Y(_3487__bF$buf3)
);

BUFX2 BUFX2_insert131 (
    .A(_3487_),
    .Y(_3487__bF$buf4)
);

BUFX2 BUFX2_insert130 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert129 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert128 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert127 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert126 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert125 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert124 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert123 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert122 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert121 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert120 (
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert119 (
    .A(selXY),
    .Y(selXY_bF$buf1)
);

BUFX2 BUFX2_insert118 (
    .A(selXY),
    .Y(selXY_bF$buf2)
);

BUFX2 BUFX2_insert117 (
    .A(selXY),
    .Y(selXY_bF$buf3)
);

BUFX2 BUFX2_insert116 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert115 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert114 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert113 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert112 (
    .A(_6562_),
    .Y(_6562__bF$buf0)
);

BUFX2 BUFX2_insert111 (
    .A(_6562_),
    .Y(_6562__bF$buf1)
);

BUFX2 BUFX2_insert110 (
    .A(_6562_),
    .Y(_6562__bF$buf2)
);

BUFX2 BUFX2_insert109 (
    .A(_6562_),
    .Y(_6562__bF$buf3)
);

BUFX2 BUFX2_insert108 (
    .A(_6562_),
    .Y(_6562__bF$buf4)
);

CLKBUF1 CLKBUF1_insert107 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert106 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert105 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert104 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert103 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert102 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert101 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert100 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert99 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert98 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert97 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert96 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert95 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert94 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert93 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert92 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert91 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert90 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert89 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert88 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert87 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert86 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert85 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert84 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert83 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert82 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert81 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert80 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert79 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert78 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert77 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert76 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert75 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert74 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert73 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert72 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert71 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert70 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert69 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert68 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert67 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert66 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert65 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert64 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert63 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert62 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert61 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert60 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert59 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert58 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert57 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert56 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert55 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert54 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert53 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert52 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert51 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert50 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert49 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf58)
);

CLKBUF1 CLKBUF1_insert48 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert47 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf60)
);

CLKBUF1 CLKBUF1_insert46 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert45 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert44 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert43 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert42 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert41 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert40 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert39 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf68)
);

CLKBUF1 CLKBUF1_insert38 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert37 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert36 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert35 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert34 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert33 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert32 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf75)
);

CLKBUF1 CLKBUF1_insert31 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert30 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert29 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf78)
);

BUFX2 BUFX2_insert28 (
    .A(_1010_),
    .Y(_1010__bF$buf0)
);

BUFX2 BUFX2_insert27 (
    .A(_1010_),
    .Y(_1010__bF$buf1)
);

BUFX2 BUFX2_insert26 (
    .A(_1010_),
    .Y(_1010__bF$buf2)
);

BUFX2 BUFX2_insert25 (
    .A(_1010_),
    .Y(_1010__bF$buf3)
);

BUFX2 BUFX2_insert24 (
    .A(_1010_),
    .Y(_1010__bF$buf4)
);

BUFX2 BUFX2_insert23 (
    .A(_1010_),
    .Y(_1010__bF$buf5)
);

BUFX2 BUFX2_insert22 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert21 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert20 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert19 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert18 (
    .A(_996_),
    .Y(_996__bF$buf0)
);

BUFX2 BUFX2_insert17 (
    .A(_996_),
    .Y(_996__bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .A(_996_),
    .Y(_996__bF$buf2)
);

BUFX2 BUFX2_insert15 (
    .A(_996_),
    .Y(_996__bF$buf3)
);

BUFX2 BUFX2_insert14 (
    .A(_996_),
    .Y(_996__bF$buf4)
);

BUFX2 BUFX2_insert13 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert12 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert11 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert10 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert9 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert8 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert7 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert6 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert5 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert4 (
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf0 )
);

BUFX2 BUFX2_insert3 (
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf1 )
);

BUFX2 BUFX2_insert2 (
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf2 )
);

BUFX2 BUFX2_insert1 (
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf3 )
);

BUFX2 BUFX2_insert0 (
    .A(\u_ot.ISreg ),
    .Y(\u_ot.ISreg_bF$buf4 )
);

INVX2 _10000_ (
    .A(_2674_),
    .Y(_2741_)
);

OAI21X1 _10001_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2741_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_2742_)
);

OAI21X1 _10002_ (
    .A(_2742_),
    .B(_2740_),
    .C(_2720_),
    .Y(_2517_)
);

INVX1 _10003_ (
    .A(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2743_)
);

INVX2 _10004_ (
    .A(_2742_),
    .Y(_2744_)
);

OAI21X1 _10005_ (
    .A(_2733_),
    .B(_2721_),
    .C(_2734_),
    .Y(_2745_)
);

INVX1 _10006_ (
    .A(_2745_),
    .Y(_2746_)
);

INVX1 _10007_ (
    .A(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2747_)
);

NAND3X1 _10008_ (
    .A(_2684_),
    .B(_2709_),
    .C(_2727_),
    .Y(_2748_)
);

INVX1 _10009_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .Y(_2749_)
);

NAND2X1 _10010_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2750_)
);

OAI21X1 _10011_ (
    .A(1'h1),
    .B(_2749_),
    .C(_2750_),
    .Y(_2751_)
);

NAND2X1 _10012_ (
    .A(_2649__bF$buf4),
    .B(_2703_),
    .Y(_2752_)
);

OAI21X1 _10013_ (
    .A(_2649__bF$buf3),
    .B(_2751_),
    .C(_2752_),
    .Y(_2753_)
);

NOR2X1 _10014_ (
    .A(1'h0),
    .B(_2649__bF$buf2),
    .Y(_2754_)
);

NOR2X1 _10015_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_2755_)
);

AOI22X1 _10016_ (
    .A(_2696_),
    .B(_2755_),
    .C(_2754_),
    .D(_2692_),
    .Y(_2756_)
);

OAI21X1 _10017_ (
    .A(_2648__bF$buf4),
    .B(_2753_),
    .C(_2756_),
    .Y(_2757_)
);

NAND3X1 _10018_ (
    .A(_2686__bF$buf5),
    .B(_2757_),
    .C(_2748_),
    .Y(_2758_)
);

INVX1 _10019_ (
    .A(_2748_),
    .Y(_2759_)
);

INVX1 _10020_ (
    .A(_2757_),
    .Y(_2760_)
);

OAI21X1 _10021_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2759_),
    .C(_2760_),
    .Y(_2761_)
);

NAND3X1 _10022_ (
    .A(_2747_),
    .B(_2758_),
    .C(_2761_),
    .Y(_2762_)
);

AOI21X1 _10023_ (
    .A(_2761_),
    .B(_2758_),
    .C(_2747_),
    .Y(_2763_)
);

INVX1 _10024_ (
    .A(_2763_),
    .Y(_2764_)
);

NAND2X1 _10025_ (
    .A(_2762_),
    .B(_2764_),
    .Y(_2765_)
);

AOI21X1 _10026_ (
    .A(_2765_),
    .B(_2746_),
    .C(_2674_),
    .Y(_2766_)
);

OAI21X1 _10027_ (
    .A(_2746_),
    .B(_2765_),
    .C(_2766_),
    .Y(_2767_)
);

AOI22X1 _10028_ (
    .A(_2743_),
    .B(_2672__bF$buf4),
    .C(_2767_),
    .D(_2744_),
    .Y(_2518_)
);

AOI21X1 _10029_ (
    .A(_2745_),
    .B(_2762_),
    .C(_2763_),
    .Y(_2768_)
);

INVX1 _10030_ (
    .A(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2769_)
);

INVX1 _10031_ (
    .A(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2770_)
);

NAND2X1 _10032_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2771_)
);

OAI21X1 _10033_ (
    .A(1'h1),
    .B(_2770_),
    .C(_2771_),
    .Y(_2772_)
);

NAND2X1 _10034_ (
    .A(_2649__bF$buf1),
    .B(_2722_),
    .Y(_2773_)
);

OAI21X1 _10035_ (
    .A(_2649__bF$buf0),
    .B(_2772_),
    .C(_2773_),
    .Y(_2774_)
);

NAND2X1 _10036_ (
    .A(_2648__bF$buf3),
    .B(_2677_),
    .Y(_2775_)
);

OAI21X1 _10037_ (
    .A(_2648__bF$buf2),
    .B(_2774_),
    .C(_2775_),
    .Y(_2776_)
);

INVX2 _10038_ (
    .A(_2776_),
    .Y(_2777_)
);

OAI21X1 _10039_ (
    .A(_2757_),
    .B(_2748_),
    .C(_2686__bF$buf4),
    .Y(_2778_)
);

OR2X2 _10040_ (
    .A(_2778_),
    .B(_2777_),
    .Y(_2779_)
);

NOR2X1 _10041_ (
    .A(_2757_),
    .B(_2748_),
    .Y(_2780_)
);

OAI21X1 _10042_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2780_),
    .C(_2777_),
    .Y(_2781_)
);

NAND3X1 _10043_ (
    .A(_2769_),
    .B(_2781_),
    .C(_2779_),
    .Y(_2782_)
);

NOR2X1 _10044_ (
    .A(_2777_),
    .B(_2778_),
    .Y(_2783_)
);

AND2X2 _10045_ (
    .A(_2778_),
    .B(_2777_),
    .Y(_2784_)
);

OAI21X1 _10046_ (
    .A(_2783_),
    .B(_2784_),
    .C(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2785_)
);

NAND2X1 _10047_ (
    .A(_2785_),
    .B(_2782_),
    .Y(_2786_)
);

AOI21X1 _10048_ (
    .A(_2768_),
    .B(_2786_),
    .C(_2674_),
    .Y(_2787_)
);

OAI21X1 _10049_ (
    .A(_2768_),
    .B(_2786_),
    .C(_2787_),
    .Y(_2788_)
);

AOI22X1 _10050_ (
    .A(_2619_),
    .B(_2672__bF$buf3),
    .C(_2788_),
    .D(_2744_),
    .Y(_2519_)
);

OAI21X1 _10051_ (
    .A(_2786_),
    .B(_2768_),
    .C(_2785_),
    .Y(_2789_)
);

INVX1 _10052_ (
    .A(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_2790_)
);

NAND3X1 _10053_ (
    .A(_2760_),
    .B(_2777_),
    .C(_2759_),
    .Y(_2791_)
);

NAND2X1 _10054_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2792_)
);

INVX1 _10055_ (
    .A(_2792_),
    .Y(_2793_)
);

AOI21X1 _10056_ (
    .A(_2751_),
    .B(_2649__bF$buf4),
    .C(_2793_),
    .Y(_2794_)
);

NAND2X1 _10057_ (
    .A(_2648__bF$buf1),
    .B(_2705_),
    .Y(_2795_)
);

OAI21X1 _10058_ (
    .A(_2648__bF$buf0),
    .B(_2794_),
    .C(_2795_),
    .Y(_2796_)
);

NAND3X1 _10059_ (
    .A(_2686__bF$buf3),
    .B(_2796_),
    .C(_2791_),
    .Y(_2797_)
);

NOR3X1 _10060_ (
    .A(_2757_),
    .B(_2776_),
    .C(_2748_),
    .Y(_2798_)
);

INVX1 _10061_ (
    .A(_2796_),
    .Y(_2799_)
);

OAI21X1 _10062_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2798_),
    .C(_2799_),
    .Y(_2800_)
);

NAND3X1 _10063_ (
    .A(_2790_),
    .B(_2797_),
    .C(_2800_),
    .Y(_2801_)
);

AOI21X1 _10064_ (
    .A(_2800_),
    .B(_2797_),
    .C(_2790_),
    .Y(_2802_)
);

INVX1 _10065_ (
    .A(_2802_),
    .Y(_2803_)
);

NAND2X1 _10066_ (
    .A(_2801_),
    .B(_2803_),
    .Y(_2804_)
);

AND2X2 _10067_ (
    .A(_2789_),
    .B(_2804_),
    .Y(_2805_)
);

OAI21X1 _10068_ (
    .A(_2804_),
    .B(_2789_),
    .C(_2741_),
    .Y(_2806_)
);

OAI21X1 _10069_ (
    .A(_2806_),
    .B(_2805_),
    .C(_2744_),
    .Y(_2807_)
);

OAI21X1 _10070_ (
    .A(_2627_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_2807_),
    .Y(_2520_)
);

INVX1 _10071_ (
    .A(\genblk1[3].u_ce.Ycalc [6]),
    .Y(_2808_)
);

INVX1 _10072_ (
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2809_)
);

NAND3X1 _10073_ (
    .A(_2777_),
    .B(_2799_),
    .C(_2780_),
    .Y(_2810_)
);

AOI21X1 _10074_ (
    .A(_2772_),
    .B(_2649__bF$buf3),
    .C(_2793_),
    .Y(_2811_)
);

NAND2X1 _10075_ (
    .A(_2648__bF$buf4),
    .B(_2723_),
    .Y(_2812_)
);

OAI21X1 _10076_ (
    .A(_2648__bF$buf3),
    .B(_2811_),
    .C(_2812_),
    .Y(_2813_)
);

NAND3X1 _10077_ (
    .A(_2686__bF$buf2),
    .B(_2813_),
    .C(_2810_),
    .Y(_2814_)
);

INVX1 _10078_ (
    .A(_2813_),
    .Y(_2815_)
);

OAI21X1 _10079_ (
    .A(_2796_),
    .B(_2791_),
    .C(_2686__bF$buf1),
    .Y(_2816_)
);

NAND2X1 _10080_ (
    .A(_2815_),
    .B(_2816_),
    .Y(_2817_)
);

NAND3X1 _10081_ (
    .A(_2809_),
    .B(_2814_),
    .C(_2817_),
    .Y(_2818_)
);

NAND3X1 _10082_ (
    .A(_2686__bF$buf0),
    .B(_2815_),
    .C(_2810_),
    .Y(_2819_)
);

NAND2X1 _10083_ (
    .A(_2813_),
    .B(_2816_),
    .Y(_2820_)
);

NAND3X1 _10084_ (
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .B(_2819_),
    .C(_2820_),
    .Y(_2821_)
);

NAND2X1 _10085_ (
    .A(_2818_),
    .B(_2821_),
    .Y(_2822_)
);

AOI21X1 _10086_ (
    .A(_2779_),
    .B(_2781_),
    .C(_2769_),
    .Y(_2823_)
);

NOR2X1 _10087_ (
    .A(_2823_),
    .B(_2802_),
    .Y(_2824_)
);

OAI21X1 _10088_ (
    .A(_2786_),
    .B(_2768_),
    .C(_2824_),
    .Y(_2825_)
);

NAND2X1 _10089_ (
    .A(_2801_),
    .B(_2825_),
    .Y(_2826_)
);

AOI21X1 _10090_ (
    .A(_2826_),
    .B(_2822_),
    .C(_2674_),
    .Y(_2827_)
);

OAI21X1 _10091_ (
    .A(_2822_),
    .B(_2826_),
    .C(_2827_),
    .Y(_2828_)
);

AOI22X1 _10092_ (
    .A(_2808_),
    .B(_2672__bF$buf2),
    .C(_2828_),
    .D(_2744_),
    .Y(_2521_)
);

INVX1 _10093_ (
    .A(\genblk1[3].u_ce.Ycalc [7]),
    .Y(_2829_)
);

AOI21X1 _10094_ (
    .A(_2817_),
    .B(_2814_),
    .C(_2809_),
    .Y(_2830_)
);

AND2X2 _10095_ (
    .A(_2782_),
    .B(_2785_),
    .Y(_2831_)
);

NAND3X1 _10096_ (
    .A(_2801_),
    .B(_2803_),
    .C(_2831_),
    .Y(_2832_)
);

AOI21X1 _10097_ (
    .A(_2823_),
    .B(_2801_),
    .C(_2802_),
    .Y(_2833_)
);

OAI21X1 _10098_ (
    .A(_2768_),
    .B(_2832_),
    .C(_2833_),
    .Y(_2834_)
);

AOI21X1 _10099_ (
    .A(_2834_),
    .B(_2818_),
    .C(_2830_),
    .Y(_2835_)
);

INVX1 _10100_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2836_)
);

NAND3X1 _10101_ (
    .A(_2799_),
    .B(_2815_),
    .C(_2798_),
    .Y(_2837_)
);

INVX1 _10102_ (
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2838_)
);

NOR2X1 _10103_ (
    .A(_2648__bF$buf2),
    .B(_2838_),
    .Y(_2839_)
);

INVX1 _10104_ (
    .A(_2839_),
    .Y(_2840_)
);

OAI21X1 _10105_ (
    .A(1'h0),
    .B(_2753_),
    .C(_2840_),
    .Y(_2841_)
);

NAND3X1 _10106_ (
    .A(_2686__bF$buf5),
    .B(_2841_),
    .C(_2837_),
    .Y(_2842_)
);

INVX1 _10107_ (
    .A(_2841_),
    .Y(_2843_)
);

OAI21X1 _10108_ (
    .A(_2813_),
    .B(_2810_),
    .C(_2686__bF$buf4),
    .Y(_2844_)
);

NAND2X1 _10109_ (
    .A(_2843_),
    .B(_2844_),
    .Y(_2845_)
);

NAND3X1 _10110_ (
    .A(_2836_),
    .B(_2842_),
    .C(_2845_),
    .Y(_2846_)
);

NAND3X1 _10111_ (
    .A(_2686__bF$buf3),
    .B(_2843_),
    .C(_2837_),
    .Y(_2847_)
);

NAND2X1 _10112_ (
    .A(_2841_),
    .B(_2844_),
    .Y(_2848_)
);

NAND3X1 _10113_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(_2847_),
    .C(_2848_),
    .Y(_2849_)
);

NAND2X1 _10114_ (
    .A(_2846_),
    .B(_2849_),
    .Y(_2850_)
);

INVX1 _10115_ (
    .A(_2850_),
    .Y(_2851_)
);

NOR2X1 _10116_ (
    .A(_2851_),
    .B(_2835_),
    .Y(_2852_)
);

OAI21X1 _10117_ (
    .A(_2822_),
    .B(_2826_),
    .C(_2821_),
    .Y(_2853_)
);

OAI21X1 _10118_ (
    .A(_2850_),
    .B(_2853_),
    .C(_2741_),
    .Y(_2854_)
);

OAI21X1 _10119_ (
    .A(_2686__bF$buf2),
    .B(_2741_),
    .C(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .Y(_2855_)
);

INVX1 _10120_ (
    .A(_2855_),
    .Y(_2856_)
);

OAI21X1 _10121_ (
    .A(_2854_),
    .B(_2852_),
    .C(_2856_),
    .Y(_2857_)
);

OAI21X1 _10122_ (
    .A(_2829_),
    .B(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .C(_2857_),
    .Y(_2522_)
);

INVX1 _10123_ (
    .A(\genblk1[3].u_ce.Ycalc [8]),
    .Y(_2858_)
);

OAI21X1 _10124_ (
    .A(_2821_),
    .B(_2850_),
    .C(_2849_),
    .Y(_2859_)
);

NOR2X1 _10125_ (
    .A(_2822_),
    .B(_2850_),
    .Y(_2860_)
);

AOI21X1 _10126_ (
    .A(_2860_),
    .B(_2834_),
    .C(_2859_),
    .Y(_2861_)
);

INVX1 _10127_ (
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_2862_)
);

OR2X2 _10128_ (
    .A(_2837_),
    .B(_2841_),
    .Y(_2863_)
);

OAI21X1 _10129_ (
    .A(1'h0),
    .B(_2774_),
    .C(_2840_),
    .Y(_2864_)
);

NAND3X1 _10130_ (
    .A(_2686__bF$buf1),
    .B(_2864_),
    .C(_2863_),
    .Y(_2865_)
);

NOR2X1 _10131_ (
    .A(_2841_),
    .B(_2837_),
    .Y(_2866_)
);

INVX1 _10132_ (
    .A(_2864_),
    .Y(_2867_)
);

OAI21X1 _10133_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2866_),
    .C(_2867_),
    .Y(_2868_)
);

NAND3X1 _10134_ (
    .A(_2862_),
    .B(_2868_),
    .C(_2865_),
    .Y(_2869_)
);

NAND3X1 _10135_ (
    .A(_2686__bF$buf0),
    .B(_2867_),
    .C(_2863_),
    .Y(_2870_)
);

OAI21X1 _10136_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2866_),
    .C(_2864_),
    .Y(_2871_)
);

NAND3X1 _10137_ (
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .B(_2871_),
    .C(_2870_),
    .Y(_2872_)
);

AND2X2 _10138_ (
    .A(_2869_),
    .B(_2872_),
    .Y(_2873_)
);

INVX1 _10139_ (
    .A(_2873_),
    .Y(_2874_)
);

AOI21X1 _10140_ (
    .A(_2861_),
    .B(_2874_),
    .C(_2674_),
    .Y(_2875_)
);

OAI21X1 _10141_ (
    .A(_2861_),
    .B(_2874_),
    .C(_2875_),
    .Y(_2876_)
);

AOI22X1 _10142_ (
    .A(_2858_),
    .B(_2672__bF$buf1),
    .C(_2876_),
    .D(_2856_),
    .Y(_2523_)
);

NAND2X1 _10143_ (
    .A(_2830_),
    .B(_2846_),
    .Y(_2877_)
);

AND2X2 _10144_ (
    .A(_2877_),
    .B(_2849_),
    .Y(_2878_)
);

AND2X2 _10145_ (
    .A(_2818_),
    .B(_2821_),
    .Y(_2879_)
);

NAND3X1 _10146_ (
    .A(_2846_),
    .B(_2849_),
    .C(_2879_),
    .Y(_2880_)
);

OAI21X1 _10147_ (
    .A(_2826_),
    .B(_2880_),
    .C(_2878_),
    .Y(_2881_)
);

INVX1 _10148_ (
    .A(_2872_),
    .Y(_2882_)
);

AOI21X1 _10149_ (
    .A(_2881_),
    .B(_2869_),
    .C(_2882_),
    .Y(_2883_)
);

INVX1 _10150_ (
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_2884_)
);

NOR3X1 _10151_ (
    .A(_2841_),
    .B(_2864_),
    .C(_2837_),
    .Y(_2885_)
);

INVX1 _10152_ (
    .A(_2885_),
    .Y(_2886_)
);

OAI21X1 _10153_ (
    .A(1'h0),
    .B(_2794_),
    .C(_2840_),
    .Y(_2887_)
);

NAND3X1 _10154_ (
    .A(_2686__bF$buf5),
    .B(_2887_),
    .C(_2886_),
    .Y(_2888_)
);

INVX1 _10155_ (
    .A(_2887_),
    .Y(_2889_)
);

OAI21X1 _10156_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2885_),
    .C(_2889_),
    .Y(_2890_)
);

NAND3X1 _10157_ (
    .A(_2884_),
    .B(_2890_),
    .C(_2888_),
    .Y(_2891_)
);

NAND3X1 _10158_ (
    .A(_2686__bF$buf4),
    .B(_2889_),
    .C(_2886_),
    .Y(_2892_)
);

OAI21X1 _10159_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2885_),
    .C(_2887_),
    .Y(_2893_)
);

NAND3X1 _10160_ (
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .B(_2893_),
    .C(_2892_),
    .Y(_2894_)
);

AND2X2 _10161_ (
    .A(_2891_),
    .B(_2894_),
    .Y(_2895_)
);

AND2X2 _10162_ (
    .A(_2883_),
    .B(_2895_),
    .Y(_2896_)
);

OAI21X1 _10163_ (
    .A(_2895_),
    .B(_2883_),
    .C(_2741_),
    .Y(_2897_)
);

OAI21X1 _10164_ (
    .A(_2897_),
    .B(_2896_),
    .C(_2744_),
    .Y(_2898_)
);

OAI21X1 _10165_ (
    .A(_2624_),
    .B(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .C(_2898_),
    .Y(_2524_)
);

INVX1 _10166_ (
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .Y(_2899_)
);

OAI21X1 _10167_ (
    .A(1'h0),
    .B(_2811_),
    .C(_2840_),
    .Y(_2900_)
);

INVX1 _10168_ (
    .A(_2900_),
    .Y(_2901_)
);

AOI21X1 _10169_ (
    .A(_2885_),
    .B(_2889_),
    .C(_2901_),
    .Y(_2902_)
);

NAND3X1 _10170_ (
    .A(_2889_),
    .B(_2901_),
    .C(_2885_),
    .Y(_2903_)
);

NAND2X1 _10171_ (
    .A(_2686__bF$buf3),
    .B(_2903_),
    .Y(_2904_)
);

NAND2X1 _10172_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2900_),
    .Y(_2905_)
);

OAI21X1 _10173_ (
    .A(_2902_),
    .B(_2904_),
    .C(_2905_),
    .Y(_2906_)
);

NAND2X1 _10174_ (
    .A(_2899_),
    .B(_2906_),
    .Y(_2907_)
);

INVX1 _10175_ (
    .A(_2902_),
    .Y(_2908_)
);

AND2X2 _10176_ (
    .A(_2903_),
    .B(_2686__bF$buf2),
    .Y(_2909_)
);

NAND2X1 _10177_ (
    .A(_2908_),
    .B(_2909_),
    .Y(_2910_)
);

NAND3X1 _10178_ (
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .B(_2905_),
    .C(_2910_),
    .Y(_2911_)
);

NAND2X1 _10179_ (
    .A(_2907_),
    .B(_2911_),
    .Y(_2912_)
);

AOI21X1 _10180_ (
    .A(_2888_),
    .B(_2890_),
    .C(_2884_),
    .Y(_2913_)
);

AOI21X1 _10181_ (
    .A(_2882_),
    .B(_2891_),
    .C(_2913_),
    .Y(_2914_)
);

NAND3X1 _10182_ (
    .A(_2873_),
    .B(_2895_),
    .C(_2881_),
    .Y(_2915_)
);

AOI21X1 _10183_ (
    .A(_2915_),
    .B(_2914_),
    .C(_2912_),
    .Y(_2916_)
);

AND2X2 _10184_ (
    .A(_2911_),
    .B(_2907_),
    .Y(_2917_)
);

NAND3X1 _10185_ (
    .A(_2891_),
    .B(_2894_),
    .C(_2873_),
    .Y(_2918_)
);

OAI21X1 _10186_ (
    .A(_2918_),
    .B(_2861_),
    .C(_2914_),
    .Y(_2919_)
);

OAI21X1 _10187_ (
    .A(_2917_),
    .B(_2919_),
    .C(_2741_),
    .Y(_2920_)
);

OR2X2 _10188_ (
    .A(_2920_),
    .B(_2916_),
    .Y(_2921_)
);

AOI22X1 _10189_ (
    .A(_2616_),
    .B(_2672__bF$buf0),
    .C(_2921_),
    .D(_2744_),
    .Y(_2525_)
);

NAND2X1 _10190_ (
    .A(\genblk1[3].u_ce.Ycalc [11]),
    .B(_2672__bF$buf4),
    .Y(_2922_)
);

INVX1 _10191_ (
    .A(_2911_),
    .Y(_2923_)
);

NAND2X1 _10192_ (
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .B(_2838_),
    .Y(_2924_)
);

INVX1 _10193_ (
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_2925_)
);

NAND2X1 _10194_ (
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .B(_2925_),
    .Y(_2926_)
);

NAND2X1 _10195_ (
    .A(_2924_),
    .B(_2926_),
    .Y(_2927_)
);

INVX1 _10196_ (
    .A(_2927_),
    .Y(_2928_)
);

NAND2X1 _10197_ (
    .A(_2928_),
    .B(_2904_),
    .Y(_2929_)
);

NAND2X1 _10198_ (
    .A(_2927_),
    .B(_2909_),
    .Y(_2930_)
);

NAND2X1 _10199_ (
    .A(_2929_),
    .B(_2930_),
    .Y(_2931_)
);

INVX1 _10200_ (
    .A(_2931_),
    .Y(_2932_)
);

NOR3X1 _10201_ (
    .A(_2923_),
    .B(_2932_),
    .C(_2916_),
    .Y(_2933_)
);

AOI21X1 _10202_ (
    .A(_2919_),
    .B(_2917_),
    .C(_2923_),
    .Y(_2934_)
);

OAI21X1 _10203_ (
    .A(_2931_),
    .B(_2934_),
    .C(_2741_),
    .Y(_2935_)
);

OAI21X1 _10204_ (
    .A(_2933_),
    .B(_2935_),
    .C(_2744_),
    .Y(_2936_)
);

NAND2X1 _10205_ (
    .A(_2922_),
    .B(_2936_),
    .Y(_2526_)
);

NAND2X1 _10206_ (
    .A(\genblk1[3].u_ce.Xcalc [0]),
    .B(_2672__bF$buf3),
    .Y(_2937_)
);

INVX1 _10207_ (
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2938_)
);

NAND2X1 _10208_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2939_)
);

OAI21X1 _10209_ (
    .A(1'h1),
    .B(_2938_),
    .C(_2939_),
    .Y(_2940_)
);

NAND2X1 _10210_ (
    .A(1'h1),
    .B(_2940_),
    .Y(_2941_)
);

NOR2X1 _10211_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_2942_)
);

NOR2X1 _10212_ (
    .A(1'h1),
    .B(_2678_),
    .Y(_2943_)
);

AOI22X1 _10213_ (
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .B(_2942_),
    .C(_2943_),
    .D(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2944_)
);

NAND3X1 _10214_ (
    .A(_2648__bF$buf1),
    .B(_2941_),
    .C(_2944_),
    .Y(_2945_)
);

NAND2X1 _10215_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2946_)
);

OAI21X1 _10216_ (
    .A(1'h1),
    .B(_2809_),
    .C(_2946_),
    .Y(_2947_)
);

NAND2X1 _10217_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_2948_)
);

OAI21X1 _10218_ (
    .A(1'h1),
    .B(_2769_),
    .C(_2948_),
    .Y(_2949_)
);

MUX2X1 _10219_ (
    .A(_2949_),
    .B(_2947_),
    .S(_2649__bF$buf2),
    .Y(_2950_)
);

NAND2X1 _10220_ (
    .A(1'h0),
    .B(_2950_),
    .Y(_2951_)
);

AND2X2 _10221_ (
    .A(_2945_),
    .B(_2951_),
    .Y(_2952_)
);

NOR2X1 _10222_ (
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .B(_2952_),
    .Y(_2953_)
);

NAND2X1 _10223_ (
    .A(_2649__bF$buf1),
    .B(_2949_),
    .Y(_2954_)
);

NAND2X1 _10224_ (
    .A(1'h1),
    .B(_2947_),
    .Y(_2955_)
);

NAND2X1 _10225_ (
    .A(_2954_),
    .B(_2955_),
    .Y(_2956_)
);

OAI21X1 _10226_ (
    .A(_2648__bF$buf0),
    .B(_2956_),
    .C(_2945_),
    .Y(_2957_)
);

OAI21X1 _10227_ (
    .A(_2660_),
    .B(_2957_),
    .C(_2670_),
    .Y(_2958_)
);

OAI21X1 _10228_ (
    .A(_2958_),
    .B(_2953_),
    .C(_2937_),
    .Y(_2527_)
);

NAND2X1 _10229_ (
    .A(\genblk1[3].u_ce.Xcalc [1]),
    .B(_2672__bF$buf2),
    .Y(_2959_)
);

NOR2X1 _10230_ (
    .A(_2660_),
    .B(_2957_),
    .Y(_2960_)
);

NAND2X1 _10231_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2961_)
);

OAI21X1 _10232_ (
    .A(1'h1),
    .B(_2747_),
    .C(_2961_),
    .Y(_2962_)
);

NAND2X1 _10233_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2963_)
);

OAI21X1 _10234_ (
    .A(1'h1),
    .B(_2685_),
    .C(_2963_),
    .Y(_2964_)
);

MUX2X1 _10235_ (
    .A(_2964_),
    .B(_2962_),
    .S(_2649__bF$buf0),
    .Y(_2965_)
);

NAND2X1 _10236_ (
    .A(_2648__bF$buf4),
    .B(_2965_),
    .Y(_2966_)
);

NAND2X1 _10237_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_2967_)
);

OAI21X1 _10238_ (
    .A(1'h1),
    .B(_2836_),
    .C(_2967_),
    .Y(_2968_)
);

INVX1 _10239_ (
    .A(_2968_),
    .Y(_2969_)
);

NAND2X1 _10240_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2970_)
);

OAI21X1 _10241_ (
    .A(1'h1),
    .B(_2790_),
    .C(_2970_),
    .Y(_2971_)
);

NAND2X1 _10242_ (
    .A(_2649__bF$buf4),
    .B(_2971_),
    .Y(_2972_)
);

OAI21X1 _10243_ (
    .A(_2649__bF$buf3),
    .B(_2969_),
    .C(_2972_),
    .Y(_2973_)
);

OAI21X1 _10244_ (
    .A(_2648__bF$buf3),
    .B(_2973_),
    .C(_2966_),
    .Y(_2974_)
);

NAND3X1 _10245_ (
    .A(_2686__bF$buf1),
    .B(_2974_),
    .C(_2952_),
    .Y(_2975_)
);

MUX2X1 _10246_ (
    .A(_2971_),
    .B(_2968_),
    .S(_2649__bF$buf2),
    .Y(_2976_)
);

MUX2X1 _10247_ (
    .A(_2976_),
    .B(_2965_),
    .S(1'h0),
    .Y(_2977_)
);

OAI21X1 _10248_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2957_),
    .C(_2977_),
    .Y(_2978_)
);

AOI21X1 _10249_ (
    .A(_2975_),
    .B(_2978_),
    .C(_2697_),
    .Y(_2979_)
);

INVX1 _10250_ (
    .A(_2979_),
    .Y(_2980_)
);

NAND3X1 _10251_ (
    .A(_2697_),
    .B(_2978_),
    .C(_2975_),
    .Y(_2981_)
);

AND2X2 _10252_ (
    .A(_2980_),
    .B(_2981_),
    .Y(_2982_)
);

NAND2X1 _10253_ (
    .A(_2960_),
    .B(_2982_),
    .Y(_2983_)
);

OR2X2 _10254_ (
    .A(_2982_),
    .B(_2960_),
    .Y(_2984_)
);

AOI21X1 _10255_ (
    .A(_2984_),
    .B(_2983_),
    .C(_2674_),
    .Y(_2985_)
);

OAI21X1 _10256_ (
    .A(_2672__bF$buf1),
    .B(_2985_),
    .C(_2959_),
    .Y(_2528_)
);

NAND2X1 _10257_ (
    .A(\genblk1[3].u_ce.Xcalc [2]),
    .B(_2672__bF$buf0),
    .Y(_2986_)
);

AOI21X1 _10258_ (
    .A(_2960_),
    .B(_2981_),
    .C(_2979_),
    .Y(_2987_)
);

NAND2X1 _10259_ (
    .A(_2957_),
    .B(_2974_),
    .Y(_2988_)
);

NAND2X1 _10260_ (
    .A(1'h1),
    .B(_2884_),
    .Y(_2989_)
);

OAI21X1 _10261_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .C(_2989_),
    .Y(_2990_)
);

NAND2X1 _10262_ (
    .A(_2649__bF$buf1),
    .B(_2947_),
    .Y(_2991_)
);

OAI21X1 _10263_ (
    .A(_2649__bF$buf0),
    .B(_2990_),
    .C(_2991_),
    .Y(_2992_)
);

NAND2X1 _10264_ (
    .A(_2755_),
    .B(_2940_),
    .Y(_2993_)
);

NAND2X1 _10265_ (
    .A(_2949_),
    .B(_2754_),
    .Y(_2994_)
);

NAND2X1 _10266_ (
    .A(_2993_),
    .B(_2994_),
    .Y(_2995_)
);

AOI21X1 _10267_ (
    .A(_2992_),
    .B(1'h0),
    .C(_2995_),
    .Y(_2996_)
);

INVX1 _10268_ (
    .A(_2996_),
    .Y(_2997_)
);

NAND3X1 _10269_ (
    .A(_2686__bF$buf0),
    .B(_2997_),
    .C(_2988_),
    .Y(_2998_)
);

AOI21X1 _10270_ (
    .A(_2945_),
    .B(_2951_),
    .C(_2977_),
    .Y(_2999_)
);

OAI21X1 _10271_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2999_),
    .C(_2996_),
    .Y(_3000_)
);

NAND3X1 _10272_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(_3000_),
    .C(_2998_),
    .Y(_3001_)
);

INVX1 _10273_ (
    .A(_3001_),
    .Y(_3002_)
);

AOI21X1 _10274_ (
    .A(_2998_),
    .B(_3000_),
    .C(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_3003_)
);

NOR2X1 _10275_ (
    .A(_3003_),
    .B(_3002_),
    .Y(_3004_)
);

AND2X2 _10276_ (
    .A(_3004_),
    .B(_2987_),
    .Y(_3005_)
);

NOR2X1 _10277_ (
    .A(_2987_),
    .B(_3004_),
    .Y(_3006_)
);

OAI21X1 _10278_ (
    .A(_3006_),
    .B(_3005_),
    .C(_2741_),
    .Y(_3007_)
);

OAI21X1 _10279_ (
    .A(_2672__bF$buf4),
    .B(_3007_),
    .C(_2986_),
    .Y(_2529_)
);

OAI21X1 _10280_ (
    .A(_3003_),
    .B(_2987_),
    .C(_3001_),
    .Y(_3008_)
);

INVX1 _10281_ (
    .A(_3008_),
    .Y(_3009_)
);

NAND2X1 _10282_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [10]),
    .Y(_3010_)
);

OAI21X1 _10283_ (
    .A(1'h1),
    .B(_2884_),
    .C(_3010_),
    .Y(_3011_)
);

MUX2X1 _10284_ (
    .A(_3011_),
    .B(_2968_),
    .S(1'h1),
    .Y(_3012_)
);

NOR2X1 _10285_ (
    .A(_2648__bF$buf2),
    .B(_3012_),
    .Y(_3013_)
);

NAND2X1 _10286_ (
    .A(_2755_),
    .B(_2962_),
    .Y(_3014_)
);

NAND2X1 _10287_ (
    .A(_2971_),
    .B(_2754_),
    .Y(_3015_)
);

NAND2X1 _10288_ (
    .A(_3014_),
    .B(_3015_),
    .Y(_3016_)
);

OR2X2 _10289_ (
    .A(_3013_),
    .B(_3016_),
    .Y(_3017_)
);

OAI21X1 _10290_ (
    .A(_2997_),
    .B(_2988_),
    .C(_2686__bF$buf5),
    .Y(_3018_)
);

OR2X2 _10291_ (
    .A(_3018_),
    .B(_3017_),
    .Y(_3019_)
);

OAI21X1 _10292_ (
    .A(_3013_),
    .B(_3016_),
    .C(_3018_),
    .Y(_3020_)
);

AOI21X1 _10293_ (
    .A(_3019_),
    .B(_3020_),
    .C(_2694_),
    .Y(_3021_)
);

INVX1 _10294_ (
    .A(_3021_),
    .Y(_3022_)
);

NAND3X1 _10295_ (
    .A(_2694_),
    .B(_3020_),
    .C(_3019_),
    .Y(_3023_)
);

NAND2X1 _10296_ (
    .A(_3023_),
    .B(_3022_),
    .Y(_3024_)
);

OR2X2 _10297_ (
    .A(_3024_),
    .B(_3009_),
    .Y(_3025_)
);

NAND2X1 _10298_ (
    .A(_3009_),
    .B(_3024_),
    .Y(_3026_)
);

NAND2X1 _10299_ (
    .A(_3026_),
    .B(_3025_),
    .Y(_3027_)
);

AOI22X1 _10300_ (
    .A(_2640_),
    .B(_2672__bF$buf3),
    .C(_3027_),
    .D(_2670_),
    .Y(_2530_)
);

AOI21X1 _10301_ (
    .A(_3008_),
    .B(_3023_),
    .C(_3021_),
    .Y(_3028_)
);

NAND2X1 _10302_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_3029_)
);

OAI21X1 _10303_ (
    .A(1'h1),
    .B(_2899_),
    .C(_3029_),
    .Y(_3030_)
);

NAND2X1 _10304_ (
    .A(1'h1),
    .B(_3030_),
    .Y(_3031_)
);

OAI21X1 _10305_ (
    .A(1'h1),
    .B(_2990_),
    .C(_3031_),
    .Y(_3032_)
);

NAND2X1 _10306_ (
    .A(1'h0),
    .B(_3032_),
    .Y(_3033_)
);

OAI21X1 _10307_ (
    .A(1'h0),
    .B(_2950_),
    .C(_3033_),
    .Y(_3034_)
);

INVX1 _10308_ (
    .A(_3034_),
    .Y(_3035_)
);

NAND3X1 _10309_ (
    .A(_2996_),
    .B(_2957_),
    .C(_2974_),
    .Y(_3036_)
);

OAI21X1 _10310_ (
    .A(_3017_),
    .B(_3036_),
    .C(_2686__bF$buf4),
    .Y(_3037_)
);

OR2X2 _10311_ (
    .A(_3037_),
    .B(_3035_),
    .Y(_3038_)
);

NOR2X1 _10312_ (
    .A(_3017_),
    .B(_3036_),
    .Y(_3039_)
);

OAI21X1 _10313_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3039_),
    .C(_3035_),
    .Y(_3040_)
);

NAND3X1 _10314_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(_3040_),
    .C(_3038_),
    .Y(_3041_)
);

OR2X2 _10315_ (
    .A(_3037_),
    .B(_3034_),
    .Y(_3042_)
);

OAI21X1 _10316_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3039_),
    .C(_3034_),
    .Y(_3043_)
);

NAND3X1 _10317_ (
    .A(_2653_),
    .B(_3043_),
    .C(_3042_),
    .Y(_3044_)
);

NAND2X1 _10318_ (
    .A(_3041_),
    .B(_3044_),
    .Y(_3045_)
);

OR2X2 _10319_ (
    .A(_3028_),
    .B(_3045_),
    .Y(_3046_)
);

NAND2X1 _10320_ (
    .A(_3045_),
    .B(_3028_),
    .Y(_3047_)
);

NAND2X1 _10321_ (
    .A(_3047_),
    .B(_3046_),
    .Y(_3048_)
);

AOI22X1 _10322_ (
    .A(_2635_),
    .B(_2672__bF$buf2),
    .C(_3048_),
    .D(_2670_),
    .Y(_2531_)
);

INVX1 _10323_ (
    .A(\genblk1[3].u_ce.Xcalc [5]),
    .Y(_3049_)
);

OAI21X1 _10324_ (
    .A(_3045_),
    .B(_3028_),
    .C(_3041_),
    .Y(_3050_)
);

NAND2X1 _10325_ (
    .A(_3035_),
    .B(_3039_),
    .Y(_3051_)
);

NOR2X1 _10326_ (
    .A(_2649__bF$buf4),
    .B(_2925_),
    .Y(_3052_)
);

AOI21X1 _10327_ (
    .A(_2649__bF$buf3),
    .B(_3011_),
    .C(_3052_),
    .Y(_3053_)
);

NAND2X1 _10328_ (
    .A(_2648__bF$buf1),
    .B(_2973_),
    .Y(_3054_)
);

OAI21X1 _10329_ (
    .A(_2648__bF$buf0),
    .B(_3053_),
    .C(_3054_),
    .Y(_3055_)
);

INVX1 _10330_ (
    .A(_3055_),
    .Y(_3056_)
);

NAND3X1 _10331_ (
    .A(_2686__bF$buf3),
    .B(_3056_),
    .C(_3051_),
    .Y(_3057_)
);

NOR2X1 _10332_ (
    .A(_3016_),
    .B(_3013_),
    .Y(_3058_)
);

NAND3X1 _10333_ (
    .A(_2996_),
    .B(_3058_),
    .C(_2999_),
    .Y(_3059_)
);

OAI21X1 _10334_ (
    .A(_3034_),
    .B(_3059_),
    .C(_2686__bF$buf2),
    .Y(_3060_)
);

NAND2X1 _10335_ (
    .A(_3055_),
    .B(_3060_),
    .Y(_3061_)
);

AOI21X1 _10336_ (
    .A(_3057_),
    .B(_3061_),
    .C(_2690_),
    .Y(_3062_)
);

INVX1 _10337_ (
    .A(_3062_),
    .Y(_3063_)
);

NAND3X1 _10338_ (
    .A(_2690_),
    .B(_3061_),
    .C(_3057_),
    .Y(_3064_)
);

NAND2X1 _10339_ (
    .A(_3064_),
    .B(_3063_),
    .Y(_3065_)
);

NOR2X1 _10340_ (
    .A(_3065_),
    .B(_3050_),
    .Y(_3066_)
);

AND2X2 _10341_ (
    .A(_3050_),
    .B(_3065_),
    .Y(_3067_)
);

OAI21X1 _10342_ (
    .A(_3066_),
    .B(_3067_),
    .C(_2670_),
    .Y(_3068_)
);

OAI21X1 _10343_ (
    .A(_3049_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_3068_),
    .Y(_2532_)
);

INVX1 _10344_ (
    .A(\genblk1[3].u_ce.Xcalc [6]),
    .Y(_3069_)
);

NAND3X1 _10345_ (
    .A(_3035_),
    .B(_3056_),
    .C(_3039_),
    .Y(_3070_)
);

AOI21X1 _10346_ (
    .A(_2649__bF$buf2),
    .B(_3030_),
    .C(_3052_),
    .Y(_3071_)
);

NAND2X1 _10347_ (
    .A(1'h0),
    .B(_3071_),
    .Y(_3072_)
);

OAI21X1 _10348_ (
    .A(1'h0),
    .B(_2992_),
    .C(_3072_),
    .Y(_3073_)
);

NAND3X1 _10349_ (
    .A(_2686__bF$buf1),
    .B(_3073_),
    .C(_3070_),
    .Y(_3074_)
);

NOR3X1 _10350_ (
    .A(_3034_),
    .B(_3055_),
    .C(_3059_),
    .Y(_3075_)
);

INVX1 _10351_ (
    .A(_3073_),
    .Y(_3076_)
);

OAI21X1 _10352_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3075_),
    .C(_3076_),
    .Y(_3077_)
);

NAND2X1 _10353_ (
    .A(_3074_),
    .B(_3077_),
    .Y(_3078_)
);

NAND2X1 _10354_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(_3078_),
    .Y(_3079_)
);

NAND3X1 _10355_ (
    .A(_2650_),
    .B(_3074_),
    .C(_3077_),
    .Y(_3080_)
);

NAND2X1 _10356_ (
    .A(_3080_),
    .B(_3079_),
    .Y(_3081_)
);

AOI21X1 _10357_ (
    .A(_3042_),
    .B(_3043_),
    .C(_2653_),
    .Y(_3082_)
);

NOR2X1 _10358_ (
    .A(_3082_),
    .B(_3062_),
    .Y(_3083_)
);

OAI21X1 _10359_ (
    .A(_3045_),
    .B(_3028_),
    .C(_3083_),
    .Y(_3084_)
);

NAND2X1 _10360_ (
    .A(_3064_),
    .B(_3084_),
    .Y(_3085_)
);

NOR2X1 _10361_ (
    .A(_3081_),
    .B(_3085_),
    .Y(_3086_)
);

AND2X2 _10362_ (
    .A(_3079_),
    .B(_3080_),
    .Y(_3087_)
);

AND2X2 _10363_ (
    .A(_3041_),
    .B(_3044_),
    .Y(_3088_)
);

NAND3X1 _10364_ (
    .A(_3064_),
    .B(_3088_),
    .C(_3063_),
    .Y(_3089_)
);

AOI21X1 _10365_ (
    .A(_3082_),
    .B(_3064_),
    .C(_3062_),
    .Y(_3090_)
);

OAI21X1 _10366_ (
    .A(_3028_),
    .B(_3089_),
    .C(_3090_),
    .Y(_3091_)
);

NOR2X1 _10367_ (
    .A(_3087_),
    .B(_3091_),
    .Y(_3092_)
);

OAI21X1 _10368_ (
    .A(_3092_),
    .B(_3086_),
    .C(_2741_),
    .Y(_3093_)
);

NAND2X1 _10369_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .B(_3093_),
    .Y(_3094_)
);

OAI21X1 _10370_ (
    .A(_3069_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3094_),
    .Y(_2533_)
);

INVX1 _10371_ (
    .A(\genblk1[3].u_ce.Xcalc [7]),
    .Y(_3095_)
);

INVX1 _10372_ (
    .A(_3079_),
    .Y(_3096_)
);

NAND2X1 _10373_ (
    .A(_3073_),
    .B(_3075_),
    .Y(_3097_)
);

NOR2X1 _10374_ (
    .A(_2648__bF$buf4),
    .B(_2925_),
    .Y(_3098_)
);

INVX1 _10375_ (
    .A(_3098_),
    .Y(_3099_)
);

OAI21X1 _10376_ (
    .A(1'h0),
    .B(_3012_),
    .C(_3099_),
    .Y(_3100_)
);

NAND3X1 _10377_ (
    .A(_2686__bF$buf0),
    .B(_3100_),
    .C(_3097_),
    .Y(_3101_)
);

INVX1 _10378_ (
    .A(_3100_),
    .Y(_3102_)
);

OAI21X1 _10379_ (
    .A(_3076_),
    .B(_3070_),
    .C(_2686__bF$buf5),
    .Y(_3103_)
);

NAND2X1 _10380_ (
    .A(_3102_),
    .B(_3103_),
    .Y(_3104_)
);

NAND3X1 _10381_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(_3101_),
    .C(_3104_),
    .Y(_3105_)
);

NAND3X1 _10382_ (
    .A(_2686__bF$buf4),
    .B(_3102_),
    .C(_3097_),
    .Y(_3106_)
);

NAND2X1 _10383_ (
    .A(_3100_),
    .B(_3103_),
    .Y(_3107_)
);

NAND3X1 _10384_ (
    .A(_2687_),
    .B(_3106_),
    .C(_3107_),
    .Y(_3108_)
);

NAND2X1 _10385_ (
    .A(_3105_),
    .B(_3108_),
    .Y(_3109_)
);

OAI21X1 _10386_ (
    .A(_3096_),
    .B(_3086_),
    .C(_3109_),
    .Y(_3110_)
);

NOR2X1 _10387_ (
    .A(_3096_),
    .B(_3086_),
    .Y(_3111_)
);

INVX1 _10388_ (
    .A(_3109_),
    .Y(_3112_)
);

AOI21X1 _10389_ (
    .A(_3111_),
    .B(_3112_),
    .C(_2669_),
    .Y(_3113_)
);

AOI22X1 _10390_ (
    .A(_3095_),
    .B(_2672__bF$buf1),
    .C(_3113_),
    .D(_3110_),
    .Y(_2534_)
);

OAI21X1 _10391_ (
    .A(_3079_),
    .B(_3109_),
    .C(_3105_),
    .Y(_3114_)
);

NOR2X1 _10392_ (
    .A(_3081_),
    .B(_3109_),
    .Y(_3115_)
);

AOI21X1 _10393_ (
    .A(_3115_),
    .B(_3091_),
    .C(_3114_),
    .Y(_3116_)
);

INVX1 _10394_ (
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3117_)
);

NAND3X1 _10395_ (
    .A(_3073_),
    .B(_3102_),
    .C(_3075_),
    .Y(_3118_)
);

INVX1 _10396_ (
    .A(_3032_),
    .Y(_3119_)
);

OAI21X1 _10397_ (
    .A(1'h0),
    .B(_3119_),
    .C(_3099_),
    .Y(_3120_)
);

INVX1 _10398_ (
    .A(_3120_),
    .Y(_3121_)
);

NAND3X1 _10399_ (
    .A(_2686__bF$buf3),
    .B(_3121_),
    .C(_3118_),
    .Y(_3122_)
);

OAI21X1 _10400_ (
    .A(_3100_),
    .B(_3097_),
    .C(_2686__bF$buf2),
    .Y(_3123_)
);

NAND2X1 _10401_ (
    .A(_3120_),
    .B(_3123_),
    .Y(_3124_)
);

AOI21X1 _10402_ (
    .A(_3124_),
    .B(_3122_),
    .C(_3117_),
    .Y(_3125_)
);

NAND3X1 _10403_ (
    .A(_2686__bF$buf1),
    .B(_3120_),
    .C(_3118_),
    .Y(_3126_)
);

NAND2X1 _10404_ (
    .A(_3121_),
    .B(_3123_),
    .Y(_3127_)
);

AOI21X1 _10405_ (
    .A(_3127_),
    .B(_3126_),
    .C(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3128_)
);

OAI21X1 _10406_ (
    .A(_3125_),
    .B(_3128_),
    .C(_3116_),
    .Y(_3129_)
);

INVX1 _10407_ (
    .A(_3129_),
    .Y(_3130_)
);

OR2X2 _10408_ (
    .A(_3125_),
    .B(_3128_),
    .Y(_3131_)
);

OAI21X1 _10409_ (
    .A(_3131_),
    .B(_3116_),
    .C(_2670_),
    .Y(_3132_)
);

OAI22X1 _10410_ (
    .A(_2632_),
    .B(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .C(_3132_),
    .D(_3130_),
    .Y(_2535_)
);

NAND2X1 _10411_ (
    .A(\genblk1[3].u_ce.Xcalc [9]),
    .B(_2672__bF$buf0),
    .Y(_3133_)
);

NOR2X1 _10412_ (
    .A(_3131_),
    .B(_3116_),
    .Y(_3134_)
);

NOR2X1 _10413_ (
    .A(_3125_),
    .B(_3134_),
    .Y(_3135_)
);

OAI21X1 _10414_ (
    .A(1'h0),
    .B(_3053_),
    .C(_3099_),
    .Y(_3136_)
);

INVX1 _10415_ (
    .A(_3136_),
    .Y(_3137_)
);

OAI21X1 _10416_ (
    .A(_3120_),
    .B(_3118_),
    .C(_2686__bF$buf0),
    .Y(_3138_)
);

NAND2X1 _10417_ (
    .A(_3137_),
    .B(_3138_),
    .Y(_3139_)
);

OR2X2 _10418_ (
    .A(_3138_),
    .B(_3137_),
    .Y(_3140_)
);

NAND3X1 _10419_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(_3139_),
    .C(_3140_),
    .Y(_3141_)
);

NAND2X1 _10420_ (
    .A(_3139_),
    .B(_3140_),
    .Y(_3142_)
);

NAND2X1 _10421_ (
    .A(_2749_),
    .B(_3142_),
    .Y(_3143_)
);

NAND2X1 _10422_ (
    .A(_3141_),
    .B(_3143_),
    .Y(_3144_)
);

AND2X2 _10423_ (
    .A(_3135_),
    .B(_3144_),
    .Y(_3145_)
);

OAI21X1 _10424_ (
    .A(_3144_),
    .B(_3135_),
    .C(_2670_),
    .Y(_3146_)
);

OAI21X1 _10425_ (
    .A(_3146_),
    .B(_3145_),
    .C(_3133_),
    .Y(_2536_)
);

INVX1 _10426_ (
    .A(\genblk1[3].u_ce.Xcalc [10]),
    .Y(_3147_)
);

INVX1 _10427_ (
    .A(_3141_),
    .Y(_3148_)
);

AOI21X1 _10428_ (
    .A(_3125_),
    .B(_3143_),
    .C(_3148_),
    .Y(_3149_)
);

NOR2X1 _10429_ (
    .A(_3125_),
    .B(_3128_),
    .Y(_3150_)
);

NAND3X1 _10430_ (
    .A(_3141_),
    .B(_3143_),
    .C(_3150_),
    .Y(_3151_)
);

OAI21X1 _10431_ (
    .A(_3116_),
    .B(_3151_),
    .C(_3149_),
    .Y(_3152_)
);

OAI21X1 _10432_ (
    .A(1'h0),
    .B(_3071_),
    .C(_3099_),
    .Y(_3153_)
);

INVX1 _10433_ (
    .A(_3153_),
    .Y(_3154_)
);

OR2X2 _10434_ (
    .A(_3118_),
    .B(_3120_),
    .Y(_3155_)
);

OAI21X1 _10435_ (
    .A(_3136_),
    .B(_3155_),
    .C(_2686__bF$buf5),
    .Y(_3156_)
);

NAND2X1 _10436_ (
    .A(_3154_),
    .B(_3156_),
    .Y(_3157_)
);

OR2X2 _10437_ (
    .A(_3156_),
    .B(_3154_),
    .Y(_3158_)
);

NAND3X1 _10438_ (
    .A(\genblk1[3].u_ce.Xin12b [10]),
    .B(_3157_),
    .C(_3158_),
    .Y(_3159_)
);

AND2X2 _10439_ (
    .A(_3156_),
    .B(_3154_),
    .Y(_3160_)
);

NOR2X1 _10440_ (
    .A(_3154_),
    .B(_3156_),
    .Y(_3161_)
);

OAI21X1 _10441_ (
    .A(_3161_),
    .B(_3160_),
    .C(_2770_),
    .Y(_3162_)
);

NAND2X1 _10442_ (
    .A(_3162_),
    .B(_3159_),
    .Y(_3163_)
);

AND2X2 _10443_ (
    .A(_3152_),
    .B(_3163_),
    .Y(_3164_)
);

NOR2X1 _10444_ (
    .A(_3163_),
    .B(_3152_),
    .Y(_3165_)
);

NOR2X1 _10445_ (
    .A(_3164_),
    .B(_3165_),
    .Y(_3166_)
);

AOI22X1 _10446_ (
    .A(_3147_),
    .B(_2672__bF$buf4),
    .C(_3166_),
    .D(_2670_),
    .Y(_2537_)
);

NAND2X1 _10447_ (
    .A(\genblk1[3].u_ce.Xcalc [11]),
    .B(_2672__bF$buf3),
    .Y(_3167_)
);

INVX1 _10448_ (
    .A(_3159_),
    .Y(_3168_)
);

AOI21X1 _10449_ (
    .A(_3152_),
    .B(_3162_),
    .C(_3168_),
    .Y(_3169_)
);

NAND2X1 _10450_ (
    .A(_2686__bF$buf4),
    .B(_3157_),
    .Y(_3170_)
);

NOR2X1 _10451_ (
    .A(_2927_),
    .B(_3170_),
    .Y(_3171_)
);

AOI21X1 _10452_ (
    .A(_3157_),
    .B(_2686__bF$buf3),
    .C(_2928_),
    .Y(_3172_)
);

NOR2X1 _10453_ (
    .A(_3172_),
    .B(_3171_),
    .Y(_3173_)
);

AND2X2 _10454_ (
    .A(_3169_),
    .B(_3173_),
    .Y(_3174_)
);

OAI21X1 _10455_ (
    .A(_3173_),
    .B(_3169_),
    .C(_2670_),
    .Y(_3175_)
);

OAI21X1 _10456_ (
    .A(_3175_),
    .B(_3174_),
    .C(_3167_),
    .Y(_2538_)
);

OAI21X1 _10457_ (
    .A(1'h1),
    .B(_2649__bF$buf1),
    .C(_2668_),
    .Y(_3176_)
);

OAI21X1 _10458_ (
    .A(_2943_),
    .B(_3176_),
    .C(\genblk1[3].u_ce.Ain0 [0]),
    .Y(_3177_)
);

INVX1 _10459_ (
    .A(\genblk1[3].u_ce.Ain0 [0]),
    .Y(_3178_)
);

NOR2X1 _10460_ (
    .A(_2943_),
    .B(_3176_),
    .Y(_3179_)
);

NAND2X1 _10461_ (
    .A(_3178_),
    .B(_3179_),
    .Y(_3180_)
);

NAND2X1 _10462_ (
    .A(_3177_),
    .B(_3180_),
    .Y(_3181_)
);

NAND2X1 _10463_ (
    .A(\genblk1[3].u_ce.Acalc [0]),
    .B(_2672__bF$buf2),
    .Y(_3182_)
);

OAI21X1 _10464_ (
    .A(_2672__bF$buf1),
    .B(_3181_),
    .C(_3182_),
    .Y(_2539_)
);

NAND2X1 _10465_ (
    .A(\genblk1[3].u_ce.Acalc [1]),
    .B(_2672__bF$buf0),
    .Y(_3183_)
);

INVX1 _10466_ (
    .A(_3177_),
    .Y(_3184_)
);

NOR2X1 _10467_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_3185_)
);

AOI21X1 _10468_ (
    .A(_2943_),
    .B(1'h0),
    .C(_3185_),
    .Y(_3186_)
);

NOR2X1 _10469_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3186_),
    .Y(_3187_)
);

OAI21X1 _10470_ (
    .A(_2943_),
    .B(_3176_),
    .C(_2686__bF$buf2),
    .Y(_3188_)
);

AND2X2 _10471_ (
    .A(_3188_),
    .B(_3186_),
    .Y(_3189_)
);

OR2X2 _10472_ (
    .A(_3189_),
    .B(_3187_),
    .Y(_3190_)
);

OR2X2 _10473_ (
    .A(_3190_),
    .B(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3191_)
);

OAI21X1 _10474_ (
    .A(_3187_),
    .B(_3189_),
    .C(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3192_)
);

NAND2X1 _10475_ (
    .A(_3192_),
    .B(_3191_),
    .Y(_3193_)
);

NOR2X1 _10476_ (
    .A(_3184_),
    .B(_3193_),
    .Y(_3194_)
);

NAND2X1 _10477_ (
    .A(_3184_),
    .B(_3193_),
    .Y(_3195_)
);

NAND2X1 _10478_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_3195_),
    .Y(_3196_)
);

OAI21X1 _10479_ (
    .A(_3194_),
    .B(_3196_),
    .C(_3183_),
    .Y(_2540_)
);

INVX1 _10480_ (
    .A(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3197_)
);

OAI21X1 _10481_ (
    .A(_3197_),
    .B(_3190_),
    .C(_3195_),
    .Y(_3198_)
);

OAI21X1 _10482_ (
    .A(_2678_),
    .B(_2649__bF$buf0),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_3199_)
);

OAI21X1 _10483_ (
    .A(1'h1),
    .B(1'h1),
    .C(1'h0),
    .Y(_3200_)
);

MUX2X1 _10484_ (
    .A(_3200_),
    .B(1'h0),
    .S(_3199_),
    .Y(_3201_)
);

NAND2X1 _10485_ (
    .A(\genblk1[3].u_ce.Ain1 [0]),
    .B(_3201_),
    .Y(_3202_)
);

OR2X2 _10486_ (
    .A(_3201_),
    .B(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_3203_)
);

NAND2X1 _10487_ (
    .A(_3202_),
    .B(_3203_),
    .Y(_3204_)
);

INVX1 _10488_ (
    .A(_3204_),
    .Y(_3205_)
);

NOR2X1 _10489_ (
    .A(_3205_),
    .B(_3198_),
    .Y(_3206_)
);

NAND2X1 _10490_ (
    .A(_3205_),
    .B(_3198_),
    .Y(_3207_)
);

NAND2X1 _10491_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .B(_3207_),
    .Y(_3208_)
);

OAI22X1 _10492_ (
    .A(_2594_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3206_),
    .D(_3208_),
    .Y(_2541_)
);

NOR2X1 _10493_ (
    .A(\genblk1[3].u_ce.Acalc [3]),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .Y(_3209_)
);

NAND2X1 _10494_ (
    .A(_3202_),
    .B(_3207_),
    .Y(_3210_)
);

INVX1 _10495_ (
    .A(_3210_),
    .Y(_3211_)
);

INVX1 _10496_ (
    .A(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_3212_)
);

NOR2X1 _10497_ (
    .A(1'h1),
    .B(_2649__bF$buf4),
    .Y(_3213_)
);

OAI21X1 _10498_ (
    .A(_2648__bF$buf3),
    .B(_3213_),
    .C(_2686__bF$buf1),
    .Y(_3214_)
);

OAI21X1 _10499_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_3215_)
);

OAI21X1 _10500_ (
    .A(_2678_),
    .B(_3215_),
    .C(_3214_),
    .Y(_3216_)
);

NOR2X1 _10501_ (
    .A(_3212_),
    .B(_3216_),
    .Y(_3217_)
);

NAND2X1 _10502_ (
    .A(_3212_),
    .B(_3216_),
    .Y(_3218_)
);

INVX1 _10503_ (
    .A(_3218_),
    .Y(_3219_)
);

NOR2X1 _10504_ (
    .A(_3217_),
    .B(_3219_),
    .Y(_3220_)
);

OAI21X1 _10505_ (
    .A(_3220_),
    .B(_3211_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_3221_)
);

AOI21X1 _10506_ (
    .A(_3211_),
    .B(_3220_),
    .C(_3221_),
    .Y(_3222_)
);

NOR2X1 _10507_ (
    .A(_3209_),
    .B(_3222_),
    .Y(_2542_)
);

NAND2X1 _10508_ (
    .A(\genblk1[3].u_ce.Acalc [4]),
    .B(_2672__bF$buf4),
    .Y(_3223_)
);

INVX1 _10509_ (
    .A(\genblk1[3].u_ce.Ain12b [4]),
    .Y(_3224_)
);

AOI21X1 _10510_ (
    .A(_2943_),
    .B(1'h0),
    .C(_2686__bF$buf0),
    .Y(_3225_)
);

OAI21X1 _10511_ (
    .A(1'h0),
    .B(_2943_),
    .C(_3225_),
    .Y(_3226_)
);

OAI21X1 _10512_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3186_),
    .C(_3226_),
    .Y(_3227_)
);

OR2X2 _10513_ (
    .A(_3227_),
    .B(_3224_),
    .Y(_3228_)
);

NAND2X1 _10514_ (
    .A(_3224_),
    .B(_3227_),
    .Y(_3229_)
);

NAND2X1 _10515_ (
    .A(_3229_),
    .B(_3228_),
    .Y(_3230_)
);

AOI21X1 _10516_ (
    .A(_3210_),
    .B(_3218_),
    .C(_3217_),
    .Y(_3231_)
);

AND2X2 _10517_ (
    .A(_3231_),
    .B(_3230_),
    .Y(_3232_)
);

OAI21X1 _10518_ (
    .A(_3230_),
    .B(_3231_),
    .C(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .Y(_3233_)
);

OAI21X1 _10519_ (
    .A(_3233_),
    .B(_3232_),
    .C(_3223_),
    .Y(_2543_)
);

OAI21X1 _10520_ (
    .A(_3230_),
    .B(_3231_),
    .C(_3228_),
    .Y(_3234_)
);

INVX1 _10521_ (
    .A(\genblk1[3].u_ce.Ain12b [5]),
    .Y(_3235_)
);

OAI21X1 _10522_ (
    .A(_2942_),
    .B(_2755_),
    .C(_2686__bF$buf5),
    .Y(_3236_)
);

OAI21X1 _10523_ (
    .A(1'h1),
    .B(1'h1),
    .C(_2668_),
    .Y(_3237_)
);

OR2X2 _10524_ (
    .A(_3237_),
    .B(_2686__bF$buf4),
    .Y(_3238_)
);

NAND2X1 _10525_ (
    .A(_3236_),
    .B(_3238_),
    .Y(_3239_)
);

OR2X2 _10526_ (
    .A(_3239_),
    .B(_3235_),
    .Y(_3240_)
);

NAND2X1 _10527_ (
    .A(_3235_),
    .B(_3239_),
    .Y(_3241_)
);

NAND2X1 _10528_ (
    .A(_3241_),
    .B(_3240_),
    .Y(_3242_)
);

INVX1 _10529_ (
    .A(_3242_),
    .Y(_3243_)
);

NOR2X1 _10530_ (
    .A(_3243_),
    .B(_3234_),
    .Y(_3244_)
);

NAND2X1 _10531_ (
    .A(_3243_),
    .B(_3234_),
    .Y(_3245_)
);

NAND2X1 _10532_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .B(_3245_),
    .Y(_3246_)
);

OAI22X1 _10533_ (
    .A(_2611_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3244_),
    .D(_3246_),
    .Y(_2544_)
);

NAND2X1 _10534_ (
    .A(\genblk1[3].u_ce.Acalc [6]),
    .B(_2672__bF$buf3),
    .Y(_3247_)
);

INVX1 _10535_ (
    .A(_3230_),
    .Y(_3248_)
);

NAND2X1 _10536_ (
    .A(_3243_),
    .B(_3248_),
    .Y(_3249_)
);

OAI21X1 _10537_ (
    .A(_3228_),
    .B(_3242_),
    .C(_3240_),
    .Y(_3250_)
);

INVX1 _10538_ (
    .A(_3250_),
    .Y(_3251_)
);

OAI21X1 _10539_ (
    .A(_3249_),
    .B(_3231_),
    .C(_3251_),
    .Y(_3252_)
);

OAI21X1 _10540_ (
    .A(1'h1),
    .B(_2678_),
    .C(_2648__bF$buf2),
    .Y(_3253_)
);

NOR2X1 _10541_ (
    .A(_3253_),
    .B(_3213_),
    .Y(_3254_)
);

NAND2X1 _10542_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3254_),
    .Y(_3255_)
);

OAI21X1 _10543_ (
    .A(_3253_),
    .B(_3213_),
    .C(_2686__bF$buf3),
    .Y(_3256_)
);

NAND2X1 _10544_ (
    .A(_3256_),
    .B(_3255_),
    .Y(_3257_)
);

NAND2X1 _10545_ (
    .A(\genblk1[3].u_ce.Ain12b [6]),
    .B(_3257_),
    .Y(_3258_)
);

OR2X2 _10546_ (
    .A(_3257_),
    .B(\genblk1[3].u_ce.Ain12b [6]),
    .Y(_3259_)
);

NAND2X1 _10547_ (
    .A(_3258_),
    .B(_3259_),
    .Y(_3260_)
);

INVX1 _10548_ (
    .A(_3260_),
    .Y(_3261_)
);

NOR2X1 _10549_ (
    .A(_3261_),
    .B(_3252_),
    .Y(_3262_)
);

NAND2X1 _10550_ (
    .A(_3261_),
    .B(_3252_),
    .Y(_3263_)
);

NAND2X1 _10551_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .B(_3263_),
    .Y(_3264_)
);

OAI21X1 _10552_ (
    .A(_3262_),
    .B(_3264_),
    .C(_3247_),
    .Y(_2545_)
);

INVX1 _10553_ (
    .A(\genblk1[3].u_ce.Acalc [7]),
    .Y(_3265_)
);

NAND2X1 _10554_ (
    .A(_3258_),
    .B(_3263_),
    .Y(_3266_)
);

INVX1 _10555_ (
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .Y(_3267_)
);

NAND2X1 _10556_ (
    .A(_2686__bF$buf2),
    .B(_3185_),
    .Y(_3268_)
);

OR2X2 _10557_ (
    .A(_3185_),
    .B(_2686__bF$buf1),
    .Y(_3269_)
);

NAND2X1 _10558_ (
    .A(_3268_),
    .B(_3269_),
    .Y(_3270_)
);

NOR2X1 _10559_ (
    .A(_3267_),
    .B(_3270_),
    .Y(_3271_)
);

INVX1 _10560_ (
    .A(_3271_),
    .Y(_3272_)
);

NAND2X1 _10561_ (
    .A(_3267_),
    .B(_3270_),
    .Y(_3273_)
);

NAND2X1 _10562_ (
    .A(_3273_),
    .B(_3272_),
    .Y(_3274_)
);

OR2X2 _10563_ (
    .A(_3266_),
    .B(_3274_),
    .Y(_3275_)
);

AOI21X1 _10564_ (
    .A(_3266_),
    .B(_3274_),
    .C(_2672__bF$buf2),
    .Y(_3276_)
);

AOI22X1 _10565_ (
    .A(_3265_),
    .B(_2672__bF$buf1),
    .C(_3275_),
    .D(_3276_),
    .Y(_2546_)
);

NAND2X1 _10566_ (
    .A(\genblk1[3].u_ce.Acalc [8]),
    .B(_2672__bF$buf0),
    .Y(_3277_)
);

NOR2X1 _10567_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2668_),
    .Y(_3278_)
);

INVX1 _10568_ (
    .A(_3278_),
    .Y(_3279_)
);

NAND3X1 _10569_ (
    .A(\genblk1[3].u_ce.Ain12b [8]),
    .B(_3215_),
    .C(_3279_),
    .Y(_3280_)
);

INVX1 _10570_ (
    .A(_3280_),
    .Y(_3281_)
);

AOI21X1 _10571_ (
    .A(_3279_),
    .B(_3215_),
    .C(\genblk1[3].u_ce.Ain12b [8]),
    .Y(_3282_)
);

NOR2X1 _10572_ (
    .A(_3282_),
    .B(_3281_),
    .Y(_3283_)
);

OAI21X1 _10573_ (
    .A(_3258_),
    .B(_3274_),
    .C(_3272_),
    .Y(_3284_)
);

NOR2X1 _10574_ (
    .A(_3274_),
    .B(_3260_),
    .Y(_3285_)
);

AOI21X1 _10575_ (
    .A(_3285_),
    .B(_3250_),
    .C(_3284_),
    .Y(_3286_)
);

NAND3X1 _10576_ (
    .A(_3248_),
    .B(_3243_),
    .C(_3285_),
    .Y(_3287_)
);

OAI21X1 _10577_ (
    .A(_3287_),
    .B(_3231_),
    .C(_3286_),
    .Y(_3288_)
);

NOR2X1 _10578_ (
    .A(_3283_),
    .B(_3288_),
    .Y(_3289_)
);

NAND2X1 _10579_ (
    .A(_3283_),
    .B(_3288_),
    .Y(_3290_)
);

NAND2X1 _10580_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .B(_3290_),
    .Y(_3291_)
);

OAI21X1 _10581_ (
    .A(_3289_),
    .B(_3291_),
    .C(_3277_),
    .Y(_2547_)
);

AOI21X1 _10582_ (
    .A(_3288_),
    .B(_3283_),
    .C(_3281_),
    .Y(_3292_)
);

OR2X2 _10583_ (
    .A(_2686__bF$buf0),
    .B(\genblk1[3].u_ce.Ain12b [9]),
    .Y(_3293_)
);

NAND2X1 _10584_ (
    .A(\genblk1[3].u_ce.Ain12b [9]),
    .B(_2686__bF$buf5),
    .Y(_3294_)
);

NAND2X1 _10585_ (
    .A(_3294_),
    .B(_3293_),
    .Y(_3295_)
);

AND2X2 _10586_ (
    .A(_3292_),
    .B(_3295_),
    .Y(_3296_)
);

OAI21X1 _10587_ (
    .A(_3295_),
    .B(_3292_),
    .C(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .Y(_3297_)
);

OAI22X1 _10588_ (
    .A(_2608_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_3297_),
    .D(_3296_),
    .Y(_2548_)
);

NAND2X1 _10589_ (
    .A(\genblk1[3].u_ce.Acalc [10]),
    .B(_2672__bF$buf4),
    .Y(_3298_)
);

OAI21X1 _10590_ (
    .A(_3295_),
    .B(_3280_),
    .C(_3294_),
    .Y(_3299_)
);

NAND3X1 _10591_ (
    .A(_3293_),
    .B(_3294_),
    .C(_3283_),
    .Y(_3300_)
);

INVX1 _10592_ (
    .A(_3300_),
    .Y(_3301_)
);

AOI21X1 _10593_ (
    .A(_3288_),
    .B(_3301_),
    .C(_3299_),
    .Y(_3302_)
);

INVX1 _10594_ (
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .Y(_3303_)
);

NAND2X1 _10595_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3303_),
    .Y(_3304_)
);

NAND2X1 _10596_ (
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .B(_2686__bF$buf4),
    .Y(_3305_)
);

NAND2X1 _10597_ (
    .A(_3304_),
    .B(_3305_),
    .Y(_3306_)
);

AND2X2 _10598_ (
    .A(_3302_),
    .B(_3306_),
    .Y(_3307_)
);

OAI21X1 _10599_ (
    .A(_3306_),
    .B(_3302_),
    .C(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .Y(_3308_)
);

OAI21X1 _10600_ (
    .A(_3308_),
    .B(_3307_),
    .C(_3298_),
    .Y(_2549_)
);

NAND2X1 _10601_ (
    .A(\genblk1[3].u_ce.Acalc [11]),
    .B(_2672__bF$buf3),
    .Y(_3309_)
);

OAI21X1 _10602_ (
    .A(_3306_),
    .B(_3302_),
    .C(_3305_),
    .Y(_3310_)
);

OAI21X1 _10603_ (
    .A(_2672__bF$buf2),
    .B(_3310_),
    .C(_3309_),
    .Y(_2550_)
);

NAND2X1 _10604_ (
    .A(\genblk1[3].u_ce.LoadCtl [5]),
    .B(_2599_),
    .Y(_3311_)
);

NAND2X1 _10605_ (
    .A(_2600_),
    .B(_2606_),
    .Y(_3312_)
);

NOR2X1 _10606_ (
    .A(_3311_),
    .B(_3312_),
    .Y(_3313_)
);

NAND2X1 _10607_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3313_),
    .Y(_3314_)
);

OAI21X1 _10608_ (
    .A(_2770_),
    .B(_3313_),
    .C(_3314_),
    .Y(_2551_)
);

NAND2X1 _10609_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3313_),
    .Y(_3315_)
);

OAI21X1 _10610_ (
    .A(_2838_),
    .B(_3313_),
    .C(_3315_),
    .Y(_2552_)
);

INVX1 _10611_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .Y(_3316_)
);

OR2X2 _10612_ (
    .A(_3312_),
    .B(_2599_),
    .Y(_3317_)
);

OAI21X1 _10613_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3318_)
);

OAI21X1 _10614_ (
    .A(_3316_),
    .B(_3317_),
    .C(_3318_),
    .Y(_2553_)
);

INVX1 _10615_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .Y(_3319_)
);

OAI21X1 _10616_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Xin12b [9]),
    .Y(_3320_)
);

OAI21X1 _10617_ (
    .A(_3319_),
    .B(_3317_),
    .C(_3320_),
    .Y(_2554_)
);

NAND2X1 _10618_ (
    .A(_2606_),
    .B(_2603_),
    .Y(_3321_)
);

NAND2X1 _10619_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(_3321_),
    .Y(_3322_)
);

OAI21X1 _10620_ (
    .A(_3316_),
    .B(_3321_),
    .C(_3322_),
    .Y(_2555_)
);

NAND2X1 _10621_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(_3321_),
    .Y(_3323_)
);

OAI21X1 _10622_ (
    .A(_3319_),
    .B(_3321_),
    .C(_3323_),
    .Y(_2556_)
);

AND2X2 _10623_ (
    .A(_2606_),
    .B(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_3324_)
);

NAND2X1 _10624_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3324_),
    .Y(_3325_)
);

OAI21X1 _10625_ (
    .A(_2653_),
    .B(_3324_),
    .C(_3325_),
    .Y(_2557_)
);

NAND2X1 _10626_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3324_),
    .Y(_3326_)
);

OAI21X1 _10627_ (
    .A(_2690_),
    .B(_3324_),
    .C(_3326_),
    .Y(_2558_)
);

OAI21X1 _10628_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_3327_)
);

OAI21X1 _10629_ (
    .A(_3316_),
    .B(_2597_),
    .C(_3327_),
    .Y(_2559_)
);

OAI21X1 _10630_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_3328_)
);

OAI21X1 _10631_ (
    .A(_3319_),
    .B(_2597_),
    .C(_3328_),
    .Y(_2560_)
);

NAND2X1 _10632_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.X_ [0]),
    .Y(_3329_)
);

OAI21X1 _10633_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2660_),
    .C(_3329_),
    .Y(_2561_)
);

NAND2X1 _10634_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.X_ [1]),
    .Y(_3330_)
);

OAI21X1 _10635_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2697_),
    .C(_3330_),
    .Y(_2562_)
);

NAND2X1 _10636_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3313_),
    .Y(_3331_)
);

OAI21X1 _10637_ (
    .A(_2899_),
    .B(_3313_),
    .C(_3331_),
    .Y(_2563_)
);

NAND2X1 _10638_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3313_),
    .Y(_3332_)
);

OAI21X1 _10639_ (
    .A(_2925_),
    .B(_3313_),
    .C(_3332_),
    .Y(_2564_)
);

INVX1 _10640_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .Y(_3333_)
);

OAI21X1 _10641_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_3334_)
);

OAI21X1 _10642_ (
    .A(_3333_),
    .B(_3317_),
    .C(_3334_),
    .Y(_2565_)
);

INVX1 _10643_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .Y(_3335_)
);

OAI21X1 _10644_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_3336_)
);

OAI21X1 _10645_ (
    .A(_3335_),
    .B(_3317_),
    .C(_3336_),
    .Y(_2566_)
);

NAND2X1 _10646_ (
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .B(_3321_),
    .Y(_3337_)
);

OAI21X1 _10647_ (
    .A(_3333_),
    .B(_3321_),
    .C(_3337_),
    .Y(_2567_)
);

NAND2X1 _10648_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(_3321_),
    .Y(_3338_)
);

OAI21X1 _10649_ (
    .A(_3335_),
    .B(_3321_),
    .C(_3338_),
    .Y(_2568_)
);

NAND2X1 _10650_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3324_),
    .Y(_3339_)
);

OAI21X1 _10651_ (
    .A(_2769_),
    .B(_3324_),
    .C(_3339_),
    .Y(_2569_)
);

NAND2X1 _10652_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3324_),
    .Y(_3340_)
);

OAI21X1 _10653_ (
    .A(_2790_),
    .B(_3324_),
    .C(_3340_),
    .Y(_2570_)
);

OAI21X1 _10654_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_3341_)
);

OAI21X1 _10655_ (
    .A(_3333_),
    .B(_2597_),
    .C(_3341_),
    .Y(_2571_)
);

OAI21X1 _10656_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_3342_)
);

OAI21X1 _10657_ (
    .A(_3335_),
    .B(_2597_),
    .C(_3342_),
    .Y(_2572_)
);

NAND2X1 _10658_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[2].u_ce.Y_ [0]),
    .Y(_3343_)
);

OAI21X1 _10659_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_2647_),
    .C(_3343_),
    .Y(_2573_)
);

NAND2X1 _10660_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[2].u_ce.Y_ [1]),
    .Y(_3344_)
);

OAI21X1 _10661_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2685_),
    .C(_3344_),
    .Y(_2574_)
);

NAND2X1 _10662_ (
    .A(\a[3] [0]),
    .B(_3313_),
    .Y(_3345_)
);

OAI21X1 _10663_ (
    .A(_3303_),
    .B(_3313_),
    .C(_3345_),
    .Y(_2575_)
);

NAND2X1 _10664_ (
    .A(\a[3] [1]),
    .B(_3313_),
    .Y(_3346_)
);

OAI21X1 _10665_ (
    .A(_2686__bF$buf3),
    .B(_3313_),
    .C(_3346_),
    .Y(_2576_)
);

INVX1 _10666_ (
    .A(\a[3] [0]),
    .Y(_3347_)
);

OAI21X1 _10667_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Ain12b [8]),
    .Y(_3348_)
);

OAI21X1 _10668_ (
    .A(_3347_),
    .B(_3317_),
    .C(_3348_),
    .Y(_2577_)
);

INVX1 _10669_ (
    .A(\a[3] [1]),
    .Y(_3349_)
);

OAI21X1 _10670_ (
    .A(_2599_),
    .B(_3312_),
    .C(\genblk1[3].u_ce.Ain12b [9]),
    .Y(_3350_)
);

OAI21X1 _10671_ (
    .A(_3349_),
    .B(_3317_),
    .C(_3350_),
    .Y(_2578_)
);

NAND2X1 _10672_ (
    .A(\genblk1[3].u_ce.Ain12b [6]),
    .B(_3321_),
    .Y(_3351_)
);

OAI21X1 _10673_ (
    .A(_3347_),
    .B(_3321_),
    .C(_3351_),
    .Y(_2579_)
);

NAND2X1 _10674_ (
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .B(_3321_),
    .Y(_2587_)
);

OAI21X1 _10675_ (
    .A(_3349_),
    .B(_3321_),
    .C(_2587_),
    .Y(_2580_)
);

NAND2X1 _10676_ (
    .A(\a[3] [0]),
    .B(_3324_),
    .Y(_2588_)
);

OAI21X1 _10677_ (
    .A(_3224_),
    .B(_3324_),
    .C(_2588_),
    .Y(_2581_)
);

NAND2X1 _10678_ (
    .A(\a[3] [1]),
    .B(_3324_),
    .Y(_2589_)
);

OAI21X1 _10679_ (
    .A(_3235_),
    .B(_3324_),
    .C(_2589_),
    .Y(_2582_)
);

OAI21X1 _10680_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_2590_)
);

OAI21X1 _10681_ (
    .A(_3347_),
    .B(_2597_),
    .C(_2590_),
    .Y(_2583_)
);

OAI21X1 _10682_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2595_),
    .C(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_2591_)
);

OAI21X1 _10683_ (
    .A(_3349_),
    .B(_2597_),
    .C(_2591_),
    .Y(_2584_)
);

NAND2X1 _10684_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[3] [0]),
    .Y(_2592_)
);

OAI21X1 _10685_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3178_),
    .C(_2592_),
    .Y(_2585_)
);

NAND2X1 _10686_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\a[3] [1]),
    .Y(_2593_)
);

OAI21X1 _10687_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3197_),
    .C(_2593_),
    .Y(_2586_)
);

DFFPOSX1 _10688_ (
    .CLK(clk_bF$buf78),
    .D(_2514_),
    .Q(\genblk1[3].u_ce.Ycalc [0])
);

DFFPOSX1 _10689_ (
    .CLK(clk_bF$buf77),
    .D(_2515_),
    .Q(\genblk1[3].u_ce.Ycalc [1])
);

DFFPOSX1 _10690_ (
    .CLK(clk_bF$buf76),
    .D(_2516_),
    .Q(\genblk1[3].u_ce.ISout )
);

DFFPOSX1 _10691_ (
    .CLK(clk_bF$buf75),
    .D(_2517_),
    .Q(\genblk1[3].u_ce.Ycalc [2])
);

DFFPOSX1 _10692_ (
    .CLK(clk_bF$buf74),
    .D(_2518_),
    .Q(\genblk1[3].u_ce.Ycalc [3])
);

DFFPOSX1 _10693_ (
    .CLK(clk_bF$buf73),
    .D(_2519_),
    .Q(\genblk1[3].u_ce.Ycalc [4])
);

DFFPOSX1 _10694_ (
    .CLK(clk_bF$buf72),
    .D(_2520_),
    .Q(\genblk1[3].u_ce.Ycalc [5])
);

DFFPOSX1 _10695_ (
    .CLK(clk_bF$buf71),
    .D(_2521_),
    .Q(\genblk1[3].u_ce.Ycalc [6])
);

DFFPOSX1 _10696_ (
    .CLK(clk_bF$buf70),
    .D(_2522_),
    .Q(\genblk1[3].u_ce.Ycalc [7])
);

DFFPOSX1 _10697_ (
    .CLK(clk_bF$buf69),
    .D(_2523_),
    .Q(\genblk1[3].u_ce.Ycalc [8])
);

DFFPOSX1 _10698_ (
    .CLK(clk_bF$buf68),
    .D(_2524_),
    .Q(\genblk1[3].u_ce.Ycalc [9])
);

DFFPOSX1 _10699_ (
    .CLK(clk_bF$buf67),
    .D(_2525_),
    .Q(\genblk1[3].u_ce.Ycalc [10])
);

DFFPOSX1 _10700_ (
    .CLK(clk_bF$buf66),
    .D(_2526_),
    .Q(\genblk1[3].u_ce.Ycalc [11])
);

DFFPOSX1 _10701_ (
    .CLK(clk_bF$buf65),
    .D(_2527_),
    .Q(\genblk1[3].u_ce.Xcalc [0])
);

DFFPOSX1 _10702_ (
    .CLK(clk_bF$buf64),
    .D(_2528_),
    .Q(\genblk1[3].u_ce.Xcalc [1])
);

DFFPOSX1 _10703_ (
    .CLK(clk_bF$buf63),
    .D(_2529_),
    .Q(\genblk1[3].u_ce.Xcalc [2])
);

DFFPOSX1 _10704_ (
    .CLK(clk_bF$buf62),
    .D(_2530_),
    .Q(\genblk1[3].u_ce.Xcalc [3])
);

DFFPOSX1 _10705_ (
    .CLK(clk_bF$buf61),
    .D(_2531_),
    .Q(\genblk1[3].u_ce.Xcalc [4])
);

DFFPOSX1 _10706_ (
    .CLK(clk_bF$buf60),
    .D(_2532_),
    .Q(\genblk1[3].u_ce.Xcalc [5])
);

DFFPOSX1 _10707_ (
    .CLK(clk_bF$buf59),
    .D(_2533_),
    .Q(\genblk1[3].u_ce.Xcalc [6])
);

DFFPOSX1 _10708_ (
    .CLK(clk_bF$buf58),
    .D(_2534_),
    .Q(\genblk1[3].u_ce.Xcalc [7])
);

DFFPOSX1 _10709_ (
    .CLK(clk_bF$buf57),
    .D(_2535_),
    .Q(\genblk1[3].u_ce.Xcalc [8])
);

DFFPOSX1 _10710_ (
    .CLK(clk_bF$buf56),
    .D(_2536_),
    .Q(\genblk1[3].u_ce.Xcalc [9])
);

DFFPOSX1 _10711_ (
    .CLK(clk_bF$buf55),
    .D(_2537_),
    .Q(\genblk1[3].u_ce.Xcalc [10])
);

DFFPOSX1 _10712_ (
    .CLK(clk_bF$buf54),
    .D(_2538_),
    .Q(\genblk1[3].u_ce.Xcalc [11])
);

DFFPOSX1 _10713_ (
    .CLK(clk_bF$buf53),
    .D(_2539_),
    .Q(\genblk1[3].u_ce.Acalc [0])
);

DFFPOSX1 _10714_ (
    .CLK(clk_bF$buf52),
    .D(_2540_),
    .Q(\genblk1[3].u_ce.Acalc [1])
);

DFFPOSX1 _10715_ (
    .CLK(clk_bF$buf51),
    .D(_2541_),
    .Q(\genblk1[3].u_ce.Acalc [2])
);

DFFPOSX1 _10716_ (
    .CLK(clk_bF$buf50),
    .D(_2542_),
    .Q(\genblk1[3].u_ce.Acalc [3])
);

DFFPOSX1 _10717_ (
    .CLK(clk_bF$buf49),
    .D(_2543_),
    .Q(\genblk1[3].u_ce.Acalc [4])
);

DFFPOSX1 _10718_ (
    .CLK(clk_bF$buf48),
    .D(_2544_),
    .Q(\genblk1[3].u_ce.Acalc [5])
);

DFFPOSX1 _10719_ (
    .CLK(clk_bF$buf47),
    .D(_2545_),
    .Q(\genblk1[3].u_ce.Acalc [6])
);

DFFPOSX1 _10720_ (
    .CLK(clk_bF$buf46),
    .D(_2546_),
    .Q(\genblk1[3].u_ce.Acalc [7])
);

DFFPOSX1 _10721_ (
    .CLK(clk_bF$buf45),
    .D(_2547_),
    .Q(\genblk1[3].u_ce.Acalc [8])
);

DFFPOSX1 _10722_ (
    .CLK(clk_bF$buf44),
    .D(_2548_),
    .Q(\genblk1[3].u_ce.Acalc [9])
);

DFFPOSX1 _10723_ (
    .CLK(clk_bF$buf43),
    .D(_2549_),
    .Q(\genblk1[3].u_ce.Acalc [10])
);

DFFPOSX1 _10724_ (
    .CLK(clk_bF$buf42),
    .D(_2550_),
    .Q(\genblk1[3].u_ce.Acalc [11])
);

DFFPOSX1 _10725_ (
    .CLK(clk_bF$buf41),
    .D(_2551_),
    .Q(\genblk1[3].u_ce.Xin12b [10])
);

DFFPOSX1 _10726_ (
    .CLK(clk_bF$buf40),
    .D(_2552_),
    .Q(\genblk1[3].u_ce.Xin12b [11])
);

DFFPOSX1 _10727_ (
    .CLK(clk_bF$buf39),
    .D(_2553_),
    .Q(\genblk1[3].u_ce.Xin12b [8])
);

DFFPOSX1 _10728_ (
    .CLK(clk_bF$buf38),
    .D(_2554_),
    .Q(\genblk1[3].u_ce.Xin12b [9])
);

DFFPOSX1 _10729_ (
    .CLK(clk_bF$buf37),
    .D(_2555_),
    .Q(\genblk1[3].u_ce.Xin12b [6])
);

DFFPOSX1 _10730_ (
    .CLK(clk_bF$buf36),
    .D(_2556_),
    .Q(\genblk1[3].u_ce.Xin12b [7])
);

DFFPOSX1 _10731_ (
    .CLK(clk_bF$buf35),
    .D(_2557_),
    .Q(\genblk1[3].u_ce.Xin12b [4])
);

DFFPOSX1 _10732_ (
    .CLK(clk_bF$buf34),
    .D(_2558_),
    .Q(\genblk1[3].u_ce.Xin12b [5])
);

DFFPOSX1 _10733_ (
    .CLK(clk_bF$buf33),
    .D(_2559_),
    .Q(\genblk1[3].u_ce.Xin1 [0])
);

DFFPOSX1 _10734_ (
    .CLK(clk_bF$buf32),
    .D(_2560_),
    .Q(\genblk1[3].u_ce.Xin1 [1])
);

DFFPOSX1 _10735_ (
    .CLK(clk_bF$buf31),
    .D(_2561_),
    .Q(\genblk1[3].u_ce.Xin0 [0])
);

DFFPOSX1 _10736_ (
    .CLK(clk_bF$buf30),
    .D(_2562_),
    .Q(\genblk1[3].u_ce.Xin0 [1])
);

DFFPOSX1 _10737_ (
    .CLK(clk_bF$buf29),
    .D(_2563_),
    .Q(\genblk1[3].u_ce.Yin12b [10])
);

DFFPOSX1 _10738_ (
    .CLK(clk_bF$buf28),
    .D(_2564_),
    .Q(\genblk1[3].u_ce.Yin12b [11])
);

DFFPOSX1 _10739_ (
    .CLK(clk_bF$buf27),
    .D(_2565_),
    .Q(\genblk1[3].u_ce.Yin12b [8])
);

DFFPOSX1 _10740_ (
    .CLK(clk_bF$buf26),
    .D(_2566_),
    .Q(\genblk1[3].u_ce.Yin12b [9])
);

DFFPOSX1 _10741_ (
    .CLK(clk_bF$buf25),
    .D(_2567_),
    .Q(\genblk1[3].u_ce.Yin12b [6])
);

DFFPOSX1 _10742_ (
    .CLK(clk_bF$buf24),
    .D(_2568_),
    .Q(\genblk1[3].u_ce.Yin12b [7])
);

DFFPOSX1 _10743_ (
    .CLK(clk_bF$buf23),
    .D(_2569_),
    .Q(\genblk1[3].u_ce.Yin12b [4])
);

DFFPOSX1 _10744_ (
    .CLK(clk_bF$buf22),
    .D(_2570_),
    .Q(\genblk1[3].u_ce.Yin12b [5])
);

DFFPOSX1 _10745_ (
    .CLK(clk_bF$buf21),
    .D(_2571_),
    .Q(\genblk1[3].u_ce.Yin1 [0])
);

DFFPOSX1 _10746_ (
    .CLK(clk_bF$buf20),
    .D(_2572_),
    .Q(\genblk1[3].u_ce.Yin1 [1])
);

DFFPOSX1 _10747_ (
    .CLK(clk_bF$buf19),
    .D(_2573_),
    .Q(\genblk1[3].u_ce.Yin0 [0])
);

DFFPOSX1 _10748_ (
    .CLK(clk_bF$buf18),
    .D(_2574_),
    .Q(\genblk1[3].u_ce.Yin0 [1])
);

DFFPOSX1 _10749_ (
    .CLK(clk_bF$buf17),
    .D(_2575_),
    .Q(\genblk1[3].u_ce.Ain12b [10])
);

DFFPOSX1 _10750_ (
    .CLK(clk_bF$buf16),
    .D(_2576_),
    .Q(\genblk1[3].u_ce.Ain12b [11])
);

DFFPOSX1 _10751_ (
    .CLK(clk_bF$buf15),
    .D(_2577_),
    .Q(\genblk1[3].u_ce.Ain12b [8])
);

DFFPOSX1 _10752_ (
    .CLK(clk_bF$buf14),
    .D(_2578_),
    .Q(\genblk1[3].u_ce.Ain12b [9])
);

DFFPOSX1 _10753_ (
    .CLK(clk_bF$buf13),
    .D(_2579_),
    .Q(\genblk1[3].u_ce.Ain12b [6])
);

DFFPOSX1 _10754_ (
    .CLK(clk_bF$buf12),
    .D(_2580_),
    .Q(\genblk1[3].u_ce.Ain12b [7])
);

DFFPOSX1 _10755_ (
    .CLK(clk_bF$buf11),
    .D(_2581_),
    .Q(\genblk1[3].u_ce.Ain12b [4])
);

DFFPOSX1 _10756_ (
    .CLK(clk_bF$buf10),
    .D(_2582_),
    .Q(\genblk1[3].u_ce.Ain12b [5])
);

DFFPOSX1 _10757_ (
    .CLK(clk_bF$buf9),
    .D(_2583_),
    .Q(\genblk1[3].u_ce.Ain1 [0])
);

DFFPOSX1 _10758_ (
    .CLK(clk_bF$buf8),
    .D(_2584_),
    .Q(\genblk1[3].u_ce.Ain1 [1])
);

DFFPOSX1 _10759_ (
    .CLK(clk_bF$buf7),
    .D(_2585_),
    .Q(\genblk1[3].u_ce.Ain0 [0])
);

DFFPOSX1 _10760_ (
    .CLK(clk_bF$buf6),
    .D(_2586_),
    .Q(\genblk1[3].u_ce.Ain0 [1])
);

DFFPOSX1 _10761_ (
    .CLK(clk_bF$buf5),
    .D(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .Q(\genblk1[3].u_ce.LoadCtl [0])
);

DFFPOSX1 _10762_ (
    .CLK(clk_bF$buf4),
    .D(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .Q(\genblk1[3].u_ce.LoadCtl [1])
);

DFFPOSX1 _10763_ (
    .CLK(clk_bF$buf3),
    .D(\genblk1[3].u_ce.LoadCtl [1]),
    .Q(\genblk1[3].u_ce.LoadCtl [2])
);

DFFPOSX1 _10764_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[3].u_ce.LoadCtl [2]),
    .Q(\genblk1[3].u_ce.LoadCtl [3])
);

DFFPOSX1 _10765_ (
    .CLK(clk_bF$buf1),
    .D(\genblk1[3].u_ce.LoadCtl [3]),
    .Q(\genblk1[3].u_ce.LoadCtl [4])
);

DFFPOSX1 _10766_ (
    .CLK(clk_bF$buf0),
    .D(\genblk1[3].u_ce.LoadCtl [4]),
    .Q(\genblk1[3].u_ce.LoadCtl [5])
);

DFFPOSX1 _10767_ (
    .CLK(clk_bF$buf78),
    .D(\genblk1[3].u_ce.LoadCtl [5]),
    .Q(\genblk1[3].u_ce.Vld )
);

INVX1 _10768_ (
    .A(\genblk1[4].u_ce.Acalc [2]),
    .Y(_3432_)
);

INVX2 _10769_ (
    .A(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3433_)
);

NOR2X1 _10770_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3433_),
    .Y(_3434_)
);

INVX2 _10771_ (
    .A(_3434_),
    .Y(_3435_)
);

NOR2X1 _10772_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [10]),
    .Y(_3436_)
);

INVX4 _10773_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .Y(_3437_)
);

NOR2X1 _10774_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.LoadCtl [3]),
    .Y(_3438_)
);

OAI21X1 _10775_ (
    .A(_3437_),
    .B(\genblk1[4].u_ce.Acalc [8]),
    .C(_3438_),
    .Y(_3439_)
);

INVX2 _10776_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_3440_)
);

AND2X2 _10777_ (
    .A(_3440_),
    .B(\genblk1[4].u_ce.LoadCtl [3]),
    .Y(_3441_)
);

AOI22X1 _10778_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.Acalc [4]),
    .C(_3441_),
    .D(\genblk1[4].u_ce.Acalc [6]),
    .Y(_3442_)
);

OAI21X1 _10779_ (
    .A(_3436_),
    .B(_3439_),
    .C(_3442_),
    .Y(_3443_)
);

NOR2X1 _10780_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3444_)
);

AOI22X1 _10781_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.Acalc [0]),
    .C(_3443_),
    .D(_3444_),
    .Y(_3445_)
);

OAI21X1 _10782_ (
    .A(_3432_),
    .B(_3435_),
    .C(_3445_),
    .Y(\a[5] [0])
);

INVX1 _10783_ (
    .A(\genblk1[4].u_ce.Acalc [9]),
    .Y(_3446_)
);

OAI21X1 _10784_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [11]),
    .C(_3438_),
    .Y(_3447_)
);

AOI21X1 _10785_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3446_),
    .C(_3447_),
    .Y(_3448_)
);

INVX1 _10786_ (
    .A(\genblk1[4].u_ce.Acalc [5]),
    .Y(_3449_)
);

NAND2X1 _10787_ (
    .A(\genblk1[4].u_ce.Acalc [7]),
    .B(_3441_),
    .Y(_3450_)
);

OAI21X1 _10788_ (
    .A(_3440_),
    .B(_3449_),
    .C(_3450_),
    .Y(_3451_)
);

OAI21X1 _10789_ (
    .A(_3448_),
    .B(_3451_),
    .C(_3444_),
    .Y(_3452_)
);

AOI22X1 _10790_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.Acalc [1]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Acalc [3]),
    .Y(_3453_)
);

NAND2X1 _10791_ (
    .A(_3453_),
    .B(_3452_),
    .Y(\a[5] [1])
);

INVX1 _10792_ (
    .A(\genblk1[4].u_ce.Ycalc [10]),
    .Y(_3454_)
);

OAI21X1 _10793_ (
    .A(_3437_),
    .B(\genblk1[4].u_ce.Ycalc [8]),
    .C(_3438_),
    .Y(_3455_)
);

AOI21X1 _10794_ (
    .A(_3437_),
    .B(_3454_),
    .C(_3455_),
    .Y(_3456_)
);

INVX1 _10795_ (
    .A(\genblk1[4].u_ce.Ycalc [4]),
    .Y(_3457_)
);

NAND2X1 _10796_ (
    .A(\genblk1[4].u_ce.Ycalc [6]),
    .B(_3441_),
    .Y(_3458_)
);

OAI21X1 _10797_ (
    .A(_3440_),
    .B(_3457_),
    .C(_3458_),
    .Y(_3459_)
);

OAI21X1 _10798_ (
    .A(_3456_),
    .B(_3459_),
    .C(_3444_),
    .Y(_3460_)
);

AOI22X1 _10799_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.Ycalc [0]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Ycalc [2]),
    .Y(_3461_)
);

NAND2X1 _10800_ (
    .A(_3461_),
    .B(_3460_),
    .Y(\genblk1[4].u_ce.Y_ [0])
);

INVX1 _10801_ (
    .A(\genblk1[4].u_ce.Ycalc [9]),
    .Y(_3462_)
);

OAI21X1 _10802_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Ycalc [11]),
    .C(_3438_),
    .Y(_3463_)
);

AOI21X1 _10803_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3462_),
    .C(_3463_),
    .Y(_3464_)
);

INVX1 _10804_ (
    .A(\genblk1[4].u_ce.Ycalc [5]),
    .Y(_3465_)
);

NAND2X1 _10805_ (
    .A(\genblk1[4].u_ce.Ycalc [7]),
    .B(_3441_),
    .Y(_3466_)
);

OAI21X1 _10806_ (
    .A(_3440_),
    .B(_3465_),
    .C(_3466_),
    .Y(_3467_)
);

OAI21X1 _10807_ (
    .A(_3464_),
    .B(_3467_),
    .C(_3444_),
    .Y(_3468_)
);

AOI22X1 _10808_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.Ycalc [1]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3469_)
);

NAND2X1 _10809_ (
    .A(_3469_),
    .B(_3468_),
    .Y(\genblk1[4].u_ce.Y_ [1])
);

INVX1 _10810_ (
    .A(\genblk1[4].u_ce.Xcalc [8]),
    .Y(_3470_)
);

OAI21X1 _10811_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Xcalc [10]),
    .C(_3438_),
    .Y(_3471_)
);

AOI21X1 _10812_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3470_),
    .C(_3471_),
    .Y(_3472_)
);

INVX1 _10813_ (
    .A(\genblk1[4].u_ce.Xcalc [4]),
    .Y(_3473_)
);

NAND2X1 _10814_ (
    .A(\genblk1[4].u_ce.Xcalc [6]),
    .B(_3441_),
    .Y(_3474_)
);

OAI21X1 _10815_ (
    .A(_3440_),
    .B(_3473_),
    .C(_3474_),
    .Y(_3475_)
);

OAI21X1 _10816_ (
    .A(_3472_),
    .B(_3475_),
    .C(_3444_),
    .Y(_3476_)
);

AOI22X1 _10817_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Xcalc [0]),
    .C(_3434_),
    .D(\genblk1[4].u_ce.Xcalc [2]),
    .Y(_3477_)
);

NAND2X1 _10818_ (
    .A(_3477_),
    .B(_3476_),
    .Y(\genblk1[4].u_ce.X_ [0])
);

INVX1 _10819_ (
    .A(\genblk1[4].u_ce.Xcalc [3]),
    .Y(_3478_)
);

NOR2X1 _10820_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Xcalc [11]),
    .Y(_3479_)
);

OAI21X1 _10821_ (
    .A(_3437_),
    .B(\genblk1[4].u_ce.Xcalc [9]),
    .C(_3438_),
    .Y(_3480_)
);

AOI22X1 _10822_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.Xcalc [5]),
    .C(_3441_),
    .D(\genblk1[4].u_ce.Xcalc [7]),
    .Y(_3481_)
);

OAI21X1 _10823_ (
    .A(_3479_),
    .B(_3480_),
    .C(_3481_),
    .Y(_3482_)
);

AOI22X1 _10824_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.Xcalc [1]),
    .C(_3482_),
    .D(_3444_),
    .Y(_3483_)
);

OAI21X1 _10825_ (
    .A(_3478_),
    .B(_3435_),
    .C(_3483_),
    .Y(\genblk1[4].u_ce.X_ [1])
);

INVX1 _10826_ (
    .A(\genblk1[4].u_ce.Ycalc [0]),
    .Y(_3484_)
);

INVX1 _10827_ (
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .Y(_3485_)
);

INVX8 _10828_ (
    .A(1'h1),
    .Y(_3486_)
);

INVX8 _10829_ (
    .A(1'h0),
    .Y(_3487_)
);

INVX1 _10830_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_3488_)
);

NAND2X1 _10831_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3489_)
);

OAI21X1 _10832_ (
    .A(1'h0),
    .B(_3488_),
    .C(_3489_),
    .Y(_3490_)
);

INVX1 _10833_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .Y(_3491_)
);

NAND2X1 _10834_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3492_)
);

OAI21X1 _10835_ (
    .A(1'h0),
    .B(_3491_),
    .C(_3492_),
    .Y(_3493_)
);

MUX2X1 _10836_ (
    .A(_3493_),
    .B(_3490_),
    .S(_3487__bF$buf4),
    .Y(_3494_)
);

INVX1 _10837_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3495_)
);

NAND2X1 _10838_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3496_)
);

OAI21X1 _10839_ (
    .A(1'h0),
    .B(_3495_),
    .C(_3496_),
    .Y(_3497_)
);

INVX1 _10840_ (
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .Y(_3498_)
);

NAND2X1 _10841_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_3499_)
);

OAI21X1 _10842_ (
    .A(1'h0),
    .B(_3498_),
    .C(_3499_),
    .Y(_3500_)
);

MUX2X1 _10843_ (
    .A(_3500_),
    .B(_3497_),
    .S(_3487__bF$buf3),
    .Y(_3501_)
);

MUX2X1 _10844_ (
    .A(_3501_),
    .B(_3494_),
    .S(_3486__bF$buf4),
    .Y(_3502_)
);

NOR2X1 _10845_ (
    .A(_3485_),
    .B(_3502_),
    .Y(_3503_)
);

NAND2X1 _10846_ (
    .A(_3485_),
    .B(_3502_),
    .Y(_3504_)
);

INVX1 _10847_ (
    .A(_3504_),
    .Y(_3505_)
);

NAND2X1 _10848_ (
    .A(_3486__bF$buf3),
    .B(_3487__bF$buf2),
    .Y(_3506_)
);

OAI21X1 _10849_ (
    .A(1'h0),
    .B(_3506_),
    .C(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_3507_)
);

INVX2 _10850_ (
    .A(_3507_),
    .Y(_3508_)
);

OAI21X1 _10851_ (
    .A(_3503_),
    .B(_3505_),
    .C(_3508_),
    .Y(_3509_)
);

OAI21X1 _10852_ (
    .A(_3484_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3509_),
    .Y(_3352_)
);

INVX8 _10853_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_3510_)
);

NAND2X1 _10854_ (
    .A(\genblk1[4].u_ce.Ycalc [1]),
    .B(_3510__bF$buf4),
    .Y(_3511_)
);

NOR2X1 _10855_ (
    .A(1'h0),
    .B(_3506_),
    .Y(_3512_)
);

MUX2X1 _10856_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(\genblk1[4].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_3513_)
);

MUX2X1 _10857_ (
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .B(\genblk1[4].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_3514_)
);

MUX2X1 _10858_ (
    .A(_3514_),
    .B(_3513_),
    .S(_3487__bF$buf1),
    .Y(_3515_)
);

INVX2 _10859_ (
    .A(1'h0),
    .Y(_3516_)
);

NAND2X1 _10860_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(_3516_),
    .Y(_3517_)
);

AOI21X1 _10861_ (
    .A(_3517_),
    .B(_3496_),
    .C(_3487__bF$buf0),
    .Y(_3518_)
);

NAND3X1 _10862_ (
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .B(_3516_),
    .C(_3487__bF$buf4),
    .Y(_3519_)
);

NAND3X1 _10863_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(1'h0),
    .C(_3487__bF$buf3),
    .Y(_3520_)
);

NAND3X1 _10864_ (
    .A(_3486__bF$buf2),
    .B(_3520_),
    .C(_3519_),
    .Y(_3521_)
);

OAI22X1 _10865_ (
    .A(_3518_),
    .B(_3521_),
    .C(_3486__bF$buf1),
    .D(_3515_),
    .Y(_3522_)
);

INVX1 _10866_ (
    .A(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3523_)
);

INVX8 _10867_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_3524_)
);

INVX1 _10868_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3525_)
);

NAND2X1 _10869_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3526_)
);

OAI21X1 _10870_ (
    .A(1'h0),
    .B(_3525_),
    .C(_3526_),
    .Y(_3527_)
);

INVX1 _10871_ (
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3528_)
);

NAND2X1 _10872_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_3529_)
);

OAI21X1 _10873_ (
    .A(1'h0),
    .B(_3528_),
    .C(_3529_),
    .Y(_3530_)
);

MUX2X1 _10874_ (
    .A(_3530_),
    .B(_3527_),
    .S(_3487__bF$buf2),
    .Y(_3531_)
);

INVX1 _10875_ (
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3532_)
);

NAND2X1 _10876_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [4]),
    .Y(_3533_)
);

OAI21X1 _10877_ (
    .A(1'h0),
    .B(_3532_),
    .C(_3533_),
    .Y(_3534_)
);

INVX1 _10878_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .Y(_3535_)
);

NAND2X1 _10879_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3536_)
);

OAI21X1 _10880_ (
    .A(1'h0),
    .B(_3535_),
    .C(_3536_),
    .Y(_3537_)
);

MUX2X1 _10881_ (
    .A(_3537_),
    .B(_3534_),
    .S(_3487__bF$buf1),
    .Y(_3538_)
);

MUX2X1 _10882_ (
    .A(_3538_),
    .B(_3531_),
    .S(_3486__bF$buf0),
    .Y(_3539_)
);

NAND3X1 _10883_ (
    .A(_3524__bF$buf5),
    .B(_3502_),
    .C(_3539_),
    .Y(_3540_)
);

MUX2X1 _10884_ (
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_3541_)
);

MUX2X1 _10885_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_3542_)
);

MUX2X1 _10886_ (
    .A(_3542_),
    .B(_3541_),
    .S(_3487__bF$buf0),
    .Y(_3543_)
);

MUX2X1 _10887_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_3544_)
);

MUX2X1 _10888_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(\genblk1[4].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_3545_)
);

MUX2X1 _10889_ (
    .A(_3545_),
    .B(_3544_),
    .S(_3487__bF$buf4),
    .Y(_3546_)
);

MUX2X1 _10890_ (
    .A(_3546_),
    .B(_3543_),
    .S(_3486__bF$buf4),
    .Y(_3547_)
);

OAI21X1 _10891_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3522_),
    .C(_3547_),
    .Y(_3548_)
);

AOI21X1 _10892_ (
    .A(_3548_),
    .B(_3540_),
    .C(_3523_),
    .Y(_3549_)
);

INVX1 _10893_ (
    .A(_3549_),
    .Y(_3550_)
);

NAND3X1 _10894_ (
    .A(_3523_),
    .B(_3540_),
    .C(_3548_),
    .Y(_3551_)
);

AND2X2 _10895_ (
    .A(_3550_),
    .B(_3551_),
    .Y(_3552_)
);

OAI21X1 _10896_ (
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .B(_3522_),
    .C(_3552_),
    .Y(_3553_)
);

OR2X2 _10897_ (
    .A(_3552_),
    .B(_3504_),
    .Y(_3554_)
);

AOI21X1 _10898_ (
    .A(_3554_),
    .B(_3553_),
    .C(_3512_),
    .Y(_3555_)
);

OAI21X1 _10899_ (
    .A(_3510__bF$buf3),
    .B(_3555_),
    .C(_3511_),
    .Y(_3353_)
);

INVX1 _10900_ (
    .A(\genblk1[4].u_ce.ISout ),
    .Y(_3556_)
);

NAND2X1 _10901_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(\genblk1[3].u_ce.ISout ),
    .Y(_3557_)
);

OAI21X1 _10902_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .B(_3556_),
    .C(_3557_),
    .Y(_3354_)
);

NAND2X1 _10903_ (
    .A(\genblk1[4].u_ce.Ycalc [2]),
    .B(_3510__bF$buf2),
    .Y(_3558_)
);

AOI21X1 _10904_ (
    .A(_3504_),
    .B(_3551_),
    .C(_3549_),
    .Y(_3559_)
);

MUX2X1 _10905_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(\genblk1[4].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_3560_)
);

MUX2X1 _10906_ (
    .A(_3560_),
    .B(_3513_),
    .S(1'h0),
    .Y(_3561_)
);

MUX2X1 _10907_ (
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_3562_)
);

NAND2X1 _10908_ (
    .A(1'h0),
    .B(_3486__bF$buf3),
    .Y(_3563_)
);

OAI22X1 _10909_ (
    .A(_3563_),
    .B(_3514_),
    .C(_3562_),
    .D(_3506_),
    .Y(_3564_)
);

AOI21X1 _10910_ (
    .A(1'h1),
    .B(_3561_),
    .C(_3564_),
    .Y(_3565_)
);

AOI21X1 _10911_ (
    .A(_3547_),
    .B(_3522_),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_3566_)
);

NAND2X1 _10912_ (
    .A(_3565_),
    .B(_3566_),
    .Y(_3567_)
);

INVX1 _10913_ (
    .A(_3565_),
    .Y(_3568_)
);

OAI21X1 _10914_ (
    .A(_3502_),
    .B(_3539_),
    .C(_3524__bF$buf4),
    .Y(_3569_)
);

NAND2X1 _10915_ (
    .A(_3568_),
    .B(_3569_),
    .Y(_3570_)
);

AOI21X1 _10916_ (
    .A(_3570_),
    .B(_3567_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3571_)
);

NAND3X1 _10917_ (
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .B(_3567_),
    .C(_3570_),
    .Y(_3572_)
);

INVX1 _10918_ (
    .A(_3572_),
    .Y(_3573_)
);

OR2X2 _10919_ (
    .A(_3573_),
    .B(_3571_),
    .Y(_3574_)
);

NOR2X1 _10920_ (
    .A(_3559_),
    .B(_3574_),
    .Y(_3575_)
);

INVX1 _10921_ (
    .A(_3575_),
    .Y(_3576_)
);

OAI21X1 _10922_ (
    .A(_3571_),
    .B(_3573_),
    .C(_3559_),
    .Y(_3577_)
);

AOI21X1 _10923_ (
    .A(_3576_),
    .B(_3577_),
    .C(_3512_),
    .Y(_3578_)
);

INVX2 _10924_ (
    .A(_3512_),
    .Y(_3579_)
);

OAI21X1 _10925_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3579_),
    .C(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_3580_)
);

OAI21X1 _10926_ (
    .A(_3580_),
    .B(_3578_),
    .C(_3558_),
    .Y(_3355_)
);

INVX1 _10927_ (
    .A(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3581_)
);

INVX2 _10928_ (
    .A(_3580_),
    .Y(_3582_)
);

OAI21X1 _10929_ (
    .A(_3571_),
    .B(_3559_),
    .C(_3572_),
    .Y(_3583_)
);

INVX1 _10930_ (
    .A(_3583_),
    .Y(_3584_)
);

INVX1 _10931_ (
    .A(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3585_)
);

NAND3X1 _10932_ (
    .A(_3522_),
    .B(_3547_),
    .C(_3565_),
    .Y(_3586_)
);

INVX1 _10933_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .Y(_3587_)
);

NAND2X1 _10934_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3588_)
);

OAI21X1 _10935_ (
    .A(1'h0),
    .B(_3587_),
    .C(_3588_),
    .Y(_3589_)
);

NAND2X1 _10936_ (
    .A(_3487__bF$buf3),
    .B(_3541_),
    .Y(_3590_)
);

OAI21X1 _10937_ (
    .A(_3487__bF$buf2),
    .B(_3589_),
    .C(_3590_),
    .Y(_3591_)
);

NOR2X1 _10938_ (
    .A(1'h1),
    .B(_3487__bF$buf1),
    .Y(_3592_)
);

NOR2X1 _10939_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_3593_)
);

AOI22X1 _10940_ (
    .A(_3534_),
    .B(_3593_),
    .C(_3592_),
    .D(_3530_),
    .Y(_3594_)
);

OAI21X1 _10941_ (
    .A(_3486__bF$buf2),
    .B(_3591_),
    .C(_3594_),
    .Y(_3595_)
);

NAND3X1 _10942_ (
    .A(_3524__bF$buf3),
    .B(_3595_),
    .C(_3586_),
    .Y(_3596_)
);

INVX1 _10943_ (
    .A(_3586_),
    .Y(_3597_)
);

INVX1 _10944_ (
    .A(_3595_),
    .Y(_3598_)
);

OAI21X1 _10945_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3597_),
    .C(_3598_),
    .Y(_3599_)
);

NAND3X1 _10946_ (
    .A(_3585_),
    .B(_3596_),
    .C(_3599_),
    .Y(_3600_)
);

AOI21X1 _10947_ (
    .A(_3599_),
    .B(_3596_),
    .C(_3585_),
    .Y(_3601_)
);

INVX1 _10948_ (
    .A(_3601_),
    .Y(_3602_)
);

NAND2X1 _10949_ (
    .A(_3600_),
    .B(_3602_),
    .Y(_3603_)
);

AOI21X1 _10950_ (
    .A(_3603_),
    .B(_3584_),
    .C(_3512_),
    .Y(_3604_)
);

OAI21X1 _10951_ (
    .A(_3584_),
    .B(_3603_),
    .C(_3604_),
    .Y(_3605_)
);

AOI22X1 _10952_ (
    .A(_3581_),
    .B(_3510__bF$buf1),
    .C(_3605_),
    .D(_3582_),
    .Y(_3356_)
);

AOI21X1 _10953_ (
    .A(_3583_),
    .B(_3600_),
    .C(_3601_),
    .Y(_3606_)
);

INVX1 _10954_ (
    .A(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3607_)
);

INVX1 _10955_ (
    .A(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3608_)
);

NAND2X1 _10956_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3609_)
);

OAI21X1 _10957_ (
    .A(1'h0),
    .B(_3608_),
    .C(_3609_),
    .Y(_3610_)
);

NAND2X1 _10958_ (
    .A(_3487__bF$buf0),
    .B(_3560_),
    .Y(_3611_)
);

OAI21X1 _10959_ (
    .A(_3487__bF$buf4),
    .B(_3610_),
    .C(_3611_),
    .Y(_3612_)
);

NAND2X1 _10960_ (
    .A(_3486__bF$buf1),
    .B(_3515_),
    .Y(_3613_)
);

OAI21X1 _10961_ (
    .A(_3486__bF$buf0),
    .B(_3612_),
    .C(_3613_),
    .Y(_3614_)
);

INVX2 _10962_ (
    .A(_3614_),
    .Y(_3615_)
);

OAI21X1 _10963_ (
    .A(_3595_),
    .B(_3586_),
    .C(_3524__bF$buf2),
    .Y(_3616_)
);

OR2X2 _10964_ (
    .A(_3616_),
    .B(_3615_),
    .Y(_3617_)
);

NOR2X1 _10965_ (
    .A(_3595_),
    .B(_3586_),
    .Y(_3618_)
);

OAI21X1 _10966_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3618_),
    .C(_3615_),
    .Y(_3619_)
);

NAND3X1 _10967_ (
    .A(_3607_),
    .B(_3619_),
    .C(_3617_),
    .Y(_3620_)
);

NOR2X1 _10968_ (
    .A(_3615_),
    .B(_3616_),
    .Y(_3621_)
);

AND2X2 _10969_ (
    .A(_3616_),
    .B(_3615_),
    .Y(_3622_)
);

OAI21X1 _10970_ (
    .A(_3621_),
    .B(_3622_),
    .C(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3623_)
);

NAND2X1 _10971_ (
    .A(_3623_),
    .B(_3620_),
    .Y(_3624_)
);

AOI21X1 _10972_ (
    .A(_3606_),
    .B(_3624_),
    .C(_3512_),
    .Y(_3625_)
);

OAI21X1 _10973_ (
    .A(_3606_),
    .B(_3624_),
    .C(_3625_),
    .Y(_3626_)
);

AOI22X1 _10974_ (
    .A(_3457_),
    .B(_3510__bF$buf0),
    .C(_3626_),
    .D(_3582_),
    .Y(_3357_)
);

OAI21X1 _10975_ (
    .A(_3624_),
    .B(_3606_),
    .C(_3623_),
    .Y(_3627_)
);

INVX1 _10976_ (
    .A(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3628_)
);

NAND3X1 _10977_ (
    .A(_3598_),
    .B(_3615_),
    .C(_3597_),
    .Y(_3629_)
);

NAND2X1 _10978_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3630_)
);

INVX1 _10979_ (
    .A(_3630_),
    .Y(_3631_)
);

AOI21X1 _10980_ (
    .A(_3589_),
    .B(_3487__bF$buf3),
    .C(_3631_),
    .Y(_3632_)
);

NAND2X1 _10981_ (
    .A(_3486__bF$buf4),
    .B(_3543_),
    .Y(_3633_)
);

OAI21X1 _10982_ (
    .A(_3486__bF$buf3),
    .B(_3632_),
    .C(_3633_),
    .Y(_3634_)
);

NAND3X1 _10983_ (
    .A(_3524__bF$buf1),
    .B(_3634_),
    .C(_3629_),
    .Y(_3635_)
);

NOR3X1 _10984_ (
    .A(_3595_),
    .B(_3614_),
    .C(_3586_),
    .Y(_3636_)
);

INVX1 _10985_ (
    .A(_3634_),
    .Y(_3637_)
);

OAI21X1 _10986_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3636_),
    .C(_3637_),
    .Y(_3638_)
);

NAND3X1 _10987_ (
    .A(_3628_),
    .B(_3635_),
    .C(_3638_),
    .Y(_3639_)
);

AOI21X1 _10988_ (
    .A(_3638_),
    .B(_3635_),
    .C(_3628_),
    .Y(_3640_)
);

INVX1 _10989_ (
    .A(_3640_),
    .Y(_3641_)
);

NAND2X1 _10990_ (
    .A(_3639_),
    .B(_3641_),
    .Y(_3642_)
);

AND2X2 _10991_ (
    .A(_3627_),
    .B(_3642_),
    .Y(_3643_)
);

OAI21X1 _10992_ (
    .A(_3642_),
    .B(_3627_),
    .C(_3579_),
    .Y(_3644_)
);

OAI21X1 _10993_ (
    .A(_3644_),
    .B(_3643_),
    .C(_3582_),
    .Y(_3645_)
);

OAI21X1 _10994_ (
    .A(_3465_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_3645_),
    .Y(_3358_)
);

INVX1 _10995_ (
    .A(\genblk1[4].u_ce.Ycalc [6]),
    .Y(_3646_)
);

INVX1 _10996_ (
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3647_)
);

NAND3X1 _10997_ (
    .A(_3615_),
    .B(_3637_),
    .C(_3618_),
    .Y(_3648_)
);

AOI21X1 _10998_ (
    .A(_3610_),
    .B(_3487__bF$buf2),
    .C(_3631_),
    .Y(_3649_)
);

NAND2X1 _10999_ (
    .A(_3486__bF$buf2),
    .B(_3561_),
    .Y(_3650_)
);

OAI21X1 _11000_ (
    .A(_3486__bF$buf1),
    .B(_3649_),
    .C(_3650_),
    .Y(_3651_)
);

NAND3X1 _11001_ (
    .A(_3524__bF$buf0),
    .B(_3651_),
    .C(_3648_),
    .Y(_3652_)
);

INVX1 _11002_ (
    .A(_3651_),
    .Y(_3653_)
);

OAI21X1 _11003_ (
    .A(_3634_),
    .B(_3629_),
    .C(_3524__bF$buf5),
    .Y(_3654_)
);

NAND2X1 _11004_ (
    .A(_3653_),
    .B(_3654_),
    .Y(_3655_)
);

NAND3X1 _11005_ (
    .A(_3647_),
    .B(_3652_),
    .C(_3655_),
    .Y(_3656_)
);

NAND3X1 _11006_ (
    .A(_3524__bF$buf4),
    .B(_3653_),
    .C(_3648_),
    .Y(_3657_)
);

NAND2X1 _11007_ (
    .A(_3651_),
    .B(_3654_),
    .Y(_3658_)
);

NAND3X1 _11008_ (
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .B(_3657_),
    .C(_3658_),
    .Y(_3659_)
);

NAND2X1 _11009_ (
    .A(_3656_),
    .B(_3659_),
    .Y(_3660_)
);

AOI21X1 _11010_ (
    .A(_3617_),
    .B(_3619_),
    .C(_3607_),
    .Y(_3661_)
);

NOR2X1 _11011_ (
    .A(_3661_),
    .B(_3640_),
    .Y(_3662_)
);

OAI21X1 _11012_ (
    .A(_3624_),
    .B(_3606_),
    .C(_3662_),
    .Y(_3663_)
);

NAND2X1 _11013_ (
    .A(_3639_),
    .B(_3663_),
    .Y(_3664_)
);

AOI21X1 _11014_ (
    .A(_3664_),
    .B(_3660_),
    .C(_3512_),
    .Y(_3665_)
);

OAI21X1 _11015_ (
    .A(_3660_),
    .B(_3664_),
    .C(_3665_),
    .Y(_3666_)
);

AOI22X1 _11016_ (
    .A(_3646_),
    .B(_3510__bF$buf4),
    .C(_3666_),
    .D(_3582_),
    .Y(_3359_)
);

INVX1 _11017_ (
    .A(\genblk1[4].u_ce.Ycalc [7]),
    .Y(_3667_)
);

AOI21X1 _11018_ (
    .A(_3655_),
    .B(_3652_),
    .C(_3647_),
    .Y(_3668_)
);

AND2X2 _11019_ (
    .A(_3620_),
    .B(_3623_),
    .Y(_3669_)
);

NAND3X1 _11020_ (
    .A(_3639_),
    .B(_3641_),
    .C(_3669_),
    .Y(_3670_)
);

AOI21X1 _11021_ (
    .A(_3661_),
    .B(_3639_),
    .C(_3640_),
    .Y(_3671_)
);

OAI21X1 _11022_ (
    .A(_3606_),
    .B(_3670_),
    .C(_3671_),
    .Y(_3672_)
);

AOI21X1 _11023_ (
    .A(_3672_),
    .B(_3656_),
    .C(_3668_),
    .Y(_3673_)
);

INVX1 _11024_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3674_)
);

NAND3X1 _11025_ (
    .A(_3637_),
    .B(_3653_),
    .C(_3636_),
    .Y(_3675_)
);

INVX1 _11026_ (
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3676_)
);

NOR2X1 _11027_ (
    .A(_3486__bF$buf0),
    .B(_3676_),
    .Y(_3677_)
);

INVX1 _11028_ (
    .A(_3677_),
    .Y(_3678_)
);

OAI21X1 _11029_ (
    .A(1'h1),
    .B(_3591_),
    .C(_3678_),
    .Y(_3679_)
);

NAND3X1 _11030_ (
    .A(_3524__bF$buf3),
    .B(_3679_),
    .C(_3675_),
    .Y(_3680_)
);

INVX1 _11031_ (
    .A(_3679_),
    .Y(_3681_)
);

OAI21X1 _11032_ (
    .A(_3651_),
    .B(_3648_),
    .C(_3524__bF$buf2),
    .Y(_3682_)
);

NAND2X1 _11033_ (
    .A(_3681_),
    .B(_3682_),
    .Y(_3683_)
);

NAND3X1 _11034_ (
    .A(_3674_),
    .B(_3680_),
    .C(_3683_),
    .Y(_3684_)
);

NAND3X1 _11035_ (
    .A(_3524__bF$buf1),
    .B(_3681_),
    .C(_3675_),
    .Y(_3685_)
);

NAND2X1 _11036_ (
    .A(_3679_),
    .B(_3682_),
    .Y(_3686_)
);

NAND3X1 _11037_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(_3685_),
    .C(_3686_),
    .Y(_3687_)
);

NAND2X1 _11038_ (
    .A(_3684_),
    .B(_3687_),
    .Y(_3688_)
);

INVX1 _11039_ (
    .A(_3688_),
    .Y(_3689_)
);

NOR2X1 _11040_ (
    .A(_3689_),
    .B(_3673_),
    .Y(_3690_)
);

OAI21X1 _11041_ (
    .A(_3660_),
    .B(_3664_),
    .C(_3659_),
    .Y(_3691_)
);

OAI21X1 _11042_ (
    .A(_3688_),
    .B(_3691_),
    .C(_3579_),
    .Y(_3692_)
);

OAI21X1 _11043_ (
    .A(_3524__bF$buf0),
    .B(_3579_),
    .C(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_3693_)
);

INVX1 _11044_ (
    .A(_3693_),
    .Y(_3694_)
);

OAI21X1 _11045_ (
    .A(_3692_),
    .B(_3690_),
    .C(_3694_),
    .Y(_3695_)
);

OAI21X1 _11046_ (
    .A(_3667_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_3695_),
    .Y(_3360_)
);

INVX1 _11047_ (
    .A(\genblk1[4].u_ce.Ycalc [8]),
    .Y(_3696_)
);

OAI21X1 _11048_ (
    .A(_3659_),
    .B(_3688_),
    .C(_3687_),
    .Y(_3697_)
);

NOR2X1 _11049_ (
    .A(_3660_),
    .B(_3688_),
    .Y(_3698_)
);

AOI21X1 _11050_ (
    .A(_3698_),
    .B(_3672_),
    .C(_3697_),
    .Y(_3699_)
);

INVX1 _11051_ (
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3700_)
);

OR2X2 _11052_ (
    .A(_3675_),
    .B(_3679_),
    .Y(_3701_)
);

OAI21X1 _11053_ (
    .A(1'h1),
    .B(_3612_),
    .C(_3678_),
    .Y(_3702_)
);

NAND3X1 _11054_ (
    .A(_3524__bF$buf5),
    .B(_3702_),
    .C(_3701_),
    .Y(_3703_)
);

NOR2X1 _11055_ (
    .A(_3679_),
    .B(_3675_),
    .Y(_3704_)
);

INVX1 _11056_ (
    .A(_3702_),
    .Y(_3705_)
);

OAI21X1 _11057_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3704_),
    .C(_3705_),
    .Y(_3706_)
);

NAND3X1 _11058_ (
    .A(_3700_),
    .B(_3706_),
    .C(_3703_),
    .Y(_3707_)
);

NAND3X1 _11059_ (
    .A(_3524__bF$buf4),
    .B(_3705_),
    .C(_3701_),
    .Y(_3708_)
);

OAI21X1 _11060_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3704_),
    .C(_3702_),
    .Y(_3709_)
);

NAND3X1 _11061_ (
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .B(_3709_),
    .C(_3708_),
    .Y(_3710_)
);

AND2X2 _11062_ (
    .A(_3707_),
    .B(_3710_),
    .Y(_3711_)
);

INVX1 _11063_ (
    .A(_3711_),
    .Y(_3712_)
);

AOI21X1 _11064_ (
    .A(_3699_),
    .B(_3712_),
    .C(_3512_),
    .Y(_3713_)
);

OAI21X1 _11065_ (
    .A(_3699_),
    .B(_3712_),
    .C(_3713_),
    .Y(_3714_)
);

AOI22X1 _11066_ (
    .A(_3696_),
    .B(_3510__bF$buf3),
    .C(_3714_),
    .D(_3694_),
    .Y(_3361_)
);

NAND2X1 _11067_ (
    .A(_3668_),
    .B(_3684_),
    .Y(_3715_)
);

AND2X2 _11068_ (
    .A(_3715_),
    .B(_3687_),
    .Y(_3716_)
);

AND2X2 _11069_ (
    .A(_3656_),
    .B(_3659_),
    .Y(_3717_)
);

NAND3X1 _11070_ (
    .A(_3684_),
    .B(_3687_),
    .C(_3717_),
    .Y(_3718_)
);

OAI21X1 _11071_ (
    .A(_3664_),
    .B(_3718_),
    .C(_3716_),
    .Y(_3719_)
);

INVX1 _11072_ (
    .A(_3710_),
    .Y(_3720_)
);

AOI21X1 _11073_ (
    .A(_3719_),
    .B(_3707_),
    .C(_3720_),
    .Y(_3721_)
);

INVX1 _11074_ (
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_3722_)
);

NOR3X1 _11075_ (
    .A(_3679_),
    .B(_3702_),
    .C(_3675_),
    .Y(_3723_)
);

INVX1 _11076_ (
    .A(_3723_),
    .Y(_3724_)
);

OAI21X1 _11077_ (
    .A(1'h1),
    .B(_3632_),
    .C(_3678_),
    .Y(_3725_)
);

NAND3X1 _11078_ (
    .A(_3524__bF$buf3),
    .B(_3725_),
    .C(_3724_),
    .Y(_3726_)
);

INVX1 _11079_ (
    .A(_3725_),
    .Y(_3727_)
);

OAI21X1 _11080_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3723_),
    .C(_3727_),
    .Y(_3728_)
);

NAND3X1 _11081_ (
    .A(_3722_),
    .B(_3728_),
    .C(_3726_),
    .Y(_3729_)
);

NAND3X1 _11082_ (
    .A(_3524__bF$buf2),
    .B(_3727_),
    .C(_3724_),
    .Y(_3730_)
);

OAI21X1 _11083_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3723_),
    .C(_3725_),
    .Y(_3731_)
);

NAND3X1 _11084_ (
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .B(_3731_),
    .C(_3730_),
    .Y(_3732_)
);

AND2X2 _11085_ (
    .A(_3729_),
    .B(_3732_),
    .Y(_3733_)
);

AND2X2 _11086_ (
    .A(_3721_),
    .B(_3733_),
    .Y(_3734_)
);

OAI21X1 _11087_ (
    .A(_3733_),
    .B(_3721_),
    .C(_3579_),
    .Y(_3735_)
);

OAI21X1 _11088_ (
    .A(_3735_),
    .B(_3734_),
    .C(_3582_),
    .Y(_3736_)
);

OAI21X1 _11089_ (
    .A(_3462_),
    .B(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .C(_3736_),
    .Y(_3362_)
);

INVX1 _11090_ (
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .Y(_3737_)
);

OAI21X1 _11091_ (
    .A(1'h1),
    .B(_3649_),
    .C(_3678_),
    .Y(_3738_)
);

INVX1 _11092_ (
    .A(_3738_),
    .Y(_3739_)
);

AOI21X1 _11093_ (
    .A(_3723_),
    .B(_3727_),
    .C(_3739_),
    .Y(_3740_)
);

NAND3X1 _11094_ (
    .A(_3727_),
    .B(_3739_),
    .C(_3723_),
    .Y(_3741_)
);

NAND2X1 _11095_ (
    .A(_3524__bF$buf1),
    .B(_3741_),
    .Y(_3742_)
);

NAND2X1 _11096_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3738_),
    .Y(_3743_)
);

OAI21X1 _11097_ (
    .A(_3740_),
    .B(_3742_),
    .C(_3743_),
    .Y(_3744_)
);

NAND2X1 _11098_ (
    .A(_3737_),
    .B(_3744_),
    .Y(_3745_)
);

INVX1 _11099_ (
    .A(_3740_),
    .Y(_3746_)
);

AND2X2 _11100_ (
    .A(_3741_),
    .B(_3524__bF$buf0),
    .Y(_3747_)
);

NAND2X1 _11101_ (
    .A(_3746_),
    .B(_3747_),
    .Y(_3748_)
);

NAND3X1 _11102_ (
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .B(_3743_),
    .C(_3748_),
    .Y(_3749_)
);

NAND2X1 _11103_ (
    .A(_3745_),
    .B(_3749_),
    .Y(_3750_)
);

AOI21X1 _11104_ (
    .A(_3726_),
    .B(_3728_),
    .C(_3722_),
    .Y(_3751_)
);

AOI21X1 _11105_ (
    .A(_3720_),
    .B(_3729_),
    .C(_3751_),
    .Y(_3752_)
);

NAND3X1 _11106_ (
    .A(_3711_),
    .B(_3733_),
    .C(_3719_),
    .Y(_3753_)
);

AOI21X1 _11107_ (
    .A(_3753_),
    .B(_3752_),
    .C(_3750_),
    .Y(_3754_)
);

AND2X2 _11108_ (
    .A(_3749_),
    .B(_3745_),
    .Y(_3755_)
);

NAND3X1 _11109_ (
    .A(_3729_),
    .B(_3732_),
    .C(_3711_),
    .Y(_3756_)
);

OAI21X1 _11110_ (
    .A(_3756_),
    .B(_3699_),
    .C(_3752_),
    .Y(_3757_)
);

OAI21X1 _11111_ (
    .A(_3755_),
    .B(_3757_),
    .C(_3579_),
    .Y(_3758_)
);

OR2X2 _11112_ (
    .A(_3758_),
    .B(_3754_),
    .Y(_3759_)
);

AOI22X1 _11113_ (
    .A(_3454_),
    .B(_3510__bF$buf2),
    .C(_3759_),
    .D(_3582_),
    .Y(_3363_)
);

NAND2X1 _11114_ (
    .A(\genblk1[4].u_ce.Ycalc [11]),
    .B(_3510__bF$buf1),
    .Y(_3760_)
);

INVX1 _11115_ (
    .A(_3749_),
    .Y(_3761_)
);

NAND2X1 _11116_ (
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .B(_3676_),
    .Y(_3762_)
);

INVX1 _11117_ (
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_3763_)
);

NAND2X1 _11118_ (
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .B(_3763_),
    .Y(_3764_)
);

NAND2X1 _11119_ (
    .A(_3762_),
    .B(_3764_),
    .Y(_3765_)
);

INVX1 _11120_ (
    .A(_3765_),
    .Y(_3766_)
);

NAND2X1 _11121_ (
    .A(_3766_),
    .B(_3742_),
    .Y(_3767_)
);

NAND2X1 _11122_ (
    .A(_3765_),
    .B(_3747_),
    .Y(_3768_)
);

NAND2X1 _11123_ (
    .A(_3767_),
    .B(_3768_),
    .Y(_3769_)
);

INVX1 _11124_ (
    .A(_3769_),
    .Y(_3770_)
);

NOR3X1 _11125_ (
    .A(_3761_),
    .B(_3770_),
    .C(_3754_),
    .Y(_3771_)
);

AOI21X1 _11126_ (
    .A(_3757_),
    .B(_3755_),
    .C(_3761_),
    .Y(_3772_)
);

OAI21X1 _11127_ (
    .A(_3769_),
    .B(_3772_),
    .C(_3579_),
    .Y(_3773_)
);

OAI21X1 _11128_ (
    .A(_3771_),
    .B(_3773_),
    .C(_3582_),
    .Y(_3774_)
);

NAND2X1 _11129_ (
    .A(_3760_),
    .B(_3774_),
    .Y(_3364_)
);

NAND2X1 _11130_ (
    .A(\genblk1[4].u_ce.Xcalc [0]),
    .B(_3510__bF$buf0),
    .Y(_3775_)
);

INVX1 _11131_ (
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3776_)
);

NAND2X1 _11132_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3777_)
);

OAI21X1 _11133_ (
    .A(1'h0),
    .B(_3776_),
    .C(_3777_),
    .Y(_3778_)
);

NAND2X1 _11134_ (
    .A(1'h0),
    .B(_3778_),
    .Y(_3779_)
);

NOR2X1 _11135_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_3780_)
);

NOR2X1 _11136_ (
    .A(1'h0),
    .B(_3516_),
    .Y(_3781_)
);

AOI22X1 _11137_ (
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .B(_3780_),
    .C(_3781_),
    .D(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3782_)
);

NAND3X1 _11138_ (
    .A(_3486__bF$buf4),
    .B(_3779_),
    .C(_3782_),
    .Y(_3783_)
);

NAND2X1 _11139_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3784_)
);

OAI21X1 _11140_ (
    .A(1'h0),
    .B(_3647_),
    .C(_3784_),
    .Y(_3785_)
);

NAND2X1 _11141_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3786_)
);

OAI21X1 _11142_ (
    .A(1'h0),
    .B(_3607_),
    .C(_3786_),
    .Y(_3787_)
);

MUX2X1 _11143_ (
    .A(_3787_),
    .B(_3785_),
    .S(_3487__bF$buf1),
    .Y(_3788_)
);

NAND2X1 _11144_ (
    .A(1'h1),
    .B(_3788_),
    .Y(_3789_)
);

AND2X2 _11145_ (
    .A(_3783_),
    .B(_3789_),
    .Y(_3790_)
);

NOR2X1 _11146_ (
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .B(_3790_),
    .Y(_3791_)
);

NAND2X1 _11147_ (
    .A(_3487__bF$buf0),
    .B(_3787_),
    .Y(_3792_)
);

NAND2X1 _11148_ (
    .A(1'h0),
    .B(_3785_),
    .Y(_3793_)
);

NAND2X1 _11149_ (
    .A(_3792_),
    .B(_3793_),
    .Y(_3794_)
);

OAI21X1 _11150_ (
    .A(_3486__bF$buf3),
    .B(_3794_),
    .C(_3783_),
    .Y(_3795_)
);

OAI21X1 _11151_ (
    .A(_3498_),
    .B(_3795_),
    .C(_3508_),
    .Y(_3796_)
);

OAI21X1 _11152_ (
    .A(_3796_),
    .B(_3791_),
    .C(_3775_),
    .Y(_3365_)
);

NAND2X1 _11153_ (
    .A(\genblk1[4].u_ce.Xcalc [1]),
    .B(_3510__bF$buf4),
    .Y(_3797_)
);

NOR2X1 _11154_ (
    .A(_3498_),
    .B(_3795_),
    .Y(_3798_)
);

NAND2X1 _11155_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3799_)
);

OAI21X1 _11156_ (
    .A(1'h0),
    .B(_3585_),
    .C(_3799_),
    .Y(_3800_)
);

NAND2X1 _11157_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3801_)
);

OAI21X1 _11158_ (
    .A(1'h0),
    .B(_3523_),
    .C(_3801_),
    .Y(_3802_)
);

MUX2X1 _11159_ (
    .A(_3802_),
    .B(_3800_),
    .S(_3487__bF$buf4),
    .Y(_3803_)
);

NAND2X1 _11160_ (
    .A(_3486__bF$buf2),
    .B(_3803_),
    .Y(_3804_)
);

NAND2X1 _11161_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3805_)
);

OAI21X1 _11162_ (
    .A(1'h0),
    .B(_3674_),
    .C(_3805_),
    .Y(_3806_)
);

INVX1 _11163_ (
    .A(_3806_),
    .Y(_3807_)
);

NAND2X1 _11164_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3808_)
);

OAI21X1 _11165_ (
    .A(1'h0),
    .B(_3628_),
    .C(_3808_),
    .Y(_3809_)
);

NAND2X1 _11166_ (
    .A(_3487__bF$buf3),
    .B(_3809_),
    .Y(_3810_)
);

OAI21X1 _11167_ (
    .A(_3487__bF$buf2),
    .B(_3807_),
    .C(_3810_),
    .Y(_3811_)
);

OAI21X1 _11168_ (
    .A(_3486__bF$buf1),
    .B(_3811_),
    .C(_3804_),
    .Y(_3812_)
);

NAND3X1 _11169_ (
    .A(_3524__bF$buf5),
    .B(_3812_),
    .C(_3790_),
    .Y(_3813_)
);

MUX2X1 _11170_ (
    .A(_3809_),
    .B(_3806_),
    .S(_3487__bF$buf1),
    .Y(_3814_)
);

MUX2X1 _11171_ (
    .A(_3814_),
    .B(_3803_),
    .S(1'h1),
    .Y(_3815_)
);

OAI21X1 _11172_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3795_),
    .C(_3815_),
    .Y(_3816_)
);

AOI21X1 _11173_ (
    .A(_3813_),
    .B(_3816_),
    .C(_3535_),
    .Y(_3817_)
);

INVX1 _11174_ (
    .A(_3817_),
    .Y(_3818_)
);

NAND3X1 _11175_ (
    .A(_3535_),
    .B(_3816_),
    .C(_3813_),
    .Y(_3819_)
);

AND2X2 _11176_ (
    .A(_3818_),
    .B(_3819_),
    .Y(_3820_)
);

NAND2X1 _11177_ (
    .A(_3798_),
    .B(_3820_),
    .Y(_3821_)
);

OR2X2 _11178_ (
    .A(_3820_),
    .B(_3798_),
    .Y(_3822_)
);

AOI21X1 _11179_ (
    .A(_3822_),
    .B(_3821_),
    .C(_3512_),
    .Y(_3823_)
);

OAI21X1 _11180_ (
    .A(_3510__bF$buf3),
    .B(_3823_),
    .C(_3797_),
    .Y(_3366_)
);

NAND2X1 _11181_ (
    .A(\genblk1[4].u_ce.Xcalc [2]),
    .B(_3510__bF$buf2),
    .Y(_3824_)
);

AOI21X1 _11182_ (
    .A(_3798_),
    .B(_3819_),
    .C(_3817_),
    .Y(_3825_)
);

NAND2X1 _11183_ (
    .A(_3795_),
    .B(_3812_),
    .Y(_3826_)
);

NAND2X1 _11184_ (
    .A(1'h0),
    .B(_3722_),
    .Y(_3827_)
);

OAI21X1 _11185_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .C(_3827_),
    .Y(_3828_)
);

NAND2X1 _11186_ (
    .A(_3487__bF$buf0),
    .B(_3785_),
    .Y(_3829_)
);

OAI21X1 _11187_ (
    .A(_3487__bF$buf4),
    .B(_3828_),
    .C(_3829_),
    .Y(_3830_)
);

NAND2X1 _11188_ (
    .A(_3593_),
    .B(_3778_),
    .Y(_3831_)
);

NAND2X1 _11189_ (
    .A(_3787_),
    .B(_3592_),
    .Y(_3832_)
);

NAND2X1 _11190_ (
    .A(_3831_),
    .B(_3832_),
    .Y(_3833_)
);

AOI21X1 _11191_ (
    .A(_3830_),
    .B(1'h1),
    .C(_3833_),
    .Y(_3834_)
);

INVX1 _11192_ (
    .A(_3834_),
    .Y(_3835_)
);

NAND3X1 _11193_ (
    .A(_3524__bF$buf4),
    .B(_3835_),
    .C(_3826_),
    .Y(_3836_)
);

AOI21X1 _11194_ (
    .A(_3783_),
    .B(_3789_),
    .C(_3815_),
    .Y(_3837_)
);

OAI21X1 _11195_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3837_),
    .C(_3834_),
    .Y(_3838_)
);

NAND3X1 _11196_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(_3838_),
    .C(_3836_),
    .Y(_3839_)
);

INVX1 _11197_ (
    .A(_3839_),
    .Y(_3840_)
);

AOI21X1 _11198_ (
    .A(_3836_),
    .B(_3838_),
    .C(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3841_)
);

NOR2X1 _11199_ (
    .A(_3841_),
    .B(_3840_),
    .Y(_3842_)
);

AND2X2 _11200_ (
    .A(_3842_),
    .B(_3825_),
    .Y(_3843_)
);

NOR2X1 _11201_ (
    .A(_3825_),
    .B(_3842_),
    .Y(_3844_)
);

OAI21X1 _11202_ (
    .A(_3844_),
    .B(_3843_),
    .C(_3579_),
    .Y(_3845_)
);

OAI21X1 _11203_ (
    .A(_3510__bF$buf1),
    .B(_3845_),
    .C(_3824_),
    .Y(_3367_)
);

OAI21X1 _11204_ (
    .A(_3841_),
    .B(_3825_),
    .C(_3839_),
    .Y(_3846_)
);

INVX1 _11205_ (
    .A(_3846_),
    .Y(_3847_)
);

NAND2X1 _11206_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [10]),
    .Y(_3848_)
);

OAI21X1 _11207_ (
    .A(1'h0),
    .B(_3722_),
    .C(_3848_),
    .Y(_3849_)
);

MUX2X1 _11208_ (
    .A(_3849_),
    .B(_3806_),
    .S(1'h0),
    .Y(_3850_)
);

NOR2X1 _11209_ (
    .A(_3486__bF$buf0),
    .B(_3850_),
    .Y(_3851_)
);

NAND2X1 _11210_ (
    .A(_3593_),
    .B(_3800_),
    .Y(_3852_)
);

NAND2X1 _11211_ (
    .A(_3809_),
    .B(_3592_),
    .Y(_3853_)
);

NAND2X1 _11212_ (
    .A(_3852_),
    .B(_3853_),
    .Y(_3854_)
);

OR2X2 _11213_ (
    .A(_3851_),
    .B(_3854_),
    .Y(_3855_)
);

OAI21X1 _11214_ (
    .A(_3835_),
    .B(_3826_),
    .C(_3524__bF$buf3),
    .Y(_3856_)
);

OR2X2 _11215_ (
    .A(_3856_),
    .B(_3855_),
    .Y(_3857_)
);

OAI21X1 _11216_ (
    .A(_3851_),
    .B(_3854_),
    .C(_3856_),
    .Y(_3858_)
);

AOI21X1 _11217_ (
    .A(_3857_),
    .B(_3858_),
    .C(_3532_),
    .Y(_3859_)
);

INVX1 _11218_ (
    .A(_3859_),
    .Y(_3860_)
);

NAND3X1 _11219_ (
    .A(_3532_),
    .B(_3858_),
    .C(_3857_),
    .Y(_3861_)
);

NAND2X1 _11220_ (
    .A(_3861_),
    .B(_3860_),
    .Y(_3862_)
);

OR2X2 _11221_ (
    .A(_3862_),
    .B(_3847_),
    .Y(_3863_)
);

NAND2X1 _11222_ (
    .A(_3847_),
    .B(_3862_),
    .Y(_3864_)
);

NAND2X1 _11223_ (
    .A(_3864_),
    .B(_3863_),
    .Y(_3865_)
);

AOI22X1 _11224_ (
    .A(_3478_),
    .B(_3510__bF$buf0),
    .C(_3865_),
    .D(_3508_),
    .Y(_3368_)
);

AOI21X1 _11225_ (
    .A(_3846_),
    .B(_3861_),
    .C(_3859_),
    .Y(_3866_)
);

NAND2X1 _11226_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_3867_)
);

OAI21X1 _11227_ (
    .A(1'h0),
    .B(_3737_),
    .C(_3867_),
    .Y(_3868_)
);

NAND2X1 _11228_ (
    .A(1'h0),
    .B(_3868_),
    .Y(_3869_)
);

OAI21X1 _11229_ (
    .A(1'h0),
    .B(_3828_),
    .C(_3869_),
    .Y(_3870_)
);

NAND2X1 _11230_ (
    .A(1'h1),
    .B(_3870_),
    .Y(_3871_)
);

OAI21X1 _11231_ (
    .A(1'h1),
    .B(_3788_),
    .C(_3871_),
    .Y(_3872_)
);

INVX1 _11232_ (
    .A(_3872_),
    .Y(_3873_)
);

NAND3X1 _11233_ (
    .A(_3834_),
    .B(_3795_),
    .C(_3812_),
    .Y(_3874_)
);

OAI21X1 _11234_ (
    .A(_3855_),
    .B(_3874_),
    .C(_3524__bF$buf2),
    .Y(_3875_)
);

OR2X2 _11235_ (
    .A(_3875_),
    .B(_3873_),
    .Y(_3876_)
);

NOR2X1 _11236_ (
    .A(_3855_),
    .B(_3874_),
    .Y(_3877_)
);

OAI21X1 _11237_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3877_),
    .C(_3873_),
    .Y(_3878_)
);

NAND3X1 _11238_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(_3878_),
    .C(_3876_),
    .Y(_3879_)
);

OR2X2 _11239_ (
    .A(_3875_),
    .B(_3872_),
    .Y(_3880_)
);

OAI21X1 _11240_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3877_),
    .C(_3872_),
    .Y(_3881_)
);

NAND3X1 _11241_ (
    .A(_3491_),
    .B(_3881_),
    .C(_3880_),
    .Y(_3882_)
);

NAND2X1 _11242_ (
    .A(_3879_),
    .B(_3882_),
    .Y(_3883_)
);

OR2X2 _11243_ (
    .A(_3866_),
    .B(_3883_),
    .Y(_3884_)
);

NAND2X1 _11244_ (
    .A(_3883_),
    .B(_3866_),
    .Y(_3885_)
);

NAND2X1 _11245_ (
    .A(_3885_),
    .B(_3884_),
    .Y(_3886_)
);

AOI22X1 _11246_ (
    .A(_3473_),
    .B(_3510__bF$buf4),
    .C(_3886_),
    .D(_3508_),
    .Y(_3369_)
);

INVX1 _11247_ (
    .A(\genblk1[4].u_ce.Xcalc [5]),
    .Y(_3887_)
);

OAI21X1 _11248_ (
    .A(_3883_),
    .B(_3866_),
    .C(_3879_),
    .Y(_3888_)
);

NAND2X1 _11249_ (
    .A(_3873_),
    .B(_3877_),
    .Y(_3889_)
);

NOR2X1 _11250_ (
    .A(_3487__bF$buf3),
    .B(_3763_),
    .Y(_3890_)
);

AOI21X1 _11251_ (
    .A(_3487__bF$buf2),
    .B(_3849_),
    .C(_3890_),
    .Y(_3891_)
);

NAND2X1 _11252_ (
    .A(_3486__bF$buf4),
    .B(_3811_),
    .Y(_3892_)
);

OAI21X1 _11253_ (
    .A(_3486__bF$buf3),
    .B(_3891_),
    .C(_3892_),
    .Y(_3893_)
);

INVX1 _11254_ (
    .A(_3893_),
    .Y(_3894_)
);

NAND3X1 _11255_ (
    .A(_3524__bF$buf1),
    .B(_3894_),
    .C(_3889_),
    .Y(_3895_)
);

NOR2X1 _11256_ (
    .A(_3854_),
    .B(_3851_),
    .Y(_3896_)
);

NAND3X1 _11257_ (
    .A(_3834_),
    .B(_3896_),
    .C(_3837_),
    .Y(_3897_)
);

OAI21X1 _11258_ (
    .A(_3872_),
    .B(_3897_),
    .C(_3524__bF$buf0),
    .Y(_3898_)
);

NAND2X1 _11259_ (
    .A(_3893_),
    .B(_3898_),
    .Y(_3899_)
);

AOI21X1 _11260_ (
    .A(_3895_),
    .B(_3899_),
    .C(_3528_),
    .Y(_3900_)
);

INVX1 _11261_ (
    .A(_3900_),
    .Y(_3901_)
);

NAND3X1 _11262_ (
    .A(_3528_),
    .B(_3899_),
    .C(_3895_),
    .Y(_3902_)
);

NAND2X1 _11263_ (
    .A(_3902_),
    .B(_3901_),
    .Y(_3903_)
);

NOR2X1 _11264_ (
    .A(_3903_),
    .B(_3888_),
    .Y(_3904_)
);

AND2X2 _11265_ (
    .A(_3888_),
    .B(_3903_),
    .Y(_3905_)
);

OAI21X1 _11266_ (
    .A(_3904_),
    .B(_3905_),
    .C(_3508_),
    .Y(_3906_)
);

OAI21X1 _11267_ (
    .A(_3887_),
    .B(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .C(_3906_),
    .Y(_3370_)
);

INVX1 _11268_ (
    .A(\genblk1[4].u_ce.Xcalc [6]),
    .Y(_3907_)
);

NAND3X1 _11269_ (
    .A(_3873_),
    .B(_3894_),
    .C(_3877_),
    .Y(_3908_)
);

AOI21X1 _11270_ (
    .A(_3487__bF$buf1),
    .B(_3868_),
    .C(_3890_),
    .Y(_3909_)
);

NAND2X1 _11271_ (
    .A(1'h1),
    .B(_3909_),
    .Y(_3910_)
);

OAI21X1 _11272_ (
    .A(1'h1),
    .B(_3830_),
    .C(_3910_),
    .Y(_3911_)
);

NAND3X1 _11273_ (
    .A(_3524__bF$buf5),
    .B(_3911_),
    .C(_3908_),
    .Y(_3912_)
);

NOR3X1 _11274_ (
    .A(_3872_),
    .B(_3893_),
    .C(_3897_),
    .Y(_3913_)
);

INVX1 _11275_ (
    .A(_3911_),
    .Y(_3914_)
);

OAI21X1 _11276_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3913_),
    .C(_3914_),
    .Y(_3915_)
);

NAND2X1 _11277_ (
    .A(_3912_),
    .B(_3915_),
    .Y(_3916_)
);

NAND2X1 _11278_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(_3916_),
    .Y(_3917_)
);

NAND3X1 _11279_ (
    .A(_3488_),
    .B(_3912_),
    .C(_3915_),
    .Y(_3918_)
);

NAND2X1 _11280_ (
    .A(_3918_),
    .B(_3917_),
    .Y(_3919_)
);

AOI21X1 _11281_ (
    .A(_3880_),
    .B(_3881_),
    .C(_3491_),
    .Y(_3920_)
);

NOR2X1 _11282_ (
    .A(_3920_),
    .B(_3900_),
    .Y(_3921_)
);

OAI21X1 _11283_ (
    .A(_3883_),
    .B(_3866_),
    .C(_3921_),
    .Y(_3922_)
);

NAND2X1 _11284_ (
    .A(_3902_),
    .B(_3922_),
    .Y(_3923_)
);

NOR2X1 _11285_ (
    .A(_3919_),
    .B(_3923_),
    .Y(_3924_)
);

AND2X2 _11286_ (
    .A(_3917_),
    .B(_3918_),
    .Y(_3925_)
);

AND2X2 _11287_ (
    .A(_3879_),
    .B(_3882_),
    .Y(_3926_)
);

NAND3X1 _11288_ (
    .A(_3902_),
    .B(_3926_),
    .C(_3901_),
    .Y(_3927_)
);

AOI21X1 _11289_ (
    .A(_3920_),
    .B(_3902_),
    .C(_3900_),
    .Y(_3928_)
);

OAI21X1 _11290_ (
    .A(_3866_),
    .B(_3927_),
    .C(_3928_),
    .Y(_3929_)
);

NOR2X1 _11291_ (
    .A(_3925_),
    .B(_3929_),
    .Y(_3930_)
);

OAI21X1 _11292_ (
    .A(_3930_),
    .B(_3924_),
    .C(_3579_),
    .Y(_3931_)
);

NAND2X1 _11293_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .B(_3931_),
    .Y(_3932_)
);

OAI21X1 _11294_ (
    .A(_3907_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_3932_),
    .Y(_3371_)
);

INVX1 _11295_ (
    .A(\genblk1[4].u_ce.Xcalc [7]),
    .Y(_3933_)
);

INVX1 _11296_ (
    .A(_3917_),
    .Y(_3934_)
);

NAND2X1 _11297_ (
    .A(_3911_),
    .B(_3913_),
    .Y(_3935_)
);

NOR2X1 _11298_ (
    .A(_3486__bF$buf2),
    .B(_3763_),
    .Y(_3936_)
);

INVX1 _11299_ (
    .A(_3936_),
    .Y(_3937_)
);

OAI21X1 _11300_ (
    .A(1'h1),
    .B(_3850_),
    .C(_3937_),
    .Y(_3938_)
);

NAND3X1 _11301_ (
    .A(_3524__bF$buf4),
    .B(_3938_),
    .C(_3935_),
    .Y(_3939_)
);

INVX1 _11302_ (
    .A(_3938_),
    .Y(_3940_)
);

OAI21X1 _11303_ (
    .A(_3914_),
    .B(_3908_),
    .C(_3524__bF$buf3),
    .Y(_3941_)
);

NAND2X1 _11304_ (
    .A(_3940_),
    .B(_3941_),
    .Y(_3942_)
);

NAND3X1 _11305_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(_3939_),
    .C(_3942_),
    .Y(_3943_)
);

NAND3X1 _11306_ (
    .A(_3524__bF$buf2),
    .B(_3940_),
    .C(_3935_),
    .Y(_3944_)
);

NAND2X1 _11307_ (
    .A(_3938_),
    .B(_3941_),
    .Y(_3945_)
);

NAND3X1 _11308_ (
    .A(_3525_),
    .B(_3944_),
    .C(_3945_),
    .Y(_3946_)
);

NAND2X1 _11309_ (
    .A(_3943_),
    .B(_3946_),
    .Y(_3947_)
);

OAI21X1 _11310_ (
    .A(_3934_),
    .B(_3924_),
    .C(_3947_),
    .Y(_3948_)
);

NOR2X1 _11311_ (
    .A(_3934_),
    .B(_3924_),
    .Y(_3949_)
);

INVX1 _11312_ (
    .A(_3947_),
    .Y(_3950_)
);

AOI21X1 _11313_ (
    .A(_3949_),
    .B(_3950_),
    .C(_3507_),
    .Y(_3951_)
);

AOI22X1 _11314_ (
    .A(_3933_),
    .B(_3510__bF$buf3),
    .C(_3951_),
    .D(_3948_),
    .Y(_3372_)
);

OAI21X1 _11315_ (
    .A(_3917_),
    .B(_3947_),
    .C(_3943_),
    .Y(_3952_)
);

NOR2X1 _11316_ (
    .A(_3919_),
    .B(_3947_),
    .Y(_3953_)
);

AOI21X1 _11317_ (
    .A(_3953_),
    .B(_3929_),
    .C(_3952_),
    .Y(_3954_)
);

INVX1 _11318_ (
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3955_)
);

NAND3X1 _11319_ (
    .A(_3911_),
    .B(_3940_),
    .C(_3913_),
    .Y(_3956_)
);

INVX1 _11320_ (
    .A(_3870_),
    .Y(_3957_)
);

OAI21X1 _11321_ (
    .A(1'h1),
    .B(_3957_),
    .C(_3937_),
    .Y(_3958_)
);

INVX1 _11322_ (
    .A(_3958_),
    .Y(_3959_)
);

NAND3X1 _11323_ (
    .A(_3524__bF$buf1),
    .B(_3959_),
    .C(_3956_),
    .Y(_3960_)
);

OAI21X1 _11324_ (
    .A(_3938_),
    .B(_3935_),
    .C(_3524__bF$buf0),
    .Y(_3961_)
);

NAND2X1 _11325_ (
    .A(_3958_),
    .B(_3961_),
    .Y(_3962_)
);

AOI21X1 _11326_ (
    .A(_3962_),
    .B(_3960_),
    .C(_3955_),
    .Y(_3963_)
);

NAND3X1 _11327_ (
    .A(_3524__bF$buf5),
    .B(_3958_),
    .C(_3956_),
    .Y(_3964_)
);

NAND2X1 _11328_ (
    .A(_3959_),
    .B(_3961_),
    .Y(_3965_)
);

AOI21X1 _11329_ (
    .A(_3965_),
    .B(_3964_),
    .C(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3966_)
);

OAI21X1 _11330_ (
    .A(_3963_),
    .B(_3966_),
    .C(_3954_),
    .Y(_3967_)
);

INVX1 _11331_ (
    .A(_3967_),
    .Y(_3968_)
);

OR2X2 _11332_ (
    .A(_3963_),
    .B(_3966_),
    .Y(_3969_)
);

OAI21X1 _11333_ (
    .A(_3969_),
    .B(_3954_),
    .C(_3508_),
    .Y(_3970_)
);

OAI22X1 _11334_ (
    .A(_3470_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_3970_),
    .D(_3968_),
    .Y(_3373_)
);

NAND2X1 _11335_ (
    .A(\genblk1[4].u_ce.Xcalc [9]),
    .B(_3510__bF$buf2),
    .Y(_3971_)
);

NOR2X1 _11336_ (
    .A(_3969_),
    .B(_3954_),
    .Y(_3972_)
);

NOR2X1 _11337_ (
    .A(_3963_),
    .B(_3972_),
    .Y(_3973_)
);

OAI21X1 _11338_ (
    .A(1'h1),
    .B(_3891_),
    .C(_3937_),
    .Y(_3974_)
);

INVX1 _11339_ (
    .A(_3974_),
    .Y(_3975_)
);

OAI21X1 _11340_ (
    .A(_3958_),
    .B(_3956_),
    .C(_3524__bF$buf4),
    .Y(_3976_)
);

NAND2X1 _11341_ (
    .A(_3975_),
    .B(_3976_),
    .Y(_3977_)
);

OR2X2 _11342_ (
    .A(_3976_),
    .B(_3975_),
    .Y(_3978_)
);

NAND3X1 _11343_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(_3977_),
    .C(_3978_),
    .Y(_3979_)
);

NAND2X1 _11344_ (
    .A(_3977_),
    .B(_3978_),
    .Y(_3980_)
);

NAND2X1 _11345_ (
    .A(_3587_),
    .B(_3980_),
    .Y(_3981_)
);

NAND2X1 _11346_ (
    .A(_3979_),
    .B(_3981_),
    .Y(_3982_)
);

AND2X2 _11347_ (
    .A(_3973_),
    .B(_3982_),
    .Y(_3983_)
);

OAI21X1 _11348_ (
    .A(_3982_),
    .B(_3973_),
    .C(_3508_),
    .Y(_3984_)
);

OAI21X1 _11349_ (
    .A(_3984_),
    .B(_3983_),
    .C(_3971_),
    .Y(_3374_)
);

INVX1 _11350_ (
    .A(\genblk1[4].u_ce.Xcalc [10]),
    .Y(_3985_)
);

INVX1 _11351_ (
    .A(_3979_),
    .Y(_3986_)
);

AOI21X1 _11352_ (
    .A(_3963_),
    .B(_3981_),
    .C(_3986_),
    .Y(_3987_)
);

NOR2X1 _11353_ (
    .A(_3963_),
    .B(_3966_),
    .Y(_3988_)
);

NAND3X1 _11354_ (
    .A(_3979_),
    .B(_3981_),
    .C(_3988_),
    .Y(_3989_)
);

OAI21X1 _11355_ (
    .A(_3954_),
    .B(_3989_),
    .C(_3987_),
    .Y(_3990_)
);

OAI21X1 _11356_ (
    .A(1'h1),
    .B(_3909_),
    .C(_3937_),
    .Y(_3991_)
);

INVX1 _11357_ (
    .A(_3991_),
    .Y(_3992_)
);

OR2X2 _11358_ (
    .A(_3956_),
    .B(_3958_),
    .Y(_3993_)
);

OAI21X1 _11359_ (
    .A(_3974_),
    .B(_3993_),
    .C(_3524__bF$buf3),
    .Y(_3994_)
);

NAND2X1 _11360_ (
    .A(_3992_),
    .B(_3994_),
    .Y(_3995_)
);

OR2X2 _11361_ (
    .A(_3994_),
    .B(_3992_),
    .Y(_3996_)
);

NAND3X1 _11362_ (
    .A(\genblk1[4].u_ce.Xin12b [10]),
    .B(_3995_),
    .C(_3996_),
    .Y(_3997_)
);

AND2X2 _11363_ (
    .A(_3994_),
    .B(_3992_),
    .Y(_3998_)
);

NOR2X1 _11364_ (
    .A(_3992_),
    .B(_3994_),
    .Y(_3999_)
);

OAI21X1 _11365_ (
    .A(_3999_),
    .B(_3998_),
    .C(_3608_),
    .Y(_4000_)
);

NAND2X1 _11366_ (
    .A(_4000_),
    .B(_3997_),
    .Y(_4001_)
);

AND2X2 _11367_ (
    .A(_3990_),
    .B(_4001_),
    .Y(_4002_)
);

NOR2X1 _11368_ (
    .A(_4001_),
    .B(_3990_),
    .Y(_4003_)
);

NOR2X1 _11369_ (
    .A(_4002_),
    .B(_4003_),
    .Y(_4004_)
);

AOI22X1 _11370_ (
    .A(_3985_),
    .B(_3510__bF$buf1),
    .C(_4004_),
    .D(_3508_),
    .Y(_3375_)
);

NAND2X1 _11371_ (
    .A(\genblk1[4].u_ce.Xcalc [11]),
    .B(_3510__bF$buf0),
    .Y(_4005_)
);

INVX1 _11372_ (
    .A(_3997_),
    .Y(_4006_)
);

AOI21X1 _11373_ (
    .A(_3990_),
    .B(_4000_),
    .C(_4006_),
    .Y(_4007_)
);

NAND2X1 _11374_ (
    .A(_3524__bF$buf2),
    .B(_3995_),
    .Y(_4008_)
);

NOR2X1 _11375_ (
    .A(_3765_),
    .B(_4008_),
    .Y(_4009_)
);

AOI21X1 _11376_ (
    .A(_3995_),
    .B(_3524__bF$buf1),
    .C(_3766_),
    .Y(_4010_)
);

NOR2X1 _11377_ (
    .A(_4010_),
    .B(_4009_),
    .Y(_4011_)
);

AND2X2 _11378_ (
    .A(_4007_),
    .B(_4011_),
    .Y(_4012_)
);

OAI21X1 _11379_ (
    .A(_4011_),
    .B(_4007_),
    .C(_3508_),
    .Y(_4013_)
);

OAI21X1 _11380_ (
    .A(_4013_),
    .B(_4012_),
    .C(_4005_),
    .Y(_3376_)
);

OAI21X1 _11381_ (
    .A(1'h0),
    .B(_3487__bF$buf0),
    .C(_3506_),
    .Y(_4014_)
);

OAI21X1 _11382_ (
    .A(_3781_),
    .B(_4014_),
    .C(\genblk1[4].u_ce.Ain0 [0]),
    .Y(_4015_)
);

INVX1 _11383_ (
    .A(\genblk1[4].u_ce.Ain0 [0]),
    .Y(_4016_)
);

NOR2X1 _11384_ (
    .A(_3781_),
    .B(_4014_),
    .Y(_4017_)
);

NAND2X1 _11385_ (
    .A(_4016_),
    .B(_4017_),
    .Y(_4018_)
);

NAND2X1 _11386_ (
    .A(_4015_),
    .B(_4018_),
    .Y(_4019_)
);

NAND2X1 _11387_ (
    .A(\genblk1[4].u_ce.Acalc [0]),
    .B(_3510__bF$buf4),
    .Y(_4020_)
);

OAI21X1 _11388_ (
    .A(_3510__bF$buf3),
    .B(_4019_),
    .C(_4020_),
    .Y(_3377_)
);

NAND2X1 _11389_ (
    .A(\genblk1[4].u_ce.Acalc [1]),
    .B(_3510__bF$buf2),
    .Y(_4021_)
);

INVX1 _11390_ (
    .A(_4015_),
    .Y(_4022_)
);

NOR2X1 _11391_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_4023_)
);

AOI21X1 _11392_ (
    .A(_3781_),
    .B(1'h1),
    .C(_4023_),
    .Y(_4024_)
);

NOR2X1 _11393_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4024_),
    .Y(_4025_)
);

OAI21X1 _11394_ (
    .A(_3781_),
    .B(_4014_),
    .C(_3524__bF$buf0),
    .Y(_4026_)
);

AND2X2 _11395_ (
    .A(_4026_),
    .B(_4024_),
    .Y(_4027_)
);

OR2X2 _11396_ (
    .A(_4027_),
    .B(_4025_),
    .Y(_4028_)
);

OR2X2 _11397_ (
    .A(_4028_),
    .B(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4029_)
);

OAI21X1 _11398_ (
    .A(_4025_),
    .B(_4027_),
    .C(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4030_)
);

NAND2X1 _11399_ (
    .A(_4030_),
    .B(_4029_),
    .Y(_4031_)
);

NOR2X1 _11400_ (
    .A(_4022_),
    .B(_4031_),
    .Y(_4032_)
);

NAND2X1 _11401_ (
    .A(_4022_),
    .B(_4031_),
    .Y(_4033_)
);

NAND2X1 _11402_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .B(_4033_),
    .Y(_4034_)
);

OAI21X1 _11403_ (
    .A(_4032_),
    .B(_4034_),
    .C(_4021_),
    .Y(_3378_)
);

INVX1 _11404_ (
    .A(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4035_)
);

OAI21X1 _11405_ (
    .A(_4035_),
    .B(_4028_),
    .C(_4033_),
    .Y(_4036_)
);

OAI21X1 _11406_ (
    .A(_3516_),
    .B(_3487__bF$buf4),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4037_)
);

OAI21X1 _11407_ (
    .A(1'h0),
    .B(1'h0),
    .C(1'h1),
    .Y(_4038_)
);

MUX2X1 _11408_ (
    .A(_4038_),
    .B(1'h1),
    .S(_4037_),
    .Y(_4039_)
);

NAND2X1 _11409_ (
    .A(\genblk1[4].u_ce.Ain1 [0]),
    .B(_4039_),
    .Y(_4040_)
);

OR2X2 _11410_ (
    .A(_4039_),
    .B(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_4041_)
);

NAND2X1 _11411_ (
    .A(_4040_),
    .B(_4041_),
    .Y(_4042_)
);

INVX1 _11412_ (
    .A(_4042_),
    .Y(_4043_)
);

NOR2X1 _11413_ (
    .A(_4043_),
    .B(_4036_),
    .Y(_4044_)
);

NAND2X1 _11414_ (
    .A(_4043_),
    .B(_4036_),
    .Y(_4045_)
);

NAND2X1 _11415_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4045_),
    .Y(_4046_)
);

OAI22X1 _11416_ (
    .A(_3432_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_4044_),
    .D(_4046_),
    .Y(_3379_)
);

NOR2X1 _11417_ (
    .A(\genblk1[4].u_ce.Acalc [3]),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_4047_)
);

NAND2X1 _11418_ (
    .A(_4040_),
    .B(_4045_),
    .Y(_4048_)
);

INVX1 _11419_ (
    .A(_4048_),
    .Y(_4049_)
);

INVX1 _11420_ (
    .A(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_4050_)
);

NOR2X1 _11421_ (
    .A(1'h0),
    .B(_3487__bF$buf3),
    .Y(_4051_)
);

OAI21X1 _11422_ (
    .A(_3486__bF$buf1),
    .B(_4051_),
    .C(_3524__bF$buf5),
    .Y(_4052_)
);

OAI21X1 _11423_ (
    .A(1'h1),
    .B(1'h0),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_4053_)
);

OAI21X1 _11424_ (
    .A(_3516_),
    .B(_4053_),
    .C(_4052_),
    .Y(_4054_)
);

NOR2X1 _11425_ (
    .A(_4050_),
    .B(_4054_),
    .Y(_4055_)
);

NAND2X1 _11426_ (
    .A(_4050_),
    .B(_4054_),
    .Y(_4056_)
);

INVX1 _11427_ (
    .A(_4056_),
    .Y(_4057_)
);

NOR2X1 _11428_ (
    .A(_4055_),
    .B(_4057_),
    .Y(_4058_)
);

OAI21X1 _11429_ (
    .A(_4058_),
    .B(_4049_),
    .C(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .Y(_4059_)
);

AOI21X1 _11430_ (
    .A(_4049_),
    .B(_4058_),
    .C(_4059_),
    .Y(_4060_)
);

NOR2X1 _11431_ (
    .A(_4047_),
    .B(_4060_),
    .Y(_3380_)
);

NAND2X1 _11432_ (
    .A(\genblk1[4].u_ce.Acalc [4]),
    .B(_3510__bF$buf1),
    .Y(_4061_)
);

INVX1 _11433_ (
    .A(\genblk1[4].u_ce.Ain12b [4]),
    .Y(_4062_)
);

AOI21X1 _11434_ (
    .A(_3781_),
    .B(1'h1),
    .C(_3524__bF$buf4),
    .Y(_4063_)
);

OAI21X1 _11435_ (
    .A(1'h1),
    .B(_3781_),
    .C(_4063_),
    .Y(_4064_)
);

OAI21X1 _11436_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4024_),
    .C(_4064_),
    .Y(_4065_)
);

OR2X2 _11437_ (
    .A(_4065_),
    .B(_4062_),
    .Y(_4066_)
);

NAND2X1 _11438_ (
    .A(_4062_),
    .B(_4065_),
    .Y(_4067_)
);

NAND2X1 _11439_ (
    .A(_4067_),
    .B(_4066_),
    .Y(_4068_)
);

AOI21X1 _11440_ (
    .A(_4048_),
    .B(_4056_),
    .C(_4055_),
    .Y(_4069_)
);

AND2X2 _11441_ (
    .A(_4069_),
    .B(_4068_),
    .Y(_4070_)
);

OAI21X1 _11442_ (
    .A(_4068_),
    .B(_4069_),
    .C(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Y(_4071_)
);

OAI21X1 _11443_ (
    .A(_4071_),
    .B(_4070_),
    .C(_4061_),
    .Y(_3381_)
);

OAI21X1 _11444_ (
    .A(_4068_),
    .B(_4069_),
    .C(_4066_),
    .Y(_4072_)
);

INVX1 _11445_ (
    .A(\genblk1[4].u_ce.Ain12b [5]),
    .Y(_4073_)
);

OAI21X1 _11446_ (
    .A(_3780_),
    .B(_3593_),
    .C(_3524__bF$buf3),
    .Y(_4074_)
);

OAI21X1 _11447_ (
    .A(1'h0),
    .B(1'h0),
    .C(_3506_),
    .Y(_4075_)
);

OR2X2 _11448_ (
    .A(_4075_),
    .B(_3524__bF$buf2),
    .Y(_4076_)
);

NAND2X1 _11449_ (
    .A(_4074_),
    .B(_4076_),
    .Y(_4077_)
);

OR2X2 _11450_ (
    .A(_4077_),
    .B(_4073_),
    .Y(_4078_)
);

NAND2X1 _11451_ (
    .A(_4073_),
    .B(_4077_),
    .Y(_4079_)
);

NAND2X1 _11452_ (
    .A(_4079_),
    .B(_4078_),
    .Y(_4080_)
);

INVX1 _11453_ (
    .A(_4080_),
    .Y(_4081_)
);

NOR2X1 _11454_ (
    .A(_4081_),
    .B(_4072_),
    .Y(_4082_)
);

NAND2X1 _11455_ (
    .A(_4081_),
    .B(_4072_),
    .Y(_4083_)
);

NAND2X1 _11456_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4083_),
    .Y(_4084_)
);

OAI22X1 _11457_ (
    .A(_3449_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_4082_),
    .D(_4084_),
    .Y(_3382_)
);

NAND2X1 _11458_ (
    .A(\genblk1[4].u_ce.Acalc [6]),
    .B(_3510__bF$buf0),
    .Y(_4085_)
);

INVX1 _11459_ (
    .A(_4068_),
    .Y(_4086_)
);

NAND2X1 _11460_ (
    .A(_4081_),
    .B(_4086_),
    .Y(_4087_)
);

OAI21X1 _11461_ (
    .A(_4066_),
    .B(_4080_),
    .C(_4078_),
    .Y(_4088_)
);

INVX1 _11462_ (
    .A(_4088_),
    .Y(_4089_)
);

OAI21X1 _11463_ (
    .A(_4087_),
    .B(_4069_),
    .C(_4089_),
    .Y(_4090_)
);

OAI21X1 _11464_ (
    .A(1'h0),
    .B(_3516_),
    .C(_3486__bF$buf0),
    .Y(_4091_)
);

NOR2X1 _11465_ (
    .A(_4091_),
    .B(_4051_),
    .Y(_4092_)
);

NAND2X1 _11466_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4092_),
    .Y(_4093_)
);

OAI21X1 _11467_ (
    .A(_4091_),
    .B(_4051_),
    .C(_3524__bF$buf1),
    .Y(_4094_)
);

NAND2X1 _11468_ (
    .A(_4094_),
    .B(_4093_),
    .Y(_4095_)
);

NAND2X1 _11469_ (
    .A(\genblk1[4].u_ce.Ain12b [6]),
    .B(_4095_),
    .Y(_4096_)
);

OR2X2 _11470_ (
    .A(_4095_),
    .B(\genblk1[4].u_ce.Ain12b [6]),
    .Y(_4097_)
);

NAND2X1 _11471_ (
    .A(_4096_),
    .B(_4097_),
    .Y(_4098_)
);

INVX1 _11472_ (
    .A(_4098_),
    .Y(_4099_)
);

NOR2X1 _11473_ (
    .A(_4099_),
    .B(_4090_),
    .Y(_4100_)
);

NAND2X1 _11474_ (
    .A(_4099_),
    .B(_4090_),
    .Y(_4101_)
);

NAND2X1 _11475_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .B(_4101_),
    .Y(_4102_)
);

OAI21X1 _11476_ (
    .A(_4100_),
    .B(_4102_),
    .C(_4085_),
    .Y(_3383_)
);

INVX1 _11477_ (
    .A(\genblk1[4].u_ce.Acalc [7]),
    .Y(_4103_)
);

NAND2X1 _11478_ (
    .A(_4096_),
    .B(_4101_),
    .Y(_4104_)
);

INVX1 _11479_ (
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .Y(_4105_)
);

NAND2X1 _11480_ (
    .A(_3524__bF$buf0),
    .B(_4023_),
    .Y(_4106_)
);

OR2X2 _11481_ (
    .A(_4023_),
    .B(_3524__bF$buf5),
    .Y(_4107_)
);

NAND2X1 _11482_ (
    .A(_4106_),
    .B(_4107_),
    .Y(_4108_)
);

NOR2X1 _11483_ (
    .A(_4105_),
    .B(_4108_),
    .Y(_4109_)
);

INVX1 _11484_ (
    .A(_4109_),
    .Y(_4110_)
);

NAND2X1 _11485_ (
    .A(_4105_),
    .B(_4108_),
    .Y(_4111_)
);

NAND2X1 _11486_ (
    .A(_4111_),
    .B(_4110_),
    .Y(_4112_)
);

OR2X2 _11487_ (
    .A(_4104_),
    .B(_4112_),
    .Y(_4113_)
);

AOI21X1 _11488_ (
    .A(_4104_),
    .B(_4112_),
    .C(_3510__bF$buf4),
    .Y(_4114_)
);

AOI22X1 _11489_ (
    .A(_4103_),
    .B(_3510__bF$buf3),
    .C(_4113_),
    .D(_4114_),
    .Y(_3384_)
);

NAND2X1 _11490_ (
    .A(\genblk1[4].u_ce.Acalc [8]),
    .B(_3510__bF$buf2),
    .Y(_4115_)
);

NOR2X1 _11491_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3506_),
    .Y(_4116_)
);

INVX1 _11492_ (
    .A(_4116_),
    .Y(_4117_)
);

NAND3X1 _11493_ (
    .A(\genblk1[4].u_ce.Ain12b [8]),
    .B(_4053_),
    .C(_4117_),
    .Y(_4118_)
);

INVX1 _11494_ (
    .A(_4118_),
    .Y(_4119_)
);

AOI21X1 _11495_ (
    .A(_4117_),
    .B(_4053_),
    .C(\genblk1[4].u_ce.Ain12b [8]),
    .Y(_4120_)
);

NOR2X1 _11496_ (
    .A(_4120_),
    .B(_4119_),
    .Y(_4121_)
);

OAI21X1 _11497_ (
    .A(_4096_),
    .B(_4112_),
    .C(_4110_),
    .Y(_4122_)
);

NOR2X1 _11498_ (
    .A(_4112_),
    .B(_4098_),
    .Y(_4123_)
);

AOI21X1 _11499_ (
    .A(_4123_),
    .B(_4088_),
    .C(_4122_),
    .Y(_4124_)
);

NAND3X1 _11500_ (
    .A(_4086_),
    .B(_4081_),
    .C(_4123_),
    .Y(_4125_)
);

OAI21X1 _11501_ (
    .A(_4125_),
    .B(_4069_),
    .C(_4124_),
    .Y(_4126_)
);

NOR2X1 _11502_ (
    .A(_4121_),
    .B(_4126_),
    .Y(_4127_)
);

NAND2X1 _11503_ (
    .A(_4121_),
    .B(_4126_),
    .Y(_4128_)
);

NAND2X1 _11504_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(_4128_),
    .Y(_4129_)
);

OAI21X1 _11505_ (
    .A(_4127_),
    .B(_4129_),
    .C(_4115_),
    .Y(_3385_)
);

AOI21X1 _11506_ (
    .A(_4126_),
    .B(_4121_),
    .C(_4119_),
    .Y(_4130_)
);

OR2X2 _11507_ (
    .A(_3524__bF$buf4),
    .B(\genblk1[4].u_ce.Ain12b [9]),
    .Y(_4131_)
);

NAND2X1 _11508_ (
    .A(\genblk1[4].u_ce.Ain12b [9]),
    .B(_3524__bF$buf3),
    .Y(_4132_)
);

NAND2X1 _11509_ (
    .A(_4132_),
    .B(_4131_),
    .Y(_4133_)
);

AND2X2 _11510_ (
    .A(_4130_),
    .B(_4133_),
    .Y(_4134_)
);

OAI21X1 _11511_ (
    .A(_4133_),
    .B(_4130_),
    .C(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Y(_4135_)
);

OAI22X1 _11512_ (
    .A(_3446_),
    .B(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .C(_4135_),
    .D(_4134_),
    .Y(_3386_)
);

NAND2X1 _11513_ (
    .A(\genblk1[4].u_ce.Acalc [10]),
    .B(_3510__bF$buf1),
    .Y(_4136_)
);

OAI21X1 _11514_ (
    .A(_4133_),
    .B(_4118_),
    .C(_4132_),
    .Y(_4137_)
);

NAND3X1 _11515_ (
    .A(_4131_),
    .B(_4132_),
    .C(_4121_),
    .Y(_4138_)
);

INVX1 _11516_ (
    .A(_4138_),
    .Y(_4139_)
);

AOI21X1 _11517_ (
    .A(_4126_),
    .B(_4139_),
    .C(_4137_),
    .Y(_4140_)
);

INVX1 _11518_ (
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .Y(_4141_)
);

NAND2X1 _11519_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4141_),
    .Y(_4142_)
);

NAND2X1 _11520_ (
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .B(_3524__bF$buf2),
    .Y(_4143_)
);

NAND2X1 _11521_ (
    .A(_4142_),
    .B(_4143_),
    .Y(_4144_)
);

AND2X2 _11522_ (
    .A(_4140_),
    .B(_4144_),
    .Y(_4145_)
);

OAI21X1 _11523_ (
    .A(_4144_),
    .B(_4140_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_4146_)
);

OAI21X1 _11524_ (
    .A(_4146_),
    .B(_4145_),
    .C(_4136_),
    .Y(_3387_)
);

NAND2X1 _11525_ (
    .A(\genblk1[4].u_ce.Acalc [11]),
    .B(_3510__bF$buf0),
    .Y(_4147_)
);

OAI21X1 _11526_ (
    .A(_4144_),
    .B(_4140_),
    .C(_4143_),
    .Y(_4148_)
);

OAI21X1 _11527_ (
    .A(_3510__bF$buf4),
    .B(_4148_),
    .C(_4147_),
    .Y(_3388_)
);

NAND2X1 _11528_ (
    .A(\genblk1[4].u_ce.LoadCtl [5]),
    .B(_3437_),
    .Y(_4149_)
);

NAND2X1 _11529_ (
    .A(_3438_),
    .B(_3444_),
    .Y(_4150_)
);

NOR2X1 _11530_ (
    .A(_4149_),
    .B(_4150_),
    .Y(_4151_)
);

NAND2X1 _11531_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4151_),
    .Y(_4152_)
);

OAI21X1 _11532_ (
    .A(_3608_),
    .B(_4151_),
    .C(_4152_),
    .Y(_3389_)
);

NAND2X1 _11533_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4151_),
    .Y(_4153_)
);

OAI21X1 _11534_ (
    .A(_3676_),
    .B(_4151_),
    .C(_4153_),
    .Y(_3390_)
);

INVX1 _11535_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .Y(_4154_)
);

OR2X2 _11536_ (
    .A(_4150_),
    .B(_3437_),
    .Y(_4155_)
);

OAI21X1 _11537_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_4156_)
);

OAI21X1 _11538_ (
    .A(_4154_),
    .B(_4155_),
    .C(_4156_),
    .Y(_3391_)
);

INVX1 _11539_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .Y(_4157_)
);

OAI21X1 _11540_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Xin12b [9]),
    .Y(_4158_)
);

OAI21X1 _11541_ (
    .A(_4157_),
    .B(_4155_),
    .C(_4158_),
    .Y(_3392_)
);

NAND2X1 _11542_ (
    .A(_3444_),
    .B(_3441_),
    .Y(_4159_)
);

NAND2X1 _11543_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(_4159_),
    .Y(_4160_)
);

OAI21X1 _11544_ (
    .A(_4154_),
    .B(_4159_),
    .C(_4160_),
    .Y(_3393_)
);

NAND2X1 _11545_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(_4159_),
    .Y(_4161_)
);

OAI21X1 _11546_ (
    .A(_4157_),
    .B(_4159_),
    .C(_4161_),
    .Y(_3394_)
);

AND2X2 _11547_ (
    .A(_3444_),
    .B(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_4162_)
);

NAND2X1 _11548_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4162_),
    .Y(_4163_)
);

OAI21X1 _11549_ (
    .A(_3491_),
    .B(_4162_),
    .C(_4163_),
    .Y(_3395_)
);

NAND2X1 _11550_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4162_),
    .Y(_4164_)
);

OAI21X1 _11551_ (
    .A(_3528_),
    .B(_4162_),
    .C(_4164_),
    .Y(_3396_)
);

OAI21X1 _11552_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_4165_)
);

OAI21X1 _11553_ (
    .A(_4154_),
    .B(_3435_),
    .C(_4165_),
    .Y(_3397_)
);

OAI21X1 _11554_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_4166_)
);

OAI21X1 _11555_ (
    .A(_4157_),
    .B(_3435_),
    .C(_4166_),
    .Y(_3398_)
);

NAND2X1 _11556_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.X_ [0]),
    .Y(_4167_)
);

OAI21X1 _11557_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3498_),
    .C(_4167_),
    .Y(_3399_)
);

NAND2X1 _11558_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.X_ [1]),
    .Y(_4168_)
);

OAI21X1 _11559_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3535_),
    .C(_4168_),
    .Y(_3400_)
);

NAND2X1 _11560_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4151_),
    .Y(_4169_)
);

OAI21X1 _11561_ (
    .A(_3737_),
    .B(_4151_),
    .C(_4169_),
    .Y(_3401_)
);

NAND2X1 _11562_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4151_),
    .Y(_4170_)
);

OAI21X1 _11563_ (
    .A(_3763_),
    .B(_4151_),
    .C(_4170_),
    .Y(_3402_)
);

INVX1 _11564_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .Y(_4171_)
);

OAI21X1 _11565_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_4172_)
);

OAI21X1 _11566_ (
    .A(_4171_),
    .B(_4155_),
    .C(_4172_),
    .Y(_3403_)
);

INVX1 _11567_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .Y(_4173_)
);

OAI21X1 _11568_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_4174_)
);

OAI21X1 _11569_ (
    .A(_4173_),
    .B(_4155_),
    .C(_4174_),
    .Y(_3404_)
);

NAND2X1 _11570_ (
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .B(_4159_),
    .Y(_4175_)
);

OAI21X1 _11571_ (
    .A(_4171_),
    .B(_4159_),
    .C(_4175_),
    .Y(_3405_)
);

NAND2X1 _11572_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(_4159_),
    .Y(_4176_)
);

OAI21X1 _11573_ (
    .A(_4173_),
    .B(_4159_),
    .C(_4176_),
    .Y(_3406_)
);

NAND2X1 _11574_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4162_),
    .Y(_4177_)
);

OAI21X1 _11575_ (
    .A(_3607_),
    .B(_4162_),
    .C(_4177_),
    .Y(_3407_)
);

NAND2X1 _11576_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4162_),
    .Y(_4178_)
);

OAI21X1 _11577_ (
    .A(_3628_),
    .B(_4162_),
    .C(_4178_),
    .Y(_3408_)
);

OAI21X1 _11578_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_4179_)
);

OAI21X1 _11579_ (
    .A(_4171_),
    .B(_3435_),
    .C(_4179_),
    .Y(_3409_)
);

OAI21X1 _11580_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_4180_)
);

OAI21X1 _11581_ (
    .A(_4173_),
    .B(_3435_),
    .C(_4180_),
    .Y(_3410_)
);

NAND2X1 _11582_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.Y_ [0]),
    .Y(_4181_)
);

OAI21X1 _11583_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3485_),
    .C(_4181_),
    .Y(_3411_)
);

NAND2X1 _11584_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.Y_ [1]),
    .Y(_4182_)
);

OAI21X1 _11585_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3523_),
    .C(_4182_),
    .Y(_3412_)
);

NAND2X1 _11586_ (
    .A(\a[4] [0]),
    .B(_4151_),
    .Y(_4183_)
);

OAI21X1 _11587_ (
    .A(_4141_),
    .B(_4151_),
    .C(_4183_),
    .Y(_3413_)
);

NAND2X1 _11588_ (
    .A(\a[4] [1]),
    .B(_4151_),
    .Y(_4184_)
);

OAI21X1 _11589_ (
    .A(_3524__bF$buf1),
    .B(_4151_),
    .C(_4184_),
    .Y(_3414_)
);

INVX1 _11590_ (
    .A(\a[4] [0]),
    .Y(_4185_)
);

OAI21X1 _11591_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Ain12b [8]),
    .Y(_4186_)
);

OAI21X1 _11592_ (
    .A(_4185_),
    .B(_4155_),
    .C(_4186_),
    .Y(_3415_)
);

INVX1 _11593_ (
    .A(\a[4] [1]),
    .Y(_4187_)
);

OAI21X1 _11594_ (
    .A(_3437_),
    .B(_4150_),
    .C(\genblk1[4].u_ce.Ain12b [9]),
    .Y(_4188_)
);

OAI21X1 _11595_ (
    .A(_4187_),
    .B(_4155_),
    .C(_4188_),
    .Y(_3416_)
);

NAND2X1 _11596_ (
    .A(\genblk1[4].u_ce.Ain12b [6]),
    .B(_4159_),
    .Y(_4189_)
);

OAI21X1 _11597_ (
    .A(_4185_),
    .B(_4159_),
    .C(_4189_),
    .Y(_3417_)
);

NAND2X1 _11598_ (
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .B(_4159_),
    .Y(_3425_)
);

OAI21X1 _11599_ (
    .A(_4187_),
    .B(_4159_),
    .C(_3425_),
    .Y(_3418_)
);

NAND2X1 _11600_ (
    .A(\a[4] [0]),
    .B(_4162_),
    .Y(_3426_)
);

OAI21X1 _11601_ (
    .A(_4062_),
    .B(_4162_),
    .C(_3426_),
    .Y(_3419_)
);

NAND2X1 _11602_ (
    .A(\a[4] [1]),
    .B(_4162_),
    .Y(_3427_)
);

OAI21X1 _11603_ (
    .A(_4073_),
    .B(_4162_),
    .C(_3427_),
    .Y(_3420_)
);

OAI21X1 _11604_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_3428_)
);

OAI21X1 _11605_ (
    .A(_4185_),
    .B(_3435_),
    .C(_3428_),
    .Y(_3421_)
);

OAI21X1 _11606_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3433_),
    .C(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_3429_)
);

OAI21X1 _11607_ (
    .A(_4187_),
    .B(_3435_),
    .C(_3429_),
    .Y(_3422_)
);

NAND2X1 _11608_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[4] [0]),
    .Y(_3430_)
);

OAI21X1 _11609_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4016_),
    .C(_3430_),
    .Y(_3423_)
);

NAND2X1 _11610_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[4] [1]),
    .Y(_3431_)
);

OAI21X1 _11611_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4035_),
    .C(_3431_),
    .Y(_3424_)
);

DFFPOSX1 _11612_ (
    .CLK(clk_bF$buf77),
    .D(_3352_),
    .Q(\genblk1[4].u_ce.Ycalc [0])
);

DFFPOSX1 _11613_ (
    .CLK(clk_bF$buf76),
    .D(_3353_),
    .Q(\genblk1[4].u_ce.Ycalc [1])
);

DFFPOSX1 _11614_ (
    .CLK(clk_bF$buf75),
    .D(_3354_),
    .Q(\genblk1[4].u_ce.ISout )
);

DFFPOSX1 _11615_ (
    .CLK(clk_bF$buf74),
    .D(_3355_),
    .Q(\genblk1[4].u_ce.Ycalc [2])
);

DFFPOSX1 _11616_ (
    .CLK(clk_bF$buf73),
    .D(_3356_),
    .Q(\genblk1[4].u_ce.Ycalc [3])
);

DFFPOSX1 _11617_ (
    .CLK(clk_bF$buf72),
    .D(_3357_),
    .Q(\genblk1[4].u_ce.Ycalc [4])
);

DFFPOSX1 _11618_ (
    .CLK(clk_bF$buf71),
    .D(_3358_),
    .Q(\genblk1[4].u_ce.Ycalc [5])
);

DFFPOSX1 _11619_ (
    .CLK(clk_bF$buf70),
    .D(_3359_),
    .Q(\genblk1[4].u_ce.Ycalc [6])
);

DFFPOSX1 _11620_ (
    .CLK(clk_bF$buf69),
    .D(_3360_),
    .Q(\genblk1[4].u_ce.Ycalc [7])
);

DFFPOSX1 _11621_ (
    .CLK(clk_bF$buf68),
    .D(_3361_),
    .Q(\genblk1[4].u_ce.Ycalc [8])
);

DFFPOSX1 _11622_ (
    .CLK(clk_bF$buf67),
    .D(_3362_),
    .Q(\genblk1[4].u_ce.Ycalc [9])
);

DFFPOSX1 _11623_ (
    .CLK(clk_bF$buf66),
    .D(_3363_),
    .Q(\genblk1[4].u_ce.Ycalc [10])
);

DFFPOSX1 _11624_ (
    .CLK(clk_bF$buf65),
    .D(_3364_),
    .Q(\genblk1[4].u_ce.Ycalc [11])
);

DFFPOSX1 _11625_ (
    .CLK(clk_bF$buf64),
    .D(_3365_),
    .Q(\genblk1[4].u_ce.Xcalc [0])
);

DFFPOSX1 _11626_ (
    .CLK(clk_bF$buf63),
    .D(_3366_),
    .Q(\genblk1[4].u_ce.Xcalc [1])
);

DFFPOSX1 _11627_ (
    .CLK(clk_bF$buf62),
    .D(_3367_),
    .Q(\genblk1[4].u_ce.Xcalc [2])
);

DFFPOSX1 _11628_ (
    .CLK(clk_bF$buf61),
    .D(_3368_),
    .Q(\genblk1[4].u_ce.Xcalc [3])
);

DFFPOSX1 _11629_ (
    .CLK(clk_bF$buf60),
    .D(_3369_),
    .Q(\genblk1[4].u_ce.Xcalc [4])
);

DFFPOSX1 _11630_ (
    .CLK(clk_bF$buf59),
    .D(_3370_),
    .Q(\genblk1[4].u_ce.Xcalc [5])
);

DFFPOSX1 _11631_ (
    .CLK(clk_bF$buf58),
    .D(_3371_),
    .Q(\genblk1[4].u_ce.Xcalc [6])
);

DFFPOSX1 _11632_ (
    .CLK(clk_bF$buf57),
    .D(_3372_),
    .Q(\genblk1[4].u_ce.Xcalc [7])
);

DFFPOSX1 _11633_ (
    .CLK(clk_bF$buf56),
    .D(_3373_),
    .Q(\genblk1[4].u_ce.Xcalc [8])
);

DFFPOSX1 _11634_ (
    .CLK(clk_bF$buf55),
    .D(_3374_),
    .Q(\genblk1[4].u_ce.Xcalc [9])
);

DFFPOSX1 _11635_ (
    .CLK(clk_bF$buf54),
    .D(_3375_),
    .Q(\genblk1[4].u_ce.Xcalc [10])
);

DFFPOSX1 _11636_ (
    .CLK(clk_bF$buf53),
    .D(_3376_),
    .Q(\genblk1[4].u_ce.Xcalc [11])
);

DFFPOSX1 _11637_ (
    .CLK(clk_bF$buf52),
    .D(_3377_),
    .Q(\genblk1[4].u_ce.Acalc [0])
);

DFFPOSX1 _11638_ (
    .CLK(clk_bF$buf51),
    .D(_3378_),
    .Q(\genblk1[4].u_ce.Acalc [1])
);

DFFPOSX1 _11639_ (
    .CLK(clk_bF$buf50),
    .D(_3379_),
    .Q(\genblk1[4].u_ce.Acalc [2])
);

DFFPOSX1 _11640_ (
    .CLK(clk_bF$buf49),
    .D(_3380_),
    .Q(\genblk1[4].u_ce.Acalc [3])
);

DFFPOSX1 _11641_ (
    .CLK(clk_bF$buf48),
    .D(_3381_),
    .Q(\genblk1[4].u_ce.Acalc [4])
);

DFFPOSX1 _11642_ (
    .CLK(clk_bF$buf47),
    .D(_3382_),
    .Q(\genblk1[4].u_ce.Acalc [5])
);

DFFPOSX1 _11643_ (
    .CLK(clk_bF$buf46),
    .D(_3383_),
    .Q(\genblk1[4].u_ce.Acalc [6])
);

DFFPOSX1 _11644_ (
    .CLK(clk_bF$buf45),
    .D(_3384_),
    .Q(\genblk1[4].u_ce.Acalc [7])
);

DFFPOSX1 _11645_ (
    .CLK(clk_bF$buf44),
    .D(_3385_),
    .Q(\genblk1[4].u_ce.Acalc [8])
);

DFFPOSX1 _11646_ (
    .CLK(clk_bF$buf43),
    .D(_3386_),
    .Q(\genblk1[4].u_ce.Acalc [9])
);

DFFPOSX1 _11647_ (
    .CLK(clk_bF$buf42),
    .D(_3387_),
    .Q(\genblk1[4].u_ce.Acalc [10])
);

DFFPOSX1 _11648_ (
    .CLK(clk_bF$buf41),
    .D(_3388_),
    .Q(\genblk1[4].u_ce.Acalc [11])
);

DFFPOSX1 _11649_ (
    .CLK(clk_bF$buf40),
    .D(_3389_),
    .Q(\genblk1[4].u_ce.Xin12b [10])
);

DFFPOSX1 _11650_ (
    .CLK(clk_bF$buf39),
    .D(_3390_),
    .Q(\genblk1[4].u_ce.Xin12b [11])
);

DFFPOSX1 _11651_ (
    .CLK(clk_bF$buf38),
    .D(_3391_),
    .Q(\genblk1[4].u_ce.Xin12b [8])
);

DFFPOSX1 _11652_ (
    .CLK(clk_bF$buf37),
    .D(_3392_),
    .Q(\genblk1[4].u_ce.Xin12b [9])
);

DFFPOSX1 _11653_ (
    .CLK(clk_bF$buf36),
    .D(_3393_),
    .Q(\genblk1[4].u_ce.Xin12b [6])
);

DFFPOSX1 _11654_ (
    .CLK(clk_bF$buf35),
    .D(_3394_),
    .Q(\genblk1[4].u_ce.Xin12b [7])
);

DFFPOSX1 _11655_ (
    .CLK(clk_bF$buf34),
    .D(_3395_),
    .Q(\genblk1[4].u_ce.Xin12b [4])
);

DFFPOSX1 _11656_ (
    .CLK(clk_bF$buf33),
    .D(_3396_),
    .Q(\genblk1[4].u_ce.Xin12b [5])
);

DFFPOSX1 _11657_ (
    .CLK(clk_bF$buf32),
    .D(_3397_),
    .Q(\genblk1[4].u_ce.Xin1 [0])
);

DFFPOSX1 _11658_ (
    .CLK(clk_bF$buf31),
    .D(_3398_),
    .Q(\genblk1[4].u_ce.Xin1 [1])
);

DFFPOSX1 _11659_ (
    .CLK(clk_bF$buf30),
    .D(_3399_),
    .Q(\genblk1[4].u_ce.Xin0 [0])
);

DFFPOSX1 _11660_ (
    .CLK(clk_bF$buf29),
    .D(_3400_),
    .Q(\genblk1[4].u_ce.Xin0 [1])
);

DFFPOSX1 _11661_ (
    .CLK(clk_bF$buf28),
    .D(_3401_),
    .Q(\genblk1[4].u_ce.Yin12b [10])
);

DFFPOSX1 _11662_ (
    .CLK(clk_bF$buf27),
    .D(_3402_),
    .Q(\genblk1[4].u_ce.Yin12b [11])
);

DFFPOSX1 _11663_ (
    .CLK(clk_bF$buf26),
    .D(_3403_),
    .Q(\genblk1[4].u_ce.Yin12b [8])
);

DFFPOSX1 _11664_ (
    .CLK(clk_bF$buf25),
    .D(_3404_),
    .Q(\genblk1[4].u_ce.Yin12b [9])
);

DFFPOSX1 _11665_ (
    .CLK(clk_bF$buf24),
    .D(_3405_),
    .Q(\genblk1[4].u_ce.Yin12b [6])
);

DFFPOSX1 _11666_ (
    .CLK(clk_bF$buf23),
    .D(_3406_),
    .Q(\genblk1[4].u_ce.Yin12b [7])
);

DFFPOSX1 _11667_ (
    .CLK(clk_bF$buf22),
    .D(_3407_),
    .Q(\genblk1[4].u_ce.Yin12b [4])
);

DFFPOSX1 _11668_ (
    .CLK(clk_bF$buf21),
    .D(_3408_),
    .Q(\genblk1[4].u_ce.Yin12b [5])
);

DFFPOSX1 _11669_ (
    .CLK(clk_bF$buf20),
    .D(_3409_),
    .Q(\genblk1[4].u_ce.Yin1 [0])
);

DFFPOSX1 _11670_ (
    .CLK(clk_bF$buf19),
    .D(_3410_),
    .Q(\genblk1[4].u_ce.Yin1 [1])
);

DFFPOSX1 _11671_ (
    .CLK(clk_bF$buf18),
    .D(_3411_),
    .Q(\genblk1[4].u_ce.Yin0 [0])
);

DFFPOSX1 _11672_ (
    .CLK(clk_bF$buf17),
    .D(_3412_),
    .Q(\genblk1[4].u_ce.Yin0 [1])
);

DFFPOSX1 _11673_ (
    .CLK(clk_bF$buf16),
    .D(_3413_),
    .Q(\genblk1[4].u_ce.Ain12b [10])
);

DFFPOSX1 _11674_ (
    .CLK(clk_bF$buf15),
    .D(_3414_),
    .Q(\genblk1[4].u_ce.Ain12b [11])
);

DFFPOSX1 _11675_ (
    .CLK(clk_bF$buf14),
    .D(_3415_),
    .Q(\genblk1[4].u_ce.Ain12b [8])
);

DFFPOSX1 _11676_ (
    .CLK(clk_bF$buf13),
    .D(_3416_),
    .Q(\genblk1[4].u_ce.Ain12b [9])
);

DFFPOSX1 _11677_ (
    .CLK(clk_bF$buf12),
    .D(_3417_),
    .Q(\genblk1[4].u_ce.Ain12b [6])
);

DFFPOSX1 _11678_ (
    .CLK(clk_bF$buf11),
    .D(_3418_),
    .Q(\genblk1[4].u_ce.Ain12b [7])
);

DFFPOSX1 _11679_ (
    .CLK(clk_bF$buf10),
    .D(_3419_),
    .Q(\genblk1[4].u_ce.Ain12b [4])
);

DFFPOSX1 _11680_ (
    .CLK(clk_bF$buf9),
    .D(_3420_),
    .Q(\genblk1[4].u_ce.Ain12b [5])
);

DFFPOSX1 _11681_ (
    .CLK(clk_bF$buf8),
    .D(_3421_),
    .Q(\genblk1[4].u_ce.Ain1 [0])
);

DFFPOSX1 _11682_ (
    .CLK(clk_bF$buf7),
    .D(_3422_),
    .Q(\genblk1[4].u_ce.Ain1 [1])
);

DFFPOSX1 _11683_ (
    .CLK(clk_bF$buf6),
    .D(_3423_),
    .Q(\genblk1[4].u_ce.Ain0 [0])
);

DFFPOSX1 _11684_ (
    .CLK(clk_bF$buf5),
    .D(_3424_),
    .Q(\genblk1[4].u_ce.Ain0 [1])
);

DFFPOSX1 _11685_ (
    .CLK(clk_bF$buf4),
    .D(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[4].u_ce.LoadCtl [0])
);

DFFPOSX1 _11686_ (
    .CLK(clk_bF$buf3),
    .D(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[4].u_ce.LoadCtl [1])
);

DFFPOSX1 _11687_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[4].u_ce.LoadCtl [1]),
    .Q(\genblk1[4].u_ce.LoadCtl [2])
);

DFFPOSX1 _11688_ (
    .CLK(clk_bF$buf1),
    .D(\genblk1[4].u_ce.LoadCtl [2]),
    .Q(\genblk1[4].u_ce.LoadCtl [3])
);

DFFPOSX1 _11689_ (
    .CLK(clk_bF$buf0),
    .D(\genblk1[4].u_ce.LoadCtl [3]),
    .Q(\genblk1[4].u_ce.LoadCtl [4])
);

DFFPOSX1 _11690_ (
    .CLK(clk_bF$buf78),
    .D(\genblk1[4].u_ce.LoadCtl [4]),
    .Q(\genblk1[4].u_ce.LoadCtl [5])
);

DFFPOSX1 _11691_ (
    .CLK(clk_bF$buf77),
    .D(\genblk1[4].u_ce.LoadCtl [5]),
    .Q(\genblk1[4].u_ce.Vld )
);

INVX1 _11692_ (
    .A(\genblk1[5].u_ce.Acalc [2]),
    .Y(_4270_)
);

INVX2 _11693_ (
    .A(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4271_)
);

NOR2X1 _11694_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4271_),
    .Y(_4272_)
);

INVX2 _11695_ (
    .A(_4272_),
    .Y(_4273_)
);

NOR2X1 _11696_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Acalc [10]),
    .Y(_4274_)
);

INVX4 _11697_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .Y(_4275_)
);

NOR2X1 _11698_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.LoadCtl [3]),
    .Y(_4276_)
);

OAI21X1 _11699_ (
    .A(_4275_),
    .B(\genblk1[5].u_ce.Acalc [8]),
    .C(_4276_),
    .Y(_4277_)
);

INVX2 _11700_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_4278_)
);

AND2X2 _11701_ (
    .A(_4278_),
    .B(\genblk1[5].u_ce.LoadCtl [3]),
    .Y(_4279_)
);

AOI22X1 _11702_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.Acalc [4]),
    .C(_4279_),
    .D(\genblk1[5].u_ce.Acalc [6]),
    .Y(_4280_)
);

OAI21X1 _11703_ (
    .A(_4274_),
    .B(_4277_),
    .C(_4280_),
    .Y(_4281_)
);

NOR2X1 _11704_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4282_)
);

AOI22X1 _11705_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Acalc [0]),
    .C(_4281_),
    .D(_4282_),
    .Y(_4283_)
);

OAI21X1 _11706_ (
    .A(_4270_),
    .B(_4273_),
    .C(_4283_),
    .Y(\a[6] [0])
);

INVX1 _11707_ (
    .A(\genblk1[5].u_ce.Acalc [9]),
    .Y(_4284_)
);

OAI21X1 _11708_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Acalc [11]),
    .C(_4276_),
    .Y(_4285_)
);

AOI21X1 _11709_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4284_),
    .C(_4285_),
    .Y(_4286_)
);

INVX1 _11710_ (
    .A(\genblk1[5].u_ce.Acalc [5]),
    .Y(_4287_)
);

NAND2X1 _11711_ (
    .A(\genblk1[5].u_ce.Acalc [7]),
    .B(_4279_),
    .Y(_4288_)
);

OAI21X1 _11712_ (
    .A(_4278_),
    .B(_4287_),
    .C(_4288_),
    .Y(_4289_)
);

OAI21X1 _11713_ (
    .A(_4286_),
    .B(_4289_),
    .C(_4282_),
    .Y(_4290_)
);

AOI22X1 _11714_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[5].u_ce.Acalc [1]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Acalc [3]),
    .Y(_4291_)
);

NAND2X1 _11715_ (
    .A(_4291_),
    .B(_4290_),
    .Y(\a[6] [1])
);

INVX1 _11716_ (
    .A(\genblk1[5].u_ce.Ycalc [10]),
    .Y(_4292_)
);

OAI21X1 _11717_ (
    .A(_4275_),
    .B(\genblk1[5].u_ce.Ycalc [8]),
    .C(_4276_),
    .Y(_4293_)
);

AOI21X1 _11718_ (
    .A(_4275_),
    .B(_4292_),
    .C(_4293_),
    .Y(_4294_)
);

INVX1 _11719_ (
    .A(\genblk1[5].u_ce.Ycalc [4]),
    .Y(_4295_)
);

NAND2X1 _11720_ (
    .A(\genblk1[5].u_ce.Ycalc [6]),
    .B(_4279_),
    .Y(_4296_)
);

OAI21X1 _11721_ (
    .A(_4278_),
    .B(_4295_),
    .C(_4296_),
    .Y(_4297_)
);

OAI21X1 _11722_ (
    .A(_4294_),
    .B(_4297_),
    .C(_4282_),
    .Y(_4298_)
);

AOI22X1 _11723_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.Ycalc [0]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Ycalc [2]),
    .Y(_4299_)
);

NAND2X1 _11724_ (
    .A(_4299_),
    .B(_4298_),
    .Y(\genblk1[5].u_ce.Y_ [0])
);

INVX1 _11725_ (
    .A(\genblk1[5].u_ce.Ycalc [9]),
    .Y(_4300_)
);

OAI21X1 _11726_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Ycalc [11]),
    .C(_4276_),
    .Y(_4301_)
);

AOI21X1 _11727_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4300_),
    .C(_4301_),
    .Y(_4302_)
);

INVX1 _11728_ (
    .A(\genblk1[5].u_ce.Ycalc [5]),
    .Y(_4303_)
);

NAND2X1 _11729_ (
    .A(\genblk1[5].u_ce.Ycalc [7]),
    .B(_4279_),
    .Y(_4304_)
);

OAI21X1 _11730_ (
    .A(_4278_),
    .B(_4303_),
    .C(_4304_),
    .Y(_4305_)
);

OAI21X1 _11731_ (
    .A(_4302_),
    .B(_4305_),
    .C(_4282_),
    .Y(_4306_)
);

AOI22X1 _11732_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.Ycalc [1]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4307_)
);

NAND2X1 _11733_ (
    .A(_4307_),
    .B(_4306_),
    .Y(\genblk1[5].u_ce.Y_ [1])
);

INVX1 _11734_ (
    .A(\genblk1[5].u_ce.Xcalc [8]),
    .Y(_4308_)
);

OAI21X1 _11735_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Xcalc [10]),
    .C(_4276_),
    .Y(_4309_)
);

AOI21X1 _11736_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4308_),
    .C(_4309_),
    .Y(_4310_)
);

INVX1 _11737_ (
    .A(\genblk1[5].u_ce.Xcalc [4]),
    .Y(_4311_)
);

NAND2X1 _11738_ (
    .A(\genblk1[5].u_ce.Xcalc [6]),
    .B(_4279_),
    .Y(_4312_)
);

OAI21X1 _11739_ (
    .A(_4278_),
    .B(_4311_),
    .C(_4312_),
    .Y(_4313_)
);

OAI21X1 _11740_ (
    .A(_4310_),
    .B(_4313_),
    .C(_4282_),
    .Y(_4314_)
);

AOI22X1 _11741_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Xcalc [0]),
    .C(_4272_),
    .D(\genblk1[5].u_ce.Xcalc [2]),
    .Y(_4315_)
);

NAND2X1 _11742_ (
    .A(_4315_),
    .B(_4314_),
    .Y(\genblk1[5].u_ce.X_ [0])
);

INVX1 _11743_ (
    .A(\genblk1[5].u_ce.Xcalc [3]),
    .Y(_4316_)
);

NOR2X1 _11744_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Xcalc [11]),
    .Y(_4317_)
);

OAI21X1 _11745_ (
    .A(_4275_),
    .B(\genblk1[5].u_ce.Xcalc [9]),
    .C(_4276_),
    .Y(_4318_)
);

AOI22X1 _11746_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.Xcalc [5]),
    .C(_4279_),
    .D(\genblk1[5].u_ce.Xcalc [7]),
    .Y(_4319_)
);

OAI21X1 _11747_ (
    .A(_4317_),
    .B(_4318_),
    .C(_4319_),
    .Y(_4320_)
);

AOI22X1 _11748_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Xcalc [1]),
    .C(_4320_),
    .D(_4282_),
    .Y(_4321_)
);

OAI21X1 _11749_ (
    .A(_4316_),
    .B(_4273_),
    .C(_4321_),
    .Y(\genblk1[5].u_ce.X_ [1])
);

INVX1 _11750_ (
    .A(\genblk1[5].u_ce.Ycalc [0]),
    .Y(_4322_)
);

INVX1 _11751_ (
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .Y(_4323_)
);

INVX8 _11752_ (
    .A(1'h1),
    .Y(_4324_)
);

INVX8 _11753_ (
    .A(1'h0),
    .Y(_4325_)
);

INVX1 _11754_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_4326_)
);

NAND2X1 _11755_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4327_)
);

OAI21X1 _11756_ (
    .A(1'h1),
    .B(_4326_),
    .C(_4327_),
    .Y(_4328_)
);

INVX1 _11757_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .Y(_4329_)
);

NAND2X1 _11758_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4330_)
);

OAI21X1 _11759_ (
    .A(1'h1),
    .B(_4329_),
    .C(_4330_),
    .Y(_4331_)
);

MUX2X1 _11760_ (
    .A(_4331_),
    .B(_4328_),
    .S(_4325__bF$buf4),
    .Y(_4332_)
);

INVX1 _11761_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4333_)
);

NAND2X1 _11762_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4334_)
);

OAI21X1 _11763_ (
    .A(1'h1),
    .B(_4333_),
    .C(_4334_),
    .Y(_4335_)
);

INVX1 _11764_ (
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .Y(_4336_)
);

NAND2X1 _11765_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_4337_)
);

OAI21X1 _11766_ (
    .A(1'h1),
    .B(_4336_),
    .C(_4337_),
    .Y(_4338_)
);

MUX2X1 _11767_ (
    .A(_4338_),
    .B(_4335_),
    .S(_4325__bF$buf3),
    .Y(_4339_)
);

MUX2X1 _11768_ (
    .A(_4339_),
    .B(_4332_),
    .S(_4324__bF$buf4),
    .Y(_4340_)
);

NOR2X1 _11769_ (
    .A(_4323_),
    .B(_4340_),
    .Y(_4341_)
);

NAND2X1 _11770_ (
    .A(_4323_),
    .B(_4340_),
    .Y(_4342_)
);

INVX1 _11771_ (
    .A(_4342_),
    .Y(_4343_)
);

NAND2X1 _11772_ (
    .A(_4324__bF$buf3),
    .B(_4325__bF$buf2),
    .Y(_4344_)
);

OAI21X1 _11773_ (
    .A(1'h1),
    .B(_4344_),
    .C(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .Y(_4345_)
);

INVX2 _11774_ (
    .A(_4345_),
    .Y(_4346_)
);

OAI21X1 _11775_ (
    .A(_4341_),
    .B(_4343_),
    .C(_4346_),
    .Y(_4347_)
);

OAI21X1 _11776_ (
    .A(_4322_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4347_),
    .Y(_4190_)
);

INVX8 _11777_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4348_)
);

NAND2X1 _11778_ (
    .A(\genblk1[5].u_ce.Ycalc [1]),
    .B(_4348__bF$buf4),
    .Y(_4349_)
);

NOR2X1 _11779_ (
    .A(1'h1),
    .B(_4344_),
    .Y(_4350_)
);

MUX2X1 _11780_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(\genblk1[5].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_4351_)
);

MUX2X1 _11781_ (
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .B(\genblk1[5].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_4352_)
);

MUX2X1 _11782_ (
    .A(_4352_),
    .B(_4351_),
    .S(_4325__bF$buf1),
    .Y(_4353_)
);

INVX2 _11783_ (
    .A(1'h1),
    .Y(_4354_)
);

NAND2X1 _11784_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(_4354_),
    .Y(_4355_)
);

AOI21X1 _11785_ (
    .A(_4355_),
    .B(_4334_),
    .C(_4325__bF$buf0),
    .Y(_4356_)
);

NAND3X1 _11786_ (
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .B(_4354_),
    .C(_4325__bF$buf4),
    .Y(_4357_)
);

NAND3X1 _11787_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(1'h1),
    .C(_4325__bF$buf3),
    .Y(_4358_)
);

NAND3X1 _11788_ (
    .A(_4324__bF$buf2),
    .B(_4358_),
    .C(_4357_),
    .Y(_4359_)
);

OAI22X1 _11789_ (
    .A(_4356_),
    .B(_4359_),
    .C(_4324__bF$buf1),
    .D(_4353_),
    .Y(_4360_)
);

INVX1 _11790_ (
    .A(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4361_)
);

INVX8 _11791_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_4362_)
);

INVX1 _11792_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4363_)
);

NAND2X1 _11793_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4364_)
);

OAI21X1 _11794_ (
    .A(1'h1),
    .B(_4363_),
    .C(_4364_),
    .Y(_4365_)
);

INVX1 _11795_ (
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4366_)
);

NAND2X1 _11796_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_4367_)
);

OAI21X1 _11797_ (
    .A(1'h1),
    .B(_4366_),
    .C(_4367_),
    .Y(_4368_)
);

MUX2X1 _11798_ (
    .A(_4368_),
    .B(_4365_),
    .S(_4325__bF$buf2),
    .Y(_4369_)
);

INVX1 _11799_ (
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4370_)
);

NAND2X1 _11800_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [4]),
    .Y(_4371_)
);

OAI21X1 _11801_ (
    .A(1'h1),
    .B(_4370_),
    .C(_4371_),
    .Y(_4372_)
);

INVX1 _11802_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .Y(_4373_)
);

NAND2X1 _11803_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4374_)
);

OAI21X1 _11804_ (
    .A(1'h1),
    .B(_4373_),
    .C(_4374_),
    .Y(_4375_)
);

MUX2X1 _11805_ (
    .A(_4375_),
    .B(_4372_),
    .S(_4325__bF$buf1),
    .Y(_4376_)
);

MUX2X1 _11806_ (
    .A(_4376_),
    .B(_4369_),
    .S(_4324__bF$buf0),
    .Y(_4377_)
);

NAND3X1 _11807_ (
    .A(_4362__bF$buf5),
    .B(_4340_),
    .C(_4377_),
    .Y(_4378_)
);

MUX2X1 _11808_ (
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_4379_)
);

MUX2X1 _11809_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_4380_)
);

MUX2X1 _11810_ (
    .A(_4380_),
    .B(_4379_),
    .S(_4325__bF$buf0),
    .Y(_4381_)
);

MUX2X1 _11811_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_4382_)
);

MUX2X1 _11812_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(\genblk1[5].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_4383_)
);

MUX2X1 _11813_ (
    .A(_4383_),
    .B(_4382_),
    .S(_4325__bF$buf4),
    .Y(_4384_)
);

MUX2X1 _11814_ (
    .A(_4384_),
    .B(_4381_),
    .S(_4324__bF$buf4),
    .Y(_4385_)
);

OAI21X1 _11815_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4360_),
    .C(_4385_),
    .Y(_4386_)
);

AOI21X1 _11816_ (
    .A(_4386_),
    .B(_4378_),
    .C(_4361_),
    .Y(_4387_)
);

INVX1 _11817_ (
    .A(_4387_),
    .Y(_4388_)
);

NAND3X1 _11818_ (
    .A(_4361_),
    .B(_4378_),
    .C(_4386_),
    .Y(_4389_)
);

AND2X2 _11819_ (
    .A(_4388_),
    .B(_4389_),
    .Y(_4390_)
);

OAI21X1 _11820_ (
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .B(_4360_),
    .C(_4390_),
    .Y(_4391_)
);

OR2X2 _11821_ (
    .A(_4390_),
    .B(_4342_),
    .Y(_4392_)
);

AOI21X1 _11822_ (
    .A(_4392_),
    .B(_4391_),
    .C(_4350_),
    .Y(_4393_)
);

OAI21X1 _11823_ (
    .A(_4348__bF$buf3),
    .B(_4393_),
    .C(_4349_),
    .Y(_4191_)
);

INVX1 _11824_ (
    .A(\genblk1[5].u_ce.ISout ),
    .Y(_4394_)
);

NAND2X1 _11825_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .B(\genblk1[4].u_ce.ISout ),
    .Y(_4395_)
);

OAI21X1 _11826_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .B(_4394_),
    .C(_4395_),
    .Y(_4192_)
);

NAND2X1 _11827_ (
    .A(\genblk1[5].u_ce.Ycalc [2]),
    .B(_4348__bF$buf2),
    .Y(_4396_)
);

AOI21X1 _11828_ (
    .A(_4342_),
    .B(_4389_),
    .C(_4387_),
    .Y(_4397_)
);

MUX2X1 _11829_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(\genblk1[5].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_4398_)
);

MUX2X1 _11830_ (
    .A(_4398_),
    .B(_4351_),
    .S(1'h0),
    .Y(_4399_)
);

MUX2X1 _11831_ (
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_4400_)
);

NAND2X1 _11832_ (
    .A(1'h0),
    .B(_4324__bF$buf3),
    .Y(_4401_)
);

OAI22X1 _11833_ (
    .A(_4401_),
    .B(_4352_),
    .C(_4400_),
    .D(_4344_),
    .Y(_4402_)
);

AOI21X1 _11834_ (
    .A(1'h1),
    .B(_4399_),
    .C(_4402_),
    .Y(_4403_)
);

AOI21X1 _11835_ (
    .A(_4385_),
    .B(_4360_),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4404_)
);

NAND2X1 _11836_ (
    .A(_4403_),
    .B(_4404_),
    .Y(_4405_)
);

INVX1 _11837_ (
    .A(_4403_),
    .Y(_4406_)
);

OAI21X1 _11838_ (
    .A(_4340_),
    .B(_4377_),
    .C(_4362__bF$buf4),
    .Y(_4407_)
);

NAND2X1 _11839_ (
    .A(_4406_),
    .B(_4407_),
    .Y(_4408_)
);

AOI21X1 _11840_ (
    .A(_4408_),
    .B(_4405_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4409_)
);

NAND3X1 _11841_ (
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .B(_4405_),
    .C(_4408_),
    .Y(_4410_)
);

INVX1 _11842_ (
    .A(_4410_),
    .Y(_4411_)
);

OR2X2 _11843_ (
    .A(_4411_),
    .B(_4409_),
    .Y(_4412_)
);

NOR2X1 _11844_ (
    .A(_4397_),
    .B(_4412_),
    .Y(_4413_)
);

INVX1 _11845_ (
    .A(_4413_),
    .Y(_4414_)
);

OAI21X1 _11846_ (
    .A(_4409_),
    .B(_4411_),
    .C(_4397_),
    .Y(_4415_)
);

AOI21X1 _11847_ (
    .A(_4414_),
    .B(_4415_),
    .C(_4350_),
    .Y(_4416_)
);

INVX2 _11848_ (
    .A(_4350_),
    .Y(_4417_)
);

OAI21X1 _11849_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4417_),
    .C(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .Y(_4418_)
);

OAI21X1 _11850_ (
    .A(_4418_),
    .B(_4416_),
    .C(_4396_),
    .Y(_4193_)
);

INVX1 _11851_ (
    .A(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4419_)
);

INVX2 _11852_ (
    .A(_4418_),
    .Y(_4420_)
);

OAI21X1 _11853_ (
    .A(_4409_),
    .B(_4397_),
    .C(_4410_),
    .Y(_4421_)
);

INVX1 _11854_ (
    .A(_4421_),
    .Y(_4422_)
);

INVX1 _11855_ (
    .A(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4423_)
);

NAND3X1 _11856_ (
    .A(_4360_),
    .B(_4385_),
    .C(_4403_),
    .Y(_4424_)
);

INVX1 _11857_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .Y(_4425_)
);

NAND2X1 _11858_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4426_)
);

OAI21X1 _11859_ (
    .A(1'h1),
    .B(_4425_),
    .C(_4426_),
    .Y(_4427_)
);

NAND2X1 _11860_ (
    .A(_4325__bF$buf3),
    .B(_4379_),
    .Y(_4428_)
);

OAI21X1 _11861_ (
    .A(_4325__bF$buf2),
    .B(_4427_),
    .C(_4428_),
    .Y(_4429_)
);

NOR2X1 _11862_ (
    .A(1'h1),
    .B(_4325__bF$buf1),
    .Y(_4430_)
);

NOR2X1 _11863_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_4431_)
);

AOI22X1 _11864_ (
    .A(_4372_),
    .B(_4431_),
    .C(_4430_),
    .D(_4368_),
    .Y(_4432_)
);

OAI21X1 _11865_ (
    .A(_4324__bF$buf2),
    .B(_4429_),
    .C(_4432_),
    .Y(_4433_)
);

NAND3X1 _11866_ (
    .A(_4362__bF$buf3),
    .B(_4433_),
    .C(_4424_),
    .Y(_4434_)
);

INVX1 _11867_ (
    .A(_4424_),
    .Y(_4435_)
);

INVX1 _11868_ (
    .A(_4433_),
    .Y(_4436_)
);

OAI21X1 _11869_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4435_),
    .C(_4436_),
    .Y(_4437_)
);

NAND3X1 _11870_ (
    .A(_4423_),
    .B(_4434_),
    .C(_4437_),
    .Y(_4438_)
);

AOI21X1 _11871_ (
    .A(_4437_),
    .B(_4434_),
    .C(_4423_),
    .Y(_4439_)
);

INVX1 _11872_ (
    .A(_4439_),
    .Y(_4440_)
);

NAND2X1 _11873_ (
    .A(_4438_),
    .B(_4440_),
    .Y(_4441_)
);

AOI21X1 _11874_ (
    .A(_4441_),
    .B(_4422_),
    .C(_4350_),
    .Y(_4442_)
);

OAI21X1 _11875_ (
    .A(_4422_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4443_)
);

AOI22X1 _11876_ (
    .A(_4419_),
    .B(_4348__bF$buf1),
    .C(_4443_),
    .D(_4420_),
    .Y(_4194_)
);

AOI21X1 _11877_ (
    .A(_4421_),
    .B(_4438_),
    .C(_4439_),
    .Y(_4444_)
);

INVX1 _11878_ (
    .A(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4445_)
);

INVX1 _11879_ (
    .A(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4446_)
);

NAND2X1 _11880_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4447_)
);

OAI21X1 _11881_ (
    .A(1'h1),
    .B(_4446_),
    .C(_4447_),
    .Y(_4448_)
);

NAND2X1 _11882_ (
    .A(_4325__bF$buf0),
    .B(_4398_),
    .Y(_4449_)
);

OAI21X1 _11883_ (
    .A(_4325__bF$buf4),
    .B(_4448_),
    .C(_4449_),
    .Y(_4450_)
);

NAND2X1 _11884_ (
    .A(_4324__bF$buf1),
    .B(_4353_),
    .Y(_4451_)
);

OAI21X1 _11885_ (
    .A(_4324__bF$buf0),
    .B(_4450_),
    .C(_4451_),
    .Y(_4452_)
);

INVX2 _11886_ (
    .A(_4452_),
    .Y(_4453_)
);

OAI21X1 _11887_ (
    .A(_4433_),
    .B(_4424_),
    .C(_4362__bF$buf2),
    .Y(_4454_)
);

OR2X2 _11888_ (
    .A(_4454_),
    .B(_4453_),
    .Y(_4455_)
);

NOR2X1 _11889_ (
    .A(_4433_),
    .B(_4424_),
    .Y(_4456_)
);

OAI21X1 _11890_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4456_),
    .C(_4453_),
    .Y(_4457_)
);

NAND3X1 _11891_ (
    .A(_4445_),
    .B(_4457_),
    .C(_4455_),
    .Y(_4458_)
);

NOR2X1 _11892_ (
    .A(_4453_),
    .B(_4454_),
    .Y(_4459_)
);

AND2X2 _11893_ (
    .A(_4454_),
    .B(_4453_),
    .Y(_4460_)
);

OAI21X1 _11894_ (
    .A(_4459_),
    .B(_4460_),
    .C(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4461_)
);

NAND2X1 _11895_ (
    .A(_4461_),
    .B(_4458_),
    .Y(_4462_)
);

AOI21X1 _11896_ (
    .A(_4444_),
    .B(_4462_),
    .C(_4350_),
    .Y(_4463_)
);

OAI21X1 _11897_ (
    .A(_4444_),
    .B(_4462_),
    .C(_4463_),
    .Y(_4464_)
);

AOI22X1 _11898_ (
    .A(_4295_),
    .B(_4348__bF$buf0),
    .C(_4464_),
    .D(_4420_),
    .Y(_4195_)
);

OAI21X1 _11899_ (
    .A(_4462_),
    .B(_4444_),
    .C(_4461_),
    .Y(_4465_)
);

INVX1 _11900_ (
    .A(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4466_)
);

NAND3X1 _11901_ (
    .A(_4436_),
    .B(_4453_),
    .C(_4435_),
    .Y(_4467_)
);

NAND2X1 _11902_ (
    .A(1'h0),
    .B(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4468_)
);

INVX1 _11903_ (
    .A(_4468_),
    .Y(_4469_)
);

AOI21X1 _11904_ (
    .A(_4427_),
    .B(_4325__bF$buf3),
    .C(_4469_),
    .Y(_4470_)
);

NAND2X1 _11905_ (
    .A(_4324__bF$buf4),
    .B(_4381_),
    .Y(_4471_)
);

OAI21X1 _11906_ (
    .A(_4324__bF$buf3),
    .B(_4470_),
    .C(_4471_),
    .Y(_4472_)
);

NAND3X1 _11907_ (
    .A(_4362__bF$buf1),
    .B(_4472_),
    .C(_4467_),
    .Y(_4473_)
);

NOR3X1 _11908_ (
    .A(_4433_),
    .B(_4452_),
    .C(_4424_),
    .Y(_4474_)
);

INVX1 _11909_ (
    .A(_4472_),
    .Y(_4475_)
);

OAI21X1 _11910_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4474_),
    .C(_4475_),
    .Y(_4476_)
);

NAND3X1 _11911_ (
    .A(_4466_),
    .B(_4473_),
    .C(_4476_),
    .Y(_4477_)
);

AOI21X1 _11912_ (
    .A(_4476_),
    .B(_4473_),
    .C(_4466_),
    .Y(_4478_)
);

INVX1 _11913_ (
    .A(_4478_),
    .Y(_4479_)
);

NAND2X1 _11914_ (
    .A(_4477_),
    .B(_4479_),
    .Y(_4480_)
);

AND2X2 _11915_ (
    .A(_4465_),
    .B(_4480_),
    .Y(_4481_)
);

OAI21X1 _11916_ (
    .A(_4480_),
    .B(_4465_),
    .C(_4417_),
    .Y(_4482_)
);

OAI21X1 _11917_ (
    .A(_4482_),
    .B(_4481_),
    .C(_4420_),
    .Y(_4483_)
);

OAI21X1 _11918_ (
    .A(_4303_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4483_),
    .Y(_4196_)
);

INVX1 _11919_ (
    .A(\genblk1[5].u_ce.Ycalc [6]),
    .Y(_4484_)
);

INVX1 _11920_ (
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4485_)
);

NAND3X1 _11921_ (
    .A(_4453_),
    .B(_4475_),
    .C(_4456_),
    .Y(_4486_)
);

AOI21X1 _11922_ (
    .A(_4448_),
    .B(_4325__bF$buf2),
    .C(_4469_),
    .Y(_4487_)
);

NAND2X1 _11923_ (
    .A(_4324__bF$buf2),
    .B(_4399_),
    .Y(_4488_)
);

OAI21X1 _11924_ (
    .A(_4324__bF$buf1),
    .B(_4487_),
    .C(_4488_),
    .Y(_4489_)
);

NAND3X1 _11925_ (
    .A(_4362__bF$buf0),
    .B(_4489_),
    .C(_4486_),
    .Y(_4490_)
);

INVX1 _11926_ (
    .A(_4489_),
    .Y(_4491_)
);

OAI21X1 _11927_ (
    .A(_4472_),
    .B(_4467_),
    .C(_4362__bF$buf5),
    .Y(_4492_)
);

NAND2X1 _11928_ (
    .A(_4491_),
    .B(_4492_),
    .Y(_4493_)
);

NAND3X1 _11929_ (
    .A(_4485_),
    .B(_4490_),
    .C(_4493_),
    .Y(_4494_)
);

NAND3X1 _11930_ (
    .A(_4362__bF$buf4),
    .B(_4491_),
    .C(_4486_),
    .Y(_4495_)
);

NAND2X1 _11931_ (
    .A(_4489_),
    .B(_4492_),
    .Y(_4496_)
);

NAND3X1 _11932_ (
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .B(_4495_),
    .C(_4496_),
    .Y(_4497_)
);

NAND2X1 _11933_ (
    .A(_4494_),
    .B(_4497_),
    .Y(_4498_)
);

AOI21X1 _11934_ (
    .A(_4455_),
    .B(_4457_),
    .C(_4445_),
    .Y(_4499_)
);

NOR2X1 _11935_ (
    .A(_4499_),
    .B(_4478_),
    .Y(_4500_)
);

OAI21X1 _11936_ (
    .A(_4462_),
    .B(_4444_),
    .C(_4500_),
    .Y(_4501_)
);

NAND2X1 _11937_ (
    .A(_4477_),
    .B(_4501_),
    .Y(_4502_)
);

AOI21X1 _11938_ (
    .A(_4502_),
    .B(_4498_),
    .C(_4350_),
    .Y(_4503_)
);

OAI21X1 _11939_ (
    .A(_4498_),
    .B(_4502_),
    .C(_4503_),
    .Y(_4504_)
);

AOI22X1 _11940_ (
    .A(_4484_),
    .B(_4348__bF$buf4),
    .C(_4504_),
    .D(_4420_),
    .Y(_4197_)
);

INVX1 _11941_ (
    .A(\genblk1[5].u_ce.Ycalc [7]),
    .Y(_4505_)
);

AOI21X1 _11942_ (
    .A(_4493_),
    .B(_4490_),
    .C(_4485_),
    .Y(_4506_)
);

AND2X2 _11943_ (
    .A(_4458_),
    .B(_4461_),
    .Y(_4507_)
);

NAND3X1 _11944_ (
    .A(_4477_),
    .B(_4479_),
    .C(_4507_),
    .Y(_4508_)
);

AOI21X1 _11945_ (
    .A(_4499_),
    .B(_4477_),
    .C(_4478_),
    .Y(_4509_)
);

OAI21X1 _11946_ (
    .A(_4444_),
    .B(_4508_),
    .C(_4509_),
    .Y(_4510_)
);

AOI21X1 _11947_ (
    .A(_4510_),
    .B(_4494_),
    .C(_4506_),
    .Y(_4511_)
);

INVX1 _11948_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4512_)
);

NAND3X1 _11949_ (
    .A(_4475_),
    .B(_4491_),
    .C(_4474_),
    .Y(_4513_)
);

INVX1 _11950_ (
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4514_)
);

NOR2X1 _11951_ (
    .A(_4324__bF$buf0),
    .B(_4514_),
    .Y(_4515_)
);

INVX1 _11952_ (
    .A(_4515_),
    .Y(_4516_)
);

OAI21X1 _11953_ (
    .A(1'h1),
    .B(_4429_),
    .C(_4516_),
    .Y(_4517_)
);

NAND3X1 _11954_ (
    .A(_4362__bF$buf3),
    .B(_4517_),
    .C(_4513_),
    .Y(_4518_)
);

INVX1 _11955_ (
    .A(_4517_),
    .Y(_4519_)
);

OAI21X1 _11956_ (
    .A(_4489_),
    .B(_4486_),
    .C(_4362__bF$buf2),
    .Y(_4520_)
);

NAND2X1 _11957_ (
    .A(_4519_),
    .B(_4520_),
    .Y(_4521_)
);

NAND3X1 _11958_ (
    .A(_4512_),
    .B(_4518_),
    .C(_4521_),
    .Y(_4522_)
);

NAND3X1 _11959_ (
    .A(_4362__bF$buf1),
    .B(_4519_),
    .C(_4513_),
    .Y(_4523_)
);

NAND2X1 _11960_ (
    .A(_4517_),
    .B(_4520_),
    .Y(_4524_)
);

NAND3X1 _11961_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(_4523_),
    .C(_4524_),
    .Y(_4525_)
);

NAND2X1 _11962_ (
    .A(_4522_),
    .B(_4525_),
    .Y(_4526_)
);

INVX1 _11963_ (
    .A(_4526_),
    .Y(_4527_)
);

NOR2X1 _11964_ (
    .A(_4527_),
    .B(_4511_),
    .Y(_4528_)
);

OAI21X1 _11965_ (
    .A(_4498_),
    .B(_4502_),
    .C(_4497_),
    .Y(_4529_)
);

OAI21X1 _11966_ (
    .A(_4526_),
    .B(_4529_),
    .C(_4417_),
    .Y(_4530_)
);

OAI21X1 _11967_ (
    .A(_4362__bF$buf0),
    .B(_4417_),
    .C(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4531_)
);

INVX1 _11968_ (
    .A(_4531_),
    .Y(_4532_)
);

OAI21X1 _11969_ (
    .A(_4530_),
    .B(_4528_),
    .C(_4532_),
    .Y(_4533_)
);

OAI21X1 _11970_ (
    .A(_4505_),
    .B(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .C(_4533_),
    .Y(_4198_)
);

INVX1 _11971_ (
    .A(\genblk1[5].u_ce.Ycalc [8]),
    .Y(_4534_)
);

OAI21X1 _11972_ (
    .A(_4497_),
    .B(_4526_),
    .C(_4525_),
    .Y(_4535_)
);

NOR2X1 _11973_ (
    .A(_4498_),
    .B(_4526_),
    .Y(_4536_)
);

AOI21X1 _11974_ (
    .A(_4536_),
    .B(_4510_),
    .C(_4535_),
    .Y(_4537_)
);

INVX1 _11975_ (
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4538_)
);

OR2X2 _11976_ (
    .A(_4513_),
    .B(_4517_),
    .Y(_4539_)
);

OAI21X1 _11977_ (
    .A(1'h1),
    .B(_4450_),
    .C(_4516_),
    .Y(_4540_)
);

NAND3X1 _11978_ (
    .A(_4362__bF$buf5),
    .B(_4540_),
    .C(_4539_),
    .Y(_4541_)
);

NOR2X1 _11979_ (
    .A(_4517_),
    .B(_4513_),
    .Y(_4542_)
);

INVX1 _11980_ (
    .A(_4540_),
    .Y(_4543_)
);

OAI21X1 _11981_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4542_),
    .C(_4543_),
    .Y(_4544_)
);

NAND3X1 _11982_ (
    .A(_4538_),
    .B(_4544_),
    .C(_4541_),
    .Y(_4545_)
);

NAND3X1 _11983_ (
    .A(_4362__bF$buf4),
    .B(_4543_),
    .C(_4539_),
    .Y(_4546_)
);

OAI21X1 _11984_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4542_),
    .C(_4540_),
    .Y(_4547_)
);

NAND3X1 _11985_ (
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .B(_4547_),
    .C(_4546_),
    .Y(_4548_)
);

AND2X2 _11986_ (
    .A(_4545_),
    .B(_4548_),
    .Y(_4549_)
);

INVX1 _11987_ (
    .A(_4549_),
    .Y(_4550_)
);

AOI21X1 _11988_ (
    .A(_4537_),
    .B(_4550_),
    .C(_4350_),
    .Y(_4551_)
);

OAI21X1 _11989_ (
    .A(_4537_),
    .B(_4550_),
    .C(_4551_),
    .Y(_4552_)
);

AOI22X1 _11990_ (
    .A(_4534_),
    .B(_4348__bF$buf3),
    .C(_4552_),
    .D(_4532_),
    .Y(_4199_)
);

NAND2X1 _11991_ (
    .A(_4506_),
    .B(_4522_),
    .Y(_4553_)
);

AND2X2 _11992_ (
    .A(_4553_),
    .B(_4525_),
    .Y(_4554_)
);

AND2X2 _11993_ (
    .A(_4494_),
    .B(_4497_),
    .Y(_4555_)
);

NAND3X1 _11994_ (
    .A(_4522_),
    .B(_4525_),
    .C(_4555_),
    .Y(_4556_)
);

OAI21X1 _11995_ (
    .A(_4502_),
    .B(_4556_),
    .C(_4554_),
    .Y(_4557_)
);

INVX1 _11996_ (
    .A(_4548_),
    .Y(_4558_)
);

AOI21X1 _11997_ (
    .A(_4557_),
    .B(_4545_),
    .C(_4558_),
    .Y(_4559_)
);

INVX1 _11998_ (
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_4560_)
);

NOR3X1 _11999_ (
    .A(_4517_),
    .B(_4540_),
    .C(_4513_),
    .Y(_4561_)
);

INVX1 _12000_ (
    .A(_4561_),
    .Y(_4562_)
);

OAI21X1 _12001_ (
    .A(1'h1),
    .B(_4470_),
    .C(_4516_),
    .Y(_4563_)
);

NAND3X1 _12002_ (
    .A(_4362__bF$buf3),
    .B(_4563_),
    .C(_4562_),
    .Y(_4564_)
);

INVX1 _12003_ (
    .A(_4563_),
    .Y(_4565_)
);

OAI21X1 _12004_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4561_),
    .C(_4565_),
    .Y(_4566_)
);

NAND3X1 _12005_ (
    .A(_4560_),
    .B(_4566_),
    .C(_4564_),
    .Y(_4567_)
);

NAND3X1 _12006_ (
    .A(_4362__bF$buf2),
    .B(_4565_),
    .C(_4562_),
    .Y(_4568_)
);

OAI21X1 _12007_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4561_),
    .C(_4563_),
    .Y(_4569_)
);

NAND3X1 _12008_ (
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .B(_4569_),
    .C(_4568_),
    .Y(_4570_)
);

AND2X2 _12009_ (
    .A(_4567_),
    .B(_4570_),
    .Y(_4571_)
);

AND2X2 _12010_ (
    .A(_4559_),
    .B(_4571_),
    .Y(_4572_)
);

OAI21X1 _12011_ (
    .A(_4571_),
    .B(_4559_),
    .C(_4417_),
    .Y(_4573_)
);

OAI21X1 _12012_ (
    .A(_4573_),
    .B(_4572_),
    .C(_4420_),
    .Y(_4574_)
);

OAI21X1 _12013_ (
    .A(_4300_),
    .B(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .C(_4574_),
    .Y(_4200_)
);

INVX1 _12014_ (
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .Y(_4575_)
);

OAI21X1 _12015_ (
    .A(1'h1),
    .B(_4487_),
    .C(_4516_),
    .Y(_4576_)
);

INVX1 _12016_ (
    .A(_4576_),
    .Y(_4577_)
);

AOI21X1 _12017_ (
    .A(_4561_),
    .B(_4565_),
    .C(_4577_),
    .Y(_4578_)
);

NAND3X1 _12018_ (
    .A(_4565_),
    .B(_4577_),
    .C(_4561_),
    .Y(_4579_)
);

NAND2X1 _12019_ (
    .A(_4362__bF$buf1),
    .B(_4579_),
    .Y(_4580_)
);

NAND2X1 _12020_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4576_),
    .Y(_4581_)
);

OAI21X1 _12021_ (
    .A(_4578_),
    .B(_4580_),
    .C(_4581_),
    .Y(_4582_)
);

NAND2X1 _12022_ (
    .A(_4575_),
    .B(_4582_),
    .Y(_4583_)
);

INVX1 _12023_ (
    .A(_4578_),
    .Y(_4584_)
);

AND2X2 _12024_ (
    .A(_4579_),
    .B(_4362__bF$buf0),
    .Y(_4585_)
);

NAND2X1 _12025_ (
    .A(_4584_),
    .B(_4585_),
    .Y(_4586_)
);

NAND3X1 _12026_ (
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .B(_4581_),
    .C(_4586_),
    .Y(_4587_)
);

NAND2X1 _12027_ (
    .A(_4583_),
    .B(_4587_),
    .Y(_4588_)
);

AOI21X1 _12028_ (
    .A(_4564_),
    .B(_4566_),
    .C(_4560_),
    .Y(_4589_)
);

AOI21X1 _12029_ (
    .A(_4558_),
    .B(_4567_),
    .C(_4589_),
    .Y(_4590_)
);

NAND3X1 _12030_ (
    .A(_4549_),
    .B(_4571_),
    .C(_4557_),
    .Y(_4591_)
);

AOI21X1 _12031_ (
    .A(_4591_),
    .B(_4590_),
    .C(_4588_),
    .Y(_4592_)
);

AND2X2 _12032_ (
    .A(_4587_),
    .B(_4583_),
    .Y(_4593_)
);

NAND3X1 _12033_ (
    .A(_4567_),
    .B(_4570_),
    .C(_4549_),
    .Y(_4594_)
);

OAI21X1 _12034_ (
    .A(_4594_),
    .B(_4537_),
    .C(_4590_),
    .Y(_4595_)
);

OAI21X1 _12035_ (
    .A(_4593_),
    .B(_4595_),
    .C(_4417_),
    .Y(_4596_)
);

OR2X2 _12036_ (
    .A(_4596_),
    .B(_4592_),
    .Y(_4597_)
);

AOI22X1 _12037_ (
    .A(_4292_),
    .B(_4348__bF$buf2),
    .C(_4597_),
    .D(_4420_),
    .Y(_4201_)
);

NAND2X1 _12038_ (
    .A(\genblk1[5].u_ce.Ycalc [11]),
    .B(_4348__bF$buf1),
    .Y(_4598_)
);

INVX1 _12039_ (
    .A(_4587_),
    .Y(_4599_)
);

NAND2X1 _12040_ (
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .B(_4514_),
    .Y(_4600_)
);

INVX1 _12041_ (
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4601_)
);

NAND2X1 _12042_ (
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .B(_4601_),
    .Y(_4602_)
);

NAND2X1 _12043_ (
    .A(_4600_),
    .B(_4602_),
    .Y(_4603_)
);

INVX1 _12044_ (
    .A(_4603_),
    .Y(_4604_)
);

NAND2X1 _12045_ (
    .A(_4604_),
    .B(_4580_),
    .Y(_4605_)
);

NAND2X1 _12046_ (
    .A(_4603_),
    .B(_4585_),
    .Y(_4606_)
);

NAND2X1 _12047_ (
    .A(_4605_),
    .B(_4606_),
    .Y(_4607_)
);

INVX1 _12048_ (
    .A(_4607_),
    .Y(_4608_)
);

NOR3X1 _12049_ (
    .A(_4599_),
    .B(_4608_),
    .C(_4592_),
    .Y(_4609_)
);

AOI21X1 _12050_ (
    .A(_4595_),
    .B(_4593_),
    .C(_4599_),
    .Y(_4610_)
);

OAI21X1 _12051_ (
    .A(_4607_),
    .B(_4610_),
    .C(_4417_),
    .Y(_4611_)
);

OAI21X1 _12052_ (
    .A(_4609_),
    .B(_4611_),
    .C(_4420_),
    .Y(_4612_)
);

NAND2X1 _12053_ (
    .A(_4598_),
    .B(_4612_),
    .Y(_4202_)
);

NAND2X1 _12054_ (
    .A(\genblk1[5].u_ce.Xcalc [0]),
    .B(_4348__bF$buf0),
    .Y(_4613_)
);

INVX1 _12055_ (
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4614_)
);

NAND2X1 _12056_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4615_)
);

OAI21X1 _12057_ (
    .A(1'h1),
    .B(_4614_),
    .C(_4615_),
    .Y(_4616_)
);

NAND2X1 _12058_ (
    .A(1'h0),
    .B(_4616_),
    .Y(_4617_)
);

NOR2X1 _12059_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_4618_)
);

NOR2X1 _12060_ (
    .A(1'h0),
    .B(_4354_),
    .Y(_4619_)
);

AOI22X1 _12061_ (
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .B(_4618_),
    .C(_4619_),
    .D(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4620_)
);

NAND3X1 _12062_ (
    .A(_4324__bF$buf4),
    .B(_4617_),
    .C(_4620_),
    .Y(_4621_)
);

NAND2X1 _12063_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4622_)
);

OAI21X1 _12064_ (
    .A(1'h1),
    .B(_4485_),
    .C(_4622_),
    .Y(_4623_)
);

NAND2X1 _12065_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4624_)
);

OAI21X1 _12066_ (
    .A(1'h1),
    .B(_4445_),
    .C(_4624_),
    .Y(_4625_)
);

MUX2X1 _12067_ (
    .A(_4625_),
    .B(_4623_),
    .S(_4325__bF$buf1),
    .Y(_4626_)
);

NAND2X1 _12068_ (
    .A(1'h1),
    .B(_4626_),
    .Y(_4627_)
);

AND2X2 _12069_ (
    .A(_4621_),
    .B(_4627_),
    .Y(_4628_)
);

NOR2X1 _12070_ (
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .B(_4628_),
    .Y(_4629_)
);

NAND2X1 _12071_ (
    .A(_4325__bF$buf0),
    .B(_4625_),
    .Y(_4630_)
);

NAND2X1 _12072_ (
    .A(1'h0),
    .B(_4623_),
    .Y(_4631_)
);

NAND2X1 _12073_ (
    .A(_4630_),
    .B(_4631_),
    .Y(_4632_)
);

OAI21X1 _12074_ (
    .A(_4324__bF$buf3),
    .B(_4632_),
    .C(_4621_),
    .Y(_4633_)
);

OAI21X1 _12075_ (
    .A(_4336_),
    .B(_4633_),
    .C(_4346_),
    .Y(_4634_)
);

OAI21X1 _12076_ (
    .A(_4634_),
    .B(_4629_),
    .C(_4613_),
    .Y(_4203_)
);

NAND2X1 _12077_ (
    .A(\genblk1[5].u_ce.Xcalc [1]),
    .B(_4348__bF$buf4),
    .Y(_4635_)
);

NOR2X1 _12078_ (
    .A(_4336_),
    .B(_4633_),
    .Y(_4636_)
);

NAND2X1 _12079_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4637_)
);

OAI21X1 _12080_ (
    .A(1'h1),
    .B(_4423_),
    .C(_4637_),
    .Y(_4638_)
);

NAND2X1 _12081_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4639_)
);

OAI21X1 _12082_ (
    .A(1'h1),
    .B(_4361_),
    .C(_4639_),
    .Y(_4640_)
);

MUX2X1 _12083_ (
    .A(_4640_),
    .B(_4638_),
    .S(_4325__bF$buf4),
    .Y(_4641_)
);

NAND2X1 _12084_ (
    .A(_4324__bF$buf2),
    .B(_4641_),
    .Y(_4642_)
);

NAND2X1 _12085_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4643_)
);

OAI21X1 _12086_ (
    .A(1'h1),
    .B(_4512_),
    .C(_4643_),
    .Y(_4644_)
);

INVX1 _12087_ (
    .A(_4644_),
    .Y(_4645_)
);

NAND2X1 _12088_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4646_)
);

OAI21X1 _12089_ (
    .A(1'h1),
    .B(_4466_),
    .C(_4646_),
    .Y(_4647_)
);

NAND2X1 _12090_ (
    .A(_4325__bF$buf3),
    .B(_4647_),
    .Y(_4648_)
);

OAI21X1 _12091_ (
    .A(_4325__bF$buf2),
    .B(_4645_),
    .C(_4648_),
    .Y(_4649_)
);

OAI21X1 _12092_ (
    .A(_4324__bF$buf1),
    .B(_4649_),
    .C(_4642_),
    .Y(_4650_)
);

NAND3X1 _12093_ (
    .A(_4362__bF$buf5),
    .B(_4650_),
    .C(_4628_),
    .Y(_4651_)
);

MUX2X1 _12094_ (
    .A(_4647_),
    .B(_4644_),
    .S(_4325__bF$buf1),
    .Y(_4652_)
);

MUX2X1 _12095_ (
    .A(_4652_),
    .B(_4641_),
    .S(1'h1),
    .Y(_4653_)
);

OAI21X1 _12096_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4633_),
    .C(_4653_),
    .Y(_4654_)
);

AOI21X1 _12097_ (
    .A(_4651_),
    .B(_4654_),
    .C(_4373_),
    .Y(_4655_)
);

INVX1 _12098_ (
    .A(_4655_),
    .Y(_4656_)
);

NAND3X1 _12099_ (
    .A(_4373_),
    .B(_4654_),
    .C(_4651_),
    .Y(_4657_)
);

AND2X2 _12100_ (
    .A(_4656_),
    .B(_4657_),
    .Y(_4658_)
);

NAND2X1 _12101_ (
    .A(_4636_),
    .B(_4658_),
    .Y(_4659_)
);

OR2X2 _12102_ (
    .A(_4658_),
    .B(_4636_),
    .Y(_4660_)
);

AOI21X1 _12103_ (
    .A(_4660_),
    .B(_4659_),
    .C(_4350_),
    .Y(_4661_)
);

OAI21X1 _12104_ (
    .A(_4348__bF$buf3),
    .B(_4661_),
    .C(_4635_),
    .Y(_4204_)
);

NAND2X1 _12105_ (
    .A(\genblk1[5].u_ce.Xcalc [2]),
    .B(_4348__bF$buf2),
    .Y(_4662_)
);

AOI21X1 _12106_ (
    .A(_4636_),
    .B(_4657_),
    .C(_4655_),
    .Y(_4663_)
);

NAND2X1 _12107_ (
    .A(_4633_),
    .B(_4650_),
    .Y(_4664_)
);

NAND2X1 _12108_ (
    .A(1'h1),
    .B(_4560_),
    .Y(_4665_)
);

OAI21X1 _12109_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .C(_4665_),
    .Y(_4666_)
);

NAND2X1 _12110_ (
    .A(_4325__bF$buf0),
    .B(_4623_),
    .Y(_4667_)
);

OAI21X1 _12111_ (
    .A(_4325__bF$buf4),
    .B(_4666_),
    .C(_4667_),
    .Y(_4668_)
);

NAND2X1 _12112_ (
    .A(_4431_),
    .B(_4616_),
    .Y(_4669_)
);

NAND2X1 _12113_ (
    .A(_4625_),
    .B(_4430_),
    .Y(_4670_)
);

NAND2X1 _12114_ (
    .A(_4669_),
    .B(_4670_),
    .Y(_4671_)
);

AOI21X1 _12115_ (
    .A(_4668_),
    .B(1'h1),
    .C(_4671_),
    .Y(_4672_)
);

INVX1 _12116_ (
    .A(_4672_),
    .Y(_4673_)
);

NAND3X1 _12117_ (
    .A(_4362__bF$buf4),
    .B(_4673_),
    .C(_4664_),
    .Y(_4674_)
);

AOI21X1 _12118_ (
    .A(_4621_),
    .B(_4627_),
    .C(_4653_),
    .Y(_4675_)
);

OAI21X1 _12119_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4675_),
    .C(_4672_),
    .Y(_4676_)
);

NAND3X1 _12120_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(_4676_),
    .C(_4674_),
    .Y(_4677_)
);

INVX1 _12121_ (
    .A(_4677_),
    .Y(_4678_)
);

AOI21X1 _12122_ (
    .A(_4674_),
    .B(_4676_),
    .C(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4679_)
);

NOR2X1 _12123_ (
    .A(_4679_),
    .B(_4678_),
    .Y(_4680_)
);

AND2X2 _12124_ (
    .A(_4680_),
    .B(_4663_),
    .Y(_4681_)
);

NOR2X1 _12125_ (
    .A(_4663_),
    .B(_4680_),
    .Y(_4682_)
);

OAI21X1 _12126_ (
    .A(_4682_),
    .B(_4681_),
    .C(_4417_),
    .Y(_4683_)
);

OAI21X1 _12127_ (
    .A(_4348__bF$buf1),
    .B(_4683_),
    .C(_4662_),
    .Y(_4205_)
);

OAI21X1 _12128_ (
    .A(_4679_),
    .B(_4663_),
    .C(_4677_),
    .Y(_4684_)
);

INVX1 _12129_ (
    .A(_4684_),
    .Y(_4685_)
);

NAND2X1 _12130_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [10]),
    .Y(_4686_)
);

OAI21X1 _12131_ (
    .A(1'h1),
    .B(_4560_),
    .C(_4686_),
    .Y(_4687_)
);

MUX2X1 _12132_ (
    .A(_4687_),
    .B(_4644_),
    .S(1'h0),
    .Y(_4688_)
);

NOR2X1 _12133_ (
    .A(_4324__bF$buf0),
    .B(_4688_),
    .Y(_4689_)
);

NAND2X1 _12134_ (
    .A(_4431_),
    .B(_4638_),
    .Y(_4690_)
);

NAND2X1 _12135_ (
    .A(_4647_),
    .B(_4430_),
    .Y(_4691_)
);

NAND2X1 _12136_ (
    .A(_4690_),
    .B(_4691_),
    .Y(_4692_)
);

OR2X2 _12137_ (
    .A(_4689_),
    .B(_4692_),
    .Y(_4693_)
);

OAI21X1 _12138_ (
    .A(_4673_),
    .B(_4664_),
    .C(_4362__bF$buf3),
    .Y(_4694_)
);

OR2X2 _12139_ (
    .A(_4694_),
    .B(_4693_),
    .Y(_4695_)
);

OAI21X1 _12140_ (
    .A(_4689_),
    .B(_4692_),
    .C(_4694_),
    .Y(_4696_)
);

AOI21X1 _12141_ (
    .A(_4695_),
    .B(_4696_),
    .C(_4370_),
    .Y(_4697_)
);

INVX1 _12142_ (
    .A(_4697_),
    .Y(_4698_)
);

NAND3X1 _12143_ (
    .A(_4370_),
    .B(_4696_),
    .C(_4695_),
    .Y(_4699_)
);

NAND2X1 _12144_ (
    .A(_4699_),
    .B(_4698_),
    .Y(_4700_)
);

OR2X2 _12145_ (
    .A(_4700_),
    .B(_4685_),
    .Y(_4701_)
);

NAND2X1 _12146_ (
    .A(_4685_),
    .B(_4700_),
    .Y(_4702_)
);

NAND2X1 _12147_ (
    .A(_4702_),
    .B(_4701_),
    .Y(_4703_)
);

AOI22X1 _12148_ (
    .A(_4316_),
    .B(_4348__bF$buf0),
    .C(_4703_),
    .D(_4346_),
    .Y(_4206_)
);

AOI21X1 _12149_ (
    .A(_4684_),
    .B(_4699_),
    .C(_4697_),
    .Y(_4704_)
);

NAND2X1 _12150_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4705_)
);

OAI21X1 _12151_ (
    .A(1'h1),
    .B(_4575_),
    .C(_4705_),
    .Y(_4706_)
);

NAND2X1 _12152_ (
    .A(1'h0),
    .B(_4706_),
    .Y(_4707_)
);

OAI21X1 _12153_ (
    .A(1'h0),
    .B(_4666_),
    .C(_4707_),
    .Y(_4708_)
);

NAND2X1 _12154_ (
    .A(1'h1),
    .B(_4708_),
    .Y(_4709_)
);

OAI21X1 _12155_ (
    .A(1'h1),
    .B(_4626_),
    .C(_4709_),
    .Y(_4710_)
);

INVX1 _12156_ (
    .A(_4710_),
    .Y(_4711_)
);

NAND3X1 _12157_ (
    .A(_4672_),
    .B(_4633_),
    .C(_4650_),
    .Y(_4712_)
);

OAI21X1 _12158_ (
    .A(_4693_),
    .B(_4712_),
    .C(_4362__bF$buf2),
    .Y(_4713_)
);

OR2X2 _12159_ (
    .A(_4713_),
    .B(_4711_),
    .Y(_4714_)
);

NOR2X1 _12160_ (
    .A(_4693_),
    .B(_4712_),
    .Y(_4715_)
);

OAI21X1 _12161_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4715_),
    .C(_4711_),
    .Y(_4716_)
);

NAND3X1 _12162_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(_4716_),
    .C(_4714_),
    .Y(_4717_)
);

OR2X2 _12163_ (
    .A(_4713_),
    .B(_4710_),
    .Y(_4718_)
);

OAI21X1 _12164_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4715_),
    .C(_4710_),
    .Y(_4719_)
);

NAND3X1 _12165_ (
    .A(_4329_),
    .B(_4719_),
    .C(_4718_),
    .Y(_4720_)
);

NAND2X1 _12166_ (
    .A(_4717_),
    .B(_4720_),
    .Y(_4721_)
);

OR2X2 _12167_ (
    .A(_4704_),
    .B(_4721_),
    .Y(_4722_)
);

NAND2X1 _12168_ (
    .A(_4721_),
    .B(_4704_),
    .Y(_4723_)
);

NAND2X1 _12169_ (
    .A(_4723_),
    .B(_4722_),
    .Y(_4724_)
);

AOI22X1 _12170_ (
    .A(_4311_),
    .B(_4348__bF$buf4),
    .C(_4724_),
    .D(_4346_),
    .Y(_4207_)
);

INVX1 _12171_ (
    .A(\genblk1[5].u_ce.Xcalc [5]),
    .Y(_4725_)
);

OAI21X1 _12172_ (
    .A(_4721_),
    .B(_4704_),
    .C(_4717_),
    .Y(_4726_)
);

NAND2X1 _12173_ (
    .A(_4711_),
    .B(_4715_),
    .Y(_4727_)
);

NOR2X1 _12174_ (
    .A(_4325__bF$buf3),
    .B(_4601_),
    .Y(_4728_)
);

AOI21X1 _12175_ (
    .A(_4325__bF$buf2),
    .B(_4687_),
    .C(_4728_),
    .Y(_4729_)
);

NAND2X1 _12176_ (
    .A(_4324__bF$buf4),
    .B(_4649_),
    .Y(_4730_)
);

OAI21X1 _12177_ (
    .A(_4324__bF$buf3),
    .B(_4729_),
    .C(_4730_),
    .Y(_4731_)
);

INVX1 _12178_ (
    .A(_4731_),
    .Y(_4732_)
);

NAND3X1 _12179_ (
    .A(_4362__bF$buf1),
    .B(_4732_),
    .C(_4727_),
    .Y(_4733_)
);

NOR2X1 _12180_ (
    .A(_4692_),
    .B(_4689_),
    .Y(_4734_)
);

NAND3X1 _12181_ (
    .A(_4672_),
    .B(_4734_),
    .C(_4675_),
    .Y(_4735_)
);

OAI21X1 _12182_ (
    .A(_4710_),
    .B(_4735_),
    .C(_4362__bF$buf0),
    .Y(_4736_)
);

NAND2X1 _12183_ (
    .A(_4731_),
    .B(_4736_),
    .Y(_4737_)
);

AOI21X1 _12184_ (
    .A(_4733_),
    .B(_4737_),
    .C(_4366_),
    .Y(_4738_)
);

INVX1 _12185_ (
    .A(_4738_),
    .Y(_4739_)
);

NAND3X1 _12186_ (
    .A(_4366_),
    .B(_4737_),
    .C(_4733_),
    .Y(_4740_)
);

NAND2X1 _12187_ (
    .A(_4740_),
    .B(_4739_),
    .Y(_4741_)
);

NOR2X1 _12188_ (
    .A(_4741_),
    .B(_4726_),
    .Y(_4742_)
);

AND2X2 _12189_ (
    .A(_4726_),
    .B(_4741_),
    .Y(_4743_)
);

OAI21X1 _12190_ (
    .A(_4742_),
    .B(_4743_),
    .C(_4346_),
    .Y(_4744_)
);

OAI21X1 _12191_ (
    .A(_4725_),
    .B(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .C(_4744_),
    .Y(_4208_)
);

INVX1 _12192_ (
    .A(\genblk1[5].u_ce.Xcalc [6]),
    .Y(_4745_)
);

NAND3X1 _12193_ (
    .A(_4711_),
    .B(_4732_),
    .C(_4715_),
    .Y(_4746_)
);

AOI21X1 _12194_ (
    .A(_4325__bF$buf1),
    .B(_4706_),
    .C(_4728_),
    .Y(_4747_)
);

NAND2X1 _12195_ (
    .A(1'h1),
    .B(_4747_),
    .Y(_4748_)
);

OAI21X1 _12196_ (
    .A(1'h1),
    .B(_4668_),
    .C(_4748_),
    .Y(_4749_)
);

NAND3X1 _12197_ (
    .A(_4362__bF$buf5),
    .B(_4749_),
    .C(_4746_),
    .Y(_4750_)
);

NOR3X1 _12198_ (
    .A(_4710_),
    .B(_4731_),
    .C(_4735_),
    .Y(_4751_)
);

INVX1 _12199_ (
    .A(_4749_),
    .Y(_4752_)
);

OAI21X1 _12200_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4751_),
    .C(_4752_),
    .Y(_4753_)
);

NAND2X1 _12201_ (
    .A(_4750_),
    .B(_4753_),
    .Y(_4754_)
);

NAND2X1 _12202_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(_4754_),
    .Y(_4755_)
);

NAND3X1 _12203_ (
    .A(_4326_),
    .B(_4750_),
    .C(_4753_),
    .Y(_4756_)
);

NAND2X1 _12204_ (
    .A(_4756_),
    .B(_4755_),
    .Y(_4757_)
);

AOI21X1 _12205_ (
    .A(_4718_),
    .B(_4719_),
    .C(_4329_),
    .Y(_4758_)
);

NOR2X1 _12206_ (
    .A(_4758_),
    .B(_4738_),
    .Y(_4759_)
);

OAI21X1 _12207_ (
    .A(_4721_),
    .B(_4704_),
    .C(_4759_),
    .Y(_4760_)
);

NAND2X1 _12208_ (
    .A(_4740_),
    .B(_4760_),
    .Y(_4761_)
);

NOR2X1 _12209_ (
    .A(_4757_),
    .B(_4761_),
    .Y(_4762_)
);

AND2X2 _12210_ (
    .A(_4755_),
    .B(_4756_),
    .Y(_4763_)
);

AND2X2 _12211_ (
    .A(_4717_),
    .B(_4720_),
    .Y(_4764_)
);

NAND3X1 _12212_ (
    .A(_4740_),
    .B(_4764_),
    .C(_4739_),
    .Y(_4765_)
);

AOI21X1 _12213_ (
    .A(_4758_),
    .B(_4740_),
    .C(_4738_),
    .Y(_4766_)
);

OAI21X1 _12214_ (
    .A(_4704_),
    .B(_4765_),
    .C(_4766_),
    .Y(_4767_)
);

NOR2X1 _12215_ (
    .A(_4763_),
    .B(_4767_),
    .Y(_4768_)
);

OAI21X1 _12216_ (
    .A(_4768_),
    .B(_4762_),
    .C(_4417_),
    .Y(_4769_)
);

NAND2X1 _12217_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .B(_4769_),
    .Y(_4770_)
);

OAI21X1 _12218_ (
    .A(_4745_),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .C(_4770_),
    .Y(_4209_)
);

INVX1 _12219_ (
    .A(\genblk1[5].u_ce.Xcalc [7]),
    .Y(_4771_)
);

INVX1 _12220_ (
    .A(_4755_),
    .Y(_4772_)
);

NAND2X1 _12221_ (
    .A(_4749_),
    .B(_4751_),
    .Y(_4773_)
);

NOR2X1 _12222_ (
    .A(_4324__bF$buf2),
    .B(_4601_),
    .Y(_4774_)
);

INVX1 _12223_ (
    .A(_4774_),
    .Y(_4775_)
);

OAI21X1 _12224_ (
    .A(1'h1),
    .B(_4688_),
    .C(_4775_),
    .Y(_4776_)
);

NAND3X1 _12225_ (
    .A(_4362__bF$buf4),
    .B(_4776_),
    .C(_4773_),
    .Y(_4777_)
);

INVX1 _12226_ (
    .A(_4776_),
    .Y(_4778_)
);

OAI21X1 _12227_ (
    .A(_4752_),
    .B(_4746_),
    .C(_4362__bF$buf3),
    .Y(_4779_)
);

NAND2X1 _12228_ (
    .A(_4778_),
    .B(_4779_),
    .Y(_4780_)
);

NAND3X1 _12229_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(_4777_),
    .C(_4780_),
    .Y(_4781_)
);

NAND3X1 _12230_ (
    .A(_4362__bF$buf2),
    .B(_4778_),
    .C(_4773_),
    .Y(_4782_)
);

NAND2X1 _12231_ (
    .A(_4776_),
    .B(_4779_),
    .Y(_4783_)
);

NAND3X1 _12232_ (
    .A(_4363_),
    .B(_4782_),
    .C(_4783_),
    .Y(_4784_)
);

NAND2X1 _12233_ (
    .A(_4781_),
    .B(_4784_),
    .Y(_4785_)
);

OAI21X1 _12234_ (
    .A(_4772_),
    .B(_4762_),
    .C(_4785_),
    .Y(_4786_)
);

NOR2X1 _12235_ (
    .A(_4772_),
    .B(_4762_),
    .Y(_4787_)
);

INVX1 _12236_ (
    .A(_4785_),
    .Y(_4788_)
);

AOI21X1 _12237_ (
    .A(_4787_),
    .B(_4788_),
    .C(_4345_),
    .Y(_4789_)
);

AOI22X1 _12238_ (
    .A(_4771_),
    .B(_4348__bF$buf3),
    .C(_4789_),
    .D(_4786_),
    .Y(_4210_)
);

OAI21X1 _12239_ (
    .A(_4755_),
    .B(_4785_),
    .C(_4781_),
    .Y(_4790_)
);

NOR2X1 _12240_ (
    .A(_4757_),
    .B(_4785_),
    .Y(_4791_)
);

AOI21X1 _12241_ (
    .A(_4791_),
    .B(_4767_),
    .C(_4790_),
    .Y(_4792_)
);

INVX1 _12242_ (
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4793_)
);

NAND3X1 _12243_ (
    .A(_4749_),
    .B(_4778_),
    .C(_4751_),
    .Y(_4794_)
);

INVX1 _12244_ (
    .A(_4708_),
    .Y(_4795_)
);

OAI21X1 _12245_ (
    .A(1'h1),
    .B(_4795_),
    .C(_4775_),
    .Y(_4796_)
);

INVX1 _12246_ (
    .A(_4796_),
    .Y(_4797_)
);

NAND3X1 _12247_ (
    .A(_4362__bF$buf1),
    .B(_4797_),
    .C(_4794_),
    .Y(_4798_)
);

OAI21X1 _12248_ (
    .A(_4776_),
    .B(_4773_),
    .C(_4362__bF$buf0),
    .Y(_4799_)
);

NAND2X1 _12249_ (
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

AOI21X1 _12250_ (
    .A(_4800_),
    .B(_4798_),
    .C(_4793_),
    .Y(_4801_)
);

NAND3X1 _12251_ (
    .A(_4362__bF$buf5),
    .B(_4796_),
    .C(_4794_),
    .Y(_4802_)
);

NAND2X1 _12252_ (
    .A(_4797_),
    .B(_4799_),
    .Y(_4803_)
);

AOI21X1 _12253_ (
    .A(_4803_),
    .B(_4802_),
    .C(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4804_)
);

OAI21X1 _12254_ (
    .A(_4801_),
    .B(_4804_),
    .C(_4792_),
    .Y(_4805_)
);

INVX1 _12255_ (
    .A(_4805_),
    .Y(_4806_)
);

OR2X2 _12256_ (
    .A(_4801_),
    .B(_4804_),
    .Y(_4807_)
);

OAI21X1 _12257_ (
    .A(_4807_),
    .B(_4792_),
    .C(_4346_),
    .Y(_4808_)
);

OAI22X1 _12258_ (
    .A(_4308_),
    .B(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .C(_4808_),
    .D(_4806_),
    .Y(_4211_)
);

NAND2X1 _12259_ (
    .A(\genblk1[5].u_ce.Xcalc [9]),
    .B(_4348__bF$buf2),
    .Y(_4809_)
);

NOR2X1 _12260_ (
    .A(_4807_),
    .B(_4792_),
    .Y(_4810_)
);

NOR2X1 _12261_ (
    .A(_4801_),
    .B(_4810_),
    .Y(_4811_)
);

OAI21X1 _12262_ (
    .A(1'h1),
    .B(_4729_),
    .C(_4775_),
    .Y(_4812_)
);

INVX1 _12263_ (
    .A(_4812_),
    .Y(_4813_)
);

OAI21X1 _12264_ (
    .A(_4796_),
    .B(_4794_),
    .C(_4362__bF$buf4),
    .Y(_4814_)
);

NAND2X1 _12265_ (
    .A(_4813_),
    .B(_4814_),
    .Y(_4815_)
);

OR2X2 _12266_ (
    .A(_4814_),
    .B(_4813_),
    .Y(_4816_)
);

NAND3X1 _12267_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(_4815_),
    .C(_4816_),
    .Y(_4817_)
);

NAND2X1 _12268_ (
    .A(_4815_),
    .B(_4816_),
    .Y(_4818_)
);

NAND2X1 _12269_ (
    .A(_4425_),
    .B(_4818_),
    .Y(_4819_)
);

NAND2X1 _12270_ (
    .A(_4817_),
    .B(_4819_),
    .Y(_4820_)
);

AND2X2 _12271_ (
    .A(_4811_),
    .B(_4820_),
    .Y(_4821_)
);

OAI21X1 _12272_ (
    .A(_4820_),
    .B(_4811_),
    .C(_4346_),
    .Y(_4822_)
);

OAI21X1 _12273_ (
    .A(_4822_),
    .B(_4821_),
    .C(_4809_),
    .Y(_4212_)
);

INVX1 _12274_ (
    .A(\genblk1[5].u_ce.Xcalc [10]),
    .Y(_4823_)
);

INVX1 _12275_ (
    .A(_4817_),
    .Y(_4824_)
);

AOI21X1 _12276_ (
    .A(_4801_),
    .B(_4819_),
    .C(_4824_),
    .Y(_4825_)
);

NOR2X1 _12277_ (
    .A(_4801_),
    .B(_4804_),
    .Y(_4826_)
);

NAND3X1 _12278_ (
    .A(_4817_),
    .B(_4819_),
    .C(_4826_),
    .Y(_4827_)
);

OAI21X1 _12279_ (
    .A(_4792_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4828_)
);

OAI21X1 _12280_ (
    .A(1'h1),
    .B(_4747_),
    .C(_4775_),
    .Y(_4829_)
);

INVX1 _12281_ (
    .A(_4829_),
    .Y(_4830_)
);

OR2X2 _12282_ (
    .A(_4794_),
    .B(_4796_),
    .Y(_4831_)
);

OAI21X1 _12283_ (
    .A(_4812_),
    .B(_4831_),
    .C(_4362__bF$buf3),
    .Y(_4832_)
);

NAND2X1 _12284_ (
    .A(_4830_),
    .B(_4832_),
    .Y(_4833_)
);

OR2X2 _12285_ (
    .A(_4832_),
    .B(_4830_),
    .Y(_4834_)
);

NAND3X1 _12286_ (
    .A(\genblk1[5].u_ce.Xin12b [10]),
    .B(_4833_),
    .C(_4834_),
    .Y(_4835_)
);

AND2X2 _12287_ (
    .A(_4832_),
    .B(_4830_),
    .Y(_4836_)
);

NOR2X1 _12288_ (
    .A(_4830_),
    .B(_4832_),
    .Y(_4837_)
);

OAI21X1 _12289_ (
    .A(_4837_),
    .B(_4836_),
    .C(_4446_),
    .Y(_4838_)
);

NAND2X1 _12290_ (
    .A(_4838_),
    .B(_4835_),
    .Y(_4839_)
);

AND2X2 _12291_ (
    .A(_4828_),
    .B(_4839_),
    .Y(_4840_)
);

NOR2X1 _12292_ (
    .A(_4839_),
    .B(_4828_),
    .Y(_4841_)
);

NOR2X1 _12293_ (
    .A(_4840_),
    .B(_4841_),
    .Y(_4842_)
);

AOI22X1 _12294_ (
    .A(_4823_),
    .B(_4348__bF$buf1),
    .C(_4842_),
    .D(_4346_),
    .Y(_4213_)
);

NAND2X1 _12295_ (
    .A(\genblk1[5].u_ce.Xcalc [11]),
    .B(_4348__bF$buf0),
    .Y(_4843_)
);

INVX1 _12296_ (
    .A(_4835_),
    .Y(_4844_)
);

AOI21X1 _12297_ (
    .A(_4828_),
    .B(_4838_),
    .C(_4844_),
    .Y(_4845_)
);

NAND2X1 _12298_ (
    .A(_4362__bF$buf2),
    .B(_4833_),
    .Y(_4846_)
);

NOR2X1 _12299_ (
    .A(_4603_),
    .B(_4846_),
    .Y(_4847_)
);

AOI21X1 _12300_ (
    .A(_4833_),
    .B(_4362__bF$buf1),
    .C(_4604_),
    .Y(_4848_)
);

NOR2X1 _12301_ (
    .A(_4848_),
    .B(_4847_),
    .Y(_4849_)
);

AND2X2 _12302_ (
    .A(_4845_),
    .B(_4849_),
    .Y(_4850_)
);

OAI21X1 _12303_ (
    .A(_4849_),
    .B(_4845_),
    .C(_4346_),
    .Y(_4851_)
);

OAI21X1 _12304_ (
    .A(_4851_),
    .B(_4850_),
    .C(_4843_),
    .Y(_4214_)
);

OAI21X1 _12305_ (
    .A(1'h1),
    .B(_4325__bF$buf0),
    .C(_4344_),
    .Y(_4852_)
);

OAI21X1 _12306_ (
    .A(_4619_),
    .B(_4852_),
    .C(\genblk1[5].u_ce.Ain0 [0]),
    .Y(_4853_)
);

INVX1 _12307_ (
    .A(\genblk1[5].u_ce.Ain0 [0]),
    .Y(_4854_)
);

NOR2X1 _12308_ (
    .A(_4619_),
    .B(_4852_),
    .Y(_4855_)
);

NAND2X1 _12309_ (
    .A(_4854_),
    .B(_4855_),
    .Y(_4856_)
);

NAND2X1 _12310_ (
    .A(_4853_),
    .B(_4856_),
    .Y(_4857_)
);

NAND2X1 _12311_ (
    .A(\genblk1[5].u_ce.Acalc [0]),
    .B(_4348__bF$buf4),
    .Y(_4858_)
);

OAI21X1 _12312_ (
    .A(_4348__bF$buf3),
    .B(_4857_),
    .C(_4858_),
    .Y(_4215_)
);

NAND2X1 _12313_ (
    .A(\genblk1[5].u_ce.Acalc [1]),
    .B(_4348__bF$buf2),
    .Y(_4859_)
);

INVX1 _12314_ (
    .A(_4853_),
    .Y(_4860_)
);

NOR2X1 _12315_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_4861_)
);

AOI21X1 _12316_ (
    .A(_4619_),
    .B(1'h1),
    .C(_4861_),
    .Y(_4862_)
);

NOR2X1 _12317_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4862_),
    .Y(_4863_)
);

OAI21X1 _12318_ (
    .A(_4619_),
    .B(_4852_),
    .C(_4362__bF$buf0),
    .Y(_4864_)
);

AND2X2 _12319_ (
    .A(_4864_),
    .B(_4862_),
    .Y(_4865_)
);

OR2X2 _12320_ (
    .A(_4865_),
    .B(_4863_),
    .Y(_4866_)
);

OR2X2 _12321_ (
    .A(_4866_),
    .B(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4867_)
);

OAI21X1 _12322_ (
    .A(_4863_),
    .B(_4865_),
    .C(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4868_)
);

NAND2X1 _12323_ (
    .A(_4868_),
    .B(_4867_),
    .Y(_4869_)
);

NOR2X1 _12324_ (
    .A(_4860_),
    .B(_4869_),
    .Y(_4870_)
);

NAND2X1 _12325_ (
    .A(_4860_),
    .B(_4869_),
    .Y(_4871_)
);

NAND2X1 _12326_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .B(_4871_),
    .Y(_4872_)
);

OAI21X1 _12327_ (
    .A(_4870_),
    .B(_4872_),
    .C(_4859_),
    .Y(_4216_)
);

INVX1 _12328_ (
    .A(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4873_)
);

OAI21X1 _12329_ (
    .A(_4873_),
    .B(_4866_),
    .C(_4871_),
    .Y(_4874_)
);

OAI21X1 _12330_ (
    .A(_4354_),
    .B(_4325__bF$buf4),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_4875_)
);

OAI21X1 _12331_ (
    .A(1'h1),
    .B(1'h0),
    .C(1'h1),
    .Y(_4876_)
);

MUX2X1 _12332_ (
    .A(_4876_),
    .B(1'h1),
    .S(_4875_),
    .Y(_4877_)
);

NAND2X1 _12333_ (
    .A(\genblk1[5].u_ce.Ain1 [0]),
    .B(_4877_),
    .Y(_4878_)
);

OR2X2 _12334_ (
    .A(_4877_),
    .B(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_4879_)
);

NAND2X1 _12335_ (
    .A(_4878_),
    .B(_4879_),
    .Y(_4880_)
);

INVX1 _12336_ (
    .A(_4880_),
    .Y(_4881_)
);

NOR2X1 _12337_ (
    .A(_4881_),
    .B(_4874_),
    .Y(_4882_)
);

NAND2X1 _12338_ (
    .A(_4881_),
    .B(_4874_),
    .Y(_4883_)
);

NAND2X1 _12339_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(_4883_),
    .Y(_4884_)
);

OAI22X1 _12340_ (
    .A(_4270_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4882_),
    .D(_4884_),
    .Y(_4217_)
);

NOR2X1 _12341_ (
    .A(\genblk1[5].u_ce.Acalc [3]),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4885_)
);

NAND2X1 _12342_ (
    .A(_4878_),
    .B(_4883_),
    .Y(_4886_)
);

INVX1 _12343_ (
    .A(_4886_),
    .Y(_4887_)
);

INVX1 _12344_ (
    .A(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_4888_)
);

NOR2X1 _12345_ (
    .A(1'h1),
    .B(_4325__bF$buf3),
    .Y(_4889_)
);

OAI21X1 _12346_ (
    .A(_4324__bF$buf1),
    .B(_4889_),
    .C(_4362__bF$buf5),
    .Y(_4890_)
);

OAI21X1 _12347_ (
    .A(1'h1),
    .B(1'h0),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_4891_)
);

OAI21X1 _12348_ (
    .A(_4354_),
    .B(_4891_),
    .C(_4890_),
    .Y(_4892_)
);

NOR2X1 _12349_ (
    .A(_4888_),
    .B(_4892_),
    .Y(_4893_)
);

NAND2X1 _12350_ (
    .A(_4888_),
    .B(_4892_),
    .Y(_4894_)
);

INVX1 _12351_ (
    .A(_4894_),
    .Y(_4895_)
);

NOR2X1 _12352_ (
    .A(_4893_),
    .B(_4895_),
    .Y(_4896_)
);

OAI21X1 _12353_ (
    .A(_4896_),
    .B(_4887_),
    .C(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .Y(_4897_)
);

AOI21X1 _12354_ (
    .A(_4887_),
    .B(_4896_),
    .C(_4897_),
    .Y(_4898_)
);

NOR2X1 _12355_ (
    .A(_4885_),
    .B(_4898_),
    .Y(_4218_)
);

NAND2X1 _12356_ (
    .A(\genblk1[5].u_ce.Acalc [4]),
    .B(_4348__bF$buf1),
    .Y(_4899_)
);

INVX1 _12357_ (
    .A(\genblk1[5].u_ce.Ain12b [4]),
    .Y(_4900_)
);

AOI21X1 _12358_ (
    .A(_4619_),
    .B(1'h1),
    .C(_4362__bF$buf4),
    .Y(_4901_)
);

OAI21X1 _12359_ (
    .A(1'h1),
    .B(_4619_),
    .C(_4901_),
    .Y(_4902_)
);

OAI21X1 _12360_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4862_),
    .C(_4902_),
    .Y(_4903_)
);

OR2X2 _12361_ (
    .A(_4903_),
    .B(_4900_),
    .Y(_4904_)
);

NAND2X1 _12362_ (
    .A(_4900_),
    .B(_4903_),
    .Y(_4905_)
);

NAND2X1 _12363_ (
    .A(_4905_),
    .B(_4904_),
    .Y(_4906_)
);

AOI21X1 _12364_ (
    .A(_4886_),
    .B(_4894_),
    .C(_4893_),
    .Y(_4907_)
);

AND2X2 _12365_ (
    .A(_4907_),
    .B(_4906_),
    .Y(_4908_)
);

OAI21X1 _12366_ (
    .A(_4906_),
    .B(_4907_),
    .C(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4909_)
);

OAI21X1 _12367_ (
    .A(_4909_),
    .B(_4908_),
    .C(_4899_),
    .Y(_4219_)
);

OAI21X1 _12368_ (
    .A(_4906_),
    .B(_4907_),
    .C(_4904_),
    .Y(_4910_)
);

INVX1 _12369_ (
    .A(\genblk1[5].u_ce.Ain12b [5]),
    .Y(_4911_)
);

OAI21X1 _12370_ (
    .A(_4618_),
    .B(_4431_),
    .C(_4362__bF$buf3),
    .Y(_4912_)
);

OAI21X1 _12371_ (
    .A(1'h1),
    .B(1'h0),
    .C(_4344_),
    .Y(_4913_)
);

OR2X2 _12372_ (
    .A(_4913_),
    .B(_4362__bF$buf2),
    .Y(_4914_)
);

NAND2X1 _12373_ (
    .A(_4912_),
    .B(_4914_),
    .Y(_4915_)
);

OR2X2 _12374_ (
    .A(_4915_),
    .B(_4911_),
    .Y(_4916_)
);

NAND2X1 _12375_ (
    .A(_4911_),
    .B(_4915_),
    .Y(_4917_)
);

NAND2X1 _12376_ (
    .A(_4917_),
    .B(_4916_),
    .Y(_4918_)
);

INVX1 _12377_ (
    .A(_4918_),
    .Y(_4919_)
);

NOR2X1 _12378_ (
    .A(_4919_),
    .B(_4910_),
    .Y(_4920_)
);

NAND2X1 _12379_ (
    .A(_4919_),
    .B(_4910_),
    .Y(_4921_)
);

NAND2X1 _12380_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .B(_4921_),
    .Y(_4922_)
);

OAI22X1 _12381_ (
    .A(_4287_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4920_),
    .D(_4922_),
    .Y(_4220_)
);

NAND2X1 _12382_ (
    .A(\genblk1[5].u_ce.Acalc [6]),
    .B(_4348__bF$buf0),
    .Y(_4923_)
);

INVX1 _12383_ (
    .A(_4906_),
    .Y(_4924_)
);

NAND2X1 _12384_ (
    .A(_4919_),
    .B(_4924_),
    .Y(_4925_)
);

OAI21X1 _12385_ (
    .A(_4904_),
    .B(_4918_),
    .C(_4916_),
    .Y(_4926_)
);

INVX1 _12386_ (
    .A(_4926_),
    .Y(_4927_)
);

OAI21X1 _12387_ (
    .A(_4925_),
    .B(_4907_),
    .C(_4927_),
    .Y(_4928_)
);

OAI21X1 _12388_ (
    .A(1'h0),
    .B(_4354_),
    .C(_4324__bF$buf0),
    .Y(_4929_)
);

NOR2X1 _12389_ (
    .A(_4929_),
    .B(_4889_),
    .Y(_4930_)
);

NAND2X1 _12390_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4930_),
    .Y(_4931_)
);

OAI21X1 _12391_ (
    .A(_4929_),
    .B(_4889_),
    .C(_4362__bF$buf1),
    .Y(_4932_)
);

NAND2X1 _12392_ (
    .A(_4932_),
    .B(_4931_),
    .Y(_4933_)
);

NAND2X1 _12393_ (
    .A(\genblk1[5].u_ce.Ain12b [6]),
    .B(_4933_),
    .Y(_4934_)
);

OR2X2 _12394_ (
    .A(_4933_),
    .B(\genblk1[5].u_ce.Ain12b [6]),
    .Y(_4935_)
);

NAND2X1 _12395_ (
    .A(_4934_),
    .B(_4935_),
    .Y(_4936_)
);

INVX1 _12396_ (
    .A(_4936_),
    .Y(_4937_)
);

NOR2X1 _12397_ (
    .A(_4937_),
    .B(_4928_),
    .Y(_4938_)
);

NAND2X1 _12398_ (
    .A(_4937_),
    .B(_4928_),
    .Y(_4939_)
);

NAND2X1 _12399_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .B(_4939_),
    .Y(_4940_)
);

OAI21X1 _12400_ (
    .A(_4938_),
    .B(_4940_),
    .C(_4923_),
    .Y(_4221_)
);

INVX1 _12401_ (
    .A(\genblk1[5].u_ce.Acalc [7]),
    .Y(_4941_)
);

NAND2X1 _12402_ (
    .A(_4934_),
    .B(_4939_),
    .Y(_4942_)
);

INVX1 _12403_ (
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .Y(_4943_)
);

NAND2X1 _12404_ (
    .A(_4362__bF$buf0),
    .B(_4861_),
    .Y(_4944_)
);

OR2X2 _12405_ (
    .A(_4861_),
    .B(_4362__bF$buf5),
    .Y(_4945_)
);

NAND2X1 _12406_ (
    .A(_4944_),
    .B(_4945_),
    .Y(_4946_)
);

NOR2X1 _12407_ (
    .A(_4943_),
    .B(_4946_),
    .Y(_4947_)
);

INVX1 _12408_ (
    .A(_4947_),
    .Y(_4948_)
);

NAND2X1 _12409_ (
    .A(_4943_),
    .B(_4946_),
    .Y(_4949_)
);

NAND2X1 _12410_ (
    .A(_4949_),
    .B(_4948_),
    .Y(_4950_)
);

OR2X2 _12411_ (
    .A(_4942_),
    .B(_4950_),
    .Y(_4951_)
);

AOI21X1 _12412_ (
    .A(_4942_),
    .B(_4950_),
    .C(_4348__bF$buf4),
    .Y(_4952_)
);

AOI22X1 _12413_ (
    .A(_4941_),
    .B(_4348__bF$buf3),
    .C(_4951_),
    .D(_4952_),
    .Y(_4222_)
);

NAND2X1 _12414_ (
    .A(\genblk1[5].u_ce.Acalc [8]),
    .B(_4348__bF$buf2),
    .Y(_4953_)
);

NOR2X1 _12415_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4344_),
    .Y(_4954_)
);

INVX1 _12416_ (
    .A(_4954_),
    .Y(_4955_)
);

NAND3X1 _12417_ (
    .A(\genblk1[5].u_ce.Ain12b [8]),
    .B(_4891_),
    .C(_4955_),
    .Y(_4956_)
);

INVX1 _12418_ (
    .A(_4956_),
    .Y(_4957_)
);

AOI21X1 _12419_ (
    .A(_4955_),
    .B(_4891_),
    .C(\genblk1[5].u_ce.Ain12b [8]),
    .Y(_4958_)
);

NOR2X1 _12420_ (
    .A(_4958_),
    .B(_4957_),
    .Y(_4959_)
);

OAI21X1 _12421_ (
    .A(_4934_),
    .B(_4950_),
    .C(_4948_),
    .Y(_4960_)
);

NOR2X1 _12422_ (
    .A(_4950_),
    .B(_4936_),
    .Y(_4961_)
);

AOI21X1 _12423_ (
    .A(_4961_),
    .B(_4926_),
    .C(_4960_),
    .Y(_4962_)
);

NAND3X1 _12424_ (
    .A(_4924_),
    .B(_4919_),
    .C(_4961_),
    .Y(_4963_)
);

OAI21X1 _12425_ (
    .A(_4963_),
    .B(_4907_),
    .C(_4962_),
    .Y(_4964_)
);

NOR2X1 _12426_ (
    .A(_4959_),
    .B(_4964_),
    .Y(_4965_)
);

NAND2X1 _12427_ (
    .A(_4959_),
    .B(_4964_),
    .Y(_4966_)
);

NAND2X1 _12428_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .B(_4966_),
    .Y(_4967_)
);

OAI21X1 _12429_ (
    .A(_4965_),
    .B(_4967_),
    .C(_4953_),
    .Y(_4223_)
);

AOI21X1 _12430_ (
    .A(_4964_),
    .B(_4959_),
    .C(_4957_),
    .Y(_4968_)
);

OR2X2 _12431_ (
    .A(_4362__bF$buf4),
    .B(\genblk1[5].u_ce.Ain12b [9]),
    .Y(_4969_)
);

NAND2X1 _12432_ (
    .A(\genblk1[5].u_ce.Ain12b [9]),
    .B(_4362__bF$buf3),
    .Y(_4970_)
);

NAND2X1 _12433_ (
    .A(_4970_),
    .B(_4969_),
    .Y(_4971_)
);

AND2X2 _12434_ (
    .A(_4968_),
    .B(_4971_),
    .Y(_4972_)
);

OAI21X1 _12435_ (
    .A(_4971_),
    .B(_4968_),
    .C(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .Y(_4973_)
);

OAI22X1 _12436_ (
    .A(_4284_),
    .B(\genblk1[5].u_ce.Vld_bF$buf4 ),
    .C(_4973_),
    .D(_4972_),
    .Y(_4224_)
);

NAND2X1 _12437_ (
    .A(\genblk1[5].u_ce.Acalc [10]),
    .B(_4348__bF$buf1),
    .Y(_4974_)
);

OAI21X1 _12438_ (
    .A(_4971_),
    .B(_4956_),
    .C(_4970_),
    .Y(_4975_)
);

NAND3X1 _12439_ (
    .A(_4969_),
    .B(_4970_),
    .C(_4959_),
    .Y(_4976_)
);

INVX1 _12440_ (
    .A(_4976_),
    .Y(_4977_)
);

AOI21X1 _12441_ (
    .A(_4964_),
    .B(_4977_),
    .C(_4975_),
    .Y(_4978_)
);

INVX1 _12442_ (
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .Y(_4979_)
);

NAND2X1 _12443_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4979_),
    .Y(_4980_)
);

NAND2X1 _12444_ (
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .B(_4362__bF$buf2),
    .Y(_4981_)
);

NAND2X1 _12445_ (
    .A(_4980_),
    .B(_4981_),
    .Y(_4982_)
);

AND2X2 _12446_ (
    .A(_4978_),
    .B(_4982_),
    .Y(_4983_)
);

OAI21X1 _12447_ (
    .A(_4982_),
    .B(_4978_),
    .C(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .Y(_4984_)
);

OAI21X1 _12448_ (
    .A(_4984_),
    .B(_4983_),
    .C(_4974_),
    .Y(_4225_)
);

NAND2X1 _12449_ (
    .A(\genblk1[5].u_ce.Acalc [11]),
    .B(_4348__bF$buf0),
    .Y(_4985_)
);

OAI21X1 _12450_ (
    .A(_4982_),
    .B(_4978_),
    .C(_4981_),
    .Y(_4986_)
);

OAI21X1 _12451_ (
    .A(_4348__bF$buf4),
    .B(_4986_),
    .C(_4985_),
    .Y(_4226_)
);

NAND2X1 _12452_ (
    .A(\genblk1[5].u_ce.LoadCtl [5]),
    .B(_4275_),
    .Y(_4987_)
);

NAND2X1 _12453_ (
    .A(_4276_),
    .B(_4282_),
    .Y(_4988_)
);

NOR2X1 _12454_ (
    .A(_4987_),
    .B(_4988_),
    .Y(_4989_)
);

NAND2X1 _12455_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_4989_),
    .Y(_4990_)
);

OAI21X1 _12456_ (
    .A(_4446_),
    .B(_4989_),
    .C(_4990_),
    .Y(_4227_)
);

NAND2X1 _12457_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_4989_),
    .Y(_4991_)
);

OAI21X1 _12458_ (
    .A(_4514_),
    .B(_4989_),
    .C(_4991_),
    .Y(_4228_)
);

INVX1 _12459_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .Y(_4992_)
);

OR2X2 _12460_ (
    .A(_4988_),
    .B(_4275_),
    .Y(_4993_)
);

OAI21X1 _12461_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4994_)
);

OAI21X1 _12462_ (
    .A(_4992_),
    .B(_4993_),
    .C(_4994_),
    .Y(_4229_)
);

INVX1 _12463_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .Y(_4995_)
);

OAI21X1 _12464_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Xin12b [9]),
    .Y(_4996_)
);

OAI21X1 _12465_ (
    .A(_4995_),
    .B(_4993_),
    .C(_4996_),
    .Y(_4230_)
);

NAND2X1 _12466_ (
    .A(_4282_),
    .B(_4279_),
    .Y(_4997_)
);

NAND2X1 _12467_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(_4997_),
    .Y(_4998_)
);

OAI21X1 _12468_ (
    .A(_4992_),
    .B(_4997_),
    .C(_4998_),
    .Y(_4231_)
);

NAND2X1 _12469_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(_4997_),
    .Y(_4999_)
);

OAI21X1 _12470_ (
    .A(_4995_),
    .B(_4997_),
    .C(_4999_),
    .Y(_4232_)
);

AND2X2 _12471_ (
    .A(_4282_),
    .B(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_5000_)
);

NAND2X1 _12472_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_5000_),
    .Y(_5001_)
);

OAI21X1 _12473_ (
    .A(_4329_),
    .B(_5000_),
    .C(_5001_),
    .Y(_4233_)
);

NAND2X1 _12474_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_5000_),
    .Y(_5002_)
);

OAI21X1 _12475_ (
    .A(_4366_),
    .B(_5000_),
    .C(_5002_),
    .Y(_4234_)
);

OAI21X1 _12476_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_5003_)
);

OAI21X1 _12477_ (
    .A(_4992_),
    .B(_4273_),
    .C(_5003_),
    .Y(_4235_)
);

OAI21X1 _12478_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_5004_)
);

OAI21X1 _12479_ (
    .A(_4995_),
    .B(_4273_),
    .C(_5004_),
    .Y(_4236_)
);

NAND2X1 _12480_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.X_ [0]),
    .Y(_5005_)
);

OAI21X1 _12481_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4336_),
    .C(_5005_),
    .Y(_4237_)
);

NAND2X1 _12482_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.X_ [1]),
    .Y(_5006_)
);

OAI21X1 _12483_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4373_),
    .C(_5006_),
    .Y(_4238_)
);

NAND2X1 _12484_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_4989_),
    .Y(_5007_)
);

OAI21X1 _12485_ (
    .A(_4575_),
    .B(_4989_),
    .C(_5007_),
    .Y(_4239_)
);

NAND2X1 _12486_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_4989_),
    .Y(_5008_)
);

OAI21X1 _12487_ (
    .A(_4601_),
    .B(_4989_),
    .C(_5008_),
    .Y(_4240_)
);

INVX1 _12488_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .Y(_5009_)
);

OAI21X1 _12489_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_5010_)
);

OAI21X1 _12490_ (
    .A(_5009_),
    .B(_4993_),
    .C(_5010_),
    .Y(_4241_)
);

INVX1 _12491_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .Y(_5011_)
);

OAI21X1 _12492_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_5012_)
);

OAI21X1 _12493_ (
    .A(_5011_),
    .B(_4993_),
    .C(_5012_),
    .Y(_4242_)
);

NAND2X1 _12494_ (
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .B(_4997_),
    .Y(_5013_)
);

OAI21X1 _12495_ (
    .A(_5009_),
    .B(_4997_),
    .C(_5013_),
    .Y(_4243_)
);

NAND2X1 _12496_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(_4997_),
    .Y(_5014_)
);

OAI21X1 _12497_ (
    .A(_5011_),
    .B(_4997_),
    .C(_5014_),
    .Y(_4244_)
);

NAND2X1 _12498_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_5000_),
    .Y(_5015_)
);

OAI21X1 _12499_ (
    .A(_4445_),
    .B(_5000_),
    .C(_5015_),
    .Y(_4245_)
);

NAND2X1 _12500_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_5000_),
    .Y(_5016_)
);

OAI21X1 _12501_ (
    .A(_4466_),
    .B(_5000_),
    .C(_5016_),
    .Y(_4246_)
);

OAI21X1 _12502_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_5017_)
);

OAI21X1 _12503_ (
    .A(_5009_),
    .B(_4273_),
    .C(_5017_),
    .Y(_4247_)
);

OAI21X1 _12504_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_5018_)
);

OAI21X1 _12505_ (
    .A(_5011_),
    .B(_4273_),
    .C(_5018_),
    .Y(_4248_)
);

NAND2X1 _12506_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Y_ [0]),
    .Y(_5019_)
);

OAI21X1 _12507_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4323_),
    .C(_5019_),
    .Y(_4249_)
);

NAND2X1 _12508_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.Y_ [1]),
    .Y(_5020_)
);

OAI21X1 _12509_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4361_),
    .C(_5020_),
    .Y(_4250_)
);

NAND2X1 _12510_ (
    .A(\a[5] [0]),
    .B(_4989_),
    .Y(_5021_)
);

OAI21X1 _12511_ (
    .A(_4979_),
    .B(_4989_),
    .C(_5021_),
    .Y(_4251_)
);

NAND2X1 _12512_ (
    .A(\a[5] [1]),
    .B(_4989_),
    .Y(_5022_)
);

OAI21X1 _12513_ (
    .A(_4362__bF$buf1),
    .B(_4989_),
    .C(_5022_),
    .Y(_4252_)
);

INVX1 _12514_ (
    .A(\a[5] [0]),
    .Y(_5023_)
);

OAI21X1 _12515_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Ain12b [8]),
    .Y(_5024_)
);

OAI21X1 _12516_ (
    .A(_5023_),
    .B(_4993_),
    .C(_5024_),
    .Y(_4253_)
);

INVX1 _12517_ (
    .A(\a[5] [1]),
    .Y(_5025_)
);

OAI21X1 _12518_ (
    .A(_4275_),
    .B(_4988_),
    .C(\genblk1[5].u_ce.Ain12b [9]),
    .Y(_5026_)
);

OAI21X1 _12519_ (
    .A(_5025_),
    .B(_4993_),
    .C(_5026_),
    .Y(_4254_)
);

NAND2X1 _12520_ (
    .A(\genblk1[5].u_ce.Ain12b [6]),
    .B(_4997_),
    .Y(_5027_)
);

OAI21X1 _12521_ (
    .A(_5023_),
    .B(_4997_),
    .C(_5027_),
    .Y(_4255_)
);

NAND2X1 _12522_ (
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .B(_4997_),
    .Y(_4263_)
);

OAI21X1 _12523_ (
    .A(_5025_),
    .B(_4997_),
    .C(_4263_),
    .Y(_4256_)
);

NAND2X1 _12524_ (
    .A(\a[5] [0]),
    .B(_5000_),
    .Y(_4264_)
);

OAI21X1 _12525_ (
    .A(_4900_),
    .B(_5000_),
    .C(_4264_),
    .Y(_4257_)
);

NAND2X1 _12526_ (
    .A(\a[5] [1]),
    .B(_5000_),
    .Y(_4265_)
);

OAI21X1 _12527_ (
    .A(_4911_),
    .B(_5000_),
    .C(_4265_),
    .Y(_4258_)
);

OAI21X1 _12528_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_4266_)
);

OAI21X1 _12529_ (
    .A(_5023_),
    .B(_4273_),
    .C(_4266_),
    .Y(_4259_)
);

OAI21X1 _12530_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4271_),
    .C(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_4267_)
);

OAI21X1 _12531_ (
    .A(_5025_),
    .B(_4273_),
    .C(_4267_),
    .Y(_4260_)
);

NAND2X1 _12532_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[5] [0]),
    .Y(_4268_)
);

OAI21X1 _12533_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4854_),
    .C(_4268_),
    .Y(_4261_)
);

NAND2X1 _12534_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[5] [1]),
    .Y(_4269_)
);

OAI21X1 _12535_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4873_),
    .C(_4269_),
    .Y(_4262_)
);

DFFPOSX1 _12536_ (
    .CLK(clk_bF$buf76),
    .D(_4190_),
    .Q(\genblk1[5].u_ce.Ycalc [0])
);

DFFPOSX1 _12537_ (
    .CLK(clk_bF$buf75),
    .D(_4191_),
    .Q(\genblk1[5].u_ce.Ycalc [1])
);

DFFPOSX1 _12538_ (
    .CLK(clk_bF$buf74),
    .D(_4192_),
    .Q(\genblk1[5].u_ce.ISout )
);

DFFPOSX1 _12539_ (
    .CLK(clk_bF$buf73),
    .D(_4193_),
    .Q(\genblk1[5].u_ce.Ycalc [2])
);

DFFPOSX1 _12540_ (
    .CLK(clk_bF$buf72),
    .D(_4194_),
    .Q(\genblk1[5].u_ce.Ycalc [3])
);

DFFPOSX1 _12541_ (
    .CLK(clk_bF$buf71),
    .D(_4195_),
    .Q(\genblk1[5].u_ce.Ycalc [4])
);

DFFPOSX1 _12542_ (
    .CLK(clk_bF$buf70),
    .D(_4196_),
    .Q(\genblk1[5].u_ce.Ycalc [5])
);

DFFPOSX1 _12543_ (
    .CLK(clk_bF$buf69),
    .D(_4197_),
    .Q(\genblk1[5].u_ce.Ycalc [6])
);

DFFPOSX1 _12544_ (
    .CLK(clk_bF$buf68),
    .D(_4198_),
    .Q(\genblk1[5].u_ce.Ycalc [7])
);

DFFPOSX1 _12545_ (
    .CLK(clk_bF$buf67),
    .D(_4199_),
    .Q(\genblk1[5].u_ce.Ycalc [8])
);

DFFPOSX1 _12546_ (
    .CLK(clk_bF$buf66),
    .D(_4200_),
    .Q(\genblk1[5].u_ce.Ycalc [9])
);

DFFPOSX1 _12547_ (
    .CLK(clk_bF$buf65),
    .D(_4201_),
    .Q(\genblk1[5].u_ce.Ycalc [10])
);

DFFPOSX1 _12548_ (
    .CLK(clk_bF$buf64),
    .D(_4202_),
    .Q(\genblk1[5].u_ce.Ycalc [11])
);

DFFPOSX1 _12549_ (
    .CLK(clk_bF$buf63),
    .D(_4203_),
    .Q(\genblk1[5].u_ce.Xcalc [0])
);

DFFPOSX1 _12550_ (
    .CLK(clk_bF$buf62),
    .D(_4204_),
    .Q(\genblk1[5].u_ce.Xcalc [1])
);

DFFPOSX1 _12551_ (
    .CLK(clk_bF$buf61),
    .D(_4205_),
    .Q(\genblk1[5].u_ce.Xcalc [2])
);

DFFPOSX1 _12552_ (
    .CLK(clk_bF$buf60),
    .D(_4206_),
    .Q(\genblk1[5].u_ce.Xcalc [3])
);

DFFPOSX1 _12553_ (
    .CLK(clk_bF$buf59),
    .D(_4207_),
    .Q(\genblk1[5].u_ce.Xcalc [4])
);

DFFPOSX1 _12554_ (
    .CLK(clk_bF$buf58),
    .D(_4208_),
    .Q(\genblk1[5].u_ce.Xcalc [5])
);

DFFPOSX1 _12555_ (
    .CLK(clk_bF$buf57),
    .D(_4209_),
    .Q(\genblk1[5].u_ce.Xcalc [6])
);

DFFPOSX1 _12556_ (
    .CLK(clk_bF$buf56),
    .D(_4210_),
    .Q(\genblk1[5].u_ce.Xcalc [7])
);

DFFPOSX1 _12557_ (
    .CLK(clk_bF$buf55),
    .D(_4211_),
    .Q(\genblk1[5].u_ce.Xcalc [8])
);

DFFPOSX1 _12558_ (
    .CLK(clk_bF$buf54),
    .D(_4212_),
    .Q(\genblk1[5].u_ce.Xcalc [9])
);

DFFPOSX1 _12559_ (
    .CLK(clk_bF$buf53),
    .D(_4213_),
    .Q(\genblk1[5].u_ce.Xcalc [10])
);

DFFPOSX1 _12560_ (
    .CLK(clk_bF$buf52),
    .D(_4214_),
    .Q(\genblk1[5].u_ce.Xcalc [11])
);

DFFPOSX1 _12561_ (
    .CLK(clk_bF$buf51),
    .D(_4215_),
    .Q(\genblk1[5].u_ce.Acalc [0])
);

DFFPOSX1 _12562_ (
    .CLK(clk_bF$buf50),
    .D(_4216_),
    .Q(\genblk1[5].u_ce.Acalc [1])
);

DFFPOSX1 _12563_ (
    .CLK(clk_bF$buf49),
    .D(_4217_),
    .Q(\genblk1[5].u_ce.Acalc [2])
);

DFFPOSX1 _12564_ (
    .CLK(clk_bF$buf48),
    .D(_4218_),
    .Q(\genblk1[5].u_ce.Acalc [3])
);

DFFPOSX1 _12565_ (
    .CLK(clk_bF$buf47),
    .D(_4219_),
    .Q(\genblk1[5].u_ce.Acalc [4])
);

DFFPOSX1 _12566_ (
    .CLK(clk_bF$buf46),
    .D(_4220_),
    .Q(\genblk1[5].u_ce.Acalc [5])
);

DFFPOSX1 _12567_ (
    .CLK(clk_bF$buf45),
    .D(_4221_),
    .Q(\genblk1[5].u_ce.Acalc [6])
);

DFFPOSX1 _12568_ (
    .CLK(clk_bF$buf44),
    .D(_4222_),
    .Q(\genblk1[5].u_ce.Acalc [7])
);

DFFPOSX1 _12569_ (
    .CLK(clk_bF$buf43),
    .D(_4223_),
    .Q(\genblk1[5].u_ce.Acalc [8])
);

DFFPOSX1 _12570_ (
    .CLK(clk_bF$buf42),
    .D(_4224_),
    .Q(\genblk1[5].u_ce.Acalc [9])
);

DFFPOSX1 _12571_ (
    .CLK(clk_bF$buf41),
    .D(_4225_),
    .Q(\genblk1[5].u_ce.Acalc [10])
);

DFFPOSX1 _12572_ (
    .CLK(clk_bF$buf40),
    .D(_4226_),
    .Q(\genblk1[5].u_ce.Acalc [11])
);

DFFPOSX1 _12573_ (
    .CLK(clk_bF$buf39),
    .D(_4227_),
    .Q(\genblk1[5].u_ce.Xin12b [10])
);

DFFPOSX1 _12574_ (
    .CLK(clk_bF$buf38),
    .D(_4228_),
    .Q(\genblk1[5].u_ce.Xin12b [11])
);

DFFPOSX1 _12575_ (
    .CLK(clk_bF$buf37),
    .D(_4229_),
    .Q(\genblk1[5].u_ce.Xin12b [8])
);

DFFPOSX1 _12576_ (
    .CLK(clk_bF$buf36),
    .D(_4230_),
    .Q(\genblk1[5].u_ce.Xin12b [9])
);

DFFPOSX1 _12577_ (
    .CLK(clk_bF$buf35),
    .D(_4231_),
    .Q(\genblk1[5].u_ce.Xin12b [6])
);

DFFPOSX1 _12578_ (
    .CLK(clk_bF$buf34),
    .D(_4232_),
    .Q(\genblk1[5].u_ce.Xin12b [7])
);

DFFPOSX1 _12579_ (
    .CLK(clk_bF$buf33),
    .D(_4233_),
    .Q(\genblk1[5].u_ce.Xin12b [4])
);

DFFPOSX1 _12580_ (
    .CLK(clk_bF$buf32),
    .D(_4234_),
    .Q(\genblk1[5].u_ce.Xin12b [5])
);

DFFPOSX1 _12581_ (
    .CLK(clk_bF$buf31),
    .D(_4235_),
    .Q(\genblk1[5].u_ce.Xin1 [0])
);

DFFPOSX1 _12582_ (
    .CLK(clk_bF$buf30),
    .D(_4236_),
    .Q(\genblk1[5].u_ce.Xin1 [1])
);

DFFPOSX1 _12583_ (
    .CLK(clk_bF$buf29),
    .D(_4237_),
    .Q(\genblk1[5].u_ce.Xin0 [0])
);

DFFPOSX1 _12584_ (
    .CLK(clk_bF$buf28),
    .D(_4238_),
    .Q(\genblk1[5].u_ce.Xin0 [1])
);

DFFPOSX1 _12585_ (
    .CLK(clk_bF$buf27),
    .D(_4239_),
    .Q(\genblk1[5].u_ce.Yin12b [10])
);

DFFPOSX1 _12586_ (
    .CLK(clk_bF$buf26),
    .D(_4240_),
    .Q(\genblk1[5].u_ce.Yin12b [11])
);

DFFPOSX1 _12587_ (
    .CLK(clk_bF$buf25),
    .D(_4241_),
    .Q(\genblk1[5].u_ce.Yin12b [8])
);

DFFPOSX1 _12588_ (
    .CLK(clk_bF$buf24),
    .D(_4242_),
    .Q(\genblk1[5].u_ce.Yin12b [9])
);

DFFPOSX1 _12589_ (
    .CLK(clk_bF$buf23),
    .D(_4243_),
    .Q(\genblk1[5].u_ce.Yin12b [6])
);

DFFPOSX1 _12590_ (
    .CLK(clk_bF$buf22),
    .D(_4244_),
    .Q(\genblk1[5].u_ce.Yin12b [7])
);

DFFPOSX1 _12591_ (
    .CLK(clk_bF$buf21),
    .D(_4245_),
    .Q(\genblk1[5].u_ce.Yin12b [4])
);

DFFPOSX1 _12592_ (
    .CLK(clk_bF$buf20),
    .D(_4246_),
    .Q(\genblk1[5].u_ce.Yin12b [5])
);

DFFPOSX1 _12593_ (
    .CLK(clk_bF$buf19),
    .D(_4247_),
    .Q(\genblk1[5].u_ce.Yin1 [0])
);

DFFPOSX1 _12594_ (
    .CLK(clk_bF$buf18),
    .D(_4248_),
    .Q(\genblk1[5].u_ce.Yin1 [1])
);

DFFPOSX1 _12595_ (
    .CLK(clk_bF$buf17),
    .D(_4249_),
    .Q(\genblk1[5].u_ce.Yin0 [0])
);

DFFPOSX1 _12596_ (
    .CLK(clk_bF$buf16),
    .D(_4250_),
    .Q(\genblk1[5].u_ce.Yin0 [1])
);

DFFPOSX1 _12597_ (
    .CLK(clk_bF$buf15),
    .D(_4251_),
    .Q(\genblk1[5].u_ce.Ain12b [10])
);

DFFPOSX1 _12598_ (
    .CLK(clk_bF$buf14),
    .D(_4252_),
    .Q(\genblk1[5].u_ce.Ain12b [11])
);

DFFPOSX1 _12599_ (
    .CLK(clk_bF$buf13),
    .D(_4253_),
    .Q(\genblk1[5].u_ce.Ain12b [8])
);

DFFPOSX1 _12600_ (
    .CLK(clk_bF$buf12),
    .D(_4254_),
    .Q(\genblk1[5].u_ce.Ain12b [9])
);

DFFPOSX1 _12601_ (
    .CLK(clk_bF$buf11),
    .D(_4255_),
    .Q(\genblk1[5].u_ce.Ain12b [6])
);

DFFPOSX1 _12602_ (
    .CLK(clk_bF$buf10),
    .D(_4256_),
    .Q(\genblk1[5].u_ce.Ain12b [7])
);

DFFPOSX1 _12603_ (
    .CLK(clk_bF$buf9),
    .D(_4257_),
    .Q(\genblk1[5].u_ce.Ain12b [4])
);

DFFPOSX1 _12604_ (
    .CLK(clk_bF$buf8),
    .D(_4258_),
    .Q(\genblk1[5].u_ce.Ain12b [5])
);

DFFPOSX1 _12605_ (
    .CLK(clk_bF$buf7),
    .D(_4259_),
    .Q(\genblk1[5].u_ce.Ain1 [0])
);

DFFPOSX1 _12606_ (
    .CLK(clk_bF$buf6),
    .D(_4260_),
    .Q(\genblk1[5].u_ce.Ain1 [1])
);

DFFPOSX1 _12607_ (
    .CLK(clk_bF$buf5),
    .D(_4261_),
    .Q(\genblk1[5].u_ce.Ain0 [0])
);

DFFPOSX1 _12608_ (
    .CLK(clk_bF$buf4),
    .D(_4262_),
    .Q(\genblk1[5].u_ce.Ain0 [1])
);

DFFPOSX1 _12609_ (
    .CLK(clk_bF$buf3),
    .D(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[5].u_ce.LoadCtl [0])
);

DFFPOSX1 _12610_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[5].u_ce.LoadCtl [1])
);

DFFPOSX1 _12611_ (
    .CLK(clk_bF$buf1),
    .D(\genblk1[5].u_ce.LoadCtl [1]),
    .Q(\genblk1[5].u_ce.LoadCtl [2])
);

DFFPOSX1 _12612_ (
    .CLK(clk_bF$buf0),
    .D(\genblk1[5].u_ce.LoadCtl [2]),
    .Q(\genblk1[5].u_ce.LoadCtl [3])
);

DFFPOSX1 _12613_ (
    .CLK(clk_bF$buf78),
    .D(\genblk1[5].u_ce.LoadCtl [3]),
    .Q(\genblk1[5].u_ce.LoadCtl [4])
);

DFFPOSX1 _12614_ (
    .CLK(clk_bF$buf77),
    .D(\genblk1[5].u_ce.LoadCtl [4]),
    .Q(\genblk1[5].u_ce.LoadCtl [5])
);

DFFPOSX1 _12615_ (
    .CLK(clk_bF$buf76),
    .D(\genblk1[5].u_ce.LoadCtl [5]),
    .Q(\genblk1[5].u_ce.Vld )
);

INVX2 _12616_ (
    .A(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5102_)
);

NOR2X1 _12617_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .Y(_5103_)
);

INVX2 _12618_ (
    .A(_5103_),
    .Y(_5104_)
);

INVX4 _12619_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .Y(_5105_)
);

NOR2X1 _12620_ (
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .B(\genblk1[6].u_ce.LoadCtl [3]),
    .Y(_5106_)
);

INVX2 _12621_ (
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5107_)
);

AND2X2 _12622_ (
    .A(_5107_),
    .B(\genblk1[6].u_ce.LoadCtl [3]),
    .Y(_5108_)
);

NOR2X1 _12623_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5109_)
);

INVX1 _12624_ (
    .A(\genblk1[6].u_ce.Acalc [9]),
    .Y(_5110_)
);

OAI21X1 _12625_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Acalc [11]),
    .C(_5106_),
    .Y(_5111_)
);

AOI21X1 _12626_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5110_),
    .C(_5111_),
    .Y(_5112_)
);

INVX1 _12627_ (
    .A(\genblk1[6].u_ce.Acalc [5]),
    .Y(_5113_)
);

NAND2X1 _12628_ (
    .A(\genblk1[6].u_ce.Acalc [7]),
    .B(_5108_),
    .Y(_5114_)
);

OAI21X1 _12629_ (
    .A(_5107_),
    .B(_5113_),
    .C(_5114_),
    .Y(_5115_)
);

OAI21X1 _12630_ (
    .A(_5112_),
    .B(_5115_),
    .C(_5109_),
    .Y(_5116_)
);

AOI22X1 _12631_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Acalc [1]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Acalc [3]),
    .Y(_5117_)
);

NAND2X1 _12632_ (
    .A(_5117_),
    .B(_5116_),
    .Y(\a[7] [1])
);

INVX1 _12633_ (
    .A(\genblk1[6].u_ce.Ycalc [10]),
    .Y(_5118_)
);

OAI21X1 _12634_ (
    .A(_5105_),
    .B(\genblk1[6].u_ce.Ycalc [8]),
    .C(_5106_),
    .Y(_5119_)
);

AOI21X1 _12635_ (
    .A(_5105_),
    .B(_5118_),
    .C(_5119_),
    .Y(_5120_)
);

INVX1 _12636_ (
    .A(\genblk1[6].u_ce.Ycalc [4]),
    .Y(_5121_)
);

NAND2X1 _12637_ (
    .A(\genblk1[6].u_ce.Ycalc [6]),
    .B(_5108_),
    .Y(_5122_)
);

OAI21X1 _12638_ (
    .A(_5107_),
    .B(_5121_),
    .C(_5122_),
    .Y(_5123_)
);

OAI21X1 _12639_ (
    .A(_5120_),
    .B(_5123_),
    .C(_5109_),
    .Y(_5124_)
);

AOI22X1 _12640_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Ycalc [0]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Ycalc [2]),
    .Y(_5125_)
);

NAND2X1 _12641_ (
    .A(_5125_),
    .B(_5124_),
    .Y(\genblk1[6].u_ce.Y_ [0])
);

INVX1 _12642_ (
    .A(\genblk1[6].u_ce.Ycalc [9]),
    .Y(_5126_)
);

OAI21X1 _12643_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Ycalc [11]),
    .C(_5106_),
    .Y(_5127_)
);

AOI21X1 _12644_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5126_),
    .C(_5127_),
    .Y(_5128_)
);

INVX1 _12645_ (
    .A(\genblk1[6].u_ce.Ycalc [5]),
    .Y(_5129_)
);

NAND2X1 _12646_ (
    .A(\genblk1[6].u_ce.Ycalc [7]),
    .B(_5108_),
    .Y(_5130_)
);

OAI21X1 _12647_ (
    .A(_5107_),
    .B(_5129_),
    .C(_5130_),
    .Y(_5131_)
);

OAI21X1 _12648_ (
    .A(_5128_),
    .B(_5131_),
    .C(_5109_),
    .Y(_5132_)
);

AOI22X1 _12649_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[6].u_ce.Ycalc [1]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5133_)
);

NAND2X1 _12650_ (
    .A(_5133_),
    .B(_5132_),
    .Y(\genblk1[6].u_ce.Y_ [1])
);

INVX1 _12651_ (
    .A(\genblk1[6].u_ce.Xcalc [8]),
    .Y(_5134_)
);

OAI21X1 _12652_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Xcalc [10]),
    .C(_5106_),
    .Y(_5135_)
);

AOI21X1 _12653_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5134_),
    .C(_5135_),
    .Y(_5136_)
);

INVX1 _12654_ (
    .A(\genblk1[6].u_ce.Xcalc [4]),
    .Y(_5137_)
);

NAND2X1 _12655_ (
    .A(\genblk1[6].u_ce.Xcalc [6]),
    .B(_5108_),
    .Y(_5138_)
);

OAI21X1 _12656_ (
    .A(_5107_),
    .B(_5137_),
    .C(_5138_),
    .Y(_5139_)
);

OAI21X1 _12657_ (
    .A(_5136_),
    .B(_5139_),
    .C(_5109_),
    .Y(_5140_)
);

AOI22X1 _12658_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[6].u_ce.Xcalc [0]),
    .C(_5103_),
    .D(\genblk1[6].u_ce.Xcalc [2]),
    .Y(_5141_)
);

NAND2X1 _12659_ (
    .A(_5141_),
    .B(_5140_),
    .Y(\genblk1[6].u_ce.X_ [0])
);

INVX1 _12660_ (
    .A(\genblk1[6].u_ce.Xcalc [3]),
    .Y(_5142_)
);

NOR2X1 _12661_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Xcalc [11]),
    .Y(_5143_)
);

OAI21X1 _12662_ (
    .A(_5105_),
    .B(\genblk1[6].u_ce.Xcalc [9]),
    .C(_5106_),
    .Y(_5144_)
);

AOI22X1 _12663_ (
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .B(\genblk1[6].u_ce.Xcalc [5]),
    .C(_5108_),
    .D(\genblk1[6].u_ce.Xcalc [7]),
    .Y(_5145_)
);

OAI21X1 _12664_ (
    .A(_5143_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5146_)
);

AOI22X1 _12665_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.Xcalc [1]),
    .C(_5146_),
    .D(_5109_),
    .Y(_5147_)
);

OAI21X1 _12666_ (
    .A(_5142_),
    .B(_5104_),
    .C(_5147_),
    .Y(\genblk1[6].u_ce.X_ [1])
);

INVX1 _12667_ (
    .A(\genblk1[6].u_ce.Ycalc [0]),
    .Y(_5148_)
);

INVX1 _12668_ (
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .Y(_5149_)
);

INVX8 _12669_ (
    .A(1'h1),
    .Y(_5150_)
);

INVX8 _12670_ (
    .A(1'h1),
    .Y(_5151_)
);

INVX1 _12671_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5152_)
);

NAND2X1 _12672_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5153_)
);

OAI21X1 _12673_ (
    .A(1'h0),
    .B(_5152_),
    .C(_5153_),
    .Y(_5154_)
);

INVX1 _12674_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .Y(_5155_)
);

NAND2X1 _12675_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5156_)
);

OAI21X1 _12676_ (
    .A(1'h0),
    .B(_5155_),
    .C(_5156_),
    .Y(_5157_)
);

MUX2X1 _12677_ (
    .A(_5157_),
    .B(_5154_),
    .S(_5151__bF$buf4),
    .Y(_5158_)
);

INVX1 _12678_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5159_)
);

NAND2X1 _12679_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5160_)
);

OAI21X1 _12680_ (
    .A(1'h0),
    .B(_5159_),
    .C(_5160_),
    .Y(_5161_)
);

INVX1 _12681_ (
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .Y(_5162_)
);

NAND2X1 _12682_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_5163_)
);

OAI21X1 _12683_ (
    .A(1'h0),
    .B(_5162_),
    .C(_5163_),
    .Y(_5164_)
);

MUX2X1 _12684_ (
    .A(_5164_),
    .B(_5161_),
    .S(_5151__bF$buf3),
    .Y(_5165_)
);

MUX2X1 _12685_ (
    .A(_5165_),
    .B(_5158_),
    .S(_5150__bF$buf4),
    .Y(_5166_)
);

NOR2X1 _12686_ (
    .A(_5149_),
    .B(_5166_),
    .Y(_5167_)
);

NAND2X1 _12687_ (
    .A(_5149_),
    .B(_5166_),
    .Y(_5168_)
);

INVX1 _12688_ (
    .A(_5168_),
    .Y(_5169_)
);

NAND2X1 _12689_ (
    .A(_5150__bF$buf3),
    .B(_5151__bF$buf2),
    .Y(_5170_)
);

OAI21X1 _12690_ (
    .A(1'h0),
    .B(_5170_),
    .C(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .Y(_5171_)
);

INVX2 _12691_ (
    .A(_5171_),
    .Y(_5172_)
);

OAI21X1 _12692_ (
    .A(_5167_),
    .B(_5169_),
    .C(_5172_),
    .Y(_5173_)
);

OAI21X1 _12693_ (
    .A(_5148_),
    .B(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .C(_5173_),
    .Y(_5028_)
);

INVX8 _12694_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .Y(_5174_)
);

NAND2X1 _12695_ (
    .A(\genblk1[6].u_ce.Ycalc [1]),
    .B(_5174__bF$buf4),
    .Y(_5175_)
);

NOR2X1 _12696_ (
    .A(1'h0),
    .B(_5170_),
    .Y(_5176_)
);

MUX2X1 _12697_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(\genblk1[6].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_5177_)
);

MUX2X1 _12698_ (
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .B(\genblk1[6].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_5178_)
);

MUX2X1 _12699_ (
    .A(_5178_),
    .B(_5177_),
    .S(_5151__bF$buf1),
    .Y(_5179_)
);

INVX2 _12700_ (
    .A(1'h0),
    .Y(_5180_)
);

NAND2X1 _12701_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(_5180_),
    .Y(_5181_)
);

AOI21X1 _12702_ (
    .A(_5181_),
    .B(_5160_),
    .C(_5151__bF$buf0),
    .Y(_5182_)
);

NAND3X1 _12703_ (
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .B(_5180_),
    .C(_5151__bF$buf4),
    .Y(_5183_)
);

NAND3X1 _12704_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(1'h0),
    .C(_5151__bF$buf3),
    .Y(_5184_)
);

NAND3X1 _12705_ (
    .A(_5150__bF$buf2),
    .B(_5184_),
    .C(_5183_),
    .Y(_5185_)
);

OAI22X1 _12706_ (
    .A(_5182_),
    .B(_5185_),
    .C(_5150__bF$buf1),
    .D(_5179_),
    .Y(_5186_)
);

INVX1 _12707_ (
    .A(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5187_)
);

INVX8 _12708_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_5188_)
);

INVX1 _12709_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5189_)
);

NAND2X1 _12710_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5190_)
);

OAI21X1 _12711_ (
    .A(1'h0),
    .B(_5189_),
    .C(_5190_),
    .Y(_5191_)
);

INVX1 _12712_ (
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5192_)
);

NAND2X1 _12713_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5193_)
);

OAI21X1 _12714_ (
    .A(1'h0),
    .B(_5192_),
    .C(_5193_),
    .Y(_5194_)
);

MUX2X1 _12715_ (
    .A(_5194_),
    .B(_5191_),
    .S(_5151__bF$buf2),
    .Y(_5195_)
);

INVX1 _12716_ (
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5196_)
);

NAND2X1 _12717_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [4]),
    .Y(_5197_)
);

OAI21X1 _12718_ (
    .A(1'h0),
    .B(_5196_),
    .C(_5197_),
    .Y(_5198_)
);

INVX1 _12719_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .Y(_5199_)
);

NAND2X1 _12720_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5200_)
);

OAI21X1 _12721_ (
    .A(1'h0),
    .B(_5199_),
    .C(_5200_),
    .Y(_5201_)
);

MUX2X1 _12722_ (
    .A(_5201_),
    .B(_5198_),
    .S(_5151__bF$buf1),
    .Y(_5202_)
);

MUX2X1 _12723_ (
    .A(_5202_),
    .B(_5195_),
    .S(_5150__bF$buf0),
    .Y(_5203_)
);

NAND3X1 _12724_ (
    .A(_5188__bF$buf5),
    .B(_5166_),
    .C(_5203_),
    .Y(_5204_)
);

MUX2X1 _12725_ (
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_5205_)
);

MUX2X1 _12726_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_5206_)
);

MUX2X1 _12727_ (
    .A(_5206_),
    .B(_5205_),
    .S(_5151__bF$buf0),
    .Y(_5207_)
);

MUX2X1 _12728_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_5208_)
);

MUX2X1 _12729_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(\genblk1[6].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_5209_)
);

MUX2X1 _12730_ (
    .A(_5209_),
    .B(_5208_),
    .S(_5151__bF$buf4),
    .Y(_5210_)
);

MUX2X1 _12731_ (
    .A(_5210_),
    .B(_5207_),
    .S(_5150__bF$buf4),
    .Y(_5211_)
);

OAI21X1 _12732_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5186_),
    .C(_5211_),
    .Y(_5212_)
);

AOI21X1 _12733_ (
    .A(_5212_),
    .B(_5204_),
    .C(_5187_),
    .Y(_5213_)
);

INVX1 _12734_ (
    .A(_5213_),
    .Y(_5214_)
);

NAND3X1 _12735_ (
    .A(_5187_),
    .B(_5204_),
    .C(_5212_),
    .Y(_5215_)
);

AND2X2 _12736_ (
    .A(_5214_),
    .B(_5215_),
    .Y(_5216_)
);

OAI21X1 _12737_ (
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .B(_5186_),
    .C(_5216_),
    .Y(_5217_)
);

OR2X2 _12738_ (
    .A(_5216_),
    .B(_5168_),
    .Y(_5218_)
);

AOI21X1 _12739_ (
    .A(_5218_),
    .B(_5217_),
    .C(_5176_),
    .Y(_5219_)
);

OAI21X1 _12740_ (
    .A(_5174__bF$buf3),
    .B(_5219_),
    .C(_5175_),
    .Y(_5029_)
);

INVX1 _12741_ (
    .A(\genblk1[6].u_ce.ISout ),
    .Y(_5220_)
);

NAND2X1 _12742_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .B(\genblk1[5].u_ce.ISout ),
    .Y(_5221_)
);

OAI21X1 _12743_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .B(_5220_),
    .C(_5221_),
    .Y(_5030_)
);

NAND2X1 _12744_ (
    .A(\genblk1[6].u_ce.Ycalc [2]),
    .B(_5174__bF$buf2),
    .Y(_5222_)
);

AOI21X1 _12745_ (
    .A(_5168_),
    .B(_5215_),
    .C(_5213_),
    .Y(_5223_)
);

MUX2X1 _12746_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(\genblk1[6].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_5224_)
);

MUX2X1 _12747_ (
    .A(_5224_),
    .B(_5177_),
    .S(1'h1),
    .Y(_5225_)
);

MUX2X1 _12748_ (
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_5226_)
);

NAND2X1 _12749_ (
    .A(1'h1),
    .B(_5150__bF$buf3),
    .Y(_5227_)
);

OAI22X1 _12750_ (
    .A(_5227_),
    .B(_5178_),
    .C(_5226_),
    .D(_5170_),
    .Y(_5228_)
);

AOI21X1 _12751_ (
    .A(1'h1),
    .B(_5225_),
    .C(_5228_),
    .Y(_5229_)
);

AOI21X1 _12752_ (
    .A(_5211_),
    .B(_5186_),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5230_)
);

NAND2X1 _12753_ (
    .A(_5229_),
    .B(_5230_),
    .Y(_5231_)
);

INVX1 _12754_ (
    .A(_5229_),
    .Y(_5232_)
);

OAI21X1 _12755_ (
    .A(_5166_),
    .B(_5203_),
    .C(_5188__bF$buf4),
    .Y(_5233_)
);

NAND2X1 _12756_ (
    .A(_5232_),
    .B(_5233_),
    .Y(_5234_)
);

AOI21X1 _12757_ (
    .A(_5234_),
    .B(_5231_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5235_)
);

NAND3X1 _12758_ (
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .B(_5231_),
    .C(_5234_),
    .Y(_5236_)
);

INVX1 _12759_ (
    .A(_5236_),
    .Y(_5237_)
);

OR2X2 _12760_ (
    .A(_5237_),
    .B(_5235_),
    .Y(_5238_)
);

NOR2X1 _12761_ (
    .A(_5223_),
    .B(_5238_),
    .Y(_5239_)
);

INVX1 _12762_ (
    .A(_5239_),
    .Y(_5240_)
);

OAI21X1 _12763_ (
    .A(_5235_),
    .B(_5237_),
    .C(_5223_),
    .Y(_5241_)
);

AOI21X1 _12764_ (
    .A(_5240_),
    .B(_5241_),
    .C(_5176_),
    .Y(_5242_)
);

INVX2 _12765_ (
    .A(_5176_),
    .Y(_5243_)
);

OAI21X1 _12766_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5243_),
    .C(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .Y(_5244_)
);

OAI21X1 _12767_ (
    .A(_5244_),
    .B(_5242_),
    .C(_5222_),
    .Y(_5031_)
);

INVX1 _12768_ (
    .A(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5245_)
);

INVX2 _12769_ (
    .A(_5244_),
    .Y(_5246_)
);

OAI21X1 _12770_ (
    .A(_5235_),
    .B(_5223_),
    .C(_5236_),
    .Y(_5247_)
);

INVX1 _12771_ (
    .A(_5247_),
    .Y(_5248_)
);

INVX1 _12772_ (
    .A(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5249_)
);

NAND3X1 _12773_ (
    .A(_5186_),
    .B(_5211_),
    .C(_5229_),
    .Y(_5250_)
);

INVX1 _12774_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .Y(_5251_)
);

NAND2X1 _12775_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5252_)
);

OAI21X1 _12776_ (
    .A(1'h0),
    .B(_5251_),
    .C(_5252_),
    .Y(_5253_)
);

NAND2X1 _12777_ (
    .A(_5151__bF$buf3),
    .B(_5205_),
    .Y(_5254_)
);

OAI21X1 _12778_ (
    .A(_5151__bF$buf2),
    .B(_5253_),
    .C(_5254_),
    .Y(_5255_)
);

NOR2X1 _12779_ (
    .A(1'h1),
    .B(_5151__bF$buf1),
    .Y(_5256_)
);

NOR2X1 _12780_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_5257_)
);

AOI22X1 _12781_ (
    .A(_5198_),
    .B(_5257_),
    .C(_5256_),
    .D(_5194_),
    .Y(_5258_)
);

OAI21X1 _12782_ (
    .A(_5150__bF$buf2),
    .B(_5255_),
    .C(_5258_),
    .Y(_5259_)
);

NAND3X1 _12783_ (
    .A(_5188__bF$buf3),
    .B(_5259_),
    .C(_5250_),
    .Y(_5260_)
);

INVX1 _12784_ (
    .A(_5250_),
    .Y(_5261_)
);

INVX1 _12785_ (
    .A(_5259_),
    .Y(_5262_)
);

OAI21X1 _12786_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5261_),
    .C(_5262_),
    .Y(_5263_)
);

NAND3X1 _12787_ (
    .A(_5249_),
    .B(_5260_),
    .C(_5263_),
    .Y(_5264_)
);

AOI21X1 _12788_ (
    .A(_5263_),
    .B(_5260_),
    .C(_5249_),
    .Y(_5265_)
);

INVX1 _12789_ (
    .A(_5265_),
    .Y(_5266_)
);

NAND2X1 _12790_ (
    .A(_5264_),
    .B(_5266_),
    .Y(_5267_)
);

AOI21X1 _12791_ (
    .A(_5267_),
    .B(_5248_),
    .C(_5176_),
    .Y(_5268_)
);

OAI21X1 _12792_ (
    .A(_5248_),
    .B(_5267_),
    .C(_5268_),
    .Y(_5269_)
);

AOI22X1 _12793_ (
    .A(_5245_),
    .B(_5174__bF$buf1),
    .C(_5269_),
    .D(_5246_),
    .Y(_5032_)
);

AOI21X1 _12794_ (
    .A(_5247_),
    .B(_5264_),
    .C(_5265_),
    .Y(_5270_)
);

INVX1 _12795_ (
    .A(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5271_)
);

INVX1 _12796_ (
    .A(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5272_)
);

NAND2X1 _12797_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5273_)
);

OAI21X1 _12798_ (
    .A(1'h0),
    .B(_5272_),
    .C(_5273_),
    .Y(_5274_)
);

NAND2X1 _12799_ (
    .A(_5151__bF$buf0),
    .B(_5224_),
    .Y(_5275_)
);

OAI21X1 _12800_ (
    .A(_5151__bF$buf4),
    .B(_5274_),
    .C(_5275_),
    .Y(_5276_)
);

NAND2X1 _12801_ (
    .A(_5150__bF$buf1),
    .B(_5179_),
    .Y(_5277_)
);

OAI21X1 _12802_ (
    .A(_5150__bF$buf0),
    .B(_5276_),
    .C(_5277_),
    .Y(_5278_)
);

INVX2 _12803_ (
    .A(_5278_),
    .Y(_5279_)
);

OAI21X1 _12804_ (
    .A(_5259_),
    .B(_5250_),
    .C(_5188__bF$buf2),
    .Y(_5280_)
);

OR2X2 _12805_ (
    .A(_5280_),
    .B(_5279_),
    .Y(_5281_)
);

NOR2X1 _12806_ (
    .A(_5259_),
    .B(_5250_),
    .Y(_5282_)
);

OAI21X1 _12807_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5282_),
    .C(_5279_),
    .Y(_5283_)
);

NAND3X1 _12808_ (
    .A(_5271_),
    .B(_5283_),
    .C(_5281_),
    .Y(_5284_)
);

NOR2X1 _12809_ (
    .A(_5279_),
    .B(_5280_),
    .Y(_5285_)
);

AND2X2 _12810_ (
    .A(_5280_),
    .B(_5279_),
    .Y(_5286_)
);

OAI21X1 _12811_ (
    .A(_5285_),
    .B(_5286_),
    .C(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5287_)
);

NAND2X1 _12812_ (
    .A(_5287_),
    .B(_5284_),
    .Y(_5288_)
);

AOI21X1 _12813_ (
    .A(_5270_),
    .B(_5288_),
    .C(_5176_),
    .Y(_5289_)
);

OAI21X1 _12814_ (
    .A(_5270_),
    .B(_5288_),
    .C(_5289_),
    .Y(_5290_)
);

AOI22X1 _12815_ (
    .A(_5121_),
    .B(_5174__bF$buf0),
    .C(_5290_),
    .D(_5246_),
    .Y(_5033_)
);

OAI21X1 _12816_ (
    .A(_5288_),
    .B(_5270_),
    .C(_5287_),
    .Y(_5291_)
);

INVX1 _12817_ (
    .A(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5292_)
);

NAND3X1 _12818_ (
    .A(_5262_),
    .B(_5279_),
    .C(_5261_),
    .Y(_5293_)
);

NAND2X1 _12819_ (
    .A(1'h1),
    .B(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5294_)
);

INVX1 _12820_ (
    .A(_5294_),
    .Y(_5295_)
);

AOI21X1 _12821_ (
    .A(_5253_),
    .B(_5151__bF$buf3),
    .C(_5295_),
    .Y(_5296_)
);

NAND2X1 _12822_ (
    .A(_5150__bF$buf4),
    .B(_5207_),
    .Y(_5297_)
);

OAI21X1 _12823_ (
    .A(_5150__bF$buf3),
    .B(_5296_),
    .C(_5297_),
    .Y(_5298_)
);

NAND3X1 _12824_ (
    .A(_5188__bF$buf1),
    .B(_5298_),
    .C(_5293_),
    .Y(_5299_)
);

NOR3X1 _12825_ (
    .A(_5259_),
    .B(_5278_),
    .C(_5250_),
    .Y(_5300_)
);

INVX1 _12826_ (
    .A(_5298_),
    .Y(_5301_)
);

OAI21X1 _12827_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5300_),
    .C(_5301_),
    .Y(_5302_)
);

NAND3X1 _12828_ (
    .A(_5292_),
    .B(_5299_),
    .C(_5302_),
    .Y(_5303_)
);

AOI21X1 _12829_ (
    .A(_5302_),
    .B(_5299_),
    .C(_5292_),
    .Y(_5304_)
);

INVX1 _12830_ (
    .A(_5304_),
    .Y(_5305_)
);

NAND2X1 _12831_ (
    .A(_5303_),
    .B(_5305_),
    .Y(_5306_)
);

AND2X2 _12832_ (
    .A(_5291_),
    .B(_5306_),
    .Y(_5307_)
);

OAI21X1 _12833_ (
    .A(_5306_),
    .B(_5291_),
    .C(_5243_),
    .Y(_5308_)
);

OAI21X1 _12834_ (
    .A(_5308_),
    .B(_5307_),
    .C(_5246_),
    .Y(_5309_)
);

OAI21X1 _12835_ (
    .A(_5129_),
    .B(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .C(_5309_),
    .Y(_5034_)
);

INVX1 _12836_ (
    .A(\genblk1[6].u_ce.Ycalc [6]),
    .Y(_5310_)
);

INVX1 _12837_ (
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5311_)
);

NAND3X1 _12838_ (
    .A(_5279_),
    .B(_5301_),
    .C(_5282_),
    .Y(_5312_)
);

AOI21X1 _12839_ (
    .A(_5274_),
    .B(_5151__bF$buf2),
    .C(_5295_),
    .Y(_5313_)
);

NAND2X1 _12840_ (
    .A(_5150__bF$buf2),
    .B(_5225_),
    .Y(_5314_)
);

OAI21X1 _12841_ (
    .A(_5150__bF$buf1),
    .B(_5313_),
    .C(_5314_),
    .Y(_5315_)
);

NAND3X1 _12842_ (
    .A(_5188__bF$buf0),
    .B(_5315_),
    .C(_5312_),
    .Y(_5316_)
);

INVX1 _12843_ (
    .A(_5315_),
    .Y(_5317_)
);

OAI21X1 _12844_ (
    .A(_5298_),
    .B(_5293_),
    .C(_5188__bF$buf5),
    .Y(_5318_)
);

NAND2X1 _12845_ (
    .A(_5317_),
    .B(_5318_),
    .Y(_5319_)
);

NAND3X1 _12846_ (
    .A(_5311_),
    .B(_5316_),
    .C(_5319_),
    .Y(_5320_)
);

NAND3X1 _12847_ (
    .A(_5188__bF$buf4),
    .B(_5317_),
    .C(_5312_),
    .Y(_5321_)
);

NAND2X1 _12848_ (
    .A(_5315_),
    .B(_5318_),
    .Y(_5322_)
);

NAND3X1 _12849_ (
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .B(_5321_),
    .C(_5322_),
    .Y(_5323_)
);

NAND2X1 _12850_ (
    .A(_5320_),
    .B(_5323_),
    .Y(_5324_)
);

AOI21X1 _12851_ (
    .A(_5281_),
    .B(_5283_),
    .C(_5271_),
    .Y(_5325_)
);

NOR2X1 _12852_ (
    .A(_5325_),
    .B(_5304_),
    .Y(_5326_)
);

OAI21X1 _12853_ (
    .A(_5288_),
    .B(_5270_),
    .C(_5326_),
    .Y(_5327_)
);

NAND2X1 _12854_ (
    .A(_5303_),
    .B(_5327_),
    .Y(_5328_)
);

AOI21X1 _12855_ (
    .A(_5328_),
    .B(_5324_),
    .C(_5176_),
    .Y(_5329_)
);

OAI21X1 _12856_ (
    .A(_5324_),
    .B(_5328_),
    .C(_5329_),
    .Y(_5330_)
);

AOI22X1 _12857_ (
    .A(_5310_),
    .B(_5174__bF$buf4),
    .C(_5330_),
    .D(_5246_),
    .Y(_5035_)
);

INVX1 _12858_ (
    .A(\genblk1[6].u_ce.Ycalc [7]),
    .Y(_5331_)
);

AOI21X1 _12859_ (
    .A(_5319_),
    .B(_5316_),
    .C(_5311_),
    .Y(_5332_)
);

AND2X2 _12860_ (
    .A(_5284_),
    .B(_5287_),
    .Y(_5333_)
);

NAND3X1 _12861_ (
    .A(_5303_),
    .B(_5305_),
    .C(_5333_),
    .Y(_5334_)
);

AOI21X1 _12862_ (
    .A(_5325_),
    .B(_5303_),
    .C(_5304_),
    .Y(_5335_)
);

OAI21X1 _12863_ (
    .A(_5270_),
    .B(_5334_),
    .C(_5335_),
    .Y(_5336_)
);

AOI21X1 _12864_ (
    .A(_5336_),
    .B(_5320_),
    .C(_5332_),
    .Y(_5337_)
);

INVX1 _12865_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5338_)
);

NAND3X1 _12866_ (
    .A(_5301_),
    .B(_5317_),
    .C(_5300_),
    .Y(_5339_)
);

INVX1 _12867_ (
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5340_)
);

NOR2X1 _12868_ (
    .A(_5150__bF$buf0),
    .B(_5340_),
    .Y(_5341_)
);

INVX1 _12869_ (
    .A(_5341_),
    .Y(_5342_)
);

OAI21X1 _12870_ (
    .A(1'h1),
    .B(_5255_),
    .C(_5342_),
    .Y(_5343_)
);

NAND3X1 _12871_ (
    .A(_5188__bF$buf3),
    .B(_5343_),
    .C(_5339_),
    .Y(_5344_)
);

INVX1 _12872_ (
    .A(_5343_),
    .Y(_5345_)
);

OAI21X1 _12873_ (
    .A(_5315_),
    .B(_5312_),
    .C(_5188__bF$buf2),
    .Y(_5346_)
);

NAND2X1 _12874_ (
    .A(_5345_),
    .B(_5346_),
    .Y(_5347_)
);

NAND3X1 _12875_ (
    .A(_5338_),
    .B(_5344_),
    .C(_5347_),
    .Y(_5348_)
);

NAND3X1 _12876_ (
    .A(_5188__bF$buf1),
    .B(_5345_),
    .C(_5339_),
    .Y(_5349_)
);

NAND2X1 _12877_ (
    .A(_5343_),
    .B(_5346_),
    .Y(_5350_)
);

NAND3X1 _12878_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(_5349_),
    .C(_5350_),
    .Y(_5351_)
);

NAND2X1 _12879_ (
    .A(_5348_),
    .B(_5351_),
    .Y(_5352_)
);

INVX1 _12880_ (
    .A(_5352_),
    .Y(_5353_)
);

NOR2X1 _12881_ (
    .A(_5353_),
    .B(_5337_),
    .Y(_5354_)
);

OAI21X1 _12882_ (
    .A(_5324_),
    .B(_5328_),
    .C(_5323_),
    .Y(_5355_)
);

OAI21X1 _12883_ (
    .A(_5352_),
    .B(_5355_),
    .C(_5243_),
    .Y(_5356_)
);

OAI21X1 _12884_ (
    .A(_5188__bF$buf0),
    .B(_5243_),
    .C(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .Y(_5357_)
);

INVX1 _12885_ (
    .A(_5357_),
    .Y(_5358_)
);

OAI21X1 _12886_ (
    .A(_5356_),
    .B(_5354_),
    .C(_5358_),
    .Y(_5359_)
);

OAI21X1 _12887_ (
    .A(_5331_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5359_),
    .Y(_5036_)
);

INVX1 _12888_ (
    .A(\genblk1[6].u_ce.Ycalc [8]),
    .Y(_5360_)
);

OAI21X1 _12889_ (
    .A(_5323_),
    .B(_5352_),
    .C(_5351_),
    .Y(_5361_)
);

NOR2X1 _12890_ (
    .A(_5324_),
    .B(_5352_),
    .Y(_5362_)
);

AOI21X1 _12891_ (
    .A(_5362_),
    .B(_5336_),
    .C(_5361_),
    .Y(_5363_)
);

INVX1 _12892_ (
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5364_)
);

OR2X2 _12893_ (
    .A(_5339_),
    .B(_5343_),
    .Y(_5365_)
);

OAI21X1 _12894_ (
    .A(1'h1),
    .B(_5276_),
    .C(_5342_),
    .Y(_5366_)
);

NAND3X1 _12895_ (
    .A(_5188__bF$buf5),
    .B(_5366_),
    .C(_5365_),
    .Y(_5367_)
);

NOR2X1 _12896_ (
    .A(_5343_),
    .B(_5339_),
    .Y(_5368_)
);

INVX1 _12897_ (
    .A(_5366_),
    .Y(_5369_)
);

OAI21X1 _12898_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5368_),
    .C(_5369_),
    .Y(_5370_)
);

NAND3X1 _12899_ (
    .A(_5364_),
    .B(_5370_),
    .C(_5367_),
    .Y(_5371_)
);

NAND3X1 _12900_ (
    .A(_5188__bF$buf4),
    .B(_5369_),
    .C(_5365_),
    .Y(_5372_)
);

OAI21X1 _12901_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5368_),
    .C(_5366_),
    .Y(_5373_)
);

NAND3X1 _12902_ (
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .B(_5373_),
    .C(_5372_),
    .Y(_5374_)
);

AND2X2 _12903_ (
    .A(_5371_),
    .B(_5374_),
    .Y(_5375_)
);

INVX1 _12904_ (
    .A(_5375_),
    .Y(_5376_)
);

AOI21X1 _12905_ (
    .A(_5363_),
    .B(_5376_),
    .C(_5176_),
    .Y(_5377_)
);

OAI21X1 _12906_ (
    .A(_5363_),
    .B(_5376_),
    .C(_5377_),
    .Y(_5378_)
);

AOI22X1 _12907_ (
    .A(_5360_),
    .B(_5174__bF$buf3),
    .C(_5378_),
    .D(_5358_),
    .Y(_5037_)
);

NAND2X1 _12908_ (
    .A(_5332_),
    .B(_5348_),
    .Y(_5379_)
);

AND2X2 _12909_ (
    .A(_5379_),
    .B(_5351_),
    .Y(_5380_)
);

AND2X2 _12910_ (
    .A(_5320_),
    .B(_5323_),
    .Y(_5381_)
);

NAND3X1 _12911_ (
    .A(_5348_),
    .B(_5351_),
    .C(_5381_),
    .Y(_5382_)
);

OAI21X1 _12912_ (
    .A(_5328_),
    .B(_5382_),
    .C(_5380_),
    .Y(_5383_)
);

INVX1 _12913_ (
    .A(_5374_),
    .Y(_5384_)
);

AOI21X1 _12914_ (
    .A(_5383_),
    .B(_5371_),
    .C(_5384_),
    .Y(_5385_)
);

INVX1 _12915_ (
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5386_)
);

NOR3X1 _12916_ (
    .A(_5343_),
    .B(_5366_),
    .C(_5339_),
    .Y(_5387_)
);

INVX1 _12917_ (
    .A(_5387_),
    .Y(_5388_)
);

OAI21X1 _12918_ (
    .A(1'h1),
    .B(_5296_),
    .C(_5342_),
    .Y(_5389_)
);

NAND3X1 _12919_ (
    .A(_5188__bF$buf3),
    .B(_5389_),
    .C(_5388_),
    .Y(_5390_)
);

INVX1 _12920_ (
    .A(_5389_),
    .Y(_5391_)
);

OAI21X1 _12921_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5387_),
    .C(_5391_),
    .Y(_5392_)
);

NAND3X1 _12922_ (
    .A(_5386_),
    .B(_5392_),
    .C(_5390_),
    .Y(_5393_)
);

NAND3X1 _12923_ (
    .A(_5188__bF$buf2),
    .B(_5391_),
    .C(_5388_),
    .Y(_5394_)
);

OAI21X1 _12924_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5387_),
    .C(_5389_),
    .Y(_5395_)
);

NAND3X1 _12925_ (
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .B(_5395_),
    .C(_5394_),
    .Y(_5396_)
);

AND2X2 _12926_ (
    .A(_5393_),
    .B(_5396_),
    .Y(_5397_)
);

AND2X2 _12927_ (
    .A(_5385_),
    .B(_5397_),
    .Y(_5398_)
);

OAI21X1 _12928_ (
    .A(_5397_),
    .B(_5385_),
    .C(_5243_),
    .Y(_5399_)
);

OAI21X1 _12929_ (
    .A(_5399_),
    .B(_5398_),
    .C(_5246_),
    .Y(_5400_)
);

OAI21X1 _12930_ (
    .A(_5126_),
    .B(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .C(_5400_),
    .Y(_5038_)
);

INVX1 _12931_ (
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .Y(_5401_)
);

OAI21X1 _12932_ (
    .A(1'h1),
    .B(_5313_),
    .C(_5342_),
    .Y(_5402_)
);

INVX1 _12933_ (
    .A(_5402_),
    .Y(_5403_)
);

AOI21X1 _12934_ (
    .A(_5387_),
    .B(_5391_),
    .C(_5403_),
    .Y(_5404_)
);

NAND3X1 _12935_ (
    .A(_5391_),
    .B(_5403_),
    .C(_5387_),
    .Y(_5405_)
);

NAND2X1 _12936_ (
    .A(_5188__bF$buf1),
    .B(_5405_),
    .Y(_5406_)
);

NAND2X1 _12937_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5402_),
    .Y(_5407_)
);

OAI21X1 _12938_ (
    .A(_5404_),
    .B(_5406_),
    .C(_5407_),
    .Y(_5408_)
);

NAND2X1 _12939_ (
    .A(_5401_),
    .B(_5408_),
    .Y(_5409_)
);

INVX1 _12940_ (
    .A(_5404_),
    .Y(_5410_)
);

AND2X2 _12941_ (
    .A(_5405_),
    .B(_5188__bF$buf0),
    .Y(_5411_)
);

NAND2X1 _12942_ (
    .A(_5410_),
    .B(_5411_),
    .Y(_5412_)
);

NAND3X1 _12943_ (
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .B(_5407_),
    .C(_5412_),
    .Y(_5413_)
);

NAND2X1 _12944_ (
    .A(_5409_),
    .B(_5413_),
    .Y(_5414_)
);

AOI21X1 _12945_ (
    .A(_5390_),
    .B(_5392_),
    .C(_5386_),
    .Y(_5415_)
);

AOI21X1 _12946_ (
    .A(_5384_),
    .B(_5393_),
    .C(_5415_),
    .Y(_5416_)
);

NAND3X1 _12947_ (
    .A(_5375_),
    .B(_5397_),
    .C(_5383_),
    .Y(_5417_)
);

AOI21X1 _12948_ (
    .A(_5417_),
    .B(_5416_),
    .C(_5414_),
    .Y(_5418_)
);

AND2X2 _12949_ (
    .A(_5413_),
    .B(_5409_),
    .Y(_5419_)
);

NAND3X1 _12950_ (
    .A(_5393_),
    .B(_5396_),
    .C(_5375_),
    .Y(_5420_)
);

OAI21X1 _12951_ (
    .A(_5420_),
    .B(_5363_),
    .C(_5416_),
    .Y(_5421_)
);

OAI21X1 _12952_ (
    .A(_5419_),
    .B(_5421_),
    .C(_5243_),
    .Y(_5422_)
);

OR2X2 _12953_ (
    .A(_5422_),
    .B(_5418_),
    .Y(_5423_)
);

AOI22X1 _12954_ (
    .A(_5118_),
    .B(_5174__bF$buf2),
    .C(_5423_),
    .D(_5246_),
    .Y(_5039_)
);

NAND2X1 _12955_ (
    .A(\genblk1[6].u_ce.Ycalc [11]),
    .B(_5174__bF$buf1),
    .Y(_5424_)
);

INVX1 _12956_ (
    .A(_5413_),
    .Y(_5425_)
);

NAND2X1 _12957_ (
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .B(_5340_),
    .Y(_5426_)
);

INVX1 _12958_ (
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5427_)
);

NAND2X1 _12959_ (
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .B(_5427_),
    .Y(_5428_)
);

NAND2X1 _12960_ (
    .A(_5426_),
    .B(_5428_),
    .Y(_5429_)
);

INVX1 _12961_ (
    .A(_5429_),
    .Y(_5430_)
);

NAND2X1 _12962_ (
    .A(_5430_),
    .B(_5406_),
    .Y(_5431_)
);

NAND2X1 _12963_ (
    .A(_5429_),
    .B(_5411_),
    .Y(_5432_)
);

NAND2X1 _12964_ (
    .A(_5431_),
    .B(_5432_),
    .Y(_5433_)
);

INVX1 _12965_ (
    .A(_5433_),
    .Y(_5434_)
);

NOR3X1 _12966_ (
    .A(_5425_),
    .B(_5434_),
    .C(_5418_),
    .Y(_5435_)
);

AOI21X1 _12967_ (
    .A(_5421_),
    .B(_5419_),
    .C(_5425_),
    .Y(_5436_)
);

OAI21X1 _12968_ (
    .A(_5433_),
    .B(_5436_),
    .C(_5243_),
    .Y(_5437_)
);

OAI21X1 _12969_ (
    .A(_5435_),
    .B(_5437_),
    .C(_5246_),
    .Y(_5438_)
);

NAND2X1 _12970_ (
    .A(_5424_),
    .B(_5438_),
    .Y(_5040_)
);

NAND2X1 _12971_ (
    .A(\genblk1[6].u_ce.Xcalc [0]),
    .B(_5174__bF$buf0),
    .Y(_5439_)
);

INVX1 _12972_ (
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5440_)
);

NAND2X1 _12973_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5441_)
);

OAI21X1 _12974_ (
    .A(1'h0),
    .B(_5440_),
    .C(_5441_),
    .Y(_5442_)
);

NAND2X1 _12975_ (
    .A(1'h1),
    .B(_5442_),
    .Y(_5443_)
);

NOR2X1 _12976_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_5444_)
);

NOR2X1 _12977_ (
    .A(1'h1),
    .B(_5180_),
    .Y(_5445_)
);

AOI22X1 _12978_ (
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .B(_5444_),
    .C(_5445_),
    .D(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5446_)
);

NAND3X1 _12979_ (
    .A(_5150__bF$buf4),
    .B(_5443_),
    .C(_5446_),
    .Y(_5447_)
);

NAND2X1 _12980_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5448_)
);

OAI21X1 _12981_ (
    .A(1'h0),
    .B(_5311_),
    .C(_5448_),
    .Y(_5449_)
);

NAND2X1 _12982_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5450_)
);

OAI21X1 _12983_ (
    .A(1'h0),
    .B(_5271_),
    .C(_5450_),
    .Y(_5451_)
);

MUX2X1 _12984_ (
    .A(_5451_),
    .B(_5449_),
    .S(_5151__bF$buf1),
    .Y(_5452_)
);

NAND2X1 _12985_ (
    .A(1'h1),
    .B(_5452_),
    .Y(_5453_)
);

AND2X2 _12986_ (
    .A(_5447_),
    .B(_5453_),
    .Y(_5454_)
);

NOR2X1 _12987_ (
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .B(_5454_),
    .Y(_5455_)
);

NAND2X1 _12988_ (
    .A(_5151__bF$buf0),
    .B(_5451_),
    .Y(_5456_)
);

NAND2X1 _12989_ (
    .A(1'h1),
    .B(_5449_),
    .Y(_5457_)
);

NAND2X1 _12990_ (
    .A(_5456_),
    .B(_5457_),
    .Y(_5458_)
);

OAI21X1 _12991_ (
    .A(_5150__bF$buf3),
    .B(_5458_),
    .C(_5447_),
    .Y(_5459_)
);

OAI21X1 _12992_ (
    .A(_5162_),
    .B(_5459_),
    .C(_5172_),
    .Y(_5460_)
);

OAI21X1 _12993_ (
    .A(_5460_),
    .B(_5455_),
    .C(_5439_),
    .Y(_5041_)
);

NAND2X1 _12994_ (
    .A(\genblk1[6].u_ce.Xcalc [1]),
    .B(_5174__bF$buf4),
    .Y(_5461_)
);

NOR2X1 _12995_ (
    .A(_5162_),
    .B(_5459_),
    .Y(_5462_)
);

NAND2X1 _12996_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5463_)
);

OAI21X1 _12997_ (
    .A(1'h0),
    .B(_5249_),
    .C(_5463_),
    .Y(_5464_)
);

NAND2X1 _12998_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5465_)
);

OAI21X1 _12999_ (
    .A(1'h0),
    .B(_5187_),
    .C(_5465_),
    .Y(_5466_)
);

MUX2X1 _13000_ (
    .A(_5466_),
    .B(_5464_),
    .S(_5151__bF$buf4),
    .Y(_5467_)
);

NAND2X1 _13001_ (
    .A(_5150__bF$buf2),
    .B(_5467_),
    .Y(_5468_)
);

NAND2X1 _13002_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5469_)
);

OAI21X1 _13003_ (
    .A(1'h0),
    .B(_5338_),
    .C(_5469_),
    .Y(_5470_)
);

INVX1 _13004_ (
    .A(_5470_),
    .Y(_5471_)
);

NAND2X1 _13005_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5472_)
);

OAI21X1 _13006_ (
    .A(1'h0),
    .B(_5292_),
    .C(_5472_),
    .Y(_5473_)
);

NAND2X1 _13007_ (
    .A(_5151__bF$buf3),
    .B(_5473_),
    .Y(_5474_)
);

OAI21X1 _13008_ (
    .A(_5151__bF$buf2),
    .B(_5471_),
    .C(_5474_),
    .Y(_5475_)
);

OAI21X1 _13009_ (
    .A(_5150__bF$buf1),
    .B(_5475_),
    .C(_5468_),
    .Y(_5476_)
);

NAND3X1 _13010_ (
    .A(_5188__bF$buf5),
    .B(_5476_),
    .C(_5454_),
    .Y(_5477_)
);

MUX2X1 _13011_ (
    .A(_5473_),
    .B(_5470_),
    .S(_5151__bF$buf1),
    .Y(_5478_)
);

MUX2X1 _13012_ (
    .A(_5478_),
    .B(_5467_),
    .S(1'h1),
    .Y(_5479_)
);

OAI21X1 _13013_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5459_),
    .C(_5479_),
    .Y(_5480_)
);

AOI21X1 _13014_ (
    .A(_5477_),
    .B(_5480_),
    .C(_5199_),
    .Y(_5481_)
);

INVX1 _13015_ (
    .A(_5481_),
    .Y(_5482_)
);

NAND3X1 _13016_ (
    .A(_5199_),
    .B(_5480_),
    .C(_5477_),
    .Y(_5483_)
);

AND2X2 _13017_ (
    .A(_5482_),
    .B(_5483_),
    .Y(_5484_)
);

NAND2X1 _13018_ (
    .A(_5462_),
    .B(_5484_),
    .Y(_5485_)
);

OR2X2 _13019_ (
    .A(_5484_),
    .B(_5462_),
    .Y(_5486_)
);

AOI21X1 _13020_ (
    .A(_5486_),
    .B(_5485_),
    .C(_5176_),
    .Y(_5487_)
);

OAI21X1 _13021_ (
    .A(_5174__bF$buf3),
    .B(_5487_),
    .C(_5461_),
    .Y(_5042_)
);

NAND2X1 _13022_ (
    .A(\genblk1[6].u_ce.Xcalc [2]),
    .B(_5174__bF$buf2),
    .Y(_5488_)
);

AOI21X1 _13023_ (
    .A(_5462_),
    .B(_5483_),
    .C(_5481_),
    .Y(_5489_)
);

NAND2X1 _13024_ (
    .A(_5459_),
    .B(_5476_),
    .Y(_5490_)
);

NAND2X1 _13025_ (
    .A(1'h0),
    .B(_5386_),
    .Y(_5491_)
);

OAI21X1 _13026_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .C(_5491_),
    .Y(_5492_)
);

NAND2X1 _13027_ (
    .A(_5151__bF$buf0),
    .B(_5449_),
    .Y(_5493_)
);

OAI21X1 _13028_ (
    .A(_5151__bF$buf4),
    .B(_5492_),
    .C(_5493_),
    .Y(_5494_)
);

NAND2X1 _13029_ (
    .A(_5257_),
    .B(_5442_),
    .Y(_5495_)
);

NAND2X1 _13030_ (
    .A(_5451_),
    .B(_5256_),
    .Y(_5496_)
);

NAND2X1 _13031_ (
    .A(_5495_),
    .B(_5496_),
    .Y(_5497_)
);

AOI21X1 _13032_ (
    .A(_5494_),
    .B(1'h1),
    .C(_5497_),
    .Y(_5498_)
);

INVX1 _13033_ (
    .A(_5498_),
    .Y(_5499_)
);

NAND3X1 _13034_ (
    .A(_5188__bF$buf4),
    .B(_5499_),
    .C(_5490_),
    .Y(_5500_)
);

AOI21X1 _13035_ (
    .A(_5447_),
    .B(_5453_),
    .C(_5479_),
    .Y(_5501_)
);

OAI21X1 _13036_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5501_),
    .C(_5498_),
    .Y(_5502_)
);

NAND3X1 _13037_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(_5502_),
    .C(_5500_),
    .Y(_5503_)
);

INVX1 _13038_ (
    .A(_5503_),
    .Y(_5504_)
);

AOI21X1 _13039_ (
    .A(_5500_),
    .B(_5502_),
    .C(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5505_)
);

NOR2X1 _13040_ (
    .A(_5505_),
    .B(_5504_),
    .Y(_5506_)
);

AND2X2 _13041_ (
    .A(_5506_),
    .B(_5489_),
    .Y(_5507_)
);

NOR2X1 _13042_ (
    .A(_5489_),
    .B(_5506_),
    .Y(_5508_)
);

OAI21X1 _13043_ (
    .A(_5508_),
    .B(_5507_),
    .C(_5243_),
    .Y(_5509_)
);

OAI21X1 _13044_ (
    .A(_5174__bF$buf1),
    .B(_5509_),
    .C(_5488_),
    .Y(_5043_)
);

OAI21X1 _13045_ (
    .A(_5505_),
    .B(_5489_),
    .C(_5503_),
    .Y(_5510_)
);

INVX1 _13046_ (
    .A(_5510_),
    .Y(_5511_)
);

NAND2X1 _13047_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [10]),
    .Y(_5512_)
);

OAI21X1 _13048_ (
    .A(1'h0),
    .B(_5386_),
    .C(_5512_),
    .Y(_5513_)
);

MUX2X1 _13049_ (
    .A(_5513_),
    .B(_5470_),
    .S(1'h1),
    .Y(_5514_)
);

NOR2X1 _13050_ (
    .A(_5150__bF$buf0),
    .B(_5514_),
    .Y(_5515_)
);

NAND2X1 _13051_ (
    .A(_5257_),
    .B(_5464_),
    .Y(_5516_)
);

NAND2X1 _13052_ (
    .A(_5473_),
    .B(_5256_),
    .Y(_5517_)
);

NAND2X1 _13053_ (
    .A(_5516_),
    .B(_5517_),
    .Y(_5518_)
);

OR2X2 _13054_ (
    .A(_5515_),
    .B(_5518_),
    .Y(_5519_)
);

OAI21X1 _13055_ (
    .A(_5499_),
    .B(_5490_),
    .C(_5188__bF$buf3),
    .Y(_5520_)
);

OR2X2 _13056_ (
    .A(_5520_),
    .B(_5519_),
    .Y(_5521_)
);

OAI21X1 _13057_ (
    .A(_5515_),
    .B(_5518_),
    .C(_5520_),
    .Y(_5522_)
);

AOI21X1 _13058_ (
    .A(_5521_),
    .B(_5522_),
    .C(_5196_),
    .Y(_5523_)
);

INVX1 _13059_ (
    .A(_5523_),
    .Y(_5524_)
);

NAND3X1 _13060_ (
    .A(_5196_),
    .B(_5522_),
    .C(_5521_),
    .Y(_5525_)
);

NAND2X1 _13061_ (
    .A(_5525_),
    .B(_5524_),
    .Y(_5526_)
);

OR2X2 _13062_ (
    .A(_5526_),
    .B(_5511_),
    .Y(_5527_)
);

NAND2X1 _13063_ (
    .A(_5511_),
    .B(_5526_),
    .Y(_5528_)
);

NAND2X1 _13064_ (
    .A(_5528_),
    .B(_5527_),
    .Y(_5529_)
);

AOI22X1 _13065_ (
    .A(_5142_),
    .B(_5174__bF$buf0),
    .C(_5529_),
    .D(_5172_),
    .Y(_5044_)
);

AOI21X1 _13066_ (
    .A(_5510_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5530_)
);

NAND2X1 _13067_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5531_)
);

OAI21X1 _13068_ (
    .A(1'h0),
    .B(_5401_),
    .C(_5531_),
    .Y(_5532_)
);

NAND2X1 _13069_ (
    .A(1'h1),
    .B(_5532_),
    .Y(_5533_)
);

OAI21X1 _13070_ (
    .A(1'h1),
    .B(_5492_),
    .C(_5533_),
    .Y(_5534_)
);

NAND2X1 _13071_ (
    .A(1'h1),
    .B(_5534_),
    .Y(_5535_)
);

OAI21X1 _13072_ (
    .A(1'h1),
    .B(_5452_),
    .C(_5535_),
    .Y(_5536_)
);

INVX1 _13073_ (
    .A(_5536_),
    .Y(_5537_)
);

NAND3X1 _13074_ (
    .A(_5498_),
    .B(_5459_),
    .C(_5476_),
    .Y(_5538_)
);

OAI21X1 _13075_ (
    .A(_5519_),
    .B(_5538_),
    .C(_5188__bF$buf2),
    .Y(_5539_)
);

OR2X2 _13076_ (
    .A(_5539_),
    .B(_5537_),
    .Y(_5540_)
);

NOR2X1 _13077_ (
    .A(_5519_),
    .B(_5538_),
    .Y(_5541_)
);

OAI21X1 _13078_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5541_),
    .C(_5537_),
    .Y(_5542_)
);

NAND3X1 _13079_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(_5542_),
    .C(_5540_),
    .Y(_5543_)
);

OR2X2 _13080_ (
    .A(_5539_),
    .B(_5536_),
    .Y(_5544_)
);

OAI21X1 _13081_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5541_),
    .C(_5536_),
    .Y(_5545_)
);

NAND3X1 _13082_ (
    .A(_5155_),
    .B(_5545_),
    .C(_5544_),
    .Y(_5546_)
);

NAND2X1 _13083_ (
    .A(_5543_),
    .B(_5546_),
    .Y(_5547_)
);

OR2X2 _13084_ (
    .A(_5530_),
    .B(_5547_),
    .Y(_5548_)
);

NAND2X1 _13085_ (
    .A(_5547_),
    .B(_5530_),
    .Y(_5549_)
);

NAND2X1 _13086_ (
    .A(_5549_),
    .B(_5548_),
    .Y(_5550_)
);

AOI22X1 _13087_ (
    .A(_5137_),
    .B(_5174__bF$buf4),
    .C(_5550_),
    .D(_5172_),
    .Y(_5045_)
);

INVX1 _13088_ (
    .A(\genblk1[6].u_ce.Xcalc [5]),
    .Y(_5551_)
);

OAI21X1 _13089_ (
    .A(_5547_),
    .B(_5530_),
    .C(_5543_),
    .Y(_5552_)
);

NAND2X1 _13090_ (
    .A(_5537_),
    .B(_5541_),
    .Y(_5553_)
);

NOR2X1 _13091_ (
    .A(_5151__bF$buf3),
    .B(_5427_),
    .Y(_5554_)
);

AOI21X1 _13092_ (
    .A(_5151__bF$buf2),
    .B(_5513_),
    .C(_5554_),
    .Y(_5555_)
);

NAND2X1 _13093_ (
    .A(_5150__bF$buf4),
    .B(_5475_),
    .Y(_5556_)
);

OAI21X1 _13094_ (
    .A(_5150__bF$buf3),
    .B(_5555_),
    .C(_5556_),
    .Y(_5557_)
);

INVX1 _13095_ (
    .A(_5557_),
    .Y(_5558_)
);

NAND3X1 _13096_ (
    .A(_5188__bF$buf1),
    .B(_5558_),
    .C(_5553_),
    .Y(_5559_)
);

NOR2X1 _13097_ (
    .A(_5518_),
    .B(_5515_),
    .Y(_5560_)
);

NAND3X1 _13098_ (
    .A(_5498_),
    .B(_5560_),
    .C(_5501_),
    .Y(_5561_)
);

OAI21X1 _13099_ (
    .A(_5536_),
    .B(_5561_),
    .C(_5188__bF$buf0),
    .Y(_5562_)
);

NAND2X1 _13100_ (
    .A(_5557_),
    .B(_5562_),
    .Y(_5563_)
);

AOI21X1 _13101_ (
    .A(_5559_),
    .B(_5563_),
    .C(_5192_),
    .Y(_5564_)
);

INVX1 _13102_ (
    .A(_5564_),
    .Y(_5565_)
);

NAND3X1 _13103_ (
    .A(_5192_),
    .B(_5563_),
    .C(_5559_),
    .Y(_5566_)
);

NAND2X1 _13104_ (
    .A(_5566_),
    .B(_5565_),
    .Y(_5567_)
);

NOR2X1 _13105_ (
    .A(_5567_),
    .B(_5552_),
    .Y(_5568_)
);

AND2X2 _13106_ (
    .A(_5552_),
    .B(_5567_),
    .Y(_5569_)
);

OAI21X1 _13107_ (
    .A(_5568_),
    .B(_5569_),
    .C(_5172_),
    .Y(_5570_)
);

OAI21X1 _13108_ (
    .A(_5551_),
    .B(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .C(_5570_),
    .Y(_5046_)
);

INVX1 _13109_ (
    .A(\genblk1[6].u_ce.Xcalc [6]),
    .Y(_5571_)
);

NAND3X1 _13110_ (
    .A(_5537_),
    .B(_5558_),
    .C(_5541_),
    .Y(_5572_)
);

AOI21X1 _13111_ (
    .A(_5151__bF$buf1),
    .B(_5532_),
    .C(_5554_),
    .Y(_5573_)
);

NAND2X1 _13112_ (
    .A(1'h1),
    .B(_5573_),
    .Y(_5574_)
);

OAI21X1 _13113_ (
    .A(1'h1),
    .B(_5494_),
    .C(_5574_),
    .Y(_5575_)
);

NAND3X1 _13114_ (
    .A(_5188__bF$buf5),
    .B(_5575_),
    .C(_5572_),
    .Y(_5576_)
);

NOR3X1 _13115_ (
    .A(_5536_),
    .B(_5557_),
    .C(_5561_),
    .Y(_5577_)
);

INVX1 _13116_ (
    .A(_5575_),
    .Y(_5578_)
);

OAI21X1 _13117_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5577_),
    .C(_5578_),
    .Y(_5579_)
);

NAND2X1 _13118_ (
    .A(_5576_),
    .B(_5579_),
    .Y(_5580_)
);

NAND2X1 _13119_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(_5580_),
    .Y(_5581_)
);

NAND3X1 _13120_ (
    .A(_5152_),
    .B(_5576_),
    .C(_5579_),
    .Y(_5582_)
);

NAND2X1 _13121_ (
    .A(_5582_),
    .B(_5581_),
    .Y(_5583_)
);

AOI21X1 _13122_ (
    .A(_5544_),
    .B(_5545_),
    .C(_5155_),
    .Y(_5584_)
);

NOR2X1 _13123_ (
    .A(_5584_),
    .B(_5564_),
    .Y(_5585_)
);

OAI21X1 _13124_ (
    .A(_5547_),
    .B(_5530_),
    .C(_5585_),
    .Y(_5586_)
);

NAND2X1 _13125_ (
    .A(_5566_),
    .B(_5586_),
    .Y(_5587_)
);

NOR2X1 _13126_ (
    .A(_5583_),
    .B(_5587_),
    .Y(_5588_)
);

AND2X2 _13127_ (
    .A(_5581_),
    .B(_5582_),
    .Y(_5589_)
);

AND2X2 _13128_ (
    .A(_5543_),
    .B(_5546_),
    .Y(_5590_)
);

NAND3X1 _13129_ (
    .A(_5566_),
    .B(_5590_),
    .C(_5565_),
    .Y(_5591_)
);

AOI21X1 _13130_ (
    .A(_5584_),
    .B(_5566_),
    .C(_5564_),
    .Y(_5592_)
);

OAI21X1 _13131_ (
    .A(_5530_),
    .B(_5591_),
    .C(_5592_),
    .Y(_5593_)
);

NOR2X1 _13132_ (
    .A(_5589_),
    .B(_5593_),
    .Y(_5594_)
);

OAI21X1 _13133_ (
    .A(_5594_),
    .B(_5588_),
    .C(_5243_),
    .Y(_5595_)
);

NAND2X1 _13134_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .B(_5595_),
    .Y(_5596_)
);

OAI21X1 _13135_ (
    .A(_5571_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5596_),
    .Y(_5047_)
);

INVX1 _13136_ (
    .A(\genblk1[6].u_ce.Xcalc [7]),
    .Y(_5597_)
);

INVX1 _13137_ (
    .A(_5581_),
    .Y(_5598_)
);

NAND2X1 _13138_ (
    .A(_5575_),
    .B(_5577_),
    .Y(_5599_)
);

NOR2X1 _13139_ (
    .A(_5150__bF$buf2),
    .B(_5427_),
    .Y(_5600_)
);

INVX1 _13140_ (
    .A(_5600_),
    .Y(_5601_)
);

OAI21X1 _13141_ (
    .A(1'h1),
    .B(_5514_),
    .C(_5601_),
    .Y(_5602_)
);

NAND3X1 _13142_ (
    .A(_5188__bF$buf4),
    .B(_5602_),
    .C(_5599_),
    .Y(_5603_)
);

INVX1 _13143_ (
    .A(_5602_),
    .Y(_5604_)
);

OAI21X1 _13144_ (
    .A(_5578_),
    .B(_5572_),
    .C(_5188__bF$buf3),
    .Y(_5605_)
);

NAND2X1 _13145_ (
    .A(_5604_),
    .B(_5605_),
    .Y(_5606_)
);

NAND3X1 _13146_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(_5603_),
    .C(_5606_),
    .Y(_5607_)
);

NAND3X1 _13147_ (
    .A(_5188__bF$buf2),
    .B(_5604_),
    .C(_5599_),
    .Y(_5608_)
);

NAND2X1 _13148_ (
    .A(_5602_),
    .B(_5605_),
    .Y(_5609_)
);

NAND3X1 _13149_ (
    .A(_5189_),
    .B(_5608_),
    .C(_5609_),
    .Y(_5610_)
);

NAND2X1 _13150_ (
    .A(_5607_),
    .B(_5610_),
    .Y(_5611_)
);

OAI21X1 _13151_ (
    .A(_5598_),
    .B(_5588_),
    .C(_5611_),
    .Y(_5612_)
);

NOR2X1 _13152_ (
    .A(_5598_),
    .B(_5588_),
    .Y(_5613_)
);

INVX1 _13153_ (
    .A(_5611_),
    .Y(_5614_)
);

AOI21X1 _13154_ (
    .A(_5613_),
    .B(_5614_),
    .C(_5171_),
    .Y(_5615_)
);

AOI22X1 _13155_ (
    .A(_5597_),
    .B(_5174__bF$buf3),
    .C(_5615_),
    .D(_5612_),
    .Y(_5048_)
);

OAI21X1 _13156_ (
    .A(_5581_),
    .B(_5611_),
    .C(_5607_),
    .Y(_5616_)
);

NOR2X1 _13157_ (
    .A(_5583_),
    .B(_5611_),
    .Y(_5617_)
);

AOI21X1 _13158_ (
    .A(_5617_),
    .B(_5593_),
    .C(_5616_),
    .Y(_5618_)
);

INVX1 _13159_ (
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5619_)
);

NAND3X1 _13160_ (
    .A(_5575_),
    .B(_5604_),
    .C(_5577_),
    .Y(_5620_)
);

INVX1 _13161_ (
    .A(_5534_),
    .Y(_5621_)
);

OAI21X1 _13162_ (
    .A(1'h1),
    .B(_5621_),
    .C(_5601_),
    .Y(_5622_)
);

INVX1 _13163_ (
    .A(_5622_),
    .Y(_5623_)
);

NAND3X1 _13164_ (
    .A(_5188__bF$buf1),
    .B(_5623_),
    .C(_5620_),
    .Y(_5624_)
);

OAI21X1 _13165_ (
    .A(_5602_),
    .B(_5599_),
    .C(_5188__bF$buf0),
    .Y(_5625_)
);

NAND2X1 _13166_ (
    .A(_5622_),
    .B(_5625_),
    .Y(_5626_)
);

AOI21X1 _13167_ (
    .A(_5626_),
    .B(_5624_),
    .C(_5619_),
    .Y(_5627_)
);

NAND3X1 _13168_ (
    .A(_5188__bF$buf5),
    .B(_5622_),
    .C(_5620_),
    .Y(_5628_)
);

NAND2X1 _13169_ (
    .A(_5623_),
    .B(_5625_),
    .Y(_5629_)
);

AOI21X1 _13170_ (
    .A(_5629_),
    .B(_5628_),
    .C(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5630_)
);

OAI21X1 _13171_ (
    .A(_5627_),
    .B(_5630_),
    .C(_5618_),
    .Y(_5631_)
);

INVX1 _13172_ (
    .A(_5631_),
    .Y(_5632_)
);

OR2X2 _13173_ (
    .A(_5627_),
    .B(_5630_),
    .Y(_5633_)
);

OAI21X1 _13174_ (
    .A(_5633_),
    .B(_5618_),
    .C(_5172_),
    .Y(_5634_)
);

OAI22X1 _13175_ (
    .A(_5134_),
    .B(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .C(_5634_),
    .D(_5632_),
    .Y(_5049_)
);

NAND2X1 _13176_ (
    .A(\genblk1[6].u_ce.Xcalc [9]),
    .B(_5174__bF$buf2),
    .Y(_5635_)
);

NOR2X1 _13177_ (
    .A(_5633_),
    .B(_5618_),
    .Y(_5636_)
);

NOR2X1 _13178_ (
    .A(_5627_),
    .B(_5636_),
    .Y(_5637_)
);

OAI21X1 _13179_ (
    .A(1'h1),
    .B(_5555_),
    .C(_5601_),
    .Y(_5638_)
);

INVX1 _13180_ (
    .A(_5638_),
    .Y(_5639_)
);

OAI21X1 _13181_ (
    .A(_5622_),
    .B(_5620_),
    .C(_5188__bF$buf4),
    .Y(_5640_)
);

NAND2X1 _13182_ (
    .A(_5639_),
    .B(_5640_),
    .Y(_5641_)
);

OR2X2 _13183_ (
    .A(_5640_),
    .B(_5639_),
    .Y(_5642_)
);

NAND3X1 _13184_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(_5641_),
    .C(_5642_),
    .Y(_5643_)
);

NAND2X1 _13185_ (
    .A(_5641_),
    .B(_5642_),
    .Y(_5644_)
);

NAND2X1 _13186_ (
    .A(_5251_),
    .B(_5644_),
    .Y(_5645_)
);

NAND2X1 _13187_ (
    .A(_5643_),
    .B(_5645_),
    .Y(_5646_)
);

AND2X2 _13188_ (
    .A(_5637_),
    .B(_5646_),
    .Y(_5647_)
);

OAI21X1 _13189_ (
    .A(_5646_),
    .B(_5637_),
    .C(_5172_),
    .Y(_5648_)
);

OAI21X1 _13190_ (
    .A(_5648_),
    .B(_5647_),
    .C(_5635_),
    .Y(_5050_)
);

INVX1 _13191_ (
    .A(\genblk1[6].u_ce.Xcalc [10]),
    .Y(_5649_)
);

INVX1 _13192_ (
    .A(_5643_),
    .Y(_5650_)
);

AOI21X1 _13193_ (
    .A(_5627_),
    .B(_5645_),
    .C(_5650_),
    .Y(_5651_)
);

NOR2X1 _13194_ (
    .A(_5627_),
    .B(_5630_),
    .Y(_5652_)
);

NAND3X1 _13195_ (
    .A(_5643_),
    .B(_5645_),
    .C(_5652_),
    .Y(_5653_)
);

OAI21X1 _13196_ (
    .A(_5618_),
    .B(_5653_),
    .C(_5651_),
    .Y(_5654_)
);

OAI21X1 _13197_ (
    .A(1'h1),
    .B(_5573_),
    .C(_5601_),
    .Y(_5655_)
);

INVX1 _13198_ (
    .A(_5655_),
    .Y(_5656_)
);

OR2X2 _13199_ (
    .A(_5620_),
    .B(_5622_),
    .Y(_5657_)
);

OAI21X1 _13200_ (
    .A(_5638_),
    .B(_5657_),
    .C(_5188__bF$buf3),
    .Y(_5658_)
);

NAND2X1 _13201_ (
    .A(_5656_),
    .B(_5658_),
    .Y(_5659_)
);

OR2X2 _13202_ (
    .A(_5658_),
    .B(_5656_),
    .Y(_5660_)
);

NAND3X1 _13203_ (
    .A(\genblk1[6].u_ce.Xin12b [10]),
    .B(_5659_),
    .C(_5660_),
    .Y(_5661_)
);

AND2X2 _13204_ (
    .A(_5658_),
    .B(_5656_),
    .Y(_5662_)
);

NOR2X1 _13205_ (
    .A(_5656_),
    .B(_5658_),
    .Y(_5663_)
);

OAI21X1 _13206_ (
    .A(_5663_),
    .B(_5662_),
    .C(_5272_),
    .Y(_5664_)
);

NAND2X1 _13207_ (
    .A(_5664_),
    .B(_5661_),
    .Y(_5665_)
);

AND2X2 _13208_ (
    .A(_5654_),
    .B(_5665_),
    .Y(_5666_)
);

NOR2X1 _13209_ (
    .A(_5665_),
    .B(_5654_),
    .Y(_5667_)
);

NOR2X1 _13210_ (
    .A(_5666_),
    .B(_5667_),
    .Y(_5668_)
);

AOI22X1 _13211_ (
    .A(_5649_),
    .B(_5174__bF$buf1),
    .C(_5668_),
    .D(_5172_),
    .Y(_5051_)
);

NAND2X1 _13212_ (
    .A(\genblk1[6].u_ce.Xcalc [11]),
    .B(_5174__bF$buf0),
    .Y(_5669_)
);

INVX1 _13213_ (
    .A(_5661_),
    .Y(_5670_)
);

AOI21X1 _13214_ (
    .A(_5654_),
    .B(_5664_),
    .C(_5670_),
    .Y(_5671_)
);

NAND2X1 _13215_ (
    .A(_5188__bF$buf2),
    .B(_5659_),
    .Y(_5672_)
);

NOR2X1 _13216_ (
    .A(_5429_),
    .B(_5672_),
    .Y(_5673_)
);

AOI21X1 _13217_ (
    .A(_5659_),
    .B(_5188__bF$buf1),
    .C(_5430_),
    .Y(_5674_)
);

NOR2X1 _13218_ (
    .A(_5674_),
    .B(_5673_),
    .Y(_5675_)
);

AND2X2 _13219_ (
    .A(_5671_),
    .B(_5675_),
    .Y(_5676_)
);

OAI21X1 _13220_ (
    .A(_5675_),
    .B(_5671_),
    .C(_5172_),
    .Y(_5677_)
);

OAI21X1 _13221_ (
    .A(_5677_),
    .B(_5676_),
    .C(_5669_),
    .Y(_5052_)
);

OAI21X1 _13222_ (
    .A(1'h0),
    .B(_5151__bF$buf0),
    .C(_5170_),
    .Y(_5678_)
);

OAI21X1 _13223_ (
    .A(_5445_),
    .B(_5678_),
    .C(\genblk1[6].u_ce.Ain0 [0]),
    .Y(_5679_)
);

INVX1 _13224_ (
    .A(\genblk1[6].u_ce.Ain0 [0]),
    .Y(_5680_)
);

NAND2X1 _13225_ (
    .A(\genblk1[6].u_ce.Acalc [1]),
    .B(_5174__bF$buf4),
    .Y(_5681_)
);

INVX1 _13226_ (
    .A(_5679_),
    .Y(_5682_)
);

NOR2X1 _13227_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_5683_)
);

AOI21X1 _13228_ (
    .A(_5445_),
    .B(1'h1),
    .C(_5683_),
    .Y(_5684_)
);

NOR2X1 _13229_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5684_),
    .Y(_5685_)
);

OAI21X1 _13230_ (
    .A(_5445_),
    .B(_5678_),
    .C(_5188__bF$buf0),
    .Y(_5686_)
);

AND2X2 _13231_ (
    .A(_5686_),
    .B(_5684_),
    .Y(_5687_)
);

OR2X2 _13232_ (
    .A(_5687_),
    .B(_5685_),
    .Y(_5688_)
);

OR2X2 _13233_ (
    .A(_5688_),
    .B(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5689_)
);

OAI21X1 _13234_ (
    .A(_5685_),
    .B(_5687_),
    .C(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5690_)
);

NAND2X1 _13235_ (
    .A(_5690_),
    .B(_5689_),
    .Y(_5691_)
);

NOR2X1 _13236_ (
    .A(_5682_),
    .B(_5691_),
    .Y(_5692_)
);

NAND2X1 _13237_ (
    .A(_5682_),
    .B(_5691_),
    .Y(_5693_)
);

NAND2X1 _13238_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .B(_5693_),
    .Y(_5694_)
);

OAI21X1 _13239_ (
    .A(_5692_),
    .B(_5694_),
    .C(_5681_),
    .Y(_5053_)
);

INVX1 _13240_ (
    .A(\genblk1[6].u_ce.Ain0 [1]),
    .Y(_5695_)
);

OAI21X1 _13241_ (
    .A(_5695_),
    .B(_5688_),
    .C(_5693_),
    .Y(_5696_)
);

OAI21X1 _13242_ (
    .A(_5180_),
    .B(_5151__bF$buf4),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5697_)
);

OAI21X1 _13243_ (
    .A(1'h0),
    .B(1'h1),
    .C(1'h1),
    .Y(_5698_)
);

MUX2X1 _13244_ (
    .A(_5698_),
    .B(1'h1),
    .S(_5697_),
    .Y(_5699_)
);

NAND2X1 _13245_ (
    .A(\genblk1[6].u_ce.Ain1 [0]),
    .B(_5699_),
    .Y(_5700_)
);

OR2X2 _13246_ (
    .A(_5699_),
    .B(\genblk1[6].u_ce.Ain1 [0]),
    .Y(_5701_)
);

NAND2X1 _13247_ (
    .A(_5700_),
    .B(_5701_),
    .Y(_5702_)
);

INVX1 _13248_ (
    .A(_5702_),
    .Y(_5703_)
);

NAND2X1 _13249_ (
    .A(_5703_),
    .B(_5696_),
    .Y(_5704_)
);

NOR2X1 _13250_ (
    .A(\genblk1[6].u_ce.Acalc [3]),
    .B(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .Y(_5705_)
);

NAND2X1 _13251_ (
    .A(_5700_),
    .B(_5704_),
    .Y(_5706_)
);

INVX1 _13252_ (
    .A(_5706_),
    .Y(_5707_)
);

INVX1 _13253_ (
    .A(\genblk1[6].u_ce.Ain1 [1]),
    .Y(_5708_)
);

NOR2X1 _13254_ (
    .A(1'h0),
    .B(_5151__bF$buf3),
    .Y(_5709_)
);

OAI21X1 _13255_ (
    .A(_5150__bF$buf1),
    .B(_5709_),
    .C(_5188__bF$buf5),
    .Y(_5710_)
);

OAI21X1 _13256_ (
    .A(1'h1),
    .B(1'h1),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_5711_)
);

OAI21X1 _13257_ (
    .A(_5180_),
    .B(_5711_),
    .C(_5710_),
    .Y(_5712_)
);

NOR2X1 _13258_ (
    .A(_5708_),
    .B(_5712_),
    .Y(_5713_)
);

NAND2X1 _13259_ (
    .A(_5708_),
    .B(_5712_),
    .Y(_5714_)
);

INVX1 _13260_ (
    .A(_5714_),
    .Y(_5715_)
);

NOR2X1 _13261_ (
    .A(_5713_),
    .B(_5715_),
    .Y(_5716_)
);

OAI21X1 _13262_ (
    .A(_5716_),
    .B(_5707_),
    .C(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .Y(_5717_)
);

AOI21X1 _13263_ (
    .A(_5707_),
    .B(_5716_),
    .C(_5717_),
    .Y(_5718_)
);

NOR2X1 _13264_ (
    .A(_5705_),
    .B(_5718_),
    .Y(_5054_)
);

INVX1 _13265_ (
    .A(\genblk1[6].u_ce.Ain12b [4]),
    .Y(_5719_)
);

AOI21X1 _13266_ (
    .A(_5445_),
    .B(1'h1),
    .C(_5188__bF$buf4),
    .Y(_5720_)
);

OAI21X1 _13267_ (
    .A(1'h1),
    .B(_5445_),
    .C(_5720_),
    .Y(_5721_)
);

OAI21X1 _13268_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5684_),
    .C(_5721_),
    .Y(_5722_)
);

OR2X2 _13269_ (
    .A(_5722_),
    .B(_5719_),
    .Y(_5723_)
);

NAND2X1 _13270_ (
    .A(_5719_),
    .B(_5722_),
    .Y(_5724_)
);

NAND2X1 _13271_ (
    .A(_5724_),
    .B(_5723_),
    .Y(_5725_)
);

AOI21X1 _13272_ (
    .A(_5706_),
    .B(_5714_),
    .C(_5713_),
    .Y(_5726_)
);

OAI21X1 _13273_ (
    .A(_5725_),
    .B(_5726_),
    .C(_5723_),
    .Y(_5727_)
);

INVX1 _13274_ (
    .A(\genblk1[6].u_ce.Ain12b [5]),
    .Y(_5728_)
);

OAI21X1 _13275_ (
    .A(_5444_),
    .B(_5257_),
    .C(_5188__bF$buf3),
    .Y(_5729_)
);

OAI21X1 _13276_ (
    .A(1'h0),
    .B(1'h1),
    .C(_5170_),
    .Y(_5730_)
);

OR2X2 _13277_ (
    .A(_5730_),
    .B(_5188__bF$buf2),
    .Y(_5731_)
);

NAND2X1 _13278_ (
    .A(_5729_),
    .B(_5731_),
    .Y(_5732_)
);

OR2X2 _13279_ (
    .A(_5732_),
    .B(_5728_),
    .Y(_5733_)
);

NAND2X1 _13280_ (
    .A(_5728_),
    .B(_5732_),
    .Y(_5734_)
);

NAND2X1 _13281_ (
    .A(_5734_),
    .B(_5733_),
    .Y(_5735_)
);

INVX1 _13282_ (
    .A(_5735_),
    .Y(_5736_)
);

NOR2X1 _13283_ (
    .A(_5736_),
    .B(_5727_),
    .Y(_5737_)
);

NAND2X1 _13284_ (
    .A(_5736_),
    .B(_5727_),
    .Y(_5738_)
);

NAND2X1 _13285_ (
    .A(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .B(_5738_),
    .Y(_5739_)
);

OAI22X1 _13286_ (
    .A(_5113_),
    .B(\genblk1[6].u_ce.Vld_bF$buf1 ),
    .C(_5737_),
    .D(_5739_),
    .Y(_5055_)
);

INVX1 _13287_ (
    .A(_5725_),
    .Y(_5740_)
);

NAND2X1 _13288_ (
    .A(_5736_),
    .B(_5740_),
    .Y(_5741_)
);

OAI21X1 _13289_ (
    .A(_5723_),
    .B(_5735_),
    .C(_5733_),
    .Y(_5742_)
);

INVX1 _13290_ (
    .A(_5742_),
    .Y(_5743_)
);

OAI21X1 _13291_ (
    .A(_5741_),
    .B(_5726_),
    .C(_5743_),
    .Y(_5744_)
);

OAI21X1 _13292_ (
    .A(1'h1),
    .B(_5180_),
    .C(_5150__bF$buf0),
    .Y(_5745_)
);

NOR2X1 _13293_ (
    .A(_5745_),
    .B(_5709_),
    .Y(_5746_)
);

NAND2X1 _13294_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5746_),
    .Y(_5747_)
);

OAI21X1 _13295_ (
    .A(_5745_),
    .B(_5709_),
    .C(_5188__bF$buf1),
    .Y(_5748_)
);

NAND2X1 _13296_ (
    .A(_5748_),
    .B(_5747_),
    .Y(_5749_)
);

NAND2X1 _13297_ (
    .A(\genblk1[6].u_ce.Ain12b [6]),
    .B(_5749_),
    .Y(_5750_)
);

OR2X2 _13298_ (
    .A(_5749_),
    .B(\genblk1[6].u_ce.Ain12b [6]),
    .Y(_5751_)
);

NAND2X1 _13299_ (
    .A(_5750_),
    .B(_5751_),
    .Y(_5752_)
);

INVX1 _13300_ (
    .A(_5752_),
    .Y(_5753_)
);

NAND2X1 _13301_ (
    .A(_5753_),
    .B(_5744_),
    .Y(_5754_)
);

INVX1 _13302_ (
    .A(\genblk1[6].u_ce.Acalc [7]),
    .Y(_5755_)
);

NAND2X1 _13303_ (
    .A(_5750_),
    .B(_5754_),
    .Y(_5756_)
);

INVX1 _13304_ (
    .A(\genblk1[6].u_ce.Ain12b [7]),
    .Y(_5757_)
);

NAND2X1 _13305_ (
    .A(_5188__bF$buf0),
    .B(_5683_),
    .Y(_5758_)
);

OR2X2 _13306_ (
    .A(_5683_),
    .B(_5188__bF$buf5),
    .Y(_5759_)
);

NAND2X1 _13307_ (
    .A(_5758_),
    .B(_5759_),
    .Y(_5760_)
);

NOR2X1 _13308_ (
    .A(_5757_),
    .B(_5760_),
    .Y(_5761_)
);

INVX1 _13309_ (
    .A(_5761_),
    .Y(_5762_)
);

NAND2X1 _13310_ (
    .A(_5757_),
    .B(_5760_),
    .Y(_5763_)
);

NAND2X1 _13311_ (
    .A(_5763_),
    .B(_5762_),
    .Y(_5764_)
);

OR2X2 _13312_ (
    .A(_5756_),
    .B(_5764_),
    .Y(_5765_)
);

AOI21X1 _13313_ (
    .A(_5756_),
    .B(_5764_),
    .C(_5174__bF$buf3),
    .Y(_5766_)
);

AOI22X1 _13314_ (
    .A(_5755_),
    .B(_5174__bF$buf2),
    .C(_5765_),
    .D(_5766_),
    .Y(_5056_)
);

NOR2X1 _13315_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5170_),
    .Y(_5767_)
);

INVX1 _13316_ (
    .A(_5767_),
    .Y(_5768_)
);

NAND3X1 _13317_ (
    .A(\genblk1[6].u_ce.Ain12b [8]),
    .B(_5711_),
    .C(_5768_),
    .Y(_5769_)
);

INVX1 _13318_ (
    .A(_5769_),
    .Y(_5770_)
);

AOI21X1 _13319_ (
    .A(_5768_),
    .B(_5711_),
    .C(\genblk1[6].u_ce.Ain12b [8]),
    .Y(_5771_)
);

NOR2X1 _13320_ (
    .A(_5771_),
    .B(_5770_),
    .Y(_5772_)
);

OAI21X1 _13321_ (
    .A(_5750_),
    .B(_5764_),
    .C(_5762_),
    .Y(_5773_)
);

NOR2X1 _13322_ (
    .A(_5764_),
    .B(_5752_),
    .Y(_5774_)
);

AOI21X1 _13323_ (
    .A(_5774_),
    .B(_5742_),
    .C(_5773_),
    .Y(_5775_)
);

NAND3X1 _13324_ (
    .A(_5740_),
    .B(_5736_),
    .C(_5774_),
    .Y(_5776_)
);

OAI21X1 _13325_ (
    .A(_5776_),
    .B(_5726_),
    .C(_5775_),
    .Y(_5777_)
);

AOI21X1 _13326_ (
    .A(_5777_),
    .B(_5772_),
    .C(_5770_),
    .Y(_5778_)
);

OR2X2 _13327_ (
    .A(_5188__bF$buf4),
    .B(\genblk1[6].u_ce.Ain12b [9]),
    .Y(_5779_)
);

NAND2X1 _13328_ (
    .A(\genblk1[6].u_ce.Ain12b [9]),
    .B(_5188__bF$buf3),
    .Y(_5780_)
);

NAND2X1 _13329_ (
    .A(_5780_),
    .B(_5779_),
    .Y(_5781_)
);

AND2X2 _13330_ (
    .A(_5778_),
    .B(_5781_),
    .Y(_5782_)
);

OAI21X1 _13331_ (
    .A(_5781_),
    .B(_5778_),
    .C(\genblk1[6].u_ce.Vld_bF$buf0 ),
    .Y(_5783_)
);

OAI22X1 _13332_ (
    .A(_5110_),
    .B(\genblk1[6].u_ce.Vld_bF$buf3 ),
    .C(_5783_),
    .D(_5782_),
    .Y(_5057_)
);

OAI21X1 _13333_ (
    .A(_5781_),
    .B(_5769_),
    .C(_5780_),
    .Y(_5784_)
);

NAND3X1 _13334_ (
    .A(_5779_),
    .B(_5780_),
    .C(_5772_),
    .Y(_5785_)
);

INVX1 _13335_ (
    .A(_5785_),
    .Y(_5786_)
);

AOI21X1 _13336_ (
    .A(_5777_),
    .B(_5786_),
    .C(_5784_),
    .Y(_5787_)
);

INVX1 _13337_ (
    .A(\genblk1[6].u_ce.Ain12b [10]),
    .Y(_5788_)
);

NAND2X1 _13338_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5788_),
    .Y(_5789_)
);

NAND2X1 _13339_ (
    .A(\genblk1[6].u_ce.Ain12b [10]),
    .B(_5188__bF$buf2),
    .Y(_5790_)
);

NAND2X1 _13340_ (
    .A(_5789_),
    .B(_5790_),
    .Y(_5791_)
);

NAND2X1 _13341_ (
    .A(\genblk1[6].u_ce.Acalc [11]),
    .B(_5174__bF$buf1),
    .Y(_5792_)
);

OAI21X1 _13342_ (
    .A(_5791_),
    .B(_5787_),
    .C(_5790_),
    .Y(_5793_)
);

OAI21X1 _13343_ (
    .A(_5174__bF$buf0),
    .B(_5793_),
    .C(_5792_),
    .Y(_5058_)
);

NAND2X1 _13344_ (
    .A(\genblk1[6].u_ce.LoadCtl [5]),
    .B(_5105_),
    .Y(_5794_)
);

NAND2X1 _13345_ (
    .A(_5106_),
    .B(_5109_),
    .Y(_5795_)
);

NOR2X1 _13346_ (
    .A(_5794_),
    .B(_5795_),
    .Y(_5796_)
);

NAND2X1 _13347_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5796_),
    .Y(_5797_)
);

OAI21X1 _13348_ (
    .A(_5272_),
    .B(_5796_),
    .C(_5797_),
    .Y(_5059_)
);

NAND2X1 _13349_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5796_),
    .Y(_5798_)
);

OAI21X1 _13350_ (
    .A(_5340_),
    .B(_5796_),
    .C(_5798_),
    .Y(_5060_)
);

INVX1 _13351_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .Y(_5799_)
);

OR2X2 _13352_ (
    .A(_5795_),
    .B(_5105_),
    .Y(_5800_)
);

OAI21X1 _13353_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5801_)
);

OAI21X1 _13354_ (
    .A(_5799_),
    .B(_5800_),
    .C(_5801_),
    .Y(_5061_)
);

INVX1 _13355_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .Y(_5802_)
);

OAI21X1 _13356_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Xin12b [9]),
    .Y(_5803_)
);

OAI21X1 _13357_ (
    .A(_5802_),
    .B(_5800_),
    .C(_5803_),
    .Y(_5062_)
);

NAND2X1 _13358_ (
    .A(_5109_),
    .B(_5108_),
    .Y(_5804_)
);

NAND2X1 _13359_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(_5804_),
    .Y(_5805_)
);

OAI21X1 _13360_ (
    .A(_5799_),
    .B(_5804_),
    .C(_5805_),
    .Y(_5063_)
);

NAND2X1 _13361_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(_5804_),
    .Y(_5806_)
);

OAI21X1 _13362_ (
    .A(_5802_),
    .B(_5804_),
    .C(_5806_),
    .Y(_5064_)
);

AND2X2 _13363_ (
    .A(_5109_),
    .B(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5807_)
);

NAND2X1 _13364_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5807_),
    .Y(_5808_)
);

OAI21X1 _13365_ (
    .A(_5155_),
    .B(_5807_),
    .C(_5808_),
    .Y(_5065_)
);

NAND2X1 _13366_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5807_),
    .Y(_5809_)
);

OAI21X1 _13367_ (
    .A(_5192_),
    .B(_5807_),
    .C(_5809_),
    .Y(_5066_)
);

OAI21X1 _13368_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5810_)
);

OAI21X1 _13369_ (
    .A(_5799_),
    .B(_5104_),
    .C(_5810_),
    .Y(_5067_)
);

OAI21X1 _13370_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5811_)
);

OAI21X1 _13371_ (
    .A(_5802_),
    .B(_5104_),
    .C(_5811_),
    .Y(_5068_)
);

NAND2X1 _13372_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.X_ [0]),
    .Y(_5812_)
);

OAI21X1 _13373_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5162_),
    .C(_5812_),
    .Y(_5069_)
);

NAND2X1 _13374_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.X_ [1]),
    .Y(_5813_)
);

OAI21X1 _13375_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5199_),
    .C(_5813_),
    .Y(_5070_)
);

NAND2X1 _13376_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5796_),
    .Y(_5814_)
);

OAI21X1 _13377_ (
    .A(_5401_),
    .B(_5796_),
    .C(_5814_),
    .Y(_5071_)
);

NAND2X1 _13378_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5796_),
    .Y(_5815_)
);

OAI21X1 _13379_ (
    .A(_5427_),
    .B(_5796_),
    .C(_5815_),
    .Y(_5072_)
);

INVX1 _13380_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5816_)
);

OAI21X1 _13381_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5817_)
);

OAI21X1 _13382_ (
    .A(_5816_),
    .B(_5800_),
    .C(_5817_),
    .Y(_5073_)
);

INVX1 _13383_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5818_)
);

OAI21X1 _13384_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5819_)
);

OAI21X1 _13385_ (
    .A(_5818_),
    .B(_5800_),
    .C(_5819_),
    .Y(_5074_)
);

NAND2X1 _13386_ (
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .B(_5804_),
    .Y(_5820_)
);

OAI21X1 _13387_ (
    .A(_5816_),
    .B(_5804_),
    .C(_5820_),
    .Y(_5075_)
);

NAND2X1 _13388_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(_5804_),
    .Y(_5821_)
);

OAI21X1 _13389_ (
    .A(_5818_),
    .B(_5804_),
    .C(_5821_),
    .Y(_5076_)
);

NAND2X1 _13390_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5807_),
    .Y(_5822_)
);

OAI21X1 _13391_ (
    .A(_5271_),
    .B(_5807_),
    .C(_5822_),
    .Y(_5077_)
);

NAND2X1 _13392_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5807_),
    .Y(_5823_)
);

OAI21X1 _13393_ (
    .A(_5292_),
    .B(_5807_),
    .C(_5823_),
    .Y(_5078_)
);

OAI21X1 _13394_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5824_)
);

OAI21X1 _13395_ (
    .A(_5816_),
    .B(_5104_),
    .C(_5824_),
    .Y(_5079_)
);

OAI21X1 _13396_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5825_)
);

OAI21X1 _13397_ (
    .A(_5818_),
    .B(_5104_),
    .C(_5825_),
    .Y(_5080_)
);

NAND2X1 _13398_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5826_)
);

OAI21X1 _13399_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5149_),
    .C(_5826_),
    .Y(_5081_)
);

NAND2X1 _13400_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5827_)
);

OAI21X1 _13401_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5187_),
    .C(_5827_),
    .Y(_5082_)
);

NAND2X1 _13402_ (
    .A(\a[6] [0]),
    .B(_5796_),
    .Y(_5828_)
);

OAI21X1 _13403_ (
    .A(_5788_),
    .B(_5796_),
    .C(_5828_),
    .Y(_5083_)
);

NAND2X1 _13404_ (
    .A(\a[6] [1]),
    .B(_5796_),
    .Y(_5829_)
);

OAI21X1 _13405_ (
    .A(_5188__bF$buf1),
    .B(_5796_),
    .C(_5829_),
    .Y(_5084_)
);

INVX1 _13406_ (
    .A(\a[6] [0]),
    .Y(_5830_)
);

OAI21X1 _13407_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Ain12b [8]),
    .Y(_5831_)
);

OAI21X1 _13408_ (
    .A(_5830_),
    .B(_5800_),
    .C(_5831_),
    .Y(_5085_)
);

INVX1 _13409_ (
    .A(\a[6] [1]),
    .Y(_5832_)
);

OAI21X1 _13410_ (
    .A(_5105_),
    .B(_5795_),
    .C(\genblk1[6].u_ce.Ain12b [9]),
    .Y(_5833_)
);

OAI21X1 _13411_ (
    .A(_5832_),
    .B(_5800_),
    .C(_5833_),
    .Y(_5086_)
);

NAND2X1 _13412_ (
    .A(\genblk1[6].u_ce.Ain12b [6]),
    .B(_5804_),
    .Y(_5834_)
);

OAI21X1 _13413_ (
    .A(_5830_),
    .B(_5804_),
    .C(_5834_),
    .Y(_5087_)
);

NAND2X1 _13414_ (
    .A(\genblk1[6].u_ce.Ain12b [7]),
    .B(_5804_),
    .Y(_5095_)
);

OAI21X1 _13415_ (
    .A(_5832_),
    .B(_5804_),
    .C(_5095_),
    .Y(_5088_)
);

NAND2X1 _13416_ (
    .A(\a[6] [0]),
    .B(_5807_),
    .Y(_5096_)
);

OAI21X1 _13417_ (
    .A(_5719_),
    .B(_5807_),
    .C(_5096_),
    .Y(_5089_)
);

NAND2X1 _13418_ (
    .A(\a[6] [1]),
    .B(_5807_),
    .Y(_5097_)
);

OAI21X1 _13419_ (
    .A(_5728_),
    .B(_5807_),
    .C(_5097_),
    .Y(_5090_)
);

OAI21X1 _13420_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Ain1 [0]),
    .Y(_5098_)
);

OAI21X1 _13421_ (
    .A(_5830_),
    .B(_5104_),
    .C(_5098_),
    .Y(_5091_)
);

OAI21X1 _13422_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_5102_),
    .C(\genblk1[6].u_ce.Ain1 [1]),
    .Y(_5099_)
);

OAI21X1 _13423_ (
    .A(_5832_),
    .B(_5104_),
    .C(_5099_),
    .Y(_5092_)
);

NAND2X1 _13424_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\a[6] [0]),
    .Y(_5100_)
);

OAI21X1 _13425_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5680_),
    .C(_5100_),
    .Y(_5093_)
);

NAND2X1 _13426_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[6] [1]),
    .Y(_5101_)
);

OAI21X1 _13427_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5695_),
    .C(_5101_),
    .Y(_5094_)
);

DFFPOSX1 _13428_ (
    .CLK(clk_bF$buf75),
    .D(_5028_),
    .Q(\genblk1[6].u_ce.Ycalc [0])
);

DFFPOSX1 _13429_ (
    .CLK(clk_bF$buf74),
    .D(_5029_),
    .Q(\genblk1[6].u_ce.Ycalc [1])
);

DFFPOSX1 _13430_ (
    .CLK(clk_bF$buf73),
    .D(_5030_),
    .Q(\genblk1[6].u_ce.ISout )
);

DFFPOSX1 _13431_ (
    .CLK(clk_bF$buf72),
    .D(_5031_),
    .Q(\genblk1[6].u_ce.Ycalc [2])
);

DFFPOSX1 _13432_ (
    .CLK(clk_bF$buf71),
    .D(_5032_),
    .Q(\genblk1[6].u_ce.Ycalc [3])
);

DFFPOSX1 _13433_ (
    .CLK(clk_bF$buf70),
    .D(_5033_),
    .Q(\genblk1[6].u_ce.Ycalc [4])
);

DFFPOSX1 _13434_ (
    .CLK(clk_bF$buf69),
    .D(_5034_),
    .Q(\genblk1[6].u_ce.Ycalc [5])
);

DFFPOSX1 _13435_ (
    .CLK(clk_bF$buf68),
    .D(_5035_),
    .Q(\genblk1[6].u_ce.Ycalc [6])
);

DFFPOSX1 _13436_ (
    .CLK(clk_bF$buf67),
    .D(_5036_),
    .Q(\genblk1[6].u_ce.Ycalc [7])
);

DFFPOSX1 _13437_ (
    .CLK(clk_bF$buf66),
    .D(_5037_),
    .Q(\genblk1[6].u_ce.Ycalc [8])
);

DFFPOSX1 _13438_ (
    .CLK(clk_bF$buf65),
    .D(_5038_),
    .Q(\genblk1[6].u_ce.Ycalc [9])
);

DFFPOSX1 _13439_ (
    .CLK(clk_bF$buf64),
    .D(_5039_),
    .Q(\genblk1[6].u_ce.Ycalc [10])
);

DFFPOSX1 _13440_ (
    .CLK(clk_bF$buf63),
    .D(_5040_),
    .Q(\genblk1[6].u_ce.Ycalc [11])
);

DFFPOSX1 _13441_ (
    .CLK(clk_bF$buf62),
    .D(_5041_),
    .Q(\genblk1[6].u_ce.Xcalc [0])
);

DFFPOSX1 _13442_ (
    .CLK(clk_bF$buf61),
    .D(_5042_),
    .Q(\genblk1[6].u_ce.Xcalc [1])
);

DFFPOSX1 _13443_ (
    .CLK(clk_bF$buf60),
    .D(_5043_),
    .Q(\genblk1[6].u_ce.Xcalc [2])
);

DFFPOSX1 _13444_ (
    .CLK(clk_bF$buf59),
    .D(_5044_),
    .Q(\genblk1[6].u_ce.Xcalc [3])
);

DFFPOSX1 _13445_ (
    .CLK(clk_bF$buf58),
    .D(_5045_),
    .Q(\genblk1[6].u_ce.Xcalc [4])
);

DFFPOSX1 _13446_ (
    .CLK(clk_bF$buf57),
    .D(_5046_),
    .Q(\genblk1[6].u_ce.Xcalc [5])
);

DFFPOSX1 _13447_ (
    .CLK(clk_bF$buf56),
    .D(_5047_),
    .Q(\genblk1[6].u_ce.Xcalc [6])
);

DFFPOSX1 _13448_ (
    .CLK(clk_bF$buf55),
    .D(_5048_),
    .Q(\genblk1[6].u_ce.Xcalc [7])
);

DFFPOSX1 _13449_ (
    .CLK(clk_bF$buf54),
    .D(_5049_),
    .Q(\genblk1[6].u_ce.Xcalc [8])
);

DFFPOSX1 _13450_ (
    .CLK(clk_bF$buf53),
    .D(_5050_),
    .Q(\genblk1[6].u_ce.Xcalc [9])
);

DFFPOSX1 _13451_ (
    .CLK(clk_bF$buf52),
    .D(_5051_),
    .Q(\genblk1[6].u_ce.Xcalc [10])
);

DFFPOSX1 _13452_ (
    .CLK(clk_bF$buf51),
    .D(_5052_),
    .Q(\genblk1[6].u_ce.Xcalc [11])
);

DFFPOSX1 _13453_ (
    .CLK(clk_bF$buf50),
    .D(_5053_),
    .Q(\genblk1[6].u_ce.Acalc [1])
);

DFFPOSX1 _13454_ (
    .CLK(clk_bF$buf49),
    .D(_5054_),
    .Q(\genblk1[6].u_ce.Acalc [3])
);

DFFPOSX1 _13455_ (
    .CLK(clk_bF$buf48),
    .D(_5055_),
    .Q(\genblk1[6].u_ce.Acalc [5])
);

DFFPOSX1 _13456_ (
    .CLK(clk_bF$buf47),
    .D(_5056_),
    .Q(\genblk1[6].u_ce.Acalc [7])
);

DFFPOSX1 _13457_ (
    .CLK(clk_bF$buf46),
    .D(_5057_),
    .Q(\genblk1[6].u_ce.Acalc [9])
);

DFFPOSX1 _13458_ (
    .CLK(clk_bF$buf45),
    .D(_5058_),
    .Q(\genblk1[6].u_ce.Acalc [11])
);

DFFPOSX1 _13459_ (
    .CLK(clk_bF$buf44),
    .D(_5059_),
    .Q(\genblk1[6].u_ce.Xin12b [10])
);

DFFPOSX1 _13460_ (
    .CLK(clk_bF$buf43),
    .D(_5060_),
    .Q(\genblk1[6].u_ce.Xin12b [11])
);

DFFPOSX1 _13461_ (
    .CLK(clk_bF$buf42),
    .D(_5061_),
    .Q(\genblk1[6].u_ce.Xin12b [8])
);

DFFPOSX1 _13462_ (
    .CLK(clk_bF$buf41),
    .D(_5062_),
    .Q(\genblk1[6].u_ce.Xin12b [9])
);

DFFPOSX1 _13463_ (
    .CLK(clk_bF$buf40),
    .D(_5063_),
    .Q(\genblk1[6].u_ce.Xin12b [6])
);

DFFPOSX1 _13464_ (
    .CLK(clk_bF$buf39),
    .D(_5064_),
    .Q(\genblk1[6].u_ce.Xin12b [7])
);

DFFPOSX1 _13465_ (
    .CLK(clk_bF$buf38),
    .D(_5065_),
    .Q(\genblk1[6].u_ce.Xin12b [4])
);

DFFPOSX1 _13466_ (
    .CLK(clk_bF$buf37),
    .D(_5066_),
    .Q(\genblk1[6].u_ce.Xin12b [5])
);

DFFPOSX1 _13467_ (
    .CLK(clk_bF$buf36),
    .D(_5067_),
    .Q(\genblk1[6].u_ce.Xin1 [0])
);

DFFPOSX1 _13468_ (
    .CLK(clk_bF$buf35),
    .D(_5068_),
    .Q(\genblk1[6].u_ce.Xin1 [1])
);

DFFPOSX1 _13469_ (
    .CLK(clk_bF$buf34),
    .D(_5069_),
    .Q(\genblk1[6].u_ce.Xin0 [0])
);

DFFPOSX1 _13470_ (
    .CLK(clk_bF$buf33),
    .D(_5070_),
    .Q(\genblk1[6].u_ce.Xin0 [1])
);

DFFPOSX1 _13471_ (
    .CLK(clk_bF$buf32),
    .D(_5071_),
    .Q(\genblk1[6].u_ce.Yin12b [10])
);

DFFPOSX1 _13472_ (
    .CLK(clk_bF$buf31),
    .D(_5072_),
    .Q(\genblk1[6].u_ce.Yin12b [11])
);

DFFPOSX1 _13473_ (
    .CLK(clk_bF$buf30),
    .D(_5073_),
    .Q(\genblk1[6].u_ce.Yin12b [8])
);

DFFPOSX1 _13474_ (
    .CLK(clk_bF$buf29),
    .D(_5074_),
    .Q(\genblk1[6].u_ce.Yin12b [9])
);

DFFPOSX1 _13475_ (
    .CLK(clk_bF$buf28),
    .D(_5075_),
    .Q(\genblk1[6].u_ce.Yin12b [6])
);

DFFPOSX1 _13476_ (
    .CLK(clk_bF$buf27),
    .D(_5076_),
    .Q(\genblk1[6].u_ce.Yin12b [7])
);

DFFPOSX1 _13477_ (
    .CLK(clk_bF$buf26),
    .D(_5077_),
    .Q(\genblk1[6].u_ce.Yin12b [4])
);

DFFPOSX1 _13478_ (
    .CLK(clk_bF$buf25),
    .D(_5078_),
    .Q(\genblk1[6].u_ce.Yin12b [5])
);

DFFPOSX1 _13479_ (
    .CLK(clk_bF$buf24),
    .D(_5079_),
    .Q(\genblk1[6].u_ce.Yin1 [0])
);

DFFPOSX1 _13480_ (
    .CLK(clk_bF$buf23),
    .D(_5080_),
    .Q(\genblk1[6].u_ce.Yin1 [1])
);

DFFPOSX1 _13481_ (
    .CLK(clk_bF$buf22),
    .D(_5081_),
    .Q(\genblk1[6].u_ce.Yin0 [0])
);

DFFPOSX1 _13482_ (
    .CLK(clk_bF$buf21),
    .D(_5082_),
    .Q(\genblk1[6].u_ce.Yin0 [1])
);

DFFPOSX1 _13483_ (
    .CLK(clk_bF$buf20),
    .D(_5083_),
    .Q(\genblk1[6].u_ce.Ain12b [10])
);

DFFPOSX1 _13484_ (
    .CLK(clk_bF$buf19),
    .D(_5084_),
    .Q(\genblk1[6].u_ce.Ain12b [11])
);

DFFPOSX1 _13485_ (
    .CLK(clk_bF$buf18),
    .D(_5085_),
    .Q(\genblk1[6].u_ce.Ain12b [8])
);

DFFPOSX1 _13486_ (
    .CLK(clk_bF$buf17),
    .D(_5086_),
    .Q(\genblk1[6].u_ce.Ain12b [9])
);

DFFPOSX1 _13487_ (
    .CLK(clk_bF$buf16),
    .D(_5087_),
    .Q(\genblk1[6].u_ce.Ain12b [6])
);

DFFPOSX1 _13488_ (
    .CLK(clk_bF$buf15),
    .D(_5088_),
    .Q(\genblk1[6].u_ce.Ain12b [7])
);

DFFPOSX1 _13489_ (
    .CLK(clk_bF$buf14),
    .D(_5089_),
    .Q(\genblk1[6].u_ce.Ain12b [4])
);

DFFPOSX1 _13490_ (
    .CLK(clk_bF$buf13),
    .D(_5090_),
    .Q(\genblk1[6].u_ce.Ain12b [5])
);

DFFPOSX1 _13491_ (
    .CLK(clk_bF$buf12),
    .D(_5091_),
    .Q(\genblk1[6].u_ce.Ain1 [0])
);

DFFPOSX1 _13492_ (
    .CLK(clk_bF$buf11),
    .D(_5092_),
    .Q(\genblk1[6].u_ce.Ain1 [1])
);

DFFPOSX1 _13493_ (
    .CLK(clk_bF$buf10),
    .D(_5093_),
    .Q(\genblk1[6].u_ce.Ain0 [0])
);

DFFPOSX1 _13494_ (
    .CLK(clk_bF$buf9),
    .D(_5094_),
    .Q(\genblk1[6].u_ce.Ain0 [1])
);

DFFPOSX1 _13495_ (
    .CLK(clk_bF$buf8),
    .D(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[6].u_ce.LoadCtl [0])
);

DFFPOSX1 _13496_ (
    .CLK(clk_bF$buf7),
    .D(\genblk1[6].u_ce.LoadCtl_0_bF$buf4 ),
    .Q(\genblk1[6].u_ce.LoadCtl [1])
);

DFFPOSX1 _13497_ (
    .CLK(clk_bF$buf6),
    .D(\genblk1[6].u_ce.LoadCtl [1]),
    .Q(\genblk1[6].u_ce.LoadCtl [2])
);

DFFPOSX1 _13498_ (
    .CLK(clk_bF$buf5),
    .D(\genblk1[6].u_ce.LoadCtl [2]),
    .Q(\genblk1[6].u_ce.LoadCtl [3])
);

DFFPOSX1 _13499_ (
    .CLK(clk_bF$buf4),
    .D(\genblk1[6].u_ce.LoadCtl [3]),
    .Q(\genblk1[6].u_ce.LoadCtl [4])
);

DFFPOSX1 _13500_ (
    .CLK(clk_bF$buf3),
    .D(\genblk1[6].u_ce.LoadCtl [4]),
    .Q(\genblk1[6].u_ce.LoadCtl [5])
);

DFFPOSX1 _13501_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[6].u_ce.LoadCtl [5]),
    .Q(\genblk1[6].u_ce.Vld )
);

INVX2 _13502_ (
    .A(\genblk1[7].u_ce.LoadCtl [1]),
    .Y(_5885_)
);

NOR2X1 _13503_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5885_),
    .Y(_5886_)
);

INVX2 _13504_ (
    .A(_5886_),
    .Y(_5887_)
);

INVX2 _13505_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .Y(_5888_)
);

NOR2X1 _13506_ (
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .B(\genblk1[7].u_ce.LoadCtl [3]),
    .Y(_5889_)
);

INVX1 _13507_ (
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .Y(_5890_)
);

AND2X2 _13508_ (
    .A(_5890_),
    .B(\genblk1[7].u_ce.LoadCtl [3]),
    .Y(_5891_)
);

NOR2X1 _13509_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[7].u_ce.LoadCtl [1]),
    .Y(_5892_)
);

INVX1 _13510_ (
    .A(\genblk1[7].u_ce.Ycalc [10]),
    .Y(_5893_)
);

OAI21X1 _13511_ (
    .A(_5888_),
    .B(\genblk1[7].u_ce.Ycalc [8]),
    .C(_5889_),
    .Y(_5894_)
);

AOI21X1 _13512_ (
    .A(_5888_),
    .B(_5893_),
    .C(_5894_),
    .Y(_5895_)
);

INVX1 _13513_ (
    .A(\genblk1[7].u_ce.Ycalc [4]),
    .Y(_5896_)
);

NAND2X1 _13514_ (
    .A(\genblk1[7].u_ce.Ycalc [6]),
    .B(_5891_),
    .Y(_5897_)
);

OAI21X1 _13515_ (
    .A(_5890_),
    .B(_5896_),
    .C(_5897_),
    .Y(_5898_)
);

OAI21X1 _13516_ (
    .A(_5895_),
    .B(_5898_),
    .C(_5892_),
    .Y(_5899_)
);

AOI22X1 _13517_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[7].u_ce.Ycalc [0]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Ycalc [2]),
    .Y(_5900_)
);

NAND2X1 _13518_ (
    .A(_5900_),
    .B(_5899_),
    .Y(\genblk1[7].u_ce.Y_ [0])
);

INVX1 _13519_ (
    .A(\genblk1[7].u_ce.Ycalc [9]),
    .Y(_5901_)
);

OAI21X1 _13520_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Ycalc [11]),
    .C(_5889_),
    .Y(_5902_)
);

AOI21X1 _13521_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(_5901_),
    .C(_5902_),
    .Y(_5903_)
);

INVX1 _13522_ (
    .A(\genblk1[7].u_ce.Ycalc [5]),
    .Y(_5904_)
);

NAND2X1 _13523_ (
    .A(\genblk1[7].u_ce.Ycalc [7]),
    .B(_5891_),
    .Y(_5905_)
);

OAI21X1 _13524_ (
    .A(_5890_),
    .B(_5904_),
    .C(_5905_),
    .Y(_5906_)
);

OAI21X1 _13525_ (
    .A(_5903_),
    .B(_5906_),
    .C(_5892_),
    .Y(_5907_)
);

AOI22X1 _13526_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[7].u_ce.Ycalc [1]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Ycalc [3]),
    .Y(_5908_)
);

NAND2X1 _13527_ (
    .A(_5908_),
    .B(_5907_),
    .Y(\genblk1[7].u_ce.Y_ [1])
);

INVX1 _13528_ (
    .A(\genblk1[7].u_ce.Xcalc [8]),
    .Y(_5909_)
);

OAI21X1 _13529_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Xcalc [10]),
    .C(_5889_),
    .Y(_5910_)
);

AOI21X1 _13530_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(_5909_),
    .C(_5910_),
    .Y(_5911_)
);

INVX1 _13531_ (
    .A(\genblk1[7].u_ce.Xcalc [4]),
    .Y(_5912_)
);

NAND2X1 _13532_ (
    .A(\genblk1[7].u_ce.Xcalc [6]),
    .B(_5891_),
    .Y(_5913_)
);

OAI21X1 _13533_ (
    .A(_5890_),
    .B(_5912_),
    .C(_5913_),
    .Y(_5914_)
);

OAI21X1 _13534_ (
    .A(_5911_),
    .B(_5914_),
    .C(_5892_),
    .Y(_5915_)
);

AOI22X1 _13535_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[7].u_ce.Xcalc [0]),
    .C(_5886_),
    .D(\genblk1[7].u_ce.Xcalc [2]),
    .Y(_5916_)
);

NAND2X1 _13536_ (
    .A(_5916_),
    .B(_5915_),
    .Y(\genblk1[7].u_ce.X_ [0])
);

INVX1 _13537_ (
    .A(\genblk1[7].u_ce.Xcalc [3]),
    .Y(_5917_)
);

NOR2X1 _13538_ (
    .A(\genblk1[7].u_ce.LoadCtl [4]),
    .B(\genblk1[7].u_ce.Xcalc [11]),
    .Y(_5918_)
);

OAI21X1 _13539_ (
    .A(_5888_),
    .B(\genblk1[7].u_ce.Xcalc [9]),
    .C(_5889_),
    .Y(_5919_)
);

AOI22X1 _13540_ (
    .A(\genblk1[7].u_ce.LoadCtl [2]),
    .B(\genblk1[7].u_ce.Xcalc [5]),
    .C(_5891_),
    .D(\genblk1[7].u_ce.Xcalc [7]),
    .Y(_5920_)
);

OAI21X1 _13541_ (
    .A(_5918_),
    .B(_5919_),
    .C(_5920_),
    .Y(_5921_)
);

AOI22X1 _13542_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[7].u_ce.Xcalc [1]),
    .C(_5921_),
    .D(_5892_),
    .Y(_5922_)
);

OAI21X1 _13543_ (
    .A(_5917_),
    .B(_5887_),
    .C(_5922_),
    .Y(\genblk1[7].u_ce.X_ [1])
);

INVX1 _13544_ (
    .A(\genblk1[7].u_ce.Ycalc [0]),
    .Y(_5923_)
);

INVX1 _13545_ (
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .Y(_5924_)
);

INVX4 _13546_ (
    .A(1'h1),
    .Y(_5925_)
);

INVX8 _13547_ (
    .A(1'h1),
    .Y(_5926_)
);

INVX1 _13548_ (
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .Y(_5927_)
);

NAND2X1 _13549_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [7]),
    .Y(_5928_)
);

OAI21X1 _13550_ (
    .A(1'h1),
    .B(_5927_),
    .C(_5928_),
    .Y(_5929_)
);

INVX1 _13551_ (
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .Y(_5930_)
);

NAND2X1 _13552_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [5]),
    .Y(_5931_)
);

OAI21X1 _13553_ (
    .A(1'h1),
    .B(_5930_),
    .C(_5931_),
    .Y(_5932_)
);

MUX2X1 _13554_ (
    .A(_5932_),
    .B(_5929_),
    .S(_5926__bF$buf4),
    .Y(_5933_)
);

INVX1 _13555_ (
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_5934_)
);

NAND2X1 _13556_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_5935_)
);

OAI21X1 _13557_ (
    .A(1'h1),
    .B(_5934_),
    .C(_5935_),
    .Y(_5936_)
);

INVX1 _13558_ (
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .Y(_5937_)
);

NAND2X1 _13559_ (
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_5938_)
);

OAI21X1 _13560_ (
    .A(1'h1),
    .B(_5937_),
    .C(_5938_),
    .Y(_5939_)
);

MUX2X1 _13561_ (
    .A(_5939_),
    .B(_5936_),
    .S(_5926__bF$buf3),
    .Y(_5940_)
);

MUX2X1 _13562_ (
    .A(_5940_),
    .B(_5933_),
    .S(_5925__bF$buf3),
    .Y(_5941_)
);

NOR2X1 _13563_ (
    .A(_5924_),
    .B(_5941_),
    .Y(_5942_)
);

NAND2X1 _13564_ (
    .A(_5924_),
    .B(_5941_),
    .Y(_5943_)
);

INVX1 _13565_ (
    .A(_5943_),
    .Y(_5944_)
);

NAND2X1 _13566_ (
    .A(_5925__bF$buf2),
    .B(_5926__bF$buf2),
    .Y(_5945_)
);

OAI21X1 _13567_ (
    .A(1'h1),
    .B(_5945_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_5946_)
);

INVX2 _13568_ (
    .A(_5946_),
    .Y(_5947_)
);

OAI21X1 _13569_ (
    .A(_5942_),
    .B(_5944_),
    .C(_5947_),
    .Y(_5948_)
);

OAI21X1 _13570_ (
    .A(_5923_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_5948_),
    .Y(_5835_)
);

INVX4 _13571_ (
    .A(\genblk1[7].u_ce.Vld ),
    .Y(_5949_)
);

NAND2X1 _13572_ (
    .A(\genblk1[7].u_ce.Ycalc [1]),
    .B(_5949__bF$buf3),
    .Y(_5950_)
);

NOR2X1 _13573_ (
    .A(1'h1),
    .B(_5945_),
    .Y(_5951_)
);

MUX2X1 _13574_ (
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(\genblk1[7].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_5952_)
);

MUX2X1 _13575_ (
    .A(\genblk1[7].u_ce.Xin12b [5]),
    .B(\genblk1[7].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_5953_)
);

MUX2X1 _13576_ (
    .A(_5953_),
    .B(_5952_),
    .S(_5926__bF$buf1),
    .Y(_5954_)
);

INVX1 _13577_ (
    .A(1'h1),
    .Y(_5955_)
);

NAND2X1 _13578_ (
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(_5955_),
    .Y(_5956_)
);

AOI21X1 _13579_ (
    .A(_5956_),
    .B(_5935_),
    .C(_5926__bF$buf0),
    .Y(_5957_)
);

NAND3X1 _13580_ (
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .B(_5955_),
    .C(_5926__bF$buf4),
    .Y(_5958_)
);

NAND3X1 _13581_ (
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .B(1'h1),
    .C(_5926__bF$buf3),
    .Y(_5959_)
);

NAND3X1 _13582_ (
    .A(_5925__bF$buf1),
    .B(_5959_),
    .C(_5958_),
    .Y(_5960_)
);

OAI22X1 _13583_ (
    .A(_5957_),
    .B(_5960_),
    .C(_5925__bF$buf0),
    .D(_5954_),
    .Y(_5961_)
);

INVX1 _13584_ (
    .A(\genblk1[7].u_ce.Yin0 [1]),
    .Y(_5962_)
);

INVX8 _13585_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_5963_)
);

INVX1 _13586_ (
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .Y(_5964_)
);

NAND2X1 _13587_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_5965_)
);

OAI21X1 _13588_ (
    .A(1'h1),
    .B(_5964_),
    .C(_5965_),
    .Y(_5966_)
);

INVX1 _13589_ (
    .A(\genblk1[7].u_ce.Xin12b [5]),
    .Y(_5967_)
);

NAND2X1 _13590_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [6]),
    .Y(_5968_)
);

OAI21X1 _13591_ (
    .A(1'h1),
    .B(_5967_),
    .C(_5968_),
    .Y(_5969_)
);

MUX2X1 _13592_ (
    .A(_5969_),
    .B(_5966_),
    .S(_5926__bF$buf2),
    .Y(_5970_)
);

INVX1 _13593_ (
    .A(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_5971_)
);

NAND2X1 _13594_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [4]),
    .Y(_5972_)
);

OAI21X1 _13595_ (
    .A(1'h1),
    .B(_5971_),
    .C(_5972_),
    .Y(_5973_)
);

INVX1 _13596_ (
    .A(\genblk1[7].u_ce.Xin0 [1]),
    .Y(_5974_)
);

NAND2X1 _13597_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_5975_)
);

OAI21X1 _13598_ (
    .A(1'h1),
    .B(_5974_),
    .C(_5975_),
    .Y(_5976_)
);

MUX2X1 _13599_ (
    .A(_5976_),
    .B(_5973_),
    .S(_5926__bF$buf1),
    .Y(_5977_)
);

MUX2X1 _13600_ (
    .A(_5977_),
    .B(_5970_),
    .S(_5925__bF$buf3),
    .Y(_5978_)
);

NAND3X1 _13601_ (
    .A(_5963__bF$buf5),
    .B(_5941_),
    .C(_5978_),
    .Y(_5979_)
);

MUX2X1 _13602_ (
    .A(\genblk1[7].u_ce.Xin12b [8]),
    .B(\genblk1[7].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_5980_)
);

MUX2X1 _13603_ (
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(\genblk1[7].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_5981_)
);

MUX2X1 _13604_ (
    .A(_5981_),
    .B(_5980_),
    .S(_5926__bF$buf0),
    .Y(_5982_)
);

MUX2X1 _13605_ (
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .B(\genblk1[7].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_5983_)
);

MUX2X1 _13606_ (
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(\genblk1[7].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_5984_)
);

MUX2X1 _13607_ (
    .A(_5984_),
    .B(_5983_),
    .S(_5926__bF$buf4),
    .Y(_5985_)
);

MUX2X1 _13608_ (
    .A(_5985_),
    .B(_5982_),
    .S(_5925__bF$buf2),
    .Y(_5986_)
);

OAI21X1 _13609_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5961_),
    .C(_5986_),
    .Y(_5987_)
);

AOI21X1 _13610_ (
    .A(_5987_),
    .B(_5979_),
    .C(_5962_),
    .Y(_5988_)
);

INVX1 _13611_ (
    .A(_5988_),
    .Y(_5989_)
);

NAND3X1 _13612_ (
    .A(_5962_),
    .B(_5979_),
    .C(_5987_),
    .Y(_5990_)
);

AND2X2 _13613_ (
    .A(_5989_),
    .B(_5990_),
    .Y(_5991_)
);

OAI21X1 _13614_ (
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .B(_5961_),
    .C(_5991_),
    .Y(_5992_)
);

OR2X2 _13615_ (
    .A(_5991_),
    .B(_5943_),
    .Y(_5993_)
);

AOI21X1 _13616_ (
    .A(_5993_),
    .B(_5992_),
    .C(_5951_),
    .Y(_5994_)
);

OAI21X1 _13617_ (
    .A(_5949__bF$buf2),
    .B(_5994_),
    .C(_5950_),
    .Y(_5836_)
);

INVX1 _13618_ (
    .A(\genblk1[7].u_ce.ISout ),
    .Y(_5995_)
);

NAND2X1 _13619_ (
    .A(\genblk1[7].u_ce.Vld ),
    .B(\genblk1[6].u_ce.ISout ),
    .Y(_5996_)
);

OAI21X1 _13620_ (
    .A(\genblk1[7].u_ce.Vld ),
    .B(_5995_),
    .C(_5996_),
    .Y(_5837_)
);

NAND2X1 _13621_ (
    .A(\genblk1[7].u_ce.Ycalc [2]),
    .B(_5949__bF$buf1),
    .Y(_5997_)
);

AOI21X1 _13622_ (
    .A(_5943_),
    .B(_5990_),
    .C(_5988_),
    .Y(_5998_)
);

MUX2X1 _13623_ (
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .B(\genblk1[7].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_5999_)
);

MUX2X1 _13624_ (
    .A(_5999_),
    .B(_5952_),
    .S(1'h1),
    .Y(_6000_)
);

MUX2X1 _13625_ (
    .A(\genblk1[7].u_ce.Xin1 [1]),
    .B(\genblk1[7].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_6001_)
);

NAND2X1 _13626_ (
    .A(1'h1),
    .B(_5925__bF$buf1),
    .Y(_6002_)
);

OAI22X1 _13627_ (
    .A(_6002_),
    .B(_5953_),
    .C(_6001_),
    .D(_5945_),
    .Y(_6003_)
);

AOI21X1 _13628_ (
    .A(1'h1),
    .B(_6000_),
    .C(_6003_),
    .Y(_6004_)
);

AOI21X1 _13629_ (
    .A(_5986_),
    .B(_5961_),
    .C(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_6005_)
);

NAND2X1 _13630_ (
    .A(_6004_),
    .B(_6005_),
    .Y(_6006_)
);

INVX1 _13631_ (
    .A(_6004_),
    .Y(_6007_)
);

OAI21X1 _13632_ (
    .A(_5941_),
    .B(_5978_),
    .C(_5963__bF$buf4),
    .Y(_6008_)
);

NAND2X1 _13633_ (
    .A(_6007_),
    .B(_6008_),
    .Y(_6009_)
);

AOI21X1 _13634_ (
    .A(_6009_),
    .B(_6006_),
    .C(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6010_)
);

NAND3X1 _13635_ (
    .A(\genblk1[7].u_ce.Yin1 [0]),
    .B(_6006_),
    .C(_6009_),
    .Y(_6011_)
);

INVX1 _13636_ (
    .A(_6011_),
    .Y(_6012_)
);

OR2X2 _13637_ (
    .A(_6012_),
    .B(_6010_),
    .Y(_6013_)
);

NOR2X1 _13638_ (
    .A(_5998_),
    .B(_6013_),
    .Y(_6014_)
);

INVX1 _13639_ (
    .A(_6014_),
    .Y(_6015_)
);

OAI21X1 _13640_ (
    .A(_6010_),
    .B(_6012_),
    .C(_5998_),
    .Y(_6016_)
);

AOI21X1 _13641_ (
    .A(_6015_),
    .B(_6016_),
    .C(_5951_),
    .Y(_6017_)
);

INVX2 _13642_ (
    .A(_5951_),
    .Y(_6018_)
);

OAI21X1 _13643_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6018_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_6019_)
);

OAI21X1 _13644_ (
    .A(_6019_),
    .B(_6017_),
    .C(_5997_),
    .Y(_5838_)
);

INVX1 _13645_ (
    .A(\genblk1[7].u_ce.Ycalc [3]),
    .Y(_6020_)
);

INVX2 _13646_ (
    .A(_6019_),
    .Y(_6021_)
);

OAI21X1 _13647_ (
    .A(_6010_),
    .B(_5998_),
    .C(_6011_),
    .Y(_6022_)
);

INVX1 _13648_ (
    .A(_6022_),
    .Y(_6023_)
);

INVX1 _13649_ (
    .A(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6024_)
);

NAND3X1 _13650_ (
    .A(_5961_),
    .B(_5986_),
    .C(_6004_),
    .Y(_6025_)
);

INVX1 _13651_ (
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .Y(_6026_)
);

NAND2X1 _13652_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [10]),
    .Y(_6027_)
);

OAI21X1 _13653_ (
    .A(1'h1),
    .B(_6026_),
    .C(_6027_),
    .Y(_6028_)
);

NAND2X1 _13654_ (
    .A(_5926__bF$buf3),
    .B(_5980_),
    .Y(_6029_)
);

OAI21X1 _13655_ (
    .A(_5926__bF$buf2),
    .B(_6028_),
    .C(_6029_),
    .Y(_6030_)
);

NOR2X1 _13656_ (
    .A(1'h1),
    .B(_5926__bF$buf1),
    .Y(_6031_)
);

NOR2X1 _13657_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_6032_)
);

AOI22X1 _13658_ (
    .A(_5973_),
    .B(_6032_),
    .C(_6031_),
    .D(_5969_),
    .Y(_6033_)
);

OAI21X1 _13659_ (
    .A(_5925__bF$buf0),
    .B(_6030_),
    .C(_6033_),
    .Y(_6034_)
);

NAND3X1 _13660_ (
    .A(_5963__bF$buf3),
    .B(_6034_),
    .C(_6025_),
    .Y(_6035_)
);

INVX1 _13661_ (
    .A(_6025_),
    .Y(_6036_)
);

INVX1 _13662_ (
    .A(_6034_),
    .Y(_6037_)
);

OAI21X1 _13663_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6036_),
    .C(_6037_),
    .Y(_6038_)
);

NAND3X1 _13664_ (
    .A(_6024_),
    .B(_6035_),
    .C(_6038_),
    .Y(_6039_)
);

AOI21X1 _13665_ (
    .A(_6038_),
    .B(_6035_),
    .C(_6024_),
    .Y(_6040_)
);

INVX1 _13666_ (
    .A(_6040_),
    .Y(_6041_)
);

NAND2X1 _13667_ (
    .A(_6039_),
    .B(_6041_),
    .Y(_6042_)
);

AOI21X1 _13668_ (
    .A(_6042_),
    .B(_6023_),
    .C(_5951_),
    .Y(_6043_)
);

OAI21X1 _13669_ (
    .A(_6023_),
    .B(_6042_),
    .C(_6043_),
    .Y(_6044_)
);

AOI22X1 _13670_ (
    .A(_6020_),
    .B(_5949__bF$buf0),
    .C(_6044_),
    .D(_6021_),
    .Y(_5839_)
);

AOI21X1 _13671_ (
    .A(_6022_),
    .B(_6039_),
    .C(_6040_),
    .Y(_6045_)
);

INVX1 _13672_ (
    .A(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6046_)
);

INVX1 _13673_ (
    .A(\genblk1[7].u_ce.Xin12b [10]),
    .Y(_6047_)
);

NAND2X1 _13674_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6048_)
);

OAI21X1 _13675_ (
    .A(1'h1),
    .B(_6047_),
    .C(_6048_),
    .Y(_6049_)
);

NAND2X1 _13676_ (
    .A(_5926__bF$buf0),
    .B(_5999_),
    .Y(_6050_)
);

OAI21X1 _13677_ (
    .A(_5926__bF$buf4),
    .B(_6049_),
    .C(_6050_),
    .Y(_6051_)
);

NAND2X1 _13678_ (
    .A(_5925__bF$buf3),
    .B(_5954_),
    .Y(_6052_)
);

OAI21X1 _13679_ (
    .A(_5925__bF$buf2),
    .B(_6051_),
    .C(_6052_),
    .Y(_6053_)
);

INVX2 _13680_ (
    .A(_6053_),
    .Y(_6054_)
);

OAI21X1 _13681_ (
    .A(_6034_),
    .B(_6025_),
    .C(_5963__bF$buf2),
    .Y(_6055_)
);

OR2X2 _13682_ (
    .A(_6055_),
    .B(_6054_),
    .Y(_6056_)
);

NOR2X1 _13683_ (
    .A(_6034_),
    .B(_6025_),
    .Y(_6057_)
);

OAI21X1 _13684_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_6057_),
    .C(_6054_),
    .Y(_6058_)
);

NAND3X1 _13685_ (
    .A(_6046_),
    .B(_6058_),
    .C(_6056_),
    .Y(_6059_)
);

NOR2X1 _13686_ (
    .A(_6054_),
    .B(_6055_),
    .Y(_6060_)
);

AND2X2 _13687_ (
    .A(_6055_),
    .B(_6054_),
    .Y(_6061_)
);

OAI21X1 _13688_ (
    .A(_6060_),
    .B(_6061_),
    .C(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6062_)
);

NAND2X1 _13689_ (
    .A(_6062_),
    .B(_6059_),
    .Y(_6063_)
);

AOI21X1 _13690_ (
    .A(_6045_),
    .B(_6063_),
    .C(_5951_),
    .Y(_6064_)
);

OAI21X1 _13691_ (
    .A(_6045_),
    .B(_6063_),
    .C(_6064_),
    .Y(_6065_)
);

AOI22X1 _13692_ (
    .A(_5896_),
    .B(_5949__bF$buf3),
    .C(_6065_),
    .D(_6021_),
    .Y(_5840_)
);

OAI21X1 _13693_ (
    .A(_6063_),
    .B(_6045_),
    .C(_6062_),
    .Y(_6066_)
);

INVX1 _13694_ (
    .A(\genblk1[7].u_ce.Yin12b [5]),
    .Y(_6067_)
);

NAND3X1 _13695_ (
    .A(_6037_),
    .B(_6054_),
    .C(_6036_),
    .Y(_6068_)
);

NAND2X1 _13696_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6069_)
);

INVX1 _13697_ (
    .A(_6069_),
    .Y(_6070_)
);

AOI21X1 _13698_ (
    .A(_6028_),
    .B(_5926__bF$buf3),
    .C(_6070_),
    .Y(_6071_)
);

NAND2X1 _13699_ (
    .A(_5925__bF$buf1),
    .B(_5982_),
    .Y(_6072_)
);

OAI21X1 _13700_ (
    .A(_5925__bF$buf0),
    .B(_6071_),
    .C(_6072_),
    .Y(_6073_)
);

NAND3X1 _13701_ (
    .A(_5963__bF$buf1),
    .B(_6073_),
    .C(_6068_),
    .Y(_6074_)
);

NOR3X1 _13702_ (
    .A(_6034_),
    .B(_6053_),
    .C(_6025_),
    .Y(_6075_)
);

INVX1 _13703_ (
    .A(_6073_),
    .Y(_6076_)
);

OAI21X1 _13704_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6075_),
    .C(_6076_),
    .Y(_6077_)
);

NAND3X1 _13705_ (
    .A(_6067_),
    .B(_6074_),
    .C(_6077_),
    .Y(_6078_)
);

AOI21X1 _13706_ (
    .A(_6077_),
    .B(_6074_),
    .C(_6067_),
    .Y(_6079_)
);

INVX1 _13707_ (
    .A(_6079_),
    .Y(_6080_)
);

NAND2X1 _13708_ (
    .A(_6078_),
    .B(_6080_),
    .Y(_6081_)
);

AND2X2 _13709_ (
    .A(_6066_),
    .B(_6081_),
    .Y(_6082_)
);

OAI21X1 _13710_ (
    .A(_6081_),
    .B(_6066_),
    .C(_6018_),
    .Y(_6083_)
);

OAI21X1 _13711_ (
    .A(_6083_),
    .B(_6082_),
    .C(_6021_),
    .Y(_6084_)
);

OAI21X1 _13712_ (
    .A(_5904_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6084_),
    .Y(_5841_)
);

INVX1 _13713_ (
    .A(\genblk1[7].u_ce.Ycalc [6]),
    .Y(_6085_)
);

INVX1 _13714_ (
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .Y(_6086_)
);

NAND3X1 _13715_ (
    .A(_6054_),
    .B(_6076_),
    .C(_6057_),
    .Y(_6087_)
);

AOI21X1 _13716_ (
    .A(_6049_),
    .B(_5926__bF$buf2),
    .C(_6070_),
    .Y(_6088_)
);

NAND2X1 _13717_ (
    .A(_5925__bF$buf3),
    .B(_6000_),
    .Y(_6089_)
);

OAI21X1 _13718_ (
    .A(_5925__bF$buf2),
    .B(_6088_),
    .C(_6089_),
    .Y(_6090_)
);

NAND3X1 _13719_ (
    .A(_5963__bF$buf0),
    .B(_6090_),
    .C(_6087_),
    .Y(_6091_)
);

INVX1 _13720_ (
    .A(_6090_),
    .Y(_6092_)
);

OAI21X1 _13721_ (
    .A(_6073_),
    .B(_6068_),
    .C(_5963__bF$buf5),
    .Y(_6093_)
);

NAND2X1 _13722_ (
    .A(_6092_),
    .B(_6093_),
    .Y(_6094_)
);

NAND3X1 _13723_ (
    .A(_6086_),
    .B(_6091_),
    .C(_6094_),
    .Y(_6095_)
);

NAND3X1 _13724_ (
    .A(_5963__bF$buf4),
    .B(_6092_),
    .C(_6087_),
    .Y(_6096_)
);

NAND2X1 _13725_ (
    .A(_6090_),
    .B(_6093_),
    .Y(_6097_)
);

NAND3X1 _13726_ (
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .B(_6096_),
    .C(_6097_),
    .Y(_6098_)
);

NAND2X1 _13727_ (
    .A(_6095_),
    .B(_6098_),
    .Y(_6099_)
);

AOI21X1 _13728_ (
    .A(_6056_),
    .B(_6058_),
    .C(_6046_),
    .Y(_6100_)
);

NOR2X1 _13729_ (
    .A(_6100_),
    .B(_6079_),
    .Y(_6101_)
);

OAI21X1 _13730_ (
    .A(_6063_),
    .B(_6045_),
    .C(_6101_),
    .Y(_6102_)
);

NAND2X1 _13731_ (
    .A(_6078_),
    .B(_6102_),
    .Y(_6103_)
);

AOI21X1 _13732_ (
    .A(_6103_),
    .B(_6099_),
    .C(_5951_),
    .Y(_6104_)
);

OAI21X1 _13733_ (
    .A(_6099_),
    .B(_6103_),
    .C(_6104_),
    .Y(_6105_)
);

AOI22X1 _13734_ (
    .A(_6085_),
    .B(_5949__bF$buf2),
    .C(_6105_),
    .D(_6021_),
    .Y(_5842_)
);

INVX1 _13735_ (
    .A(\genblk1[7].u_ce.Ycalc [7]),
    .Y(_6106_)
);

AOI21X1 _13736_ (
    .A(_6094_),
    .B(_6091_),
    .C(_6086_),
    .Y(_6107_)
);

AND2X2 _13737_ (
    .A(_6059_),
    .B(_6062_),
    .Y(_6108_)
);

NAND3X1 _13738_ (
    .A(_6078_),
    .B(_6080_),
    .C(_6108_),
    .Y(_6109_)
);

AOI21X1 _13739_ (
    .A(_6100_),
    .B(_6078_),
    .C(_6079_),
    .Y(_6110_)
);

OAI21X1 _13740_ (
    .A(_6045_),
    .B(_6109_),
    .C(_6110_),
    .Y(_6111_)
);

AOI21X1 _13741_ (
    .A(_6111_),
    .B(_6095_),
    .C(_6107_),
    .Y(_6112_)
);

INVX1 _13742_ (
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .Y(_6113_)
);

NAND3X1 _13743_ (
    .A(_6076_),
    .B(_6092_),
    .C(_6075_),
    .Y(_6114_)
);

INVX1 _13744_ (
    .A(\genblk1[7].u_ce.Xin12b [11]),
    .Y(_6115_)
);

NOR2X1 _13745_ (
    .A(_5925__bF$buf1),
    .B(_6115_),
    .Y(_6116_)
);

INVX1 _13746_ (
    .A(_6116_),
    .Y(_6117_)
);

OAI21X1 _13747_ (
    .A(1'h1),
    .B(_6030_),
    .C(_6117_),
    .Y(_6118_)
);

NAND3X1 _13748_ (
    .A(_5963__bF$buf3),
    .B(_6118_),
    .C(_6114_),
    .Y(_6119_)
);

INVX1 _13749_ (
    .A(_6118_),
    .Y(_6120_)
);

OAI21X1 _13750_ (
    .A(_6090_),
    .B(_6087_),
    .C(_5963__bF$buf2),
    .Y(_6121_)
);

NAND2X1 _13751_ (
    .A(_6120_),
    .B(_6121_),
    .Y(_6122_)
);

NAND3X1 _13752_ (
    .A(_6113_),
    .B(_6119_),
    .C(_6122_),
    .Y(_6123_)
);

NAND3X1 _13753_ (
    .A(_5963__bF$buf1),
    .B(_6120_),
    .C(_6114_),
    .Y(_6124_)
);

NAND2X1 _13754_ (
    .A(_6118_),
    .B(_6121_),
    .Y(_6125_)
);

NAND3X1 _13755_ (
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .B(_6124_),
    .C(_6125_),
    .Y(_6126_)
);

NAND2X1 _13756_ (
    .A(_6123_),
    .B(_6126_),
    .Y(_6127_)
);

INVX1 _13757_ (
    .A(_6127_),
    .Y(_6128_)
);

NOR2X1 _13758_ (
    .A(_6128_),
    .B(_6112_),
    .Y(_6129_)
);

OAI21X1 _13759_ (
    .A(_6099_),
    .B(_6103_),
    .C(_6098_),
    .Y(_6130_)
);

OAI21X1 _13760_ (
    .A(_6127_),
    .B(_6130_),
    .C(_6018_),
    .Y(_6131_)
);

OAI21X1 _13761_ (
    .A(_5963__bF$buf0),
    .B(_6018_),
    .C(\genblk1[7].u_ce.Vld ),
    .Y(_6132_)
);

INVX1 _13762_ (
    .A(_6132_),
    .Y(_6133_)
);

OAI21X1 _13763_ (
    .A(_6131_),
    .B(_6129_),
    .C(_6133_),
    .Y(_6134_)
);

OAI21X1 _13764_ (
    .A(_6106_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6134_),
    .Y(_5843_)
);

INVX1 _13765_ (
    .A(\genblk1[7].u_ce.Ycalc [8]),
    .Y(_6135_)
);

OAI21X1 _13766_ (
    .A(_6098_),
    .B(_6127_),
    .C(_6126_),
    .Y(_6136_)
);

NOR2X1 _13767_ (
    .A(_6099_),
    .B(_6127_),
    .Y(_6137_)
);

AOI21X1 _13768_ (
    .A(_6137_),
    .B(_6111_),
    .C(_6136_),
    .Y(_6138_)
);

INVX1 _13769_ (
    .A(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6139_)
);

OR2X2 _13770_ (
    .A(_6114_),
    .B(_6118_),
    .Y(_6140_)
);

OAI21X1 _13771_ (
    .A(1'h1),
    .B(_6051_),
    .C(_6117_),
    .Y(_6141_)
);

NAND3X1 _13772_ (
    .A(_5963__bF$buf5),
    .B(_6141_),
    .C(_6140_),
    .Y(_6142_)
);

NOR2X1 _13773_ (
    .A(_6118_),
    .B(_6114_),
    .Y(_6143_)
);

INVX1 _13774_ (
    .A(_6141_),
    .Y(_6144_)
);

OAI21X1 _13775_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6143_),
    .C(_6144_),
    .Y(_6145_)
);

NAND3X1 _13776_ (
    .A(_6139_),
    .B(_6145_),
    .C(_6142_),
    .Y(_6146_)
);

NAND3X1 _13777_ (
    .A(_5963__bF$buf4),
    .B(_6144_),
    .C(_6140_),
    .Y(_6147_)
);

OAI21X1 _13778_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6143_),
    .C(_6141_),
    .Y(_6148_)
);

NAND3X1 _13779_ (
    .A(\genblk1[7].u_ce.Yin12b [8]),
    .B(_6148_),
    .C(_6147_),
    .Y(_6149_)
);

AND2X2 _13780_ (
    .A(_6146_),
    .B(_6149_),
    .Y(_6150_)
);

INVX1 _13781_ (
    .A(_6150_),
    .Y(_6151_)
);

AOI21X1 _13782_ (
    .A(_6138_),
    .B(_6151_),
    .C(_5951_),
    .Y(_6152_)
);

OAI21X1 _13783_ (
    .A(_6138_),
    .B(_6151_),
    .C(_6152_),
    .Y(_6153_)
);

AOI22X1 _13784_ (
    .A(_6135_),
    .B(_5949__bF$buf1),
    .C(_6153_),
    .D(_6133_),
    .Y(_5844_)
);

NAND2X1 _13785_ (
    .A(_6107_),
    .B(_6123_),
    .Y(_6154_)
);

AND2X2 _13786_ (
    .A(_6154_),
    .B(_6126_),
    .Y(_6155_)
);

AND2X2 _13787_ (
    .A(_6095_),
    .B(_6098_),
    .Y(_6156_)
);

NAND3X1 _13788_ (
    .A(_6123_),
    .B(_6126_),
    .C(_6156_),
    .Y(_6157_)
);

OAI21X1 _13789_ (
    .A(_6103_),
    .B(_6157_),
    .C(_6155_),
    .Y(_6158_)
);

INVX1 _13790_ (
    .A(_6149_),
    .Y(_6159_)
);

AOI21X1 _13791_ (
    .A(_6158_),
    .B(_6146_),
    .C(_6159_),
    .Y(_6160_)
);

INVX1 _13792_ (
    .A(\genblk1[7].u_ce.Yin12b [9]),
    .Y(_6161_)
);

NOR3X1 _13793_ (
    .A(_6118_),
    .B(_6141_),
    .C(_6114_),
    .Y(_6162_)
);

INVX1 _13794_ (
    .A(_6162_),
    .Y(_6163_)
);

OAI21X1 _13795_ (
    .A(1'h1),
    .B(_6071_),
    .C(_6117_),
    .Y(_6164_)
);

NAND3X1 _13796_ (
    .A(_5963__bF$buf3),
    .B(_6164_),
    .C(_6163_),
    .Y(_6165_)
);

INVX1 _13797_ (
    .A(_6164_),
    .Y(_6166_)
);

OAI21X1 _13798_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_6162_),
    .C(_6166_),
    .Y(_6167_)
);

NAND3X1 _13799_ (
    .A(_6161_),
    .B(_6167_),
    .C(_6165_),
    .Y(_6168_)
);

NAND3X1 _13800_ (
    .A(_5963__bF$buf2),
    .B(_6166_),
    .C(_6163_),
    .Y(_6169_)
);

OAI21X1 _13801_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6162_),
    .C(_6164_),
    .Y(_6170_)
);

NAND3X1 _13802_ (
    .A(\genblk1[7].u_ce.Yin12b [9]),
    .B(_6170_),
    .C(_6169_),
    .Y(_6171_)
);

AND2X2 _13803_ (
    .A(_6168_),
    .B(_6171_),
    .Y(_6172_)
);

AND2X2 _13804_ (
    .A(_6160_),
    .B(_6172_),
    .Y(_6173_)
);

OAI21X1 _13805_ (
    .A(_6172_),
    .B(_6160_),
    .C(_6018_),
    .Y(_6174_)
);

OAI21X1 _13806_ (
    .A(_6174_),
    .B(_6173_),
    .C(_6021_),
    .Y(_6175_)
);

OAI21X1 _13807_ (
    .A(_5901_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6175_),
    .Y(_5845_)
);

INVX1 _13808_ (
    .A(\genblk1[7].u_ce.Yin12b [10]),
    .Y(_6176_)
);

OAI21X1 _13809_ (
    .A(1'h1),
    .B(_6088_),
    .C(_6117_),
    .Y(_6177_)
);

INVX1 _13810_ (
    .A(_6177_),
    .Y(_6178_)
);

AOI21X1 _13811_ (
    .A(_6162_),
    .B(_6166_),
    .C(_6178_),
    .Y(_6179_)
);

NAND3X1 _13812_ (
    .A(_6166_),
    .B(_6178_),
    .C(_6162_),
    .Y(_6180_)
);

NAND2X1 _13813_ (
    .A(_5963__bF$buf1),
    .B(_6180_),
    .Y(_6181_)
);

NAND2X1 _13814_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6177_),
    .Y(_6182_)
);

OAI21X1 _13815_ (
    .A(_6179_),
    .B(_6181_),
    .C(_6182_),
    .Y(_6183_)
);

NAND2X1 _13816_ (
    .A(_6176_),
    .B(_6183_),
    .Y(_6184_)
);

INVX1 _13817_ (
    .A(_6179_),
    .Y(_6185_)
);

AND2X2 _13818_ (
    .A(_6180_),
    .B(_5963__bF$buf0),
    .Y(_6186_)
);

NAND2X1 _13819_ (
    .A(_6185_),
    .B(_6186_),
    .Y(_6187_)
);

NAND3X1 _13820_ (
    .A(\genblk1[7].u_ce.Yin12b [10]),
    .B(_6182_),
    .C(_6187_),
    .Y(_6188_)
);

NAND2X1 _13821_ (
    .A(_6184_),
    .B(_6188_),
    .Y(_6189_)
);

AOI21X1 _13822_ (
    .A(_6165_),
    .B(_6167_),
    .C(_6161_),
    .Y(_6190_)
);

AOI21X1 _13823_ (
    .A(_6159_),
    .B(_6168_),
    .C(_6190_),
    .Y(_6191_)
);

NAND3X1 _13824_ (
    .A(_6150_),
    .B(_6172_),
    .C(_6158_),
    .Y(_6192_)
);

AOI21X1 _13825_ (
    .A(_6192_),
    .B(_6191_),
    .C(_6189_),
    .Y(_6193_)
);

AND2X2 _13826_ (
    .A(_6188_),
    .B(_6184_),
    .Y(_6194_)
);

NAND3X1 _13827_ (
    .A(_6168_),
    .B(_6171_),
    .C(_6150_),
    .Y(_6195_)
);

OAI21X1 _13828_ (
    .A(_6195_),
    .B(_6138_),
    .C(_6191_),
    .Y(_6196_)
);

OAI21X1 _13829_ (
    .A(_6194_),
    .B(_6196_),
    .C(_6018_),
    .Y(_6197_)
);

OR2X2 _13830_ (
    .A(_6197_),
    .B(_6193_),
    .Y(_6198_)
);

AOI22X1 _13831_ (
    .A(_5893_),
    .B(_5949__bF$buf0),
    .C(_6198_),
    .D(_6021_),
    .Y(_5846_)
);

NAND2X1 _13832_ (
    .A(\genblk1[7].u_ce.Ycalc [11]),
    .B(_5949__bF$buf3),
    .Y(_6199_)
);

INVX1 _13833_ (
    .A(_6188_),
    .Y(_6200_)
);

NAND2X1 _13834_ (
    .A(\genblk1[7].u_ce.Yin12b [11]),
    .B(_6115_),
    .Y(_6201_)
);

INVX1 _13835_ (
    .A(\genblk1[7].u_ce.Yin12b [11]),
    .Y(_6202_)
);

NAND2X1 _13836_ (
    .A(\genblk1[7].u_ce.Xin12b [11]),
    .B(_6202_),
    .Y(_6203_)
);

NAND2X1 _13837_ (
    .A(_6201_),
    .B(_6203_),
    .Y(_6204_)
);

INVX1 _13838_ (
    .A(_6204_),
    .Y(_6205_)
);

NAND2X1 _13839_ (
    .A(_6205_),
    .B(_6181_),
    .Y(_6206_)
);

NAND2X1 _13840_ (
    .A(_6204_),
    .B(_6186_),
    .Y(_6207_)
);

NAND2X1 _13841_ (
    .A(_6206_),
    .B(_6207_),
    .Y(_6208_)
);

INVX1 _13842_ (
    .A(_6208_),
    .Y(_6209_)
);

NOR3X1 _13843_ (
    .A(_6200_),
    .B(_6209_),
    .C(_6193_),
    .Y(_6210_)
);

AOI21X1 _13844_ (
    .A(_6196_),
    .B(_6194_),
    .C(_6200_),
    .Y(_6211_)
);

OAI21X1 _13845_ (
    .A(_6208_),
    .B(_6211_),
    .C(_6018_),
    .Y(_6212_)
);

OAI21X1 _13846_ (
    .A(_6210_),
    .B(_6212_),
    .C(_6021_),
    .Y(_6213_)
);

NAND2X1 _13847_ (
    .A(_6199_),
    .B(_6213_),
    .Y(_5847_)
);

NAND2X1 _13848_ (
    .A(\genblk1[7].u_ce.Xcalc [0]),
    .B(_5949__bF$buf2),
    .Y(_6214_)
);

INVX1 _13849_ (
    .A(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6215_)
);

NAND2X1 _13850_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6216_)
);

OAI21X1 _13851_ (
    .A(1'h1),
    .B(_6215_),
    .C(_6216_),
    .Y(_6217_)
);

NAND2X1 _13852_ (
    .A(1'h1),
    .B(_6217_),
    .Y(_6218_)
);

NOR2X1 _13853_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_6219_)
);

NOR2X1 _13854_ (
    .A(1'h1),
    .B(_5955_),
    .Y(_6220_)
);

AOI22X1 _13855_ (
    .A(\genblk1[7].u_ce.Yin0 [0]),
    .B(_6219_),
    .C(_6220_),
    .D(\genblk1[7].u_ce.Yin0 [1]),
    .Y(_6221_)
);

NAND3X1 _13856_ (
    .A(_5925__bF$buf0),
    .B(_6218_),
    .C(_6221_),
    .Y(_6222_)
);

NAND2X1 _13857_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [7]),
    .Y(_6223_)
);

OAI21X1 _13858_ (
    .A(1'h1),
    .B(_6086_),
    .C(_6223_),
    .Y(_6224_)
);

NAND2X1 _13859_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [5]),
    .Y(_6225_)
);

OAI21X1 _13860_ (
    .A(1'h1),
    .B(_6046_),
    .C(_6225_),
    .Y(_6226_)
);

MUX2X1 _13861_ (
    .A(_6226_),
    .B(_6224_),
    .S(_5926__bF$buf1),
    .Y(_6227_)
);

NAND2X1 _13862_ (
    .A(1'h1),
    .B(_6227_),
    .Y(_6228_)
);

AND2X2 _13863_ (
    .A(_6222_),
    .B(_6228_),
    .Y(_6229_)
);

NOR2X1 _13864_ (
    .A(\genblk1[7].u_ce.Xin0 [0]),
    .B(_6229_),
    .Y(_6230_)
);

NAND2X1 _13865_ (
    .A(_5926__bF$buf0),
    .B(_6226_),
    .Y(_6231_)
);

NAND2X1 _13866_ (
    .A(1'h1),
    .B(_6224_),
    .Y(_6232_)
);

NAND2X1 _13867_ (
    .A(_6231_),
    .B(_6232_),
    .Y(_6233_)
);

OAI21X1 _13868_ (
    .A(_5925__bF$buf3),
    .B(_6233_),
    .C(_6222_),
    .Y(_6234_)
);

OAI21X1 _13869_ (
    .A(_5937_),
    .B(_6234_),
    .C(_5947_),
    .Y(_6235_)
);

OAI21X1 _13870_ (
    .A(_6235_),
    .B(_6230_),
    .C(_6214_),
    .Y(_5848_)
);

NAND2X1 _13871_ (
    .A(\genblk1[7].u_ce.Xcalc [1]),
    .B(_5949__bF$buf1),
    .Y(_6236_)
);

NOR2X1 _13872_ (
    .A(_5937_),
    .B(_6234_),
    .Y(_6237_)
);

NAND2X1 _13873_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [4]),
    .Y(_6238_)
);

OAI21X1 _13874_ (
    .A(1'h1),
    .B(_6024_),
    .C(_6238_),
    .Y(_6239_)
);

NAND2X1 _13875_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6240_)
);

OAI21X1 _13876_ (
    .A(1'h1),
    .B(_5962_),
    .C(_6240_),
    .Y(_6241_)
);

MUX2X1 _13877_ (
    .A(_6241_),
    .B(_6239_),
    .S(_5926__bF$buf4),
    .Y(_6242_)
);

NAND2X1 _13878_ (
    .A(_5925__bF$buf2),
    .B(_6242_),
    .Y(_6243_)
);

NAND2X1 _13879_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6244_)
);

OAI21X1 _13880_ (
    .A(1'h1),
    .B(_6113_),
    .C(_6244_),
    .Y(_6245_)
);

INVX1 _13881_ (
    .A(_6245_),
    .Y(_6246_)
);

NAND2X1 _13882_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [6]),
    .Y(_6247_)
);

OAI21X1 _13883_ (
    .A(1'h1),
    .B(_6067_),
    .C(_6247_),
    .Y(_6248_)
);

NAND2X1 _13884_ (
    .A(_5926__bF$buf3),
    .B(_6248_),
    .Y(_6249_)
);

OAI21X1 _13885_ (
    .A(_5926__bF$buf2),
    .B(_6246_),
    .C(_6249_),
    .Y(_6250_)
);

OAI21X1 _13886_ (
    .A(_5925__bF$buf1),
    .B(_6250_),
    .C(_6243_),
    .Y(_6251_)
);

NAND3X1 _13887_ (
    .A(_5963__bF$buf5),
    .B(_6251_),
    .C(_6229_),
    .Y(_6252_)
);

MUX2X1 _13888_ (
    .A(_6248_),
    .B(_6245_),
    .S(_5926__bF$buf1),
    .Y(_6253_)
);

MUX2X1 _13889_ (
    .A(_6253_),
    .B(_6242_),
    .S(1'h1),
    .Y(_6254_)
);

OAI21X1 _13890_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6234_),
    .C(_6254_),
    .Y(_6255_)
);

AOI21X1 _13891_ (
    .A(_6252_),
    .B(_6255_),
    .C(_5974_),
    .Y(_6256_)
);

INVX1 _13892_ (
    .A(_6256_),
    .Y(_6257_)
);

NAND3X1 _13893_ (
    .A(_5974_),
    .B(_6255_),
    .C(_6252_),
    .Y(_6258_)
);

AND2X2 _13894_ (
    .A(_6257_),
    .B(_6258_),
    .Y(_6259_)
);

NAND2X1 _13895_ (
    .A(_6237_),
    .B(_6259_),
    .Y(_6260_)
);

OR2X2 _13896_ (
    .A(_6259_),
    .B(_6237_),
    .Y(_6261_)
);

AOI21X1 _13897_ (
    .A(_6261_),
    .B(_6260_),
    .C(_5951_),
    .Y(_6262_)
);

OAI21X1 _13898_ (
    .A(_5949__bF$buf0),
    .B(_6262_),
    .C(_6236_),
    .Y(_5849_)
);

NAND2X1 _13899_ (
    .A(\genblk1[7].u_ce.Xcalc [2]),
    .B(_5949__bF$buf3),
    .Y(_6263_)
);

AOI21X1 _13900_ (
    .A(_6237_),
    .B(_6258_),
    .C(_6256_),
    .Y(_6264_)
);

NAND2X1 _13901_ (
    .A(_6234_),
    .B(_6251_),
    .Y(_6265_)
);

NAND2X1 _13902_ (
    .A(1'h1),
    .B(_6161_),
    .Y(_6266_)
);

OAI21X1 _13903_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [8]),
    .C(_6266_),
    .Y(_6267_)
);

NAND2X1 _13904_ (
    .A(_5926__bF$buf0),
    .B(_6224_),
    .Y(_6268_)
);

OAI21X1 _13905_ (
    .A(_5926__bF$buf4),
    .B(_6267_),
    .C(_6268_),
    .Y(_6269_)
);

NAND2X1 _13906_ (
    .A(_6032_),
    .B(_6217_),
    .Y(_6270_)
);

NAND2X1 _13907_ (
    .A(_6226_),
    .B(_6031_),
    .Y(_6271_)
);

NAND2X1 _13908_ (
    .A(_6270_),
    .B(_6271_),
    .Y(_6272_)
);

AOI21X1 _13909_ (
    .A(_6269_),
    .B(1'h1),
    .C(_6272_),
    .Y(_6273_)
);

INVX1 _13910_ (
    .A(_6273_),
    .Y(_6274_)
);

NAND3X1 _13911_ (
    .A(_5963__bF$buf4),
    .B(_6274_),
    .C(_6265_),
    .Y(_6275_)
);

AOI21X1 _13912_ (
    .A(_6222_),
    .B(_6228_),
    .C(_6254_),
    .Y(_6276_)
);

OAI21X1 _13913_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf2 ),
    .B(_6276_),
    .C(_6273_),
    .Y(_6277_)
);

NAND3X1 _13914_ (
    .A(\genblk1[7].u_ce.Xin1 [0]),
    .B(_6277_),
    .C(_6275_),
    .Y(_6278_)
);

INVX1 _13915_ (
    .A(_6278_),
    .Y(_6279_)
);

AOI21X1 _13916_ (
    .A(_6275_),
    .B(_6277_),
    .C(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_6280_)
);

NOR2X1 _13917_ (
    .A(_6280_),
    .B(_6279_),
    .Y(_6281_)
);

AND2X2 _13918_ (
    .A(_6281_),
    .B(_6264_),
    .Y(_6282_)
);

NOR2X1 _13919_ (
    .A(_6264_),
    .B(_6281_),
    .Y(_6283_)
);

OAI21X1 _13920_ (
    .A(_6283_),
    .B(_6282_),
    .C(_6018_),
    .Y(_6284_)
);

OAI21X1 _13921_ (
    .A(_5949__bF$buf2),
    .B(_6284_),
    .C(_6263_),
    .Y(_5850_)
);

OAI21X1 _13922_ (
    .A(_6280_),
    .B(_6264_),
    .C(_6278_),
    .Y(_6285_)
);

INVX1 _13923_ (
    .A(_6285_),
    .Y(_6286_)
);

NAND2X1 _13924_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [10]),
    .Y(_6287_)
);

OAI21X1 _13925_ (
    .A(1'h1),
    .B(_6161_),
    .C(_6287_),
    .Y(_6288_)
);

MUX2X1 _13926_ (
    .A(_6288_),
    .B(_6245_),
    .S(1'h1),
    .Y(_6289_)
);

NOR2X1 _13927_ (
    .A(_5925__bF$buf0),
    .B(_6289_),
    .Y(_6290_)
);

NAND2X1 _13928_ (
    .A(_6032_),
    .B(_6239_),
    .Y(_6291_)
);

NAND2X1 _13929_ (
    .A(_6248_),
    .B(_6031_),
    .Y(_6292_)
);

NAND2X1 _13930_ (
    .A(_6291_),
    .B(_6292_),
    .Y(_6293_)
);

OR2X2 _13931_ (
    .A(_6290_),
    .B(_6293_),
    .Y(_6294_)
);

OAI21X1 _13932_ (
    .A(_6274_),
    .B(_6265_),
    .C(_5963__bF$buf3),
    .Y(_6295_)
);

OR2X2 _13933_ (
    .A(_6295_),
    .B(_6294_),
    .Y(_6296_)
);

OAI21X1 _13934_ (
    .A(_6290_),
    .B(_6293_),
    .C(_6295_),
    .Y(_6297_)
);

AOI21X1 _13935_ (
    .A(_6296_),
    .B(_6297_),
    .C(_5971_),
    .Y(_6298_)
);

INVX1 _13936_ (
    .A(_6298_),
    .Y(_6299_)
);

NAND3X1 _13937_ (
    .A(_5971_),
    .B(_6297_),
    .C(_6296_),
    .Y(_6300_)
);

NAND2X1 _13938_ (
    .A(_6300_),
    .B(_6299_),
    .Y(_6301_)
);

OR2X2 _13939_ (
    .A(_6301_),
    .B(_6286_),
    .Y(_6302_)
);

NAND2X1 _13940_ (
    .A(_6286_),
    .B(_6301_),
    .Y(_6303_)
);

NAND2X1 _13941_ (
    .A(_6303_),
    .B(_6302_),
    .Y(_6304_)
);

AOI22X1 _13942_ (
    .A(_5917_),
    .B(_5949__bF$buf1),
    .C(_6304_),
    .D(_5947_),
    .Y(_5851_)
);

AOI21X1 _13943_ (
    .A(_6285_),
    .B(_6300_),
    .C(_6298_),
    .Y(_6305_)
);

NAND2X1 _13944_ (
    .A(1'h1),
    .B(\genblk1[7].u_ce.Yin12b [11]),
    .Y(_6306_)
);

OAI21X1 _13945_ (
    .A(1'h1),
    .B(_6176_),
    .C(_6306_),
    .Y(_6307_)
);

NAND2X1 _13946_ (
    .A(1'h1),
    .B(_6307_),
    .Y(_6308_)
);

OAI21X1 _13947_ (
    .A(1'h1),
    .B(_6267_),
    .C(_6308_),
    .Y(_6309_)
);

NAND2X1 _13948_ (
    .A(1'h1),
    .B(_6309_),
    .Y(_6310_)
);

OAI21X1 _13949_ (
    .A(1'h1),
    .B(_6227_),
    .C(_6310_),
    .Y(_6311_)
);

INVX1 _13950_ (
    .A(_6311_),
    .Y(_6312_)
);

NAND3X1 _13951_ (
    .A(_6273_),
    .B(_6234_),
    .C(_6251_),
    .Y(_6313_)
);

OAI21X1 _13952_ (
    .A(_6294_),
    .B(_6313_),
    .C(_5963__bF$buf2),
    .Y(_6314_)
);

OR2X2 _13953_ (
    .A(_6314_),
    .B(_6312_),
    .Y(_6315_)
);

NOR2X1 _13954_ (
    .A(_6294_),
    .B(_6313_),
    .Y(_6316_)
);

OAI21X1 _13955_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf1 ),
    .B(_6316_),
    .C(_6312_),
    .Y(_6317_)
);

NAND3X1 _13956_ (
    .A(\genblk1[7].u_ce.Xin12b [4]),
    .B(_6317_),
    .C(_6315_),
    .Y(_6318_)
);

OR2X2 _13957_ (
    .A(_6314_),
    .B(_6311_),
    .Y(_6319_)
);

OAI21X1 _13958_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf0 ),
    .B(_6316_),
    .C(_6311_),
    .Y(_6320_)
);

NAND3X1 _13959_ (
    .A(_5930_),
    .B(_6320_),
    .C(_6319_),
    .Y(_6321_)
);

NAND2X1 _13960_ (
    .A(_6318_),
    .B(_6321_),
    .Y(_6322_)
);

OR2X2 _13961_ (
    .A(_6305_),
    .B(_6322_),
    .Y(_6323_)
);

NAND2X1 _13962_ (
    .A(_6322_),
    .B(_6305_),
    .Y(_6324_)
);

NAND2X1 _13963_ (
    .A(_6324_),
    .B(_6323_),
    .Y(_6325_)
);

AOI22X1 _13964_ (
    .A(_5912_),
    .B(_5949__bF$buf0),
    .C(_6325_),
    .D(_5947_),
    .Y(_5852_)
);

INVX1 _13965_ (
    .A(\genblk1[7].u_ce.Xcalc [5]),
    .Y(_6326_)
);

OAI21X1 _13966_ (
    .A(_6322_),
    .B(_6305_),
    .C(_6318_),
    .Y(_6327_)
);

NAND2X1 _13967_ (
    .A(_6312_),
    .B(_6316_),
    .Y(_6328_)
);

NOR2X1 _13968_ (
    .A(_5926__bF$buf3),
    .B(_6202_),
    .Y(_6329_)
);

AOI21X1 _13969_ (
    .A(_5926__bF$buf2),
    .B(_6288_),
    .C(_6329_),
    .Y(_6330_)
);

NAND2X1 _13970_ (
    .A(_5925__bF$buf3),
    .B(_6250_),
    .Y(_6331_)
);

OAI21X1 _13971_ (
    .A(_5925__bF$buf2),
    .B(_6330_),
    .C(_6331_),
    .Y(_6332_)
);

INVX1 _13972_ (
    .A(_6332_),
    .Y(_6333_)
);

NAND3X1 _13973_ (
    .A(_5963__bF$buf1),
    .B(_6333_),
    .C(_6328_),
    .Y(_6334_)
);

NOR2X1 _13974_ (
    .A(_6293_),
    .B(_6290_),
    .Y(_6335_)
);

NAND3X1 _13975_ (
    .A(_6273_),
    .B(_6335_),
    .C(_6276_),
    .Y(_6336_)
);

OAI21X1 _13976_ (
    .A(_6311_),
    .B(_6336_),
    .C(_5963__bF$buf0),
    .Y(_6337_)
);

NAND2X1 _13977_ (
    .A(_6332_),
    .B(_6337_),
    .Y(_6338_)
);

AOI21X1 _13978_ (
    .A(_6334_),
    .B(_6338_),
    .C(_5967_),
    .Y(_6339_)
);

INVX1 _13979_ (
    .A(_6339_),
    .Y(_6340_)
);

NAND3X1 _13980_ (
    .A(_5967_),
    .B(_6338_),
    .C(_6334_),
    .Y(_6341_)
);

NAND2X1 _13981_ (
    .A(_6341_),
    .B(_6340_),
    .Y(_6342_)
);

NOR2X1 _13982_ (
    .A(_6342_),
    .B(_6327_),
    .Y(_6343_)
);

AND2X2 _13983_ (
    .A(_6327_),
    .B(_6342_),
    .Y(_6344_)
);

OAI21X1 _13984_ (
    .A(_6343_),
    .B(_6344_),
    .C(_5947_),
    .Y(_6345_)
);

OAI21X1 _13985_ (
    .A(_6326_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6345_),
    .Y(_5853_)
);

INVX1 _13986_ (
    .A(\genblk1[7].u_ce.Xcalc [6]),
    .Y(_6346_)
);

NAND3X1 _13987_ (
    .A(_6312_),
    .B(_6333_),
    .C(_6316_),
    .Y(_6347_)
);

AOI21X1 _13988_ (
    .A(_5926__bF$buf1),
    .B(_6307_),
    .C(_6329_),
    .Y(_6348_)
);

NAND2X1 _13989_ (
    .A(1'h1),
    .B(_6348_),
    .Y(_6349_)
);

OAI21X1 _13990_ (
    .A(1'h1),
    .B(_6269_),
    .C(_6349_),
    .Y(_6350_)
);

NAND3X1 _13991_ (
    .A(_5963__bF$buf5),
    .B(_6350_),
    .C(_6347_),
    .Y(_6351_)
);

NOR3X1 _13992_ (
    .A(_6311_),
    .B(_6332_),
    .C(_6336_),
    .Y(_6352_)
);

INVX1 _13993_ (
    .A(_6350_),
    .Y(_6353_)
);

OAI21X1 _13994_ (
    .A(\genblk1[7].u_ce.Ain12b_11_bF$buf3 ),
    .B(_6352_),
    .C(_6353_),
    .Y(_6354_)
);

NAND2X1 _13995_ (
    .A(_6351_),
    .B(_6354_),
    .Y(_6355_)
);

NAND2X1 _13996_ (
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(_6355_),
    .Y(_6356_)
);

NAND3X1 _13997_ (
    .A(_5927_),
    .B(_6351_),
    .C(_6354_),
    .Y(_6357_)
);

NAND2X1 _13998_ (
    .A(_6357_),
    .B(_6356_),
    .Y(_6358_)
);

AOI21X1 _13999_ (
    .A(_6319_),
    .B(_6320_),
    .C(_5930_),
    .Y(_6359_)
);

NOR2X1 _14000_ (
    .A(_6359_),
    .B(_6339_),
    .Y(_6360_)
);

OAI21X1 _14001_ (
    .A(_6322_),
    .B(_6305_),
    .C(_6360_),
    .Y(_6361_)
);

NAND2X1 _14002_ (
    .A(_6341_),
    .B(_6361_),
    .Y(_6362_)
);

NOR2X1 _14003_ (
    .A(_6358_),
    .B(_6362_),
    .Y(_6363_)
);

AND2X2 _14004_ (
    .A(_6356_),
    .B(_6357_),
    .Y(_6364_)
);

AND2X2 _14005_ (
    .A(_6318_),
    .B(_6321_),
    .Y(_6365_)
);

NAND3X1 _14006_ (
    .A(_6341_),
    .B(_6365_),
    .C(_6340_),
    .Y(_6366_)
);

AOI21X1 _14007_ (
    .A(_6359_),
    .B(_6341_),
    .C(_6339_),
    .Y(_6367_)
);

OAI21X1 _14008_ (
    .A(_6305_),
    .B(_6366_),
    .C(_6367_),
    .Y(_6368_)
);

NOR2X1 _14009_ (
    .A(_6364_),
    .B(_6368_),
    .Y(_6369_)
);

OAI21X1 _14010_ (
    .A(_6369_),
    .B(_6363_),
    .C(_6018_),
    .Y(_6370_)
);

NAND2X1 _14011_ (
    .A(\genblk1[7].u_ce.Vld ),
    .B(_6370_),
    .Y(_6371_)
);

OAI21X1 _14012_ (
    .A(_6346_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6371_),
    .Y(_5854_)
);

INVX1 _14013_ (
    .A(\genblk1[7].u_ce.Xcalc [7]),
    .Y(_6372_)
);

INVX1 _14014_ (
    .A(_6356_),
    .Y(_6373_)
);

NAND2X1 _14015_ (
    .A(_6350_),
    .B(_6352_),
    .Y(_6374_)
);

NOR2X1 _14016_ (
    .A(_5925__bF$buf1),
    .B(_6202_),
    .Y(_6375_)
);

INVX1 _14017_ (
    .A(_6375_),
    .Y(_6376_)
);

OAI21X1 _14018_ (
    .A(1'h1),
    .B(_6289_),
    .C(_6376_),
    .Y(_6377_)
);

NAND3X1 _14019_ (
    .A(_5963__bF$buf4),
    .B(_6377_),
    .C(_6374_),
    .Y(_6378_)
);

INVX1 _14020_ (
    .A(_6377_),
    .Y(_6379_)
);

OAI21X1 _14021_ (
    .A(_6353_),
    .B(_6347_),
    .C(_5963__bF$buf3),
    .Y(_6380_)
);

NAND2X1 _14022_ (
    .A(_6379_),
    .B(_6380_),
    .Y(_6381_)
);

NAND3X1 _14023_ (
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(_6378_),
    .C(_6381_),
    .Y(_6382_)
);

NAND3X1 _14024_ (
    .A(_5963__bF$buf2),
    .B(_6379_),
    .C(_6374_),
    .Y(_6383_)
);

NAND2X1 _14025_ (
    .A(_6377_),
    .B(_6380_),
    .Y(_6384_)
);

NAND3X1 _14026_ (
    .A(_5964_),
    .B(_6383_),
    .C(_6384_),
    .Y(_6385_)
);

NAND2X1 _14027_ (
    .A(_6382_),
    .B(_6385_),
    .Y(_6386_)
);

OAI21X1 _14028_ (
    .A(_6373_),
    .B(_6363_),
    .C(_6386_),
    .Y(_6387_)
);

NOR2X1 _14029_ (
    .A(_6373_),
    .B(_6363_),
    .Y(_6388_)
);

INVX1 _14030_ (
    .A(_6386_),
    .Y(_6389_)
);

AOI21X1 _14031_ (
    .A(_6388_),
    .B(_6389_),
    .C(_5946_),
    .Y(_6390_)
);

AOI22X1 _14032_ (
    .A(_6372_),
    .B(_5949__bF$buf3),
    .C(_6390_),
    .D(_6387_),
    .Y(_5855_)
);

OAI21X1 _14033_ (
    .A(_6356_),
    .B(_6386_),
    .C(_6382_),
    .Y(_6391_)
);

NOR2X1 _14034_ (
    .A(_6358_),
    .B(_6386_),
    .Y(_6392_)
);

AOI21X1 _14035_ (
    .A(_6392_),
    .B(_6368_),
    .C(_6391_),
    .Y(_6393_)
);

INVX1 _14036_ (
    .A(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6394_)
);

NAND3X1 _14037_ (
    .A(_6350_),
    .B(_6379_),
    .C(_6352_),
    .Y(_6395_)
);

INVX1 _14038_ (
    .A(_6309_),
    .Y(_6396_)
);

OAI21X1 _14039_ (
    .A(1'h1),
    .B(_6396_),
    .C(_6376_),
    .Y(_6397_)
);

INVX1 _14040_ (
    .A(_6397_),
    .Y(_6398_)
);

NAND3X1 _14041_ (
    .A(_5963__bF$buf1),
    .B(_6398_),
    .C(_6395_),
    .Y(_6399_)
);

OAI21X1 _14042_ (
    .A(_6377_),
    .B(_6374_),
    .C(_5963__bF$buf0),
    .Y(_6400_)
);

NAND2X1 _14043_ (
    .A(_6397_),
    .B(_6400_),
    .Y(_6401_)
);

AOI21X1 _14044_ (
    .A(_6401_),
    .B(_6399_),
    .C(_6394_),
    .Y(_6402_)
);

NAND3X1 _14045_ (
    .A(_5963__bF$buf5),
    .B(_6397_),
    .C(_6395_),
    .Y(_6403_)
);

NAND2X1 _14046_ (
    .A(_6398_),
    .B(_6400_),
    .Y(_6404_)
);

AOI21X1 _14047_ (
    .A(_6404_),
    .B(_6403_),
    .C(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6405_)
);

OAI21X1 _14048_ (
    .A(_6402_),
    .B(_6405_),
    .C(_6393_),
    .Y(_6406_)
);

INVX1 _14049_ (
    .A(_6406_),
    .Y(_6407_)
);

OR2X2 _14050_ (
    .A(_6402_),
    .B(_6405_),
    .Y(_6408_)
);

OAI21X1 _14051_ (
    .A(_6408_),
    .B(_6393_),
    .C(_5947_),
    .Y(_6409_)
);

OAI22X1 _14052_ (
    .A(_5909_),
    .B(\genblk1[7].u_ce.Vld ),
    .C(_6409_),
    .D(_6407_),
    .Y(_5856_)
);

NAND2X1 _14053_ (
    .A(\genblk1[7].u_ce.Xcalc [9]),
    .B(_5949__bF$buf2),
    .Y(_6410_)
);

NOR2X1 _14054_ (
    .A(_6408_),
    .B(_6393_),
    .Y(_6411_)
);

NOR2X1 _14055_ (
    .A(_6402_),
    .B(_6411_),
    .Y(_6412_)
);

OAI21X1 _14056_ (
    .A(1'h1),
    .B(_6330_),
    .C(_6376_),
    .Y(_6413_)
);

INVX1 _14057_ (
    .A(_6413_),
    .Y(_6414_)
);

OAI21X1 _14058_ (
    .A(_6397_),
    .B(_6395_),
    .C(_5963__bF$buf4),
    .Y(_6415_)
);

NAND2X1 _14059_ (
    .A(_6414_),
    .B(_6415_),
    .Y(_6416_)
);

OR2X2 _14060_ (
    .A(_6415_),
    .B(_6414_),
    .Y(_6417_)
);

NAND3X1 _14061_ (
    .A(\genblk1[7].u_ce.Xin12b [9]),
    .B(_6416_),
    .C(_6417_),
    .Y(_6418_)
);

NAND2X1 _14062_ (
    .A(_6416_),
    .B(_6417_),
    .Y(_6419_)
);

NAND2X1 _14063_ (
    .A(_6026_),
    .B(_6419_),
    .Y(_6420_)
);

NAND2X1 _14064_ (
    .A(_6418_),
    .B(_6420_),
    .Y(_6421_)
);

AND2X2 _14065_ (
    .A(_6412_),
    .B(_6421_),
    .Y(_6422_)
);

OAI21X1 _14066_ (
    .A(_6421_),
    .B(_6412_),
    .C(_5947_),
    .Y(_6423_)
);

OAI21X1 _14067_ (
    .A(_6423_),
    .B(_6422_),
    .C(_6410_),
    .Y(_5857_)
);

INVX1 _14068_ (
    .A(\genblk1[7].u_ce.Xcalc [10]),
    .Y(_6424_)
);

INVX1 _14069_ (
    .A(_6418_),
    .Y(_6425_)
);

AOI21X1 _14070_ (
    .A(_6402_),
    .B(_6420_),
    .C(_6425_),
    .Y(_6426_)
);

NOR2X1 _14071_ (
    .A(_6402_),
    .B(_6405_),
    .Y(_6427_)
);

NAND3X1 _14072_ (
    .A(_6418_),
    .B(_6420_),
    .C(_6427_),
    .Y(_6428_)
);

OAI21X1 _14073_ (
    .A(_6393_),
    .B(_6428_),
    .C(_6426_),
    .Y(_6429_)
);

OAI21X1 _14074_ (
    .A(1'h1),
    .B(_6348_),
    .C(_6376_),
    .Y(_6430_)
);

INVX1 _14075_ (
    .A(_6430_),
    .Y(_6431_)
);

OR2X2 _14076_ (
    .A(_6395_),
    .B(_6397_),
    .Y(_6432_)
);

OAI21X1 _14077_ (
    .A(_6413_),
    .B(_6432_),
    .C(_5963__bF$buf3),
    .Y(_6433_)
);

NAND2X1 _14078_ (
    .A(_6431_),
    .B(_6433_),
    .Y(_6434_)
);

OR2X2 _14079_ (
    .A(_6433_),
    .B(_6431_),
    .Y(_6435_)
);

NAND3X1 _14080_ (
    .A(\genblk1[7].u_ce.Xin12b [10]),
    .B(_6434_),
    .C(_6435_),
    .Y(_6436_)
);

AND2X2 _14081_ (
    .A(_6433_),
    .B(_6431_),
    .Y(_6437_)
);

NOR2X1 _14082_ (
    .A(_6431_),
    .B(_6433_),
    .Y(_6438_)
);

OAI21X1 _14083_ (
    .A(_6438_),
    .B(_6437_),
    .C(_6047_),
    .Y(_6439_)
);

NAND2X1 _14084_ (
    .A(_6439_),
    .B(_6436_),
    .Y(_6440_)
);

AND2X2 _14085_ (
    .A(_6429_),
    .B(_6440_),
    .Y(_6441_)
);

NOR2X1 _14086_ (
    .A(_6440_),
    .B(_6429_),
    .Y(_6442_)
);

NOR2X1 _14087_ (
    .A(_6441_),
    .B(_6442_),
    .Y(_6443_)
);

AOI22X1 _14088_ (
    .A(_6424_),
    .B(_5949__bF$buf1),
    .C(_6443_),
    .D(_5947_),
    .Y(_5858_)
);

NAND2X1 _14089_ (
    .A(\genblk1[7].u_ce.Xcalc [11]),
    .B(_5949__bF$buf0),
    .Y(_6444_)
);

INVX1 _14090_ (
    .A(_6436_),
    .Y(_6445_)
);

AOI21X1 _14091_ (
    .A(_6429_),
    .B(_6439_),
    .C(_6445_),
    .Y(_6446_)
);

NAND2X1 _14092_ (
    .A(_5963__bF$buf2),
    .B(_6434_),
    .Y(_6447_)
);

NOR2X1 _14093_ (
    .A(_6204_),
    .B(_6447_),
    .Y(_6448_)
);

AOI21X1 _14094_ (
    .A(_6434_),
    .B(_5963__bF$buf1),
    .C(_6205_),
    .Y(_6449_)
);

NOR2X1 _14095_ (
    .A(_6449_),
    .B(_6448_),
    .Y(_6450_)
);

AND2X2 _14096_ (
    .A(_6446_),
    .B(_6450_),
    .Y(_6451_)
);

OAI21X1 _14097_ (
    .A(_6450_),
    .B(_6446_),
    .C(_5947_),
    .Y(_6452_)
);

OAI21X1 _14098_ (
    .A(_6452_),
    .B(_6451_),
    .C(_6444_),
    .Y(_5859_)
);

NAND2X1 _14099_ (
    .A(\genblk1[7].u_ce.LoadCtl [5]),
    .B(_5888_),
    .Y(_6453_)
);

NAND2X1 _14100_ (
    .A(_5889_),
    .B(_5892_),
    .Y(_6454_)
);

NOR2X1 _14101_ (
    .A(_6453_),
    .B(_6454_),
    .Y(_6455_)
);

NAND2X1 _14102_ (
    .A(\genblk1[6].u_ce.X_ [0]),
    .B(_6455_),
    .Y(_6456_)
);

OAI21X1 _14103_ (
    .A(_6047_),
    .B(_6455_),
    .C(_6456_),
    .Y(_5860_)
);

NAND2X1 _14104_ (
    .A(\genblk1[6].u_ce.X_ [1]),
    .B(_6455_),
    .Y(_6457_)
);

OAI21X1 _14105_ (
    .A(_6115_),
    .B(_6455_),
    .C(_6457_),
    .Y(_5861_)
);

INVX1 _14106_ (
    .A(\genblk1[6].u_ce.X_ [0]),
    .Y(_6458_)
);

OR2X2 _14107_ (
    .A(_6454_),
    .B(_5888_),
    .Y(_6459_)
);

OAI21X1 _14108_ (
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Xin12b [8]),
    .Y(_6460_)
);

OAI21X1 _14109_ (
    .A(_6458_),
    .B(_6459_),
    .C(_6460_),
    .Y(_5862_)
);

INVX1 _14110_ (
    .A(\genblk1[6].u_ce.X_ [1]),
    .Y(_6461_)
);

OAI21X1 _14111_ (
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Xin12b [9]),
    .Y(_6462_)
);

OAI21X1 _14112_ (
    .A(_6461_),
    .B(_6459_),
    .C(_6462_),
    .Y(_5863_)
);

NAND2X1 _14113_ (
    .A(_5892_),
    .B(_5891_),
    .Y(_6463_)
);

NAND2X1 _14114_ (
    .A(\genblk1[7].u_ce.Xin12b [6]),
    .B(_6463_),
    .Y(_6464_)
);

OAI21X1 _14115_ (
    .A(_6458_),
    .B(_6463_),
    .C(_6464_),
    .Y(_5864_)
);

NAND2X1 _14116_ (
    .A(\genblk1[7].u_ce.Xin12b [7]),
    .B(_6463_),
    .Y(_6465_)
);

OAI21X1 _14117_ (
    .A(_6461_),
    .B(_6463_),
    .C(_6465_),
    .Y(_5865_)
);

AND2X2 _14118_ (
    .A(_5892_),
    .B(\genblk1[7].u_ce.LoadCtl [2]),
    .Y(_6466_)
);

NAND2X1 _14119_ (
    .A(\genblk1[6].u_ce.X_ [0]),
    .B(_6466_),
    .Y(_6467_)
);

OAI21X1 _14120_ (
    .A(_5930_),
    .B(_6466_),
    .C(_6467_),
    .Y(_5866_)
);

NAND2X1 _14121_ (
    .A(\genblk1[6].u_ce.X_ [1]),
    .B(_6466_),
    .Y(_6468_)
);

OAI21X1 _14122_ (
    .A(_5967_),
    .B(_6466_),
    .C(_6468_),
    .Y(_5867_)
);

OAI21X1 _14123_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Xin1 [0]),
    .Y(_6469_)
);

OAI21X1 _14124_ (
    .A(_6458_),
    .B(_5887_),
    .C(_6469_),
    .Y(_5868_)
);

OAI21X1 _14125_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Xin1 [1]),
    .Y(_6470_)
);

OAI21X1 _14126_ (
    .A(_6461_),
    .B(_5887_),
    .C(_6470_),
    .Y(_5869_)
);

NAND2X1 _14127_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.X_ [0]),
    .Y(_6471_)
);

OAI21X1 _14128_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5937_),
    .C(_6471_),
    .Y(_5870_)
);

NAND2X1 _14129_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.X_ [1]),
    .Y(_6472_)
);

OAI21X1 _14130_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5974_),
    .C(_6472_),
    .Y(_5871_)
);

NAND2X1 _14131_ (
    .A(\genblk1[6].u_ce.Y_ [0]),
    .B(_6455_),
    .Y(_6473_)
);

OAI21X1 _14132_ (
    .A(_6176_),
    .B(_6455_),
    .C(_6473_),
    .Y(_5872_)
);

NAND2X1 _14133_ (
    .A(\genblk1[6].u_ce.Y_ [1]),
    .B(_6455_),
    .Y(_6474_)
);

OAI21X1 _14134_ (
    .A(_6202_),
    .B(_6455_),
    .C(_6474_),
    .Y(_5873_)
);

INVX1 _14135_ (
    .A(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6475_)
);

OAI21X1 _14136_ (
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Yin12b [8]),
    .Y(_6476_)
);

OAI21X1 _14137_ (
    .A(_6475_),
    .B(_6459_),
    .C(_6476_),
    .Y(_5874_)
);

INVX1 _14138_ (
    .A(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6477_)
);

OAI21X1 _14139_ (
    .A(_5888_),
    .B(_6454_),
    .C(\genblk1[7].u_ce.Yin12b [9]),
    .Y(_6478_)
);

OAI21X1 _14140_ (
    .A(_6477_),
    .B(_6459_),
    .C(_6478_),
    .Y(_5875_)
);

NAND2X1 _14141_ (
    .A(\genblk1[7].u_ce.Yin12b [6]),
    .B(_6463_),
    .Y(_6479_)
);

OAI21X1 _14142_ (
    .A(_6475_),
    .B(_6463_),
    .C(_6479_),
    .Y(_5876_)
);

NAND2X1 _14143_ (
    .A(\genblk1[7].u_ce.Yin12b [7]),
    .B(_6463_),
    .Y(_6480_)
);

OAI21X1 _14144_ (
    .A(_6477_),
    .B(_6463_),
    .C(_6480_),
    .Y(_5877_)
);

NAND2X1 _14145_ (
    .A(\genblk1[6].u_ce.Y_ [0]),
    .B(_6466_),
    .Y(_6481_)
);

OAI21X1 _14146_ (
    .A(_6046_),
    .B(_6466_),
    .C(_6481_),
    .Y(_5878_)
);

NAND2X1 _14147_ (
    .A(\genblk1[6].u_ce.Y_ [1]),
    .B(_6466_),
    .Y(_6482_)
);

OAI21X1 _14148_ (
    .A(_6067_),
    .B(_6466_),
    .C(_6482_),
    .Y(_5879_)
);

OAI21X1 _14149_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Yin1 [0]),
    .Y(_6483_)
);

OAI21X1 _14150_ (
    .A(_6475_),
    .B(_5887_),
    .C(_6483_),
    .Y(_5880_)
);

OAI21X1 _14151_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5885_),
    .C(\genblk1[7].u_ce.Yin1 [1]),
    .Y(_6484_)
);

OAI21X1 _14152_ (
    .A(_6477_),
    .B(_5887_),
    .C(_6484_),
    .Y(_5881_)
);

NAND2X1 _14153_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6485_)
);

OAI21X1 _14154_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5924_),
    .C(_6485_),
    .Y(_5882_)
);

NAND2X1 _14155_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6486_)
);

OAI21X1 _14156_ (
    .A(\genblk1[7].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5962_),
    .C(_6486_),
    .Y(_5883_)
);

NAND2X1 _14157_ (
    .A(\a[7] [1]),
    .B(_6455_),
    .Y(_6487_)
);

OAI21X1 _14158_ (
    .A(_5963__bF$buf0),
    .B(_6455_),
    .C(_6487_),
    .Y(_5884_)
);

DFFPOSX1 _14159_ (
    .CLK(clk_bF$buf1),
    .D(_5835_),
    .Q(\genblk1[7].u_ce.Ycalc [0])
);

DFFPOSX1 _14160_ (
    .CLK(clk_bF$buf0),
    .D(_5836_),
    .Q(\genblk1[7].u_ce.Ycalc [1])
);

DFFPOSX1 _14161_ (
    .CLK(clk_bF$buf78),
    .D(_5837_),
    .Q(\genblk1[7].u_ce.ISout )
);

DFFPOSX1 _14162_ (
    .CLK(clk_bF$buf77),
    .D(_5838_),
    .Q(\genblk1[7].u_ce.Ycalc [2])
);

DFFPOSX1 _14163_ (
    .CLK(clk_bF$buf76),
    .D(_5839_),
    .Q(\genblk1[7].u_ce.Ycalc [3])
);

DFFPOSX1 _14164_ (
    .CLK(clk_bF$buf75),
    .D(_5840_),
    .Q(\genblk1[7].u_ce.Ycalc [4])
);

DFFPOSX1 _14165_ (
    .CLK(clk_bF$buf74),
    .D(_5841_),
    .Q(\genblk1[7].u_ce.Ycalc [5])
);

DFFPOSX1 _14166_ (
    .CLK(clk_bF$buf73),
    .D(_5842_),
    .Q(\genblk1[7].u_ce.Ycalc [6])
);

DFFPOSX1 _14167_ (
    .CLK(clk_bF$buf72),
    .D(_5843_),
    .Q(\genblk1[7].u_ce.Ycalc [7])
);

DFFPOSX1 _14168_ (
    .CLK(clk_bF$buf71),
    .D(_5844_),
    .Q(\genblk1[7].u_ce.Ycalc [8])
);

DFFPOSX1 _14169_ (
    .CLK(clk_bF$buf70),
    .D(_5845_),
    .Q(\genblk1[7].u_ce.Ycalc [9])
);

DFFPOSX1 _14170_ (
    .CLK(clk_bF$buf69),
    .D(_5846_),
    .Q(\genblk1[7].u_ce.Ycalc [10])
);

DFFPOSX1 _14171_ (
    .CLK(clk_bF$buf68),
    .D(_5847_),
    .Q(\genblk1[7].u_ce.Ycalc [11])
);

DFFPOSX1 _14172_ (
    .CLK(clk_bF$buf67),
    .D(_5848_),
    .Q(\genblk1[7].u_ce.Xcalc [0])
);

DFFPOSX1 _14173_ (
    .CLK(clk_bF$buf66),
    .D(_5849_),
    .Q(\genblk1[7].u_ce.Xcalc [1])
);

DFFPOSX1 _14174_ (
    .CLK(clk_bF$buf65),
    .D(_5850_),
    .Q(\genblk1[7].u_ce.Xcalc [2])
);

DFFPOSX1 _14175_ (
    .CLK(clk_bF$buf64),
    .D(_5851_),
    .Q(\genblk1[7].u_ce.Xcalc [3])
);

DFFPOSX1 _14176_ (
    .CLK(clk_bF$buf63),
    .D(_5852_),
    .Q(\genblk1[7].u_ce.Xcalc [4])
);

DFFPOSX1 _14177_ (
    .CLK(clk_bF$buf62),
    .D(_5853_),
    .Q(\genblk1[7].u_ce.Xcalc [5])
);

DFFPOSX1 _14178_ (
    .CLK(clk_bF$buf61),
    .D(_5854_),
    .Q(\genblk1[7].u_ce.Xcalc [6])
);

DFFPOSX1 _14179_ (
    .CLK(clk_bF$buf60),
    .D(_5855_),
    .Q(\genblk1[7].u_ce.Xcalc [7])
);

DFFPOSX1 _14180_ (
    .CLK(clk_bF$buf59),
    .D(_5856_),
    .Q(\genblk1[7].u_ce.Xcalc [8])
);

DFFPOSX1 _14181_ (
    .CLK(clk_bF$buf58),
    .D(_5857_),
    .Q(\genblk1[7].u_ce.Xcalc [9])
);

DFFPOSX1 _14182_ (
    .CLK(clk_bF$buf57),
    .D(_5858_),
    .Q(\genblk1[7].u_ce.Xcalc [10])
);

DFFPOSX1 _14183_ (
    .CLK(clk_bF$buf56),
    .D(_5859_),
    .Q(\genblk1[7].u_ce.Xcalc [11])
);

DFFPOSX1 _14184_ (
    .CLK(clk_bF$buf55),
    .D(_5860_),
    .Q(\genblk1[7].u_ce.Xin12b [10])
);

DFFPOSX1 _14185_ (
    .CLK(clk_bF$buf54),
    .D(_5861_),
    .Q(\genblk1[7].u_ce.Xin12b [11])
);

DFFPOSX1 _14186_ (
    .CLK(clk_bF$buf53),
    .D(_5862_),
    .Q(\genblk1[7].u_ce.Xin12b [8])
);

DFFPOSX1 _14187_ (
    .CLK(clk_bF$buf52),
    .D(_5863_),
    .Q(\genblk1[7].u_ce.Xin12b [9])
);

DFFPOSX1 _14188_ (
    .CLK(clk_bF$buf51),
    .D(_5864_),
    .Q(\genblk1[7].u_ce.Xin12b [6])
);

DFFPOSX1 _14189_ (
    .CLK(clk_bF$buf50),
    .D(_5865_),
    .Q(\genblk1[7].u_ce.Xin12b [7])
);

DFFPOSX1 _14190_ (
    .CLK(clk_bF$buf49),
    .D(_5866_),
    .Q(\genblk1[7].u_ce.Xin12b [4])
);

DFFPOSX1 _14191_ (
    .CLK(clk_bF$buf48),
    .D(_5867_),
    .Q(\genblk1[7].u_ce.Xin12b [5])
);

DFFPOSX1 _14192_ (
    .CLK(clk_bF$buf47),
    .D(_5868_),
    .Q(\genblk1[7].u_ce.Xin1 [0])
);

DFFPOSX1 _14193_ (
    .CLK(clk_bF$buf46),
    .D(_5869_),
    .Q(\genblk1[7].u_ce.Xin1 [1])
);

DFFPOSX1 _14194_ (
    .CLK(clk_bF$buf45),
    .D(_5870_),
    .Q(\genblk1[7].u_ce.Xin0 [0])
);

DFFPOSX1 _14195_ (
    .CLK(clk_bF$buf44),
    .D(_5871_),
    .Q(\genblk1[7].u_ce.Xin0 [1])
);

DFFPOSX1 _14196_ (
    .CLK(clk_bF$buf43),
    .D(_5872_),
    .Q(\genblk1[7].u_ce.Yin12b [10])
);

DFFPOSX1 _14197_ (
    .CLK(clk_bF$buf42),
    .D(_5873_),
    .Q(\genblk1[7].u_ce.Yin12b [11])
);

DFFPOSX1 _14198_ (
    .CLK(clk_bF$buf41),
    .D(_5874_),
    .Q(\genblk1[7].u_ce.Yin12b [8])
);

DFFPOSX1 _14199_ (
    .CLK(clk_bF$buf40),
    .D(_5875_),
    .Q(\genblk1[7].u_ce.Yin12b [9])
);

DFFPOSX1 _14200_ (
    .CLK(clk_bF$buf39),
    .D(_5876_),
    .Q(\genblk1[7].u_ce.Yin12b [6])
);

DFFPOSX1 _14201_ (
    .CLK(clk_bF$buf38),
    .D(_5877_),
    .Q(\genblk1[7].u_ce.Yin12b [7])
);

DFFPOSX1 _14202_ (
    .CLK(clk_bF$buf37),
    .D(_5878_),
    .Q(\genblk1[7].u_ce.Yin12b [4])
);

DFFPOSX1 _14203_ (
    .CLK(clk_bF$buf36),
    .D(_5879_),
    .Q(\genblk1[7].u_ce.Yin12b [5])
);

DFFPOSX1 _14204_ (
    .CLK(clk_bF$buf35),
    .D(_5880_),
    .Q(\genblk1[7].u_ce.Yin1 [0])
);

DFFPOSX1 _14205_ (
    .CLK(clk_bF$buf34),
    .D(_5881_),
    .Q(\genblk1[7].u_ce.Yin1 [1])
);

DFFPOSX1 _14206_ (
    .CLK(clk_bF$buf33),
    .D(_5882_),
    .Q(\genblk1[7].u_ce.Yin0 [0])
);

DFFPOSX1 _14207_ (
    .CLK(clk_bF$buf32),
    .D(_5883_),
    .Q(\genblk1[7].u_ce.Yin0 [1])
);

DFFPOSX1 _14208_ (
    .CLK(clk_bF$buf31),
    .D(_5884_),
    .Q(\genblk1[7].u_ce.Ain12b [11])
);

DFFPOSX1 _14209_ (
    .CLK(clk_bF$buf30),
    .D(\genblk1[6].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[7].u_ce.LoadCtl [0])
);

DFFPOSX1 _14210_ (
    .CLK(clk_bF$buf29),
    .D(\genblk1[7].u_ce.LoadCtl_0_bF$buf1 ),
    .Q(\genblk1[7].u_ce.LoadCtl [1])
);

DFFPOSX1 _14211_ (
    .CLK(clk_bF$buf28),
    .D(\genblk1[7].u_ce.LoadCtl [1]),
    .Q(\genblk1[7].u_ce.LoadCtl [2])
);

DFFPOSX1 _14212_ (
    .CLK(clk_bF$buf27),
    .D(\genblk1[7].u_ce.LoadCtl [2]),
    .Q(\genblk1[7].u_ce.LoadCtl [3])
);

DFFPOSX1 _14213_ (
    .CLK(clk_bF$buf26),
    .D(\genblk1[7].u_ce.LoadCtl [3]),
    .Q(\genblk1[7].u_ce.LoadCtl [4])
);

DFFPOSX1 _14214_ (
    .CLK(clk_bF$buf25),
    .D(\genblk1[7].u_ce.LoadCtl [4]),
    .Q(\genblk1[7].u_ce.LoadCtl [5])
);

DFFPOSX1 _14215_ (
    .CLK(clk_bF$buf24),
    .D(\genblk1[7].u_ce.LoadCtl [5]),
    .Q(\genblk1[7].u_ce.Vld )
);

INVX1 _14216_ (
    .A(\u_ot.Ycalc [0]),
    .Y(_6537_)
);

NAND2X1 _14217_ (
    .A(\u_ot.Xcalc [0]),
    .B(selXY_bF$buf3),
    .Y(_6538_)
);

OAI21X1 _14218_ (
    .A(selXY_bF$buf2),
    .B(_6537_),
    .C(_6538_),
    .Y(_7071_[0])
);

INVX1 _14219_ (
    .A(\u_ot.Ycalc [1]),
    .Y(_6539_)
);

NAND2X1 _14220_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [1]),
    .Y(_6540_)
);

OAI21X1 _14221_ (
    .A(selXY_bF$buf0),
    .B(_6539_),
    .C(_6540_),
    .Y(_7071_[1])
);

INVX1 _14222_ (
    .A(\u_ot.Ycalc [2]),
    .Y(_6541_)
);

NAND2X1 _14223_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [2]),
    .Y(_6542_)
);

OAI21X1 _14224_ (
    .A(selXY_bF$buf2),
    .B(_6541_),
    .C(_6542_),
    .Y(_7071_[2])
);

INVX1 _14225_ (
    .A(\u_ot.Ycalc [3]),
    .Y(_6543_)
);

NAND2X1 _14226_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [3]),
    .Y(_6544_)
);

OAI21X1 _14227_ (
    .A(selXY_bF$buf0),
    .B(_6543_),
    .C(_6544_),
    .Y(_7071_[3])
);

INVX1 _14228_ (
    .A(\u_ot.Ycalc [4]),
    .Y(_6545_)
);

NAND2X1 _14229_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [4]),
    .Y(_6546_)
);

OAI21X1 _14230_ (
    .A(selXY_bF$buf2),
    .B(_6545_),
    .C(_6546_),
    .Y(_7071_[4])
);

INVX1 _14231_ (
    .A(\u_ot.Ycalc [5]),
    .Y(_6547_)
);

NAND2X1 _14232_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [5]),
    .Y(_6548_)
);

OAI21X1 _14233_ (
    .A(selXY_bF$buf0),
    .B(_6547_),
    .C(_6548_),
    .Y(_7071_[5])
);

INVX1 _14234_ (
    .A(\u_ot.Ycalc [6]),
    .Y(_6549_)
);

NAND2X1 _14235_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [6]),
    .Y(_6550_)
);

OAI21X1 _14236_ (
    .A(selXY_bF$buf2),
    .B(_6549_),
    .C(_6550_),
    .Y(_7071_[6])
);

INVX1 _14237_ (
    .A(\u_ot.Ycalc [7]),
    .Y(_6551_)
);

NAND2X1 _14238_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [7]),
    .Y(_6552_)
);

OAI21X1 _14239_ (
    .A(selXY_bF$buf0),
    .B(_6551_),
    .C(_6552_),
    .Y(_7071_[7])
);

INVX1 _14240_ (
    .A(\u_ot.Ycalc [8]),
    .Y(_6553_)
);

NAND2X1 _14241_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [8]),
    .Y(_6554_)
);

OAI21X1 _14242_ (
    .A(selXY_bF$buf2),
    .B(_6553_),
    .C(_6554_),
    .Y(_7071_[8])
);

INVX1 _14243_ (
    .A(\u_ot.Ycalc [9]),
    .Y(_6555_)
);

NAND2X1 _14244_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [9]),
    .Y(_6556_)
);

OAI21X1 _14245_ (
    .A(selXY_bF$buf0),
    .B(_6555_),
    .C(_6556_),
    .Y(_7071_[9])
);

INVX1 _14246_ (
    .A(\u_ot.Ycalc [10]),
    .Y(_6557_)
);

NAND2X1 _14247_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [10]),
    .Y(_6558_)
);

OAI21X1 _14248_ (
    .A(selXY_bF$buf2),
    .B(_6557_),
    .C(_6558_),
    .Y(_7071_[10])
);

INVX1 _14249_ (
    .A(\u_ot.Ycalc [11]),
    .Y(_6559_)
);

NAND2X1 _14250_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [11]),
    .Y(_6560_)
);

OAI21X1 _14251_ (
    .A(selXY_bF$buf0),
    .B(_6559_),
    .C(_6560_),
    .Y(_7071_[11])
);

INVX1 _14252_ (
    .A(\u_ot.Xin0 [0]),
    .Y(_6561_)
);

INVX8 _14253_ (
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .Y(_6562_)
);

NAND2X1 _14254_ (
    .A(\u_ot.Xcalc [0]),
    .B(_6562__bF$buf4),
    .Y(_6563_)
);

OAI21X1 _14255_ (
    .A(_6561_),
    .B(_6562__bF$buf3),
    .C(_6563_),
    .Y(_6488_)
);

NAND3X1 _14256_ (
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Xin0 [0]),
    .C(\u_ot.Xin0 [1]),
    .Y(_6564_)
);

INVX4 _14257_ (
    .A(\u_ot.ISreg_bF$buf3 ),
    .Y(_6565_)
);

INVX1 _14258_ (
    .A(\u_ot.Xin0 [1]),
    .Y(_6566_)
);

OAI21X1 _14259_ (
    .A(_6565_),
    .B(_6561_),
    .C(_6566_),
    .Y(_6567_)
);

NAND2X1 _14260_ (
    .A(_6564_),
    .B(_6567_),
    .Y(_6568_)
);

NAND2X1 _14261_ (
    .A(\u_ot.Xcalc [1]),
    .B(_6562__bF$buf2),
    .Y(_6569_)
);

OAI21X1 _14262_ (
    .A(_6562__bF$buf1),
    .B(_6568_),
    .C(_6569_),
    .Y(_6489_)
);

INVX1 _14263_ (
    .A(\u_ot.Xin1 [0]),
    .Y(_6570_)
);

OAI21X1 _14264_ (
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .C(\u_ot.ISreg_bF$buf2 ),
    .Y(_6571_)
);

OR2X2 _14265_ (
    .A(_6571_),
    .B(_6570_),
    .Y(_6572_)
);

NOR2X1 _14266_ (
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .Y(_6573_)
);

OAI21X1 _14267_ (
    .A(_6565_),
    .B(_6573_),
    .C(_6570_),
    .Y(_6574_)
);

NAND2X1 _14268_ (
    .A(_6574_),
    .B(_6572_),
    .Y(_6575_)
);

NAND2X1 _14269_ (
    .A(\u_ot.Xcalc [2]),
    .B(_6562__bF$buf0),
    .Y(_6576_)
);

OAI21X1 _14270_ (
    .A(_6562__bF$buf4),
    .B(_6575_),
    .C(_6576_),
    .Y(_6490_)
);

OAI21X1 _14271_ (
    .A(_6565_),
    .B(_6570_),
    .C(_6571_),
    .Y(_6577_)
);

NAND2X1 _14272_ (
    .A(\u_ot.Xin1 [1]),
    .B(_6577_),
    .Y(_6578_)
);

OR2X2 _14273_ (
    .A(_6577_),
    .B(\u_ot.Xin1 [1]),
    .Y(_6579_)
);

NAND2X1 _14274_ (
    .A(_6578_),
    .B(_6579_),
    .Y(_6580_)
);

NAND2X1 _14275_ (
    .A(\u_ot.Xcalc [3]),
    .B(_6562__bF$buf3),
    .Y(_6581_)
);

OAI21X1 _14276_ (
    .A(_6562__bF$buf2),
    .B(_6580_),
    .C(_6581_),
    .Y(_6491_)
);

NOR2X1 _14277_ (
    .A(\u_ot.Xin1 [0]),
    .B(\u_ot.Xin1 [1]),
    .Y(_6582_)
);

NAND2X1 _14278_ (
    .A(_6573_),
    .B(_6582_),
    .Y(_6583_)
);

NAND3X1 _14279_ (
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(\u_ot.Xin12b [4]),
    .C(_6583_),
    .Y(_6584_)
);

INVX1 _14280_ (
    .A(\u_ot.Xin12b [4]),
    .Y(_6585_)
);

AND2X2 _14281_ (
    .A(_6573_),
    .B(_6582_),
    .Y(_6586_)
);

OAI21X1 _14282_ (
    .A(_6565_),
    .B(_6586_),
    .C(_6585_),
    .Y(_6587_)
);

NAND2X1 _14283_ (
    .A(_6584_),
    .B(_6587_),
    .Y(_6588_)
);

NAND2X1 _14284_ (
    .A(\u_ot.Xcalc [4]),
    .B(_6562__bF$buf1),
    .Y(_6589_)
);

OAI21X1 _14285_ (
    .A(_6562__bF$buf0),
    .B(_6588_),
    .C(_6589_),
    .Y(_6492_)
);

INVX1 _14286_ (
    .A(\u_ot.Xcalc [5]),
    .Y(_6590_)
);

OAI21X1 _14287_ (
    .A(\u_ot.Xin12b [4]),
    .B(_6583_),
    .C(\u_ot.ISreg_bF$buf0 ),
    .Y(_6591_)
);

NAND2X1 _14288_ (
    .A(\u_ot.Xin12b [5]),
    .B(_6591_),
    .Y(_6592_)
);

NOR2X1 _14289_ (
    .A(\u_ot.Xin12b [5]),
    .B(_6591_),
    .Y(_6593_)
);

NOR2X1 _14290_ (
    .A(_6562__bF$buf4),
    .B(_6593_),
    .Y(_6594_)
);

AOI22X1 _14291_ (
    .A(_6590_),
    .B(_6562__bF$buf3),
    .C(_6594_),
    .D(_6592_),
    .Y(_6493_)
);

NOR2X1 _14292_ (
    .A(\u_ot.Xin12b [4]),
    .B(\u_ot.Xin12b [5]),
    .Y(_6595_)
);

NAND2X1 _14293_ (
    .A(_6595_),
    .B(_6586_),
    .Y(_6596_)
);

NAND3X1 _14294_ (
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Xin12b [6]),
    .C(_6596_),
    .Y(_6597_)
);

INVX1 _14295_ (
    .A(\u_ot.Xin12b [6]),
    .Y(_6598_)
);

NAND2X1 _14296_ (
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(_6596_),
    .Y(_6599_)
);

NAND2X1 _14297_ (
    .A(_6598_),
    .B(_6599_),
    .Y(_6600_)
);

NAND2X1 _14298_ (
    .A(_6597_),
    .B(_6600_),
    .Y(_6601_)
);

NAND2X1 _14299_ (
    .A(\u_ot.Xcalc [6]),
    .B(_6562__bF$buf2),
    .Y(_6602_)
);

OAI21X1 _14300_ (
    .A(_6562__bF$buf1),
    .B(_6601_),
    .C(_6602_),
    .Y(_6494_)
);

INVX1 _14301_ (
    .A(\u_ot.Xcalc [7]),
    .Y(_6603_)
);

NAND3X1 _14302_ (
    .A(_6598_),
    .B(_6595_),
    .C(_6586_),
    .Y(_6604_)
);

NAND3X1 _14303_ (
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Xin12b [7]),
    .C(_6604_),
    .Y(_6605_)
);

INVX1 _14304_ (
    .A(\u_ot.Xin12b [7]),
    .Y(_6606_)
);

NAND2X1 _14305_ (
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(\u_ot.Xin12b [6]),
    .Y(_6607_)
);

NAND3X1 _14306_ (
    .A(_6606_),
    .B(_6607_),
    .C(_6599_),
    .Y(_6608_)
);

NAND3X1 _14307_ (
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6605_),
    .C(_6608_),
    .Y(_6609_)
);

OAI21X1 _14308_ (
    .A(_6603_),
    .B(\u_ot.LoadCtl_6_bF$buf2 ),
    .C(_6609_),
    .Y(_6495_)
);

INVX1 _14309_ (
    .A(\u_ot.Xin12b [8]),
    .Y(_6610_)
);

NOR2X1 _14310_ (
    .A(\u_ot.Xin12b [6]),
    .B(\u_ot.Xin12b [7]),
    .Y(_6611_)
);

NAND2X1 _14311_ (
    .A(_6595_),
    .B(_6611_),
    .Y(_6612_)
);

OAI21X1 _14312_ (
    .A(_6583_),
    .B(_6612_),
    .C(\u_ot.ISreg_bF$buf0 ),
    .Y(_6613_)
);

OR2X2 _14313_ (
    .A(_6613_),
    .B(_6610_),
    .Y(_6614_)
);

NAND2X1 _14314_ (
    .A(_6610_),
    .B(_6613_),
    .Y(_6615_)
);

NAND2X1 _14315_ (
    .A(_6615_),
    .B(_6614_),
    .Y(_6616_)
);

NAND2X1 _14316_ (
    .A(\u_ot.Xcalc [8]),
    .B(_6562__bF$buf0),
    .Y(_6617_)
);

OAI21X1 _14317_ (
    .A(_6562__bF$buf4),
    .B(_6616_),
    .C(_6617_),
    .Y(_6496_)
);

INVX1 _14318_ (
    .A(\u_ot.Xcalc [9]),
    .Y(_6618_)
);

INVX1 _14319_ (
    .A(\u_ot.Xin12b [9]),
    .Y(_6619_)
);

OAI21X1 _14320_ (
    .A(_6565_),
    .B(_6610_),
    .C(_6613_),
    .Y(_6620_)
);

OR2X2 _14321_ (
    .A(_6620_),
    .B(_6619_),
    .Y(_6621_)
);

AOI21X1 _14322_ (
    .A(_6620_),
    .B(_6619_),
    .C(_6562__bF$buf3),
    .Y(_6622_)
);

AOI22X1 _14323_ (
    .A(_6618_),
    .B(_6562__bF$buf2),
    .C(_6621_),
    .D(_6622_),
    .Y(_6497_)
);

INVX1 _14324_ (
    .A(\u_ot.Xcalc [10]),
    .Y(_6623_)
);

AND2X2 _14325_ (
    .A(_6595_),
    .B(_6611_),
    .Y(_6624_)
);

NOR2X1 _14326_ (
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .Y(_6625_)
);

NAND3X1 _14327_ (
    .A(_6625_),
    .B(_6586_),
    .C(_6624_),
    .Y(_6626_)
);

NAND3X1 _14328_ (
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Xin12b [10]),
    .C(_6626_),
    .Y(_6627_)
);

INVX1 _14329_ (
    .A(\u_ot.Xin12b [10]),
    .Y(_6628_)
);

NAND2X1 _14330_ (
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(_6626_),
    .Y(_6629_)
);

NAND2X1 _14331_ (
    .A(_6628_),
    .B(_6629_),
    .Y(_6630_)
);

NAND3X1 _14332_ (
    .A(\u_ot.LoadCtl_6_bF$buf1 ),
    .B(_6627_),
    .C(_6630_),
    .Y(_6631_)
);

OAI21X1 _14333_ (
    .A(_6623_),
    .B(\u_ot.LoadCtl_6_bF$buf0 ),
    .C(_6631_),
    .Y(_6498_)
);

NAND2X1 _14334_ (
    .A(\u_ot.Xcalc [11]),
    .B(_6562__bF$buf1),
    .Y(_6632_)
);

INVX1 _14335_ (
    .A(\u_ot.Xin12b [11]),
    .Y(_6633_)
);

NAND2X1 _14336_ (
    .A(selSign),
    .B(_6633_),
    .Y(_6634_)
);

INVX1 _14337_ (
    .A(selSign),
    .Y(_6635_)
);

NAND2X1 _14338_ (
    .A(\u_ot.Xin12b [11]),
    .B(_6635_),
    .Y(_6636_)
);

NAND2X1 _14339_ (
    .A(_6634_),
    .B(_6636_),
    .Y(_6637_)
);

INVX1 _14340_ (
    .A(_6637_),
    .Y(_6638_)
);

NAND2X1 _14341_ (
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Xin12b [10]),
    .Y(_6639_)
);

NAND3X1 _14342_ (
    .A(_6638_),
    .B(_6639_),
    .C(_6629_),
    .Y(_6640_)
);

OAI21X1 _14343_ (
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .C(\u_ot.ISreg_bF$buf1 ),
    .Y(_6641_)
);

NAND3X1 _14344_ (
    .A(_6641_),
    .B(_6639_),
    .C(_6613_),
    .Y(_6642_)
);

NAND2X1 _14345_ (
    .A(_6637_),
    .B(_6642_),
    .Y(_6643_)
);

NAND3X1 _14346_ (
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .B(_6643_),
    .C(_6640_),
    .Y(_6644_)
);

NAND2X1 _14347_ (
    .A(_6632_),
    .B(_6644_),
    .Y(_6499_)
);

NAND2X1 _14348_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.LoadCtl_6_bF$buf3 ),
    .Y(_6645_)
);

OAI21X1 _14349_ (
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6537_),
    .C(_6645_),
    .Y(_6500_)
);

NAND3X1 _14350_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .C(\u_ot.ISreg_bF$buf0 ),
    .Y(_6646_)
);

INVX1 _14351_ (
    .A(\u_ot.Yin0 [0]),
    .Y(_6647_)
);

INVX1 _14352_ (
    .A(\u_ot.Yin0 [1]),
    .Y(_6648_)
);

OAI21X1 _14353_ (
    .A(_6647_),
    .B(_6565_),
    .C(_6648_),
    .Y(_6649_)
);

NAND3X1 _14354_ (
    .A(\u_ot.LoadCtl_6_bF$buf1 ),
    .B(_6646_),
    .C(_6649_),
    .Y(_6650_)
);

OAI21X1 _14355_ (
    .A(_6539_),
    .B(\u_ot.LoadCtl_6_bF$buf0 ),
    .C(_6650_),
    .Y(_6501_)
);

INVX1 _14356_ (
    .A(\u_ot.Yin1 [0]),
    .Y(_6651_)
);

OAI21X1 _14357_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .C(\u_ot.ISreg_bF$buf4 ),
    .Y(_6652_)
);

OR2X2 _14358_ (
    .A(_6652_),
    .B(_6651_),
    .Y(_6653_)
);

NOR2X1 _14359_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .Y(_6654_)
);

OAI21X1 _14360_ (
    .A(_6565_),
    .B(_6654_),
    .C(_6651_),
    .Y(_6655_)
);

NAND3X1 _14361_ (
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .B(_6655_),
    .C(_6653_),
    .Y(_6656_)
);

OAI21X1 _14362_ (
    .A(_6541_),
    .B(\u_ot.LoadCtl_6_bF$buf3 ),
    .C(_6656_),
    .Y(_6502_)
);

OAI21X1 _14363_ (
    .A(_6565_),
    .B(_6651_),
    .C(_6652_),
    .Y(_6657_)
);

NAND2X1 _14364_ (
    .A(\u_ot.Yin1 [1]),
    .B(_6657_),
    .Y(_6658_)
);

OR2X2 _14365_ (
    .A(_6657_),
    .B(\u_ot.Yin1 [1]),
    .Y(_6659_)
);

NAND3X1 _14366_ (
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6658_),
    .C(_6659_),
    .Y(_6660_)
);

OAI21X1 _14367_ (
    .A(_6543_),
    .B(\u_ot.LoadCtl_6_bF$buf1 ),
    .C(_6660_),
    .Y(_6503_)
);

INVX1 _14368_ (
    .A(\u_ot.Yin12b [4]),
    .Y(_6661_)
);

NOR2X1 _14369_ (
    .A(\u_ot.Yin1 [0]),
    .B(\u_ot.Yin1 [1]),
    .Y(_6662_)
);

NAND2X1 _14370_ (
    .A(_6654_),
    .B(_6662_),
    .Y(_6663_)
);

NAND2X1 _14371_ (
    .A(\u_ot.ISreg_bF$buf3 ),
    .B(_6663_),
    .Y(_6664_)
);

OR2X2 _14372_ (
    .A(_6664_),
    .B(_6661_),
    .Y(_6665_)
);

AND2X2 _14373_ (
    .A(_6654_),
    .B(_6662_),
    .Y(_6666_)
);

OAI21X1 _14374_ (
    .A(_6565_),
    .B(_6666_),
    .C(_6661_),
    .Y(_6667_)
);

NAND3X1 _14375_ (
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6667_),
    .C(_6665_),
    .Y(_6668_)
);

OAI21X1 _14376_ (
    .A(_6545_),
    .B(\u_ot.LoadCtl_6_bF$buf4 ),
    .C(_6668_),
    .Y(_6504_)
);

INVX1 _14377_ (
    .A(\u_ot.Yin12b [5]),
    .Y(_6669_)
);

OAI21X1 _14378_ (
    .A(_6565_),
    .B(_6661_),
    .C(_6664_),
    .Y(_6670_)
);

OR2X2 _14379_ (
    .A(_6670_),
    .B(_6669_),
    .Y(_6671_)
);

AOI21X1 _14380_ (
    .A(_6670_),
    .B(_6669_),
    .C(_6562__bF$buf0),
    .Y(_6672_)
);

AOI22X1 _14381_ (
    .A(_6547_),
    .B(_6562__bF$buf4),
    .C(_6671_),
    .D(_6672_),
    .Y(_6505_)
);

NOR2X1 _14382_ (
    .A(\u_ot.Yin12b [4]),
    .B(\u_ot.Yin12b [5]),
    .Y(_6673_)
);

NAND2X1 _14383_ (
    .A(_6673_),
    .B(_6666_),
    .Y(_6674_)
);

NAND3X1 _14384_ (
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Yin12b [6]),
    .C(_6674_),
    .Y(_6675_)
);

INVX1 _14385_ (
    .A(\u_ot.Yin12b [6]),
    .Y(_6676_)
);

NAND2X1 _14386_ (
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(_6674_),
    .Y(_6677_)
);

NAND2X1 _14387_ (
    .A(_6676_),
    .B(_6677_),
    .Y(_6678_)
);

NAND3X1 _14388_ (
    .A(\u_ot.LoadCtl_6_bF$buf3 ),
    .B(_6675_),
    .C(_6678_),
    .Y(_6679_)
);

OAI21X1 _14389_ (
    .A(_6549_),
    .B(\u_ot.LoadCtl_6_bF$buf2 ),
    .C(_6679_),
    .Y(_6506_)
);

NAND3X1 _14390_ (
    .A(_6676_),
    .B(_6673_),
    .C(_6666_),
    .Y(_6680_)
);

NAND3X1 _14391_ (
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(\u_ot.Yin12b [7]),
    .C(_6680_),
    .Y(_6681_)
);

INVX1 _14392_ (
    .A(\u_ot.Yin12b [7]),
    .Y(_6682_)
);

NAND2X1 _14393_ (
    .A(\u_ot.ISreg_bF$buf4 ),
    .B(\u_ot.Yin12b [6]),
    .Y(_6683_)
);

NAND3X1 _14394_ (
    .A(_6682_),
    .B(_6683_),
    .C(_6677_),
    .Y(_6684_)
);

NAND3X1 _14395_ (
    .A(\u_ot.LoadCtl_6_bF$buf1 ),
    .B(_6681_),
    .C(_6684_),
    .Y(_6685_)
);

OAI21X1 _14396_ (
    .A(_6551_),
    .B(\u_ot.LoadCtl_6_bF$buf0 ),
    .C(_6685_),
    .Y(_6507_)
);

INVX1 _14397_ (
    .A(\u_ot.Yin12b [8]),
    .Y(_6686_)
);

NOR2X1 _14398_ (
    .A(\u_ot.Yin12b [6]),
    .B(\u_ot.Yin12b [7]),
    .Y(_6687_)
);

NAND2X1 _14399_ (
    .A(_6673_),
    .B(_6687_),
    .Y(_6688_)
);

OAI21X1 _14400_ (
    .A(_6663_),
    .B(_6688_),
    .C(\u_ot.ISreg_bF$buf3 ),
    .Y(_6689_)
);

OR2X2 _14401_ (
    .A(_6689_),
    .B(_6686_),
    .Y(_6690_)
);

NAND2X1 _14402_ (
    .A(_6686_),
    .B(_6689_),
    .Y(_6691_)
);

NAND2X1 _14403_ (
    .A(_6691_),
    .B(_6690_),
    .Y(_6692_)
);

NAND2X1 _14404_ (
    .A(\u_ot.Ycalc [8]),
    .B(_6562__bF$buf3),
    .Y(_6693_)
);

OAI21X1 _14405_ (
    .A(_6562__bF$buf2),
    .B(_6692_),
    .C(_6693_),
    .Y(_6508_)
);

INVX1 _14406_ (
    .A(\u_ot.Yin12b [9]),
    .Y(_6694_)
);

OAI21X1 _14407_ (
    .A(_6565_),
    .B(_6686_),
    .C(_6689_),
    .Y(_6695_)
);

OR2X2 _14408_ (
    .A(_6695_),
    .B(_6694_),
    .Y(_6696_)
);

AOI21X1 _14409_ (
    .A(_6695_),
    .B(_6694_),
    .C(_6562__bF$buf1),
    .Y(_6697_)
);

AOI22X1 _14410_ (
    .A(_6555_),
    .B(_6562__bF$buf0),
    .C(_6696_),
    .D(_6697_),
    .Y(_6509_)
);

AND2X2 _14411_ (
    .A(_6673_),
    .B(_6687_),
    .Y(_6698_)
);

NOR2X1 _14412_ (
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .Y(_6699_)
);

NAND3X1 _14413_ (
    .A(_6699_),
    .B(_6666_),
    .C(_6698_),
    .Y(_6700_)
);

NAND3X1 _14414_ (
    .A(\u_ot.ISreg_bF$buf2 ),
    .B(\u_ot.Yin12b [10]),
    .C(_6700_),
    .Y(_6701_)
);

INVX1 _14415_ (
    .A(\u_ot.Yin12b [10]),
    .Y(_6702_)
);

NAND2X1 _14416_ (
    .A(\u_ot.ISreg_bF$buf1 ),
    .B(_6700_),
    .Y(_6703_)
);

NAND2X1 _14417_ (
    .A(_6702_),
    .B(_6703_),
    .Y(_6704_)
);

NAND3X1 _14418_ (
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .B(_6701_),
    .C(_6704_),
    .Y(_6705_)
);

OAI21X1 _14419_ (
    .A(_6557_),
    .B(\u_ot.LoadCtl_6_bF$buf3 ),
    .C(_6705_),
    .Y(_6510_)
);

NAND2X1 _14420_ (
    .A(\u_ot.Ycalc [11]),
    .B(_6562__bF$buf4),
    .Y(_6706_)
);

INVX1 _14421_ (
    .A(\u_ot.Yin12b [11]),
    .Y(_6707_)
);

NAND2X1 _14422_ (
    .A(selSign),
    .B(_6707_),
    .Y(_6708_)
);

NAND2X1 _14423_ (
    .A(\u_ot.Yin12b [11]),
    .B(_6635_),
    .Y(_6709_)
);

NAND2X1 _14424_ (
    .A(_6708_),
    .B(_6709_),
    .Y(_6710_)
);

INVX1 _14425_ (
    .A(_6710_),
    .Y(_6711_)
);

NAND2X1 _14426_ (
    .A(\u_ot.ISreg_bF$buf0 ),
    .B(\u_ot.Yin12b [10]),
    .Y(_6712_)
);

NAND3X1 _14427_ (
    .A(_6711_),
    .B(_6712_),
    .C(_6703_),
    .Y(_6713_)
);

OAI21X1 _14428_ (
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .C(\u_ot.ISreg_bF$buf4 ),
    .Y(_6714_)
);

NAND3X1 _14429_ (
    .A(_6714_),
    .B(_6712_),
    .C(_6689_),
    .Y(_6715_)
);

NAND2X1 _14430_ (
    .A(_6710_),
    .B(_6715_),
    .Y(_6716_)
);

NAND3X1 _14431_ (
    .A(\u_ot.LoadCtl_6_bF$buf2 ),
    .B(_6716_),
    .C(_6713_),
    .Y(_6717_)
);

NAND2X1 _14432_ (
    .A(_6706_),
    .B(_6717_),
    .Y(_6511_)
);

INVX2 _14433_ (
    .A(\u_ot.LoadCtl [1]),
    .Y(_6718_)
);

NOR2X1 _14434_ (
    .A(\u_ot.LoadCtl [2]),
    .B(\u_ot.LoadCtl [0]),
    .Y(_6719_)
);

AND2X2 _14435_ (
    .A(_6719_),
    .B(_6718_),
    .Y(_6720_)
);

INVX1 _14436_ (
    .A(\u_ot.LoadCtl [4]),
    .Y(_6721_)
);

NAND2X1 _14437_ (
    .A(\u_ot.LoadCtl [5]),
    .B(_6721_),
    .Y(_6722_)
);

NOR2X1 _14438_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6722_),
    .Y(_6723_)
);

AND2X2 _14439_ (
    .A(_6723_),
    .B(_6720_),
    .Y(_6724_)
);

NAND2X1 _14440_ (
    .A(\genblk1[7].u_ce.X_ [0]),
    .B(_6724_),
    .Y(_6725_)
);

OAI21X1 _14441_ (
    .A(_6628_),
    .B(_6724_),
    .C(_6725_),
    .Y(_6512_)
);

NAND2X1 _14442_ (
    .A(\genblk1[7].u_ce.X_ [1]),
    .B(_6724_),
    .Y(_6726_)
);

OAI21X1 _14443_ (
    .A(_6633_),
    .B(_6724_),
    .C(_6726_),
    .Y(_6513_)
);

INVX1 _14444_ (
    .A(\genblk1[7].u_ce.X_ [0]),
    .Y(_6727_)
);

NOR2X1 _14445_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6721_),
    .Y(_6728_)
);

NAND2X1 _14446_ (
    .A(_6728_),
    .B(_6720_),
    .Y(_6729_)
);

NAND2X1 _14447_ (
    .A(\u_ot.Xin12b [8]),
    .B(_6729_),
    .Y(_6730_)
);

OAI21X1 _14448_ (
    .A(_6727_),
    .B(_6729_),
    .C(_6730_),
    .Y(_6514_)
);

INVX1 _14449_ (
    .A(\genblk1[7].u_ce.X_ [1]),
    .Y(_6731_)
);

NAND2X1 _14450_ (
    .A(\u_ot.Xin12b [9]),
    .B(_6729_),
    .Y(_6732_)
);

OAI21X1 _14451_ (
    .A(_6731_),
    .B(_6729_),
    .C(_6732_),
    .Y(_6515_)
);

NAND2X1 _14452_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6720_),
    .Y(_6733_)
);

NAND2X1 _14453_ (
    .A(\u_ot.Xin12b [6]),
    .B(_6733_),
    .Y(_6734_)
);

OAI21X1 _14454_ (
    .A(_6727_),
    .B(_6733_),
    .C(_6734_),
    .Y(_6516_)
);

NAND2X1 _14455_ (
    .A(\u_ot.Xin12b [7]),
    .B(_6733_),
    .Y(_6735_)
);

OAI21X1 _14456_ (
    .A(_6731_),
    .B(_6733_),
    .C(_6735_),
    .Y(_6517_)
);

INVX1 _14457_ (
    .A(\u_ot.LoadCtl [0]),
    .Y(_6736_)
);

NAND3X1 _14458_ (
    .A(\u_ot.LoadCtl [2]),
    .B(_6718_),
    .C(_6736_),
    .Y(_6737_)
);

NAND2X1 _14459_ (
    .A(\u_ot.Xin12b [4]),
    .B(_6737_),
    .Y(_6738_)
);

OAI21X1 _14460_ (
    .A(_6727_),
    .B(_6737_),
    .C(_6738_),
    .Y(_6518_)
);

NAND2X1 _14461_ (
    .A(\u_ot.Xin12b [5]),
    .B(_6737_),
    .Y(_6739_)
);

OAI21X1 _14462_ (
    .A(_6731_),
    .B(_6737_),
    .C(_6739_),
    .Y(_6519_)
);

NAND2X1 _14463_ (
    .A(\u_ot.LoadCtl [1]),
    .B(_6736_),
    .Y(_6740_)
);

OAI21X1 _14464_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Xin1 [0]),
    .Y(_6741_)
);

OAI21X1 _14465_ (
    .A(_6727_),
    .B(_6740_),
    .C(_6741_),
    .Y(_6520_)
);

OAI21X1 _14466_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Xin1 [1]),
    .Y(_6742_)
);

OAI21X1 _14467_ (
    .A(_6731_),
    .B(_6740_),
    .C(_6742_),
    .Y(_6521_)
);

NAND2X1 _14468_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.X_ [0]),
    .Y(_6743_)
);

OAI21X1 _14469_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6561_),
    .C(_6743_),
    .Y(_6522_)
);

NAND2X1 _14470_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.X_ [1]),
    .Y(_6744_)
);

OAI21X1 _14471_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6566_),
    .C(_6744_),
    .Y(_6523_)
);

NAND2X1 _14472_ (
    .A(\genblk1[7].u_ce.Y_ [0]),
    .B(_6724_),
    .Y(_6745_)
);

OAI21X1 _14473_ (
    .A(_6702_),
    .B(_6724_),
    .C(_6745_),
    .Y(_6524_)
);

NAND2X1 _14474_ (
    .A(\genblk1[7].u_ce.Y_ [1]),
    .B(_6724_),
    .Y(_6746_)
);

OAI21X1 _14475_ (
    .A(_6707_),
    .B(_6724_),
    .C(_6746_),
    .Y(_6525_)
);

INVX1 _14476_ (
    .A(\genblk1[7].u_ce.Y_ [0]),
    .Y(_6747_)
);

NAND2X1 _14477_ (
    .A(\u_ot.Yin12b [8]),
    .B(_6729_),
    .Y(_6748_)
);

OAI21X1 _14478_ (
    .A(_6747_),
    .B(_6729_),
    .C(_6748_),
    .Y(_6526_)
);

INVX1 _14479_ (
    .A(\genblk1[7].u_ce.Y_ [1]),
    .Y(_6749_)
);

NAND2X1 _14480_ (
    .A(\u_ot.Yin12b [9]),
    .B(_6729_),
    .Y(_6750_)
);

OAI21X1 _14481_ (
    .A(_6749_),
    .B(_6729_),
    .C(_6750_),
    .Y(_6527_)
);

NAND2X1 _14482_ (
    .A(\u_ot.Yin12b [6]),
    .B(_6733_),
    .Y(_6751_)
);

OAI21X1 _14483_ (
    .A(_6747_),
    .B(_6733_),
    .C(_6751_),
    .Y(_6528_)
);

NAND2X1 _14484_ (
    .A(\u_ot.Yin12b [7]),
    .B(_6733_),
    .Y(_6752_)
);

OAI21X1 _14485_ (
    .A(_6749_),
    .B(_6733_),
    .C(_6752_),
    .Y(_6529_)
);

NAND2X1 _14486_ (
    .A(\u_ot.Yin12b [4]),
    .B(_6737_),
    .Y(_6753_)
);

OAI21X1 _14487_ (
    .A(_6747_),
    .B(_6737_),
    .C(_6753_),
    .Y(_6530_)
);

NAND2X1 _14488_ (
    .A(\u_ot.Yin12b [5]),
    .B(_6737_),
    .Y(_6754_)
);

OAI21X1 _14489_ (
    .A(_6749_),
    .B(_6737_),
    .C(_6754_),
    .Y(_6531_)
);

OAI21X1 _14490_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Yin1 [0]),
    .Y(_6755_)
);

OAI21X1 _14491_ (
    .A(_6747_),
    .B(_6740_),
    .C(_6755_),
    .Y(_6532_)
);

OAI21X1 _14492_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6718_),
    .C(\u_ot.Yin1 [1]),
    .Y(_6756_)
);

OAI21X1 _14493_ (
    .A(_6749_),
    .B(_6740_),
    .C(_6756_),
    .Y(_6533_)
);

NAND2X1 _14494_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.Y_ [0]),
    .Y(_6757_)
);

OAI21X1 _14495_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6647_),
    .C(_6757_),
    .Y(_6534_)
);

NAND2X1 _14496_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[7].u_ce.Y_ [1]),
    .Y(_6758_)
);

OAI21X1 _14497_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6648_),
    .C(_6758_),
    .Y(_6535_)
);

NAND2X1 _14498_ (
    .A(\u_ot.LoadCtl_6_bF$buf1 ),
    .B(\genblk1[7].u_ce.ISout ),
    .Y(_6759_)
);

OAI21X1 _14499_ (
    .A(\u_ot.LoadCtl_6_bF$buf0 ),
    .B(_6565_),
    .C(_6759_),
    .Y(_6536_)
);

DFFPOSX1 _14500_ (
    .CLK(clk_bF$buf23),
    .D(_6488_),
    .Q(\u_ot.Xcalc [0])
);

DFFPOSX1 _14501_ (
    .CLK(clk_bF$buf22),
    .D(_6489_),
    .Q(\u_ot.Xcalc [1])
);

DFFPOSX1 _14502_ (
    .CLK(clk_bF$buf21),
    .D(_6490_),
    .Q(\u_ot.Xcalc [2])
);

DFFPOSX1 _14503_ (
    .CLK(clk_bF$buf20),
    .D(_6491_),
    .Q(\u_ot.Xcalc [3])
);

DFFPOSX1 _14504_ (
    .CLK(clk_bF$buf19),
    .D(_6492_),
    .Q(\u_ot.Xcalc [4])
);

DFFPOSX1 _14505_ (
    .CLK(clk_bF$buf18),
    .D(_6493_),
    .Q(\u_ot.Xcalc [5])
);

DFFPOSX1 _14506_ (
    .CLK(clk_bF$buf17),
    .D(_6494_),
    .Q(\u_ot.Xcalc [6])
);

DFFPOSX1 _14507_ (
    .CLK(clk_bF$buf16),
    .D(_6495_),
    .Q(\u_ot.Xcalc [7])
);

DFFPOSX1 _14508_ (
    .CLK(clk_bF$buf15),
    .D(_6496_),
    .Q(\u_ot.Xcalc [8])
);

DFFPOSX1 _14509_ (
    .CLK(clk_bF$buf14),
    .D(_6497_),
    .Q(\u_ot.Xcalc [9])
);

DFFPOSX1 _14510_ (
    .CLK(clk_bF$buf13),
    .D(_6498_),
    .Q(\u_ot.Xcalc [10])
);

DFFPOSX1 _14511_ (
    .CLK(clk_bF$buf12),
    .D(_6499_),
    .Q(\u_ot.Xcalc [11])
);

DFFPOSX1 _14512_ (
    .CLK(clk_bF$buf11),
    .D(_6500_),
    .Q(\u_ot.Ycalc [0])
);

DFFPOSX1 _14513_ (
    .CLK(clk_bF$buf10),
    .D(_6501_),
    .Q(\u_ot.Ycalc [1])
);

DFFPOSX1 _14514_ (
    .CLK(clk_bF$buf9),
    .D(_6502_),
    .Q(\u_ot.Ycalc [2])
);

DFFPOSX1 _14515_ (
    .CLK(clk_bF$buf8),
    .D(_6503_),
    .Q(\u_ot.Ycalc [3])
);

DFFPOSX1 _14516_ (
    .CLK(clk_bF$buf7),
    .D(_6504_),
    .Q(\u_ot.Ycalc [4])
);

DFFPOSX1 _14517_ (
    .CLK(clk_bF$buf6),
    .D(_6505_),
    .Q(\u_ot.Ycalc [5])
);

DFFPOSX1 _14518_ (
    .CLK(clk_bF$buf5),
    .D(_6506_),
    .Q(\u_ot.Ycalc [6])
);

DFFPOSX1 _14519_ (
    .CLK(clk_bF$buf4),
    .D(_6507_),
    .Q(\u_ot.Ycalc [7])
);

DFFPOSX1 _14520_ (
    .CLK(clk_bF$buf3),
    .D(_6508_),
    .Q(\u_ot.Ycalc [8])
);

DFFPOSX1 _14521_ (
    .CLK(clk_bF$buf2),
    .D(_6509_),
    .Q(\u_ot.Ycalc [9])
);

DFFPOSX1 _14522_ (
    .CLK(clk_bF$buf1),
    .D(_6510_),
    .Q(\u_ot.Ycalc [10])
);

DFFPOSX1 _14523_ (
    .CLK(clk_bF$buf0),
    .D(_6511_),
    .Q(\u_ot.Ycalc [11])
);

DFFPOSX1 _14524_ (
    .CLK(clk_bF$buf78),
    .D(_6512_),
    .Q(\u_ot.Xin12b [10])
);

DFFPOSX1 _14525_ (
    .CLK(clk_bF$buf77),
    .D(_6513_),
    .Q(\u_ot.Xin12b [11])
);

DFFPOSX1 _14526_ (
    .CLK(clk_bF$buf76),
    .D(_6514_),
    .Q(\u_ot.Xin12b [8])
);

DFFPOSX1 _14527_ (
    .CLK(clk_bF$buf75),
    .D(_6515_),
    .Q(\u_ot.Xin12b [9])
);

DFFPOSX1 _14528_ (
    .CLK(clk_bF$buf74),
    .D(_6516_),
    .Q(\u_ot.Xin12b [6])
);

DFFPOSX1 _14529_ (
    .CLK(clk_bF$buf73),
    .D(_6517_),
    .Q(\u_ot.Xin12b [7])
);

DFFPOSX1 _14530_ (
    .CLK(clk_bF$buf72),
    .D(_6518_),
    .Q(\u_ot.Xin12b [4])
);

DFFPOSX1 _14531_ (
    .CLK(clk_bF$buf71),
    .D(_6519_),
    .Q(\u_ot.Xin12b [5])
);

DFFPOSX1 _14532_ (
    .CLK(clk_bF$buf70),
    .D(_6520_),
    .Q(\u_ot.Xin1 [0])
);

DFFPOSX1 _14533_ (
    .CLK(clk_bF$buf69),
    .D(_6521_),
    .Q(\u_ot.Xin1 [1])
);

DFFPOSX1 _14534_ (
    .CLK(clk_bF$buf68),
    .D(_6522_),
    .Q(\u_ot.Xin0 [0])
);

DFFPOSX1 _14535_ (
    .CLK(clk_bF$buf67),
    .D(_6523_),
    .Q(\u_ot.Xin0 [1])
);

DFFPOSX1 _14536_ (
    .CLK(clk_bF$buf66),
    .D(_6524_),
    .Q(\u_ot.Yin12b [10])
);

DFFPOSX1 _14537_ (
    .CLK(clk_bF$buf65),
    .D(_6525_),
    .Q(\u_ot.Yin12b [11])
);

DFFPOSX1 _14538_ (
    .CLK(clk_bF$buf64),
    .D(_6526_),
    .Q(\u_ot.Yin12b [8])
);

DFFPOSX1 _14539_ (
    .CLK(clk_bF$buf63),
    .D(_6527_),
    .Q(\u_ot.Yin12b [9])
);

DFFPOSX1 _14540_ (
    .CLK(clk_bF$buf62),
    .D(_6528_),
    .Q(\u_ot.Yin12b [6])
);

DFFPOSX1 _14541_ (
    .CLK(clk_bF$buf61),
    .D(_6529_),
    .Q(\u_ot.Yin12b [7])
);

DFFPOSX1 _14542_ (
    .CLK(clk_bF$buf60),
    .D(_6530_),
    .Q(\u_ot.Yin12b [4])
);

DFFPOSX1 _14543_ (
    .CLK(clk_bF$buf59),
    .D(_6531_),
    .Q(\u_ot.Yin12b [5])
);

DFFPOSX1 _14544_ (
    .CLK(clk_bF$buf58),
    .D(_6532_),
    .Q(\u_ot.Yin1 [0])
);

DFFPOSX1 _14545_ (
    .CLK(clk_bF$buf57),
    .D(_6533_),
    .Q(\u_ot.Yin1 [1])
);

DFFPOSX1 _14546_ (
    .CLK(clk_bF$buf56),
    .D(_6534_),
    .Q(\u_ot.Yin0 [0])
);

DFFPOSX1 _14547_ (
    .CLK(clk_bF$buf55),
    .D(_6535_),
    .Q(\u_ot.Yin0 [1])
);

DFFPOSX1 _14548_ (
    .CLK(clk_bF$buf54),
    .D(\genblk1[7].u_ce.Vld ),
    .Q(\u_ot.LoadCtl [0])
);

DFFPOSX1 _14549_ (
    .CLK(clk_bF$buf53),
    .D(\u_ot.LoadCtl [0]),
    .Q(\u_ot.LoadCtl [1])
);

DFFPOSX1 _14550_ (
    .CLK(clk_bF$buf52),
    .D(\u_ot.LoadCtl [1]),
    .Q(\u_ot.LoadCtl [2])
);

DFFPOSX1 _14551_ (
    .CLK(clk_bF$buf51),
    .D(\u_ot.LoadCtl [2]),
    .Q(\u_ot.LoadCtl [3])
);

DFFPOSX1 _14552_ (
    .CLK(clk_bF$buf50),
    .D(\u_ot.LoadCtl [3]),
    .Q(\u_ot.LoadCtl [4])
);

DFFPOSX1 _14553_ (
    .CLK(clk_bF$buf49),
    .D(\u_ot.LoadCtl [4]),
    .Q(\u_ot.LoadCtl [5])
);

DFFPOSX1 _14554_ (
    .CLK(clk_bF$buf48),
    .D(\u_ot.LoadCtl [5]),
    .Q(\u_ot.LoadCtl [6])
);

DFFPOSX1 _14555_ (
    .CLK(clk_bF$buf47),
    .D(_6536_),
    .Q(\u_ot.ISreg )
);

INVX1 _14556_ (
    .A(\u_pa.Atmp [4]),
    .Y(_6799_)
);

INVX1 _14557_ (
    .A(\u_pa.RdyCtl [2]),
    .Y(_6800_)
);

INVX1 _14558_ (
    .A(\u_pa.Atmp [6]),
    .Y(_6801_)
);

INVX1 _14559_ (
    .A(\u_pa.RdyCtl [3]),
    .Y(_6802_)
);

INVX1 _14560_ (
    .A(\u_pa.Atmp [8]),
    .Y(_6803_)
);

INVX1 _14561_ (
    .A(\u_pa.RdyCtl [4]),
    .Y(_6804_)
);

NAND2X1 _14562_ (
    .A(\u_pa.Atmp [11]),
    .B(_6804_),
    .Y(_6805_)
);

OAI21X1 _14563_ (
    .A(_6803_),
    .B(_6804_),
    .C(_6805_),
    .Y(_6806_)
);

NAND2X1 _14564_ (
    .A(_6802_),
    .B(_6806_),
    .Y(_6807_)
);

OAI21X1 _14565_ (
    .A(_6801_),
    .B(_6802_),
    .C(_6807_),
    .Y(_6808_)
);

NAND2X1 _14566_ (
    .A(_6800_),
    .B(_6808_),
    .Y(_6809_)
);

OAI21X1 _14567_ (
    .A(_6799_),
    .B(_6800_),
    .C(_6809_),
    .Y(_6810_)
);

INVX1 _14568_ (
    .A(\u_pa.Atmp [2]),
    .Y(_6811_)
);

NAND2X1 _14569_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6811_),
    .Y(_6812_)
);

OAI21X1 _14570_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6810_),
    .C(_6812_),
    .Y(_6813_)
);

NAND2X1 _14571_ (
    .A(\u_pa.Atmp [0]),
    .B(\u_pa.RdyCtl [0]),
    .Y(_6814_)
);

OAI21X1 _14572_ (
    .A(\u_pa.RdyCtl [0]),
    .B(_6813_),
    .C(_6814_),
    .Y(\a[0] [0])
);

INVX1 _14573_ (
    .A(\u_pa.Atmp [5]),
    .Y(_6815_)
);

INVX1 _14574_ (
    .A(\u_pa.Atmp [9]),
    .Y(_6816_)
);

OAI21X1 _14575_ (
    .A(_6804_),
    .B(_6816_),
    .C(_6805_),
    .Y(_6817_)
);

INVX1 _14576_ (
    .A(\u_pa.Atmp [7]),
    .Y(_6818_)
);

AOI21X1 _14577_ (
    .A(_6818_),
    .B(\u_pa.RdyCtl [3]),
    .C(\u_pa.RdyCtl [2]),
    .Y(_6819_)
);

OAI21X1 _14578_ (
    .A(\u_pa.RdyCtl [3]),
    .B(_6817_),
    .C(_6819_),
    .Y(_6820_)
);

OAI21X1 _14579_ (
    .A(_6800_),
    .B(_6815_),
    .C(_6820_),
    .Y(_6821_)
);

INVX1 _14580_ (
    .A(\u_pa.Atmp [3]),
    .Y(_6822_)
);

NAND2X1 _14581_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6822_),
    .Y(_6823_)
);

OAI21X1 _14582_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6821_),
    .C(_6823_),
    .Y(_6824_)
);

NAND2X1 _14583_ (
    .A(\u_pa.RdyCtl [0]),
    .B(\u_pa.Atmp [1]),
    .Y(_6825_)
);

OAI21X1 _14584_ (
    .A(\u_pa.RdyCtl [0]),
    .B(_6824_),
    .C(_6825_),
    .Y(\a[0] [1])
);

INVX1 _14585_ (
    .A(\u_pa.RdyCtl [5]),
    .Y(_6826_)
);

NAND2X1 _14586_ (
    .A(\u_pa.acc_reg [18]),
    .B(\u_pa.acc_reg [19]),
    .Y(_6827_)
);

INVX1 _14587_ (
    .A(\u_pa.acc_reg [18]),
    .Y(_6828_)
);

INVX1 _14588_ (
    .A(\u_pa.acc_reg [19]),
    .Y(_6829_)
);

NAND2X1 _14589_ (
    .A(_6828_),
    .B(_6829_),
    .Y(_6830_)
);

NAND2X1 _14590_ (
    .A(_6827_),
    .B(_6830_),
    .Y(_6831_)
);

NAND2X1 _14591_ (
    .A(\genblk1[0].u_ce.ISin ),
    .B(_6826_),
    .Y(_6832_)
);

OAI21X1 _14592_ (
    .A(_6826_),
    .B(_6831_),
    .C(_6832_),
    .Y(_6798_)
);

INVX8 _14593_ (
    .A(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .Y(_6833_)
);

INVX2 _14594_ (
    .A(En_bF$buf4),
    .Y(_6834_)
);

NOR2X1 _14595_ (
    .A(_6833__bF$buf4),
    .B(_6834_),
    .Y(_6760_)
);

AND2X2 _14596_ (
    .A(\u_pa.RdyCtl [0]),
    .B(En_bF$buf3),
    .Y(_6761_)
);

AND2X2 _14597_ (
    .A(\u_pa.RdyCtl [1]),
    .B(En_bF$buf2),
    .Y(_6762_)
);

NOR2X1 _14598_ (
    .A(_6800_),
    .B(_6834_),
    .Y(_6763_)
);

NOR2X1 _14599_ (
    .A(_6802_),
    .B(_6834_),
    .Y(_6764_)
);

NAND2X1 _14600_ (
    .A(En_bF$buf1),
    .B(_6804_),
    .Y(_6765_)
);

NOR2X1 _14601_ (
    .A(_6826_),
    .B(_6834_),
    .Y(_6766_)
);

INVX1 _14602_ (
    .A(\u_pa.acc_reg [0]),
    .Y(_6835_)
);

NAND2X1 _14603_ (
    .A(FCW[0]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .Y(_6836_)
);

OAI21X1 _14604_ (
    .A(_6835_),
    .B(_6836_),
    .C(En_bF$buf0),
    .Y(_6837_)
);

AOI21X1 _14605_ (
    .A(_6835_),
    .B(_6836_),
    .C(_6837_),
    .Y(_6767_)
);

NAND2X1 _14606_ (
    .A(FCW[0]),
    .B(\u_pa.acc_reg [0]),
    .Y(_6838_)
);

NAND2X1 _14607_ (
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6839_)
);

INVX1 _14608_ (
    .A(_6839_),
    .Y(_6840_)
);

NOR2X1 _14609_ (
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6841_)
);

OAI21X1 _14610_ (
    .A(_6841_),
    .B(_6840_),
    .C(_6838_),
    .Y(_6842_)
);

OR2X2 _14611_ (
    .A(_6840_),
    .B(_6841_),
    .Y(_6843_)
);

NOR2X1 _14612_ (
    .A(_6838_),
    .B(_6843_),
    .Y(_6844_)
);

INVX1 _14613_ (
    .A(_6844_),
    .Y(_6845_)
);

NAND2X1 _14614_ (
    .A(_6842_),
    .B(_6845_),
    .Y(_6846_)
);

OAI21X1 _14615_ (
    .A(\u_pa.acc_reg [1]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf4),
    .Y(_6847_)
);

AOI21X1 _14616_ (
    .A(_6846_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(_6847_),
    .Y(_6768_)
);

OAI21X1 _14617_ (
    .A(_6838_),
    .B(_6841_),
    .C(_6839_),
    .Y(_6848_)
);

AND2X2 _14618_ (
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6849_)
);

NOR2X1 _14619_ (
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6850_)
);

NOR2X1 _14620_ (
    .A(_6850_),
    .B(_6849_),
    .Y(_6851_)
);

AND2X2 _14621_ (
    .A(_6851_),
    .B(_6848_),
    .Y(_6852_)
);

NOR2X1 _14622_ (
    .A(_6833__bF$buf3),
    .B(_6852_),
    .Y(_6853_)
);

OAI21X1 _14623_ (
    .A(_6848_),
    .B(_6851_),
    .C(_6853_),
    .Y(_6854_)
);

NAND2X1 _14624_ (
    .A(\u_pa.acc_reg [2]),
    .B(_6833__bF$buf2),
    .Y(_6855_)
);

AOI21X1 _14625_ (
    .A(_6854_),
    .B(_6855_),
    .C(_6834_),
    .Y(_6769_)
);

OAI21X1 _14626_ (
    .A(\u_pa.acc_reg [3]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf3),
    .Y(_6856_)
);

AND2X2 _14627_ (
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6857_)
);

NOR2X1 _14628_ (
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6858_)
);

NOR2X1 _14629_ (
    .A(_6858_),
    .B(_6857_),
    .Y(_6859_)
);

OAI21X1 _14630_ (
    .A(_6849_),
    .B(_6852_),
    .C(_6859_),
    .Y(_6860_)
);

NOR2X1 _14631_ (
    .A(_6849_),
    .B(_6852_),
    .Y(_6861_)
);

OAI21X1 _14632_ (
    .A(_6857_),
    .B(_6858_),
    .C(_6861_),
    .Y(_6862_)
);

NAND2X1 _14633_ (
    .A(_6860_),
    .B(_6862_),
    .Y(_6863_)
);

AOI21X1 _14634_ (
    .A(_6863_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(_6856_),
    .Y(_6770_)
);

NAND3X1 _14635_ (
    .A(_6848_),
    .B(_6851_),
    .C(_6859_),
    .Y(_6864_)
);

INVX1 _14636_ (
    .A(_6858_),
    .Y(_6865_)
);

AOI21X1 _14637_ (
    .A(_6865_),
    .B(_6849_),
    .C(_6857_),
    .Y(_6866_)
);

AND2X2 _14638_ (
    .A(_6864_),
    .B(_6866_),
    .Y(_6867_)
);

AND2X2 _14639_ (
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6868_)
);

NOR2X1 _14640_ (
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6869_)
);

OAI21X1 _14641_ (
    .A(_6868_),
    .B(_6869_),
    .C(_6867_),
    .Y(_6870_)
);

NAND2X1 _14642_ (
    .A(_6866_),
    .B(_6864_),
    .Y(_6871_)
);

NOR2X1 _14643_ (
    .A(_6869_),
    .B(_6868_),
    .Y(_6872_)
);

NAND2X1 _14644_ (
    .A(_6872_),
    .B(_6871_),
    .Y(_6873_)
);

NAND2X1 _14645_ (
    .A(_6873_),
    .B(_6870_),
    .Y(_6874_)
);

OAI21X1 _14646_ (
    .A(\u_pa.acc_reg [4]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf2),
    .Y(_6875_)
);

AOI21X1 _14647_ (
    .A(_6874_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(_6875_),
    .Y(_6771_)
);

AOI21X1 _14648_ (
    .A(_6871_),
    .B(_6872_),
    .C(_6868_),
    .Y(_6876_)
);

AND2X2 _14649_ (
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6877_)
);

NOR2X1 _14650_ (
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6878_)
);

NOR2X1 _14651_ (
    .A(_6878_),
    .B(_6877_),
    .Y(_6879_)
);

NAND2X1 _14652_ (
    .A(_6879_),
    .B(_6876_),
    .Y(_6880_)
);

NOR2X1 _14653_ (
    .A(_6879_),
    .B(_6876_),
    .Y(_6881_)
);

NOR2X1 _14654_ (
    .A(_6833__bF$buf1),
    .B(_6881_),
    .Y(_6882_)
);

OAI21X1 _14655_ (
    .A(\u_pa.acc_reg [5]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(En_bF$buf1),
    .Y(_6883_)
);

AOI21X1 _14656_ (
    .A(_6882_),
    .B(_6880_),
    .C(_6883_),
    .Y(_6772_)
);

INVX1 _14657_ (
    .A(_6868_),
    .Y(_6884_)
);

INVX1 _14658_ (
    .A(_6877_),
    .Y(_6885_)
);

OAI21X1 _14659_ (
    .A(_6878_),
    .B(_6884_),
    .C(_6885_),
    .Y(_6886_)
);

AND2X2 _14660_ (
    .A(_6872_),
    .B(_6879_),
    .Y(_6887_)
);

AOI21X1 _14661_ (
    .A(_6871_),
    .B(_6887_),
    .C(_6886_),
    .Y(_6888_)
);

NAND2X1 _14662_ (
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6889_)
);

OR2X2 _14663_ (
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6890_)
);

NAND2X1 _14664_ (
    .A(_6889_),
    .B(_6890_),
    .Y(_6891_)
);

OR2X2 _14665_ (
    .A(_6888_),
    .B(_6891_),
    .Y(_6892_)
);

INVX1 _14666_ (
    .A(_6889_),
    .Y(_6893_)
);

INVX1 _14667_ (
    .A(_6890_),
    .Y(_6894_)
);

OAI21X1 _14668_ (
    .A(_6893_),
    .B(_6894_),
    .C(_6888_),
    .Y(_6895_)
);

NAND2X1 _14669_ (
    .A(_6895_),
    .B(_6892_),
    .Y(_6896_)
);

OAI21X1 _14670_ (
    .A(\u_pa.acc_reg [6]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf0),
    .Y(_6897_)
);

AOI21X1 _14671_ (
    .A(_6896_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(_6897_),
    .Y(_6773_)
);

OAI21X1 _14672_ (
    .A(_6894_),
    .B(_6888_),
    .C(_6889_),
    .Y(_6898_)
);

NAND2X1 _14673_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6899_)
);

OR2X2 _14674_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6900_)
);

NAND2X1 _14675_ (
    .A(_6899_),
    .B(_6900_),
    .Y(_6901_)
);

OR2X2 _14676_ (
    .A(_6898_),
    .B(_6901_),
    .Y(_6902_)
);

AOI21X1 _14677_ (
    .A(_6898_),
    .B(_6901_),
    .C(_6833__bF$buf0),
    .Y(_6903_)
);

OAI21X1 _14678_ (
    .A(\u_pa.acc_reg [7]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf4),
    .Y(_6904_)
);

AOI21X1 _14679_ (
    .A(_6902_),
    .B(_6903_),
    .C(_6904_),
    .Y(_6774_)
);

NAND2X1 _14680_ (
    .A(_6872_),
    .B(_6879_),
    .Y(_6905_)
);

AND2X2 _14681_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6906_)
);

NOR2X1 _14682_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6907_)
);

NOR2X1 _14683_ (
    .A(_6907_),
    .B(_6906_),
    .Y(_6908_)
);

NAND3X1 _14684_ (
    .A(_6889_),
    .B(_6890_),
    .C(_6908_),
    .Y(_6909_)
);

NOR2X1 _14685_ (
    .A(_6905_),
    .B(_6909_),
    .Y(_6910_)
);

INVX1 _14686_ (
    .A(_6878_),
    .Y(_6911_)
);

AOI21X1 _14687_ (
    .A(_6911_),
    .B(_6868_),
    .C(_6877_),
    .Y(_6912_)
);

OAI21X1 _14688_ (
    .A(_6889_),
    .B(_6907_),
    .C(_6899_),
    .Y(_6913_)
);

INVX1 _14689_ (
    .A(_6913_),
    .Y(_6914_)
);

OAI21X1 _14690_ (
    .A(_6912_),
    .B(_6909_),
    .C(_6914_),
    .Y(_6915_)
);

AOI21X1 _14691_ (
    .A(_6910_),
    .B(_6871_),
    .C(_6915_),
    .Y(_6916_)
);

NAND2X1 _14692_ (
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6917_)
);

OR2X2 _14693_ (
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6918_)
);

NAND2X1 _14694_ (
    .A(_6917_),
    .B(_6918_),
    .Y(_6919_)
);

OR2X2 _14695_ (
    .A(_6916_),
    .B(_6919_),
    .Y(_6920_)
);

NAND2X1 _14696_ (
    .A(_6919_),
    .B(_6916_),
    .Y(_6921_)
);

NAND2X1 _14697_ (
    .A(_6921_),
    .B(_6920_),
    .Y(_6922_)
);

OAI21X1 _14698_ (
    .A(\u_pa.acc_reg [8]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf3),
    .Y(_6923_)
);

AOI21X1 _14699_ (
    .A(_6922_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(_6923_),
    .Y(_6775_)
);

OAI21X1 _14700_ (
    .A(_6919_),
    .B(_6916_),
    .C(_6917_),
    .Y(_6924_)
);

NAND2X1 _14701_ (
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6925_)
);

INVX1 _14702_ (
    .A(FCW[9]),
    .Y(_6926_)
);

INVX1 _14703_ (
    .A(\u_pa.acc_reg [9]),
    .Y(_6927_)
);

NAND2X1 _14704_ (
    .A(_6926_),
    .B(_6927_),
    .Y(_6928_)
);

NAND2X1 _14705_ (
    .A(_6925_),
    .B(_6928_),
    .Y(_6929_)
);

NAND2X1 _14706_ (
    .A(_6929_),
    .B(_6924_),
    .Y(_6930_)
);

NOR2X1 _14707_ (
    .A(_6929_),
    .B(_6924_),
    .Y(_6931_)
);

NOR2X1 _14708_ (
    .A(_6833__bF$buf4),
    .B(_6931_),
    .Y(_6932_)
);

OAI21X1 _14709_ (
    .A(\u_pa.acc_reg [9]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf2),
    .Y(_6933_)
);

AOI21X1 _14710_ (
    .A(_6932_),
    .B(_6930_),
    .C(_6933_),
    .Y(_6776_)
);

NOR2X1 _14711_ (
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6934_)
);

OAI21X1 _14712_ (
    .A(_6917_),
    .B(_6934_),
    .C(_6925_),
    .Y(_6935_)
);

INVX1 _14713_ (
    .A(_6935_),
    .Y(_6936_)
);

OR2X2 _14714_ (
    .A(_6929_),
    .B(_6919_),
    .Y(_6937_)
);

OAI21X1 _14715_ (
    .A(_6937_),
    .B(_6916_),
    .C(_6936_),
    .Y(_6938_)
);

AND2X2 _14716_ (
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6939_)
);

NOR2X1 _14717_ (
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6940_)
);

NOR2X1 _14718_ (
    .A(_6940_),
    .B(_6939_),
    .Y(_6941_)
);

NAND2X1 _14719_ (
    .A(_6941_),
    .B(_6938_),
    .Y(_6942_)
);

OR2X2 _14720_ (
    .A(_6938_),
    .B(_6941_),
    .Y(_6943_)
);

NAND2X1 _14721_ (
    .A(_6942_),
    .B(_6943_),
    .Y(_6944_)
);

OAI21X1 _14722_ (
    .A(\u_pa.acc_reg [10]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf1),
    .Y(_6945_)
);

AOI21X1 _14723_ (
    .A(_6944_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(_6945_),
    .Y(_6777_)
);

NAND2X1 _14724_ (
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6946_)
);

NAND2X1 _14725_ (
    .A(_6946_),
    .B(_6942_),
    .Y(_6947_)
);

AND2X2 _14726_ (
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6948_)
);

NOR2X1 _14727_ (
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6949_)
);

NOR2X1 _14728_ (
    .A(_6949_),
    .B(_6948_),
    .Y(_6950_)
);

INVX1 _14729_ (
    .A(_6950_),
    .Y(_6951_)
);

OR2X2 _14730_ (
    .A(_6947_),
    .B(_6951_),
    .Y(_6952_)
);

AOI21X1 _14731_ (
    .A(_6947_),
    .B(_6951_),
    .C(_6833__bF$buf3),
    .Y(_6953_)
);

OAI21X1 _14732_ (
    .A(\u_pa.acc_reg [11]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf0),
    .Y(_6954_)
);

AOI21X1 _14733_ (
    .A(_6952_),
    .B(_6953_),
    .C(_6954_),
    .Y(_6778_)
);

NAND2X1 _14734_ (
    .A(\u_pa.acc_reg [12]),
    .B(_6833__bF$buf2),
    .Y(_6955_)
);

NOR2X1 _14735_ (
    .A(_6919_),
    .B(_6929_),
    .Y(_6956_)
);

NAND3X1 _14736_ (
    .A(_6941_),
    .B(_6950_),
    .C(_6956_),
    .Y(_6957_)
);

NAND3X1 _14737_ (
    .A(_6935_),
    .B(_6941_),
    .C(_6950_),
    .Y(_6958_)
);

INVX1 _14738_ (
    .A(_6949_),
    .Y(_6959_)
);

AOI21X1 _14739_ (
    .A(_6959_),
    .B(_6939_),
    .C(_6948_),
    .Y(_6960_)
);

AND2X2 _14740_ (
    .A(_6958_),
    .B(_6960_),
    .Y(_6961_)
);

OAI21X1 _14741_ (
    .A(_6957_),
    .B(_6916_),
    .C(_6961_),
    .Y(_6962_)
);

NAND2X1 _14742_ (
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6963_)
);

OR2X2 _14743_ (
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6964_)
);

NAND2X1 _14744_ (
    .A(_6963_),
    .B(_6964_),
    .Y(_6965_)
);

NOR2X1 _14745_ (
    .A(_6965_),
    .B(_6962_),
    .Y(_6966_)
);

AND2X2 _14746_ (
    .A(_6962_),
    .B(_6965_),
    .Y(_6967_)
);

OAI21X1 _14747_ (
    .A(_6966_),
    .B(_6967_),
    .C(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .Y(_6968_)
);

AOI21X1 _14748_ (
    .A(_6968_),
    .B(_6955_),
    .C(_6834_),
    .Y(_6779_)
);

INVX1 _14749_ (
    .A(_6962_),
    .Y(_6969_)
);

OAI21X1 _14750_ (
    .A(_6965_),
    .B(_6969_),
    .C(_6963_),
    .Y(_6970_)
);

NAND2X1 _14751_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6971_)
);

OR2X2 _14752_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6972_)
);

NAND2X1 _14753_ (
    .A(_6971_),
    .B(_6972_),
    .Y(_6973_)
);

OR2X2 _14754_ (
    .A(_6970_),
    .B(_6973_),
    .Y(_6974_)
);

AOI21X1 _14755_ (
    .A(_6970_),
    .B(_6973_),
    .C(_6833__bF$buf1),
    .Y(_6975_)
);

OAI21X1 _14756_ (
    .A(\u_pa.acc_reg [13]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(En_bF$buf4),
    .Y(_6976_)
);

AOI21X1 _14757_ (
    .A(_6974_),
    .B(_6975_),
    .C(_6976_),
    .Y(_6780_)
);

NOR2X1 _14758_ (
    .A(_6965_),
    .B(_6973_),
    .Y(_6977_)
);

NOR2X1 _14759_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6978_)
);

OAI21X1 _14760_ (
    .A(_6963_),
    .B(_6978_),
    .C(_6971_),
    .Y(_6979_)
);

AOI21X1 _14761_ (
    .A(_6962_),
    .B(_6977_),
    .C(_6979_),
    .Y(_6980_)
);

AND2X2 _14762_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6981_)
);

NOR2X1 _14763_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6982_)
);

OR2X2 _14764_ (
    .A(_6981_),
    .B(_6982_),
    .Y(_6983_)
);

OR2X2 _14765_ (
    .A(_6980_),
    .B(_6983_),
    .Y(_6984_)
);

OAI21X1 _14766_ (
    .A(_6981_),
    .B(_6982_),
    .C(_6980_),
    .Y(_6985_)
);

NAND2X1 _14767_ (
    .A(_6985_),
    .B(_6984_),
    .Y(_6986_)
);

OAI21X1 _14768_ (
    .A(\u_pa.acc_reg [14]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf3),
    .Y(_6987_)
);

AOI21X1 _14769_ (
    .A(_6986_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(_6987_),
    .Y(_6781_)
);

NAND2X1 _14770_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6988_)
);

NAND2X1 _14771_ (
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6989_)
);

INVX1 _14772_ (
    .A(_6989_),
    .Y(_6990_)
);

NOR2X1 _14773_ (
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6991_)
);

NOR2X1 _14774_ (
    .A(_6991_),
    .B(_6990_),
    .Y(_6992_)
);

NAND3X1 _14775_ (
    .A(_6988_),
    .B(_6992_),
    .C(_6984_),
    .Y(_6993_)
);

OAI21X1 _14776_ (
    .A(_6983_),
    .B(_6980_),
    .C(_6988_),
    .Y(_6994_)
);

INVX1 _14777_ (
    .A(_6991_),
    .Y(_6995_)
);

NAND2X1 _14778_ (
    .A(_6989_),
    .B(_6995_),
    .Y(_6996_)
);

AOI21X1 _14779_ (
    .A(_6994_),
    .B(_6996_),
    .C(_6833__bF$buf0),
    .Y(_6997_)
);

OAI21X1 _14780_ (
    .A(\u_pa.acc_reg [15]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(En_bF$buf2),
    .Y(_6998_)
);

AOI21X1 _14781_ (
    .A(_6993_),
    .B(_6997_),
    .C(_6998_),
    .Y(_6782_)
);

NOR2X1 _14782_ (
    .A(_6982_),
    .B(_6981_),
    .Y(_6999_)
);

NAND3X1 _14783_ (
    .A(_6999_),
    .B(_6992_),
    .C(_6977_),
    .Y(_7000_)
);

OR2X2 _14784_ (
    .A(_6957_),
    .B(_7000_),
    .Y(_7001_)
);

NAND2X1 _14785_ (
    .A(_6960_),
    .B(_6958_),
    .Y(_7002_)
);

NOR2X1 _14786_ (
    .A(_6983_),
    .B(_6996_),
    .Y(_7003_)
);

AND2X2 _14787_ (
    .A(_7003_),
    .B(_6977_),
    .Y(_7004_)
);

NAND3X1 _14788_ (
    .A(_6979_),
    .B(_6999_),
    .C(_6992_),
    .Y(_7005_)
);

AOI21X1 _14789_ (
    .A(_6995_),
    .B(_6981_),
    .C(_6990_),
    .Y(_7006_)
);

NAND2X1 _14790_ (
    .A(_7006_),
    .B(_7005_),
    .Y(_7007_)
);

AOI21X1 _14791_ (
    .A(_7004_),
    .B(_7002_),
    .C(_7007_),
    .Y(_7008_)
);

OAI21X1 _14792_ (
    .A(_6916_),
    .B(_7001_),
    .C(_7008_),
    .Y(_7009_)
);

AND2X2 _14793_ (
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_7010_)
);

NOR2X1 _14794_ (
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_7011_)
);

NOR2X1 _14795_ (
    .A(_7011_),
    .B(_7010_),
    .Y(_7012_)
);

NAND2X1 _14796_ (
    .A(_7012_),
    .B(_7009_),
    .Y(_7013_)
);

NOR2X1 _14797_ (
    .A(_6901_),
    .B(_6891_),
    .Y(_7014_)
);

NAND2X1 _14798_ (
    .A(_7014_),
    .B(_6887_),
    .Y(_7015_)
);

AOI21X1 _14799_ (
    .A(_7014_),
    .B(_6886_),
    .C(_6913_),
    .Y(_7016_)
);

OAI21X1 _14800_ (
    .A(_7015_),
    .B(_6867_),
    .C(_7016_),
    .Y(_7017_)
);

NOR2X1 _14801_ (
    .A(_6957_),
    .B(_7000_),
    .Y(_7018_)
);

AND2X2 _14802_ (
    .A(_7005_),
    .B(_7006_),
    .Y(_7019_)
);

OAI21X1 _14803_ (
    .A(_7000_),
    .B(_6961_),
    .C(_7019_),
    .Y(_7020_)
);

AOI21X1 _14804_ (
    .A(_7017_),
    .B(_7018_),
    .C(_7020_),
    .Y(_7021_)
);

OAI21X1 _14805_ (
    .A(_7010_),
    .B(_7011_),
    .C(_7021_),
    .Y(_7022_)
);

NAND2X1 _14806_ (
    .A(_7022_),
    .B(_7013_),
    .Y(_7023_)
);

OAI21X1 _14807_ (
    .A(\u_pa.acc_reg [16]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .C(En_bF$buf1),
    .Y(_7024_)
);

AOI21X1 _14808_ (
    .A(_7023_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .C(_7024_),
    .Y(_6783_)
);

AOI21X1 _14809_ (
    .A(_7009_),
    .B(_7012_),
    .C(_7010_),
    .Y(_7025_)
);

AND2X2 _14810_ (
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_7026_)
);

NOR2X1 _14811_ (
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_7027_)
);

NOR2X1 _14812_ (
    .A(_7027_),
    .B(_7026_),
    .Y(_7028_)
);

OR2X2 _14813_ (
    .A(_7025_),
    .B(_7028_),
    .Y(_7029_)
);

AOI21X1 _14814_ (
    .A(_7025_),
    .B(_7028_),
    .C(_6833__bF$buf4),
    .Y(_7030_)
);

OAI21X1 _14815_ (
    .A(\u_pa.acc_reg [17]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .C(En_bF$buf0),
    .Y(_7031_)
);

AOI21X1 _14816_ (
    .A(_7029_),
    .B(_7030_),
    .C(_7031_),
    .Y(_6784_)
);

NAND2X1 _14817_ (
    .A(_7012_),
    .B(_7028_),
    .Y(_7032_)
);

AOI21X1 _14818_ (
    .A(_7028_),
    .B(_7010_),
    .C(_7026_),
    .Y(_7033_)
);

OAI21X1 _14819_ (
    .A(_7032_),
    .B(_7021_),
    .C(_7033_),
    .Y(_7034_)
);

INVX1 _14820_ (
    .A(FCW[18]),
    .Y(_7035_)
);

NOR2X1 _14821_ (
    .A(_6828_),
    .B(_7035_),
    .Y(_7036_)
);

NOR2X1 _14822_ (
    .A(\u_pa.acc_reg [18]),
    .B(FCW[18]),
    .Y(_7037_)
);

NOR2X1 _14823_ (
    .A(_7037_),
    .B(_7036_),
    .Y(_7038_)
);

NAND2X1 _14824_ (
    .A(_7038_),
    .B(_7034_),
    .Y(_7039_)
);

INVX1 _14825_ (
    .A(_7032_),
    .Y(_7040_)
);

INVX1 _14826_ (
    .A(_7033_),
    .Y(_7041_)
);

AOI21X1 _14827_ (
    .A(_7009_),
    .B(_7040_),
    .C(_7041_),
    .Y(_7042_)
);

OAI21X1 _14828_ (
    .A(_7036_),
    .B(_7037_),
    .C(_7042_),
    .Y(_7043_)
);

NAND2X1 _14829_ (
    .A(_7039_),
    .B(_7043_),
    .Y(_7044_)
);

OAI21X1 _14830_ (
    .A(\u_pa.acc_reg [18]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .C(En_bF$buf4),
    .Y(_7045_)
);

AOI21X1 _14831_ (
    .A(_7044_),
    .B(\genblk1[0].u_ce.Rdy_bF$buf2 ),
    .C(_7045_),
    .Y(_6785_)
);

INVX1 _14832_ (
    .A(_6760_),
    .Y(_7046_)
);

NAND2X1 _14833_ (
    .A(\u_pa.acc_reg [19]),
    .B(En_bF$buf3),
    .Y(_7047_)
);

INVX1 _14834_ (
    .A(_7036_),
    .Y(_7048_)
);

OAI21X1 _14835_ (
    .A(_7037_),
    .B(_7042_),
    .C(_7048_),
    .Y(_7049_)
);

NAND2X1 _14836_ (
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_7050_)
);

OR2X2 _14837_ (
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_7051_)
);

NAND2X1 _14838_ (
    .A(_7050_),
    .B(_7051_),
    .Y(_7052_)
);

NAND2X1 _14839_ (
    .A(_7052_),
    .B(_7049_),
    .Y(_7053_)
);

AOI21X1 _14840_ (
    .A(_7034_),
    .B(_7038_),
    .C(_7036_),
    .Y(_7054_)
);

INVX1 _14841_ (
    .A(_7052_),
    .Y(_7055_)
);

AOI21X1 _14842_ (
    .A(_7054_),
    .B(_7055_),
    .C(_6833__bF$buf3),
    .Y(_7056_)
);

AOI22X1 _14843_ (
    .A(_7046_),
    .B(_7047_),
    .C(_7056_),
    .D(_7053_),
    .Y(_6786_)
);

NOR2X1 _14844_ (
    .A(\u_pa.Atmp [0]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf1 ),
    .Y(_7057_)
);

OAI21X1 _14845_ (
    .A(\u_pa.acc_reg [8]),
    .B(_6833__bF$buf2),
    .C(En_bF$buf2),
    .Y(_7058_)
);

NOR2X1 _14846_ (
    .A(_7057_),
    .B(_7058_),
    .Y(_6787_)
);

NOR2X1 _14847_ (
    .A(\u_pa.Atmp [1]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf0 ),
    .Y(_7059_)
);

OAI21X1 _14848_ (
    .A(\u_pa.acc_reg [9]),
    .B(_6833__bF$buf1),
    .C(En_bF$buf1),
    .Y(_7060_)
);

NOR2X1 _14849_ (
    .A(_7059_),
    .B(_7060_),
    .Y(_6788_)
);

OAI21X1 _14850_ (
    .A(\u_pa.acc_reg [10]),
    .B(_6833__bF$buf0),
    .C(En_bF$buf0),
    .Y(_7061_)
);

AOI21X1 _14851_ (
    .A(_6811_),
    .B(_6833__bF$buf4),
    .C(_7061_),
    .Y(_6789_)
);

OAI21X1 _14852_ (
    .A(\u_pa.acc_reg [11]),
    .B(_6833__bF$buf3),
    .C(En_bF$buf4),
    .Y(_7062_)
);

AOI21X1 _14853_ (
    .A(_6822_),
    .B(_6833__bF$buf2),
    .C(_7062_),
    .Y(_6790_)
);

OAI21X1 _14854_ (
    .A(\u_pa.acc_reg [12]),
    .B(_6833__bF$buf1),
    .C(En_bF$buf3),
    .Y(_7063_)
);

AOI21X1 _14855_ (
    .A(_6799_),
    .B(_6833__bF$buf0),
    .C(_7063_),
    .Y(_6791_)
);

OAI21X1 _14856_ (
    .A(\u_pa.acc_reg [13]),
    .B(_6833__bF$buf4),
    .C(En_bF$buf2),
    .Y(_7064_)
);

AOI21X1 _14857_ (
    .A(_6815_),
    .B(_6833__bF$buf3),
    .C(_7064_),
    .Y(_6792_)
);

OAI21X1 _14858_ (
    .A(\u_pa.acc_reg [14]),
    .B(_6833__bF$buf2),
    .C(En_bF$buf1),
    .Y(_7065_)
);

AOI21X1 _14859_ (
    .A(_6801_),
    .B(_6833__bF$buf1),
    .C(_7065_),
    .Y(_6793_)
);

OAI21X1 _14860_ (
    .A(\u_pa.acc_reg [15]),
    .B(_6833__bF$buf0),
    .C(En_bF$buf0),
    .Y(_7066_)
);

AOI21X1 _14861_ (
    .A(_6818_),
    .B(_6833__bF$buf4),
    .C(_7066_),
    .Y(_6794_)
);

OAI21X1 _14862_ (
    .A(\u_pa.acc_reg [16]),
    .B(_6833__bF$buf3),
    .C(En_bF$buf4),
    .Y(_7067_)
);

AOI21X1 _14863_ (
    .A(_6803_),
    .B(_6833__bF$buf2),
    .C(_7067_),
    .Y(_6795_)
);

OAI21X1 _14864_ (
    .A(\u_pa.acc_reg [17]),
    .B(_6833__bF$buf1),
    .C(En_bF$buf3),
    .Y(_7068_)
);

AOI21X1 _14865_ (
    .A(_6816_),
    .B(_6833__bF$buf0),
    .C(_7068_),
    .Y(_6796_)
);

NOR2X1 _14866_ (
    .A(\u_pa.Atmp [11]),
    .B(\genblk1[0].u_ce.Rdy_bF$buf4 ),
    .Y(_7069_)
);

OAI21X1 _14867_ (
    .A(\u_pa.acc_reg [18]),
    .B(_6833__bF$buf4),
    .C(En_bF$buf2),
    .Y(_7070_)
);

NOR2X1 _14868_ (
    .A(_7069_),
    .B(_7070_),
    .Y(_6797_)
);

DFFPOSX1 _14869_ (
    .CLK(clk_bF$buf46),
    .D(_6760_),
    .Q(\u_pa.RdyCtl [0])
);

DFFPOSX1 _14870_ (
    .CLK(clk_bF$buf45),
    .D(_6761_),
    .Q(\u_pa.RdyCtl [1])
);

DFFPOSX1 _14871_ (
    .CLK(clk_bF$buf44),
    .D(_6762_),
    .Q(\u_pa.RdyCtl [2])
);

DFFPOSX1 _14872_ (
    .CLK(clk_bF$buf43),
    .D(_6763_),
    .Q(\u_pa.RdyCtl [3])
);

DFFPOSX1 _14873_ (
    .CLK(clk_bF$buf42),
    .D(_6764_),
    .Q(\u_pa.RdyCtl [4])
);

DFFPOSX1 _14874_ (
    .CLK(clk_bF$buf41),
    .D(_6765_),
    .Q(\u_pa.RdyCtl [5])
);

DFFPOSX1 _14875_ (
    .CLK(clk_bF$buf40),
    .D(_6766_),
    .Q(\genblk1[0].u_ce.Rdy )
);

DFFPOSX1 _14876_ (
    .CLK(clk_bF$buf39),
    .D(_6767_),
    .Q(\u_pa.acc_reg [0])
);

DFFPOSX1 _14877_ (
    .CLK(clk_bF$buf38),
    .D(_6768_),
    .Q(\u_pa.acc_reg [1])
);

DFFPOSX1 _14878_ (
    .CLK(clk_bF$buf37),
    .D(_6769_),
    .Q(\u_pa.acc_reg [2])
);

DFFPOSX1 _14879_ (
    .CLK(clk_bF$buf36),
    .D(_6770_),
    .Q(\u_pa.acc_reg [3])
);

DFFPOSX1 _14880_ (
    .CLK(clk_bF$buf35),
    .D(_6771_),
    .Q(\u_pa.acc_reg [4])
);

DFFPOSX1 _14881_ (
    .CLK(clk_bF$buf34),
    .D(_6772_),
    .Q(\u_pa.acc_reg [5])
);

DFFPOSX1 _14882_ (
    .CLK(clk_bF$buf33),
    .D(_6773_),
    .Q(\u_pa.acc_reg [6])
);

DFFPOSX1 _14883_ (
    .CLK(clk_bF$buf32),
    .D(_6774_),
    .Q(\u_pa.acc_reg [7])
);

DFFPOSX1 _14884_ (
    .CLK(clk_bF$buf31),
    .D(_6775_),
    .Q(\u_pa.acc_reg [8])
);

DFFPOSX1 _14885_ (
    .CLK(clk_bF$buf30),
    .D(_6776_),
    .Q(\u_pa.acc_reg [9])
);

DFFPOSX1 _14886_ (
    .CLK(clk_bF$buf29),
    .D(_6777_),
    .Q(\u_pa.acc_reg [10])
);

DFFPOSX1 _14887_ (
    .CLK(clk_bF$buf28),
    .D(_6778_),
    .Q(\u_pa.acc_reg [11])
);

DFFPOSX1 _14888_ (
    .CLK(clk_bF$buf27),
    .D(_6779_),
    .Q(\u_pa.acc_reg [12])
);

DFFPOSX1 _14889_ (
    .CLK(clk_bF$buf26),
    .D(_6780_),
    .Q(\u_pa.acc_reg [13])
);

DFFPOSX1 _14890_ (
    .CLK(clk_bF$buf25),
    .D(_6781_),
    .Q(\u_pa.acc_reg [14])
);

DFFPOSX1 _14891_ (
    .CLK(clk_bF$buf24),
    .D(_6782_),
    .Q(\u_pa.acc_reg [15])
);

DFFPOSX1 _14892_ (
    .CLK(clk_bF$buf23),
    .D(_6783_),
    .Q(\u_pa.acc_reg [16])
);

DFFPOSX1 _14893_ (
    .CLK(clk_bF$buf22),
    .D(_6784_),
    .Q(\u_pa.acc_reg [17])
);

DFFPOSX1 _14894_ (
    .CLK(clk_bF$buf21),
    .D(_6785_),
    .Q(\u_pa.acc_reg [18])
);

DFFPOSX1 _14895_ (
    .CLK(clk_bF$buf20),
    .D(_6786_),
    .Q(\u_pa.acc_reg [19])
);

DFFPOSX1 _14896_ (
    .CLK(clk_bF$buf19),
    .D(_6787_),
    .Q(\u_pa.Atmp [0])
);

DFFPOSX1 _14897_ (
    .CLK(clk_bF$buf18),
    .D(_6788_),
    .Q(\u_pa.Atmp [1])
);

DFFPOSX1 _14898_ (
    .CLK(clk_bF$buf17),
    .D(_6789_),
    .Q(\u_pa.Atmp [2])
);

DFFPOSX1 _14899_ (
    .CLK(clk_bF$buf16),
    .D(_6790_),
    .Q(\u_pa.Atmp [3])
);

DFFPOSX1 _14900_ (
    .CLK(clk_bF$buf15),
    .D(_6791_),
    .Q(\u_pa.Atmp [4])
);

DFFPOSX1 _14901_ (
    .CLK(clk_bF$buf14),
    .D(_6792_),
    .Q(\u_pa.Atmp [5])
);

DFFPOSX1 _14902_ (
    .CLK(clk_bF$buf13),
    .D(_6793_),
    .Q(\u_pa.Atmp [6])
);

DFFPOSX1 _14903_ (
    .CLK(clk_bF$buf12),
    .D(_6794_),
    .Q(\u_pa.Atmp [7])
);

DFFPOSX1 _14904_ (
    .CLK(clk_bF$buf11),
    .D(_6795_),
    .Q(\u_pa.Atmp [8])
);

DFFPOSX1 _14905_ (
    .CLK(clk_bF$buf10),
    .D(_6796_),
    .Q(\u_pa.Atmp [9])
);

DFFPOSX1 _14906_ (
    .CLK(clk_bF$buf9),
    .D(_6797_),
    .Q(\u_pa.Atmp [11])
);

DFFPOSX1 _14907_ (
    .CLK(clk_bF$buf8),
    .D(_6798_),
    .Q(\genblk1[0].u_ce.ISin )
);

BUFX2 _14908_ (
    .A(_7071_[0]),
    .Y(Dout[0])
);

BUFX2 _14909_ (
    .A(_7071_[1]),
    .Y(Dout[1])
);

BUFX2 _14910_ (
    .A(_7071_[10]),
    .Y(Dout[10])
);

BUFX2 _14911_ (
    .A(_7071_[11]),
    .Y(Dout[11])
);

BUFX2 _14912_ (
    .A(_7071_[2]),
    .Y(Dout[2])
);

BUFX2 _14913_ (
    .A(_7071_[3]),
    .Y(Dout[3])
);

BUFX2 _14914_ (
    .A(_7071_[4]),
    .Y(Dout[4])
);

BUFX2 _14915_ (
    .A(_7071_[5]),
    .Y(Dout[5])
);

BUFX2 _14916_ (
    .A(_7071_[6]),
    .Y(Dout[6])
);

BUFX2 _14917_ (
    .A(_7071_[7]),
    .Y(Dout[7])
);

BUFX2 _14918_ (
    .A(_7071_[8]),
    .Y(Dout[8])
);

BUFX2 _14919_ (
    .A(_7071_[9]),
    .Y(Dout[9])
);

BUFX2 _14920_ (
    .A(\u_ot.LoadCtl_6_bF$buf4 ),
    .Y(Vld)
);

INVX1 _7072_ (
    .A(\genblk1[0].u_ce.Acalc [2]),
    .Y(_80_)
);

INVX2 _7073_ (
    .A(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_81_)
);

NOR2X1 _7074_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_81_),
    .Y(_82_)
);

INVX2 _7075_ (
    .A(_82_),
    .Y(_83_)
);

NOR2X1 _7076_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [10]),
    .Y(_84_)
);

INVX4 _7077_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .Y(_85_)
);

NOR2X1 _7078_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.LoadCtl [3]),
    .Y(_86_)
);

OAI21X1 _7079_ (
    .A(_85_),
    .B(\genblk1[0].u_ce.Acalc [8]),
    .C(_86_),
    .Y(_87_)
);

INVX2 _7080_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_88_)
);

AND2X2 _7081_ (
    .A(_88_),
    .B(\genblk1[0].u_ce.LoadCtl [3]),
    .Y(_89_)
);

AOI22X1 _7082_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.Acalc [4]),
    .C(_89_),
    .D(\genblk1[0].u_ce.Acalc [6]),
    .Y(_90_)
);

OAI21X1 _7083_ (
    .A(_84_),
    .B(_87_),
    .C(_90_),
    .Y(_91_)
);

NOR2X1 _7084_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_92_)
);

AOI22X1 _7085_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Acalc [0]),
    .C(_91_),
    .D(_92_),
    .Y(_93_)
);

OAI21X1 _7086_ (
    .A(_80_),
    .B(_83_),
    .C(_93_),
    .Y(\a[1] [0])
);

INVX1 _7087_ (
    .A(\genblk1[0].u_ce.Acalc [9]),
    .Y(_94_)
);

OAI21X1 _7088_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [11]),
    .C(_86_),
    .Y(_95_)
);

AOI21X1 _7089_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_94_),
    .C(_95_),
    .Y(_96_)
);

INVX1 _7090_ (
    .A(\genblk1[0].u_ce.Acalc [5]),
    .Y(_97_)
);

NAND2X1 _7091_ (
    .A(\genblk1[0].u_ce.Acalc [7]),
    .B(_89_),
    .Y(_98_)
);

OAI21X1 _7092_ (
    .A(_88_),
    .B(_97_),
    .C(_98_),
    .Y(_99_)
);

OAI21X1 _7093_ (
    .A(_96_),
    .B(_99_),
    .C(_92_),
    .Y(_100_)
);

AOI22X1 _7094_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.Acalc [1]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Acalc [3]),
    .Y(_101_)
);

NAND2X1 _7095_ (
    .A(_101_),
    .B(_100_),
    .Y(\a[1] [1])
);

INVX1 _7096_ (
    .A(\genblk1[0].u_ce.Ycalc [10]),
    .Y(_102_)
);

OAI21X1 _7097_ (
    .A(_85_),
    .B(\genblk1[0].u_ce.Ycalc [8]),
    .C(_86_),
    .Y(_103_)
);

AOI21X1 _7098_ (
    .A(_85_),
    .B(_102_),
    .C(_103_),
    .Y(_104_)
);

INVX1 _7099_ (
    .A(\genblk1[0].u_ce.Ycalc [4]),
    .Y(_105_)
);

NAND2X1 _7100_ (
    .A(\genblk1[0].u_ce.Ycalc [6]),
    .B(_89_),
    .Y(_106_)
);

OAI21X1 _7101_ (
    .A(_88_),
    .B(_105_),
    .C(_106_),
    .Y(_107_)
);

OAI21X1 _7102_ (
    .A(_104_),
    .B(_107_),
    .C(_92_),
    .Y(_108_)
);

AOI22X1 _7103_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[0].u_ce.Ycalc [0]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Ycalc [2]),
    .Y(_109_)
);

NAND2X1 _7104_ (
    .A(_109_),
    .B(_108_),
    .Y(\genblk1[0].u_ce.Y_ [0])
);

INVX1 _7105_ (
    .A(\genblk1[0].u_ce.Ycalc [9]),
    .Y(_110_)
);

OAI21X1 _7106_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Ycalc [11]),
    .C(_86_),
    .Y(_111_)
);

AOI21X1 _7107_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_110_),
    .C(_111_),
    .Y(_112_)
);

INVX1 _7108_ (
    .A(\genblk1[0].u_ce.Ycalc [5]),
    .Y(_113_)
);

NAND2X1 _7109_ (
    .A(\genblk1[0].u_ce.Ycalc [7]),
    .B(_89_),
    .Y(_114_)
);

OAI21X1 _7110_ (
    .A(_88_),
    .B(_113_),
    .C(_114_),
    .Y(_115_)
);

OAI21X1 _7111_ (
    .A(_112_),
    .B(_115_),
    .C(_92_),
    .Y(_116_)
);

AOI22X1 _7112_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.Ycalc [1]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_117_)
);

NAND2X1 _7113_ (
    .A(_117_),
    .B(_116_),
    .Y(\genblk1[0].u_ce.Y_ [1])
);

INVX1 _7114_ (
    .A(\genblk1[0].u_ce.Xcalc [8]),
    .Y(_118_)
);

OAI21X1 _7115_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Xcalc [10]),
    .C(_86_),
    .Y(_119_)
);

AOI21X1 _7116_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_118_),
    .C(_119_),
    .Y(_120_)
);

INVX1 _7117_ (
    .A(\genblk1[0].u_ce.Xcalc [4]),
    .Y(_121_)
);

NAND2X1 _7118_ (
    .A(\genblk1[0].u_ce.Xcalc [6]),
    .B(_89_),
    .Y(_122_)
);

OAI21X1 _7119_ (
    .A(_88_),
    .B(_121_),
    .C(_122_),
    .Y(_123_)
);

OAI21X1 _7120_ (
    .A(_120_),
    .B(_123_),
    .C(_92_),
    .Y(_124_)
);

AOI22X1 _7121_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.Xcalc [0]),
    .C(_82_),
    .D(\genblk1[0].u_ce.Xcalc [2]),
    .Y(_125_)
);

NAND2X1 _7122_ (
    .A(_125_),
    .B(_124_),
    .Y(\genblk1[0].u_ce.X_ [0])
);

INVX1 _7123_ (
    .A(\genblk1[0].u_ce.Xcalc [3]),
    .Y(_126_)
);

NOR2X1 _7124_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Xcalc [11]),
    .Y(_127_)
);

OAI21X1 _7125_ (
    .A(_85_),
    .B(\genblk1[0].u_ce.Xcalc [9]),
    .C(_86_),
    .Y(_128_)
);

AOI22X1 _7126_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.Xcalc [5]),
    .C(_89_),
    .D(\genblk1[0].u_ce.Xcalc [7]),
    .Y(_129_)
);

OAI21X1 _7127_ (
    .A(_127_),
    .B(_128_),
    .C(_129_),
    .Y(_130_)
);

AOI22X1 _7128_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Xcalc [1]),
    .C(_130_),
    .D(_92_),
    .Y(_131_)
);

OAI21X1 _7129_ (
    .A(_126_),
    .B(_83_),
    .C(_131_),
    .Y(\genblk1[0].u_ce.X_ [1])
);

INVX1 _7130_ (
    .A(\genblk1[0].u_ce.Ycalc [0]),
    .Y(_132_)
);

INVX1 _7131_ (
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .Y(_133_)
);

INVX8 _7132_ (
    .A(1'h0),
    .Y(_134_)
);

INVX8 _7133_ (
    .A(1'h0),
    .Y(_135_)
);

INVX1 _7134_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_136_)
);

NAND2X1 _7135_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_137_)
);

OAI21X1 _7136_ (
    .A(1'h0),
    .B(_136_),
    .C(_137_),
    .Y(_138_)
);

INVX1 _7137_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .Y(_139_)
);

NAND2X1 _7138_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_140_)
);

OAI21X1 _7139_ (
    .A(1'h0),
    .B(_139_),
    .C(_140_),
    .Y(_141_)
);

MUX2X1 _7140_ (
    .A(_141_),
    .B(_138_),
    .S(_135__bF$buf4),
    .Y(_142_)
);

INVX1 _7141_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_143_)
);

NAND2X1 _7142_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_144_)
);

OAI21X1 _7143_ (
    .A(1'h0),
    .B(_143_),
    .C(_144_),
    .Y(_145_)
);

INVX1 _7144_ (
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .Y(_146_)
);

NAND2X1 _7145_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_147_)
);

OAI21X1 _7146_ (
    .A(1'h0),
    .B(_146_),
    .C(_147_),
    .Y(_148_)
);

MUX2X1 _7147_ (
    .A(_148_),
    .B(_145_),
    .S(_135__bF$buf3),
    .Y(_149_)
);

MUX2X1 _7148_ (
    .A(_149_),
    .B(_142_),
    .S(_134__bF$buf4),
    .Y(_150_)
);

NOR2X1 _7149_ (
    .A(_133_),
    .B(_150_),
    .Y(_151_)
);

NAND2X1 _7150_ (
    .A(_133_),
    .B(_150_),
    .Y(_152_)
);

INVX1 _7151_ (
    .A(_152_),
    .Y(_153_)
);

NAND2X1 _7152_ (
    .A(_134__bF$buf3),
    .B(_135__bF$buf2),
    .Y(_154_)
);

OAI21X1 _7153_ (
    .A(1'h0),
    .B(_154_),
    .C(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .Y(_155_)
);

INVX2 _7154_ (
    .A(_155_),
    .Y(_156_)
);

OAI21X1 _7155_ (
    .A(_151_),
    .B(_153_),
    .C(_156_),
    .Y(_157_)
);

OAI21X1 _7156_ (
    .A(_132_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_157_),
    .Y(_0_)
);

INVX8 _7157_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_158_)
);

NAND2X1 _7158_ (
    .A(\genblk1[0].u_ce.Ycalc [1]),
    .B(_158__bF$buf4),
    .Y(_159_)
);

NOR2X1 _7159_ (
    .A(1'h0),
    .B(_154_),
    .Y(_160_)
);

MUX2X1 _7160_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(\genblk1[0].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_161_)
);

MUX2X1 _7161_ (
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .B(\genblk1[0].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_162_)
);

MUX2X1 _7162_ (
    .A(_162_),
    .B(_161_),
    .S(_135__bF$buf1),
    .Y(_163_)
);

INVX2 _7163_ (
    .A(1'h0),
    .Y(_164_)
);

NAND2X1 _7164_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(_164_),
    .Y(_165_)
);

AOI21X1 _7165_ (
    .A(_165_),
    .B(_144_),
    .C(_135__bF$buf0),
    .Y(_166_)
);

NAND3X1 _7166_ (
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .B(_164_),
    .C(_135__bF$buf4),
    .Y(_167_)
);

NAND3X1 _7167_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(1'h0),
    .C(_135__bF$buf3),
    .Y(_168_)
);

NAND3X1 _7168_ (
    .A(_134__bF$buf2),
    .B(_168_),
    .C(_167_),
    .Y(_169_)
);

OAI22X1 _7169_ (
    .A(_166_),
    .B(_169_),
    .C(_134__bF$buf1),
    .D(_163_),
    .Y(_170_)
);

INVX1 _7170_ (
    .A(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_171_)
);

INVX8 _7171_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_172_)
);

INVX1 _7172_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_173_)
);

NAND2X1 _7173_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_174_)
);

OAI21X1 _7174_ (
    .A(1'h0),
    .B(_173_),
    .C(_174_),
    .Y(_175_)
);

INVX1 _7175_ (
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_176_)
);

NAND2X1 _7176_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_177_)
);

OAI21X1 _7177_ (
    .A(1'h0),
    .B(_176_),
    .C(_177_),
    .Y(_178_)
);

MUX2X1 _7178_ (
    .A(_178_),
    .B(_175_),
    .S(_135__bF$buf2),
    .Y(_179_)
);

INVX1 _7179_ (
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_180_)
);

NAND2X1 _7180_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [4]),
    .Y(_181_)
);

OAI21X1 _7181_ (
    .A(1'h0),
    .B(_180_),
    .C(_181_),
    .Y(_182_)
);

INVX1 _7182_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .Y(_183_)
);

NAND2X1 _7183_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_184_)
);

OAI21X1 _7184_ (
    .A(1'h0),
    .B(_183_),
    .C(_184_),
    .Y(_185_)
);

MUX2X1 _7185_ (
    .A(_185_),
    .B(_182_),
    .S(_135__bF$buf1),
    .Y(_186_)
);

MUX2X1 _7186_ (
    .A(_186_),
    .B(_179_),
    .S(_134__bF$buf0),
    .Y(_187_)
);

NAND3X1 _7187_ (
    .A(_172__bF$buf5),
    .B(_150_),
    .C(_187_),
    .Y(_188_)
);

MUX2X1 _7188_ (
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_189_)
);

MUX2X1 _7189_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_190_)
);

MUX2X1 _7190_ (
    .A(_190_),
    .B(_189_),
    .S(_135__bF$buf0),
    .Y(_191_)
);

MUX2X1 _7191_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_192_)
);

MUX2X1 _7192_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(\genblk1[0].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_193_)
);

MUX2X1 _7193_ (
    .A(_193_),
    .B(_192_),
    .S(_135__bF$buf4),
    .Y(_194_)
);

MUX2X1 _7194_ (
    .A(_194_),
    .B(_191_),
    .S(_134__bF$buf4),
    .Y(_195_)
);

OAI21X1 _7195_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_170_),
    .C(_195_),
    .Y(_196_)
);

AOI21X1 _7196_ (
    .A(_196_),
    .B(_188_),
    .C(_171_),
    .Y(_197_)
);

INVX1 _7197_ (
    .A(_197_),
    .Y(_198_)
);

NAND3X1 _7198_ (
    .A(_171_),
    .B(_188_),
    .C(_196_),
    .Y(_199_)
);

AND2X2 _7199_ (
    .A(_198_),
    .B(_199_),
    .Y(_200_)
);

OAI21X1 _7200_ (
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .B(_170_),
    .C(_200_),
    .Y(_201_)
);

OR2X2 _7201_ (
    .A(_200_),
    .B(_152_),
    .Y(_202_)
);

AOI21X1 _7202_ (
    .A(_202_),
    .B(_201_),
    .C(_160_),
    .Y(_203_)
);

OAI21X1 _7203_ (
    .A(_158__bF$buf3),
    .B(_203_),
    .C(_159_),
    .Y(_1_)
);

INVX1 _7204_ (
    .A(\genblk1[0].u_ce.ISout ),
    .Y(_204_)
);

NAND2X1 _7205_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .B(\genblk1[0].u_ce.ISin ),
    .Y(_205_)
);

OAI21X1 _7206_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .B(_204_),
    .C(_205_),
    .Y(_2_)
);

NAND2X1 _7207_ (
    .A(\genblk1[0].u_ce.Ycalc [2]),
    .B(_158__bF$buf2),
    .Y(_206_)
);

AOI21X1 _7208_ (
    .A(_152_),
    .B(_199_),
    .C(_197_),
    .Y(_207_)
);

MUX2X1 _7209_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(\genblk1[0].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_208_)
);

MUX2X1 _7210_ (
    .A(_208_),
    .B(_161_),
    .S(1'h0),
    .Y(_209_)
);

MUX2X1 _7211_ (
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_210_)
);

NAND2X1 _7212_ (
    .A(1'h0),
    .B(_134__bF$buf3),
    .Y(_211_)
);

OAI22X1 _7213_ (
    .A(_211_),
    .B(_162_),
    .C(_210_),
    .D(_154_),
    .Y(_212_)
);

AOI21X1 _7214_ (
    .A(1'h0),
    .B(_209_),
    .C(_212_),
    .Y(_213_)
);

AOI21X1 _7215_ (
    .A(_195_),
    .B(_170_),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_214_)
);

NAND2X1 _7216_ (
    .A(_213_),
    .B(_214_),
    .Y(_215_)
);

INVX1 _7217_ (
    .A(_213_),
    .Y(_216_)
);

OAI21X1 _7218_ (
    .A(_150_),
    .B(_187_),
    .C(_172__bF$buf4),
    .Y(_217_)
);

NAND2X1 _7219_ (
    .A(_216_),
    .B(_217_),
    .Y(_218_)
);

AOI21X1 _7220_ (
    .A(_218_),
    .B(_215_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_219_)
);

NAND3X1 _7221_ (
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .B(_215_),
    .C(_218_),
    .Y(_220_)
);

INVX1 _7222_ (
    .A(_220_),
    .Y(_221_)
);

OR2X2 _7223_ (
    .A(_221_),
    .B(_219_),
    .Y(_222_)
);

NOR2X1 _7224_ (
    .A(_207_),
    .B(_222_),
    .Y(_223_)
);

INVX1 _7225_ (
    .A(_223_),
    .Y(_224_)
);

OAI21X1 _7226_ (
    .A(_219_),
    .B(_221_),
    .C(_207_),
    .Y(_225_)
);

AOI21X1 _7227_ (
    .A(_224_),
    .B(_225_),
    .C(_160_),
    .Y(_226_)
);

INVX2 _7228_ (
    .A(_160_),
    .Y(_227_)
);

OAI21X1 _7229_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_227_),
    .C(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .Y(_228_)
);

OAI21X1 _7230_ (
    .A(_228_),
    .B(_226_),
    .C(_206_),
    .Y(_3_)
);

INVX1 _7231_ (
    .A(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_229_)
);

INVX2 _7232_ (
    .A(_228_),
    .Y(_230_)
);

OAI21X1 _7233_ (
    .A(_219_),
    .B(_207_),
    .C(_220_),
    .Y(_231_)
);

INVX1 _7234_ (
    .A(_231_),
    .Y(_232_)
);

INVX1 _7235_ (
    .A(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_233_)
);

NAND3X1 _7236_ (
    .A(_170_),
    .B(_195_),
    .C(_213_),
    .Y(_234_)
);

INVX1 _7237_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .Y(_235_)
);

NAND2X1 _7238_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_236_)
);

OAI21X1 _7239_ (
    .A(1'h0),
    .B(_235_),
    .C(_236_),
    .Y(_237_)
);

NAND2X1 _7240_ (
    .A(_135__bF$buf3),
    .B(_189_),
    .Y(_238_)
);

OAI21X1 _7241_ (
    .A(_135__bF$buf2),
    .B(_237_),
    .C(_238_),
    .Y(_239_)
);

NOR2X1 _7242_ (
    .A(1'h0),
    .B(_135__bF$buf1),
    .Y(_240_)
);

NOR2X1 _7243_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_241_)
);

AOI22X1 _7244_ (
    .A(_182_),
    .B(_241_),
    .C(_240_),
    .D(_178_),
    .Y(_242_)
);

OAI21X1 _7245_ (
    .A(_134__bF$buf2),
    .B(_239_),
    .C(_242_),
    .Y(_243_)
);

NAND3X1 _7246_ (
    .A(_172__bF$buf3),
    .B(_243_),
    .C(_234_),
    .Y(_244_)
);

INVX1 _7247_ (
    .A(_234_),
    .Y(_245_)
);

INVX1 _7248_ (
    .A(_243_),
    .Y(_246_)
);

OAI21X1 _7249_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_245_),
    .C(_246_),
    .Y(_247_)
);

NAND3X1 _7250_ (
    .A(_233_),
    .B(_244_),
    .C(_247_),
    .Y(_248_)
);

AOI21X1 _7251_ (
    .A(_247_),
    .B(_244_),
    .C(_233_),
    .Y(_249_)
);

INVX1 _7252_ (
    .A(_249_),
    .Y(_250_)
);

NAND2X1 _7253_ (
    .A(_248_),
    .B(_250_),
    .Y(_251_)
);

AOI21X1 _7254_ (
    .A(_251_),
    .B(_232_),
    .C(_160_),
    .Y(_252_)
);

OAI21X1 _7255_ (
    .A(_232_),
    .B(_251_),
    .C(_252_),
    .Y(_253_)
);

AOI22X1 _7256_ (
    .A(_229_),
    .B(_158__bF$buf1),
    .C(_253_),
    .D(_230_),
    .Y(_4_)
);

AOI21X1 _7257_ (
    .A(_231_),
    .B(_248_),
    .C(_249_),
    .Y(_254_)
);

INVX1 _7258_ (
    .A(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_255_)
);

INVX1 _7259_ (
    .A(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_256_)
);

NAND2X1 _7260_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_257_)
);

OAI21X1 _7261_ (
    .A(1'h0),
    .B(_256_),
    .C(_257_),
    .Y(_258_)
);

NAND2X1 _7262_ (
    .A(_135__bF$buf0),
    .B(_208_),
    .Y(_259_)
);

OAI21X1 _7263_ (
    .A(_135__bF$buf4),
    .B(_258_),
    .C(_259_),
    .Y(_260_)
);

NAND2X1 _7264_ (
    .A(_134__bF$buf1),
    .B(_163_),
    .Y(_261_)
);

OAI21X1 _7265_ (
    .A(_134__bF$buf0),
    .B(_260_),
    .C(_261_),
    .Y(_262_)
);

INVX2 _7266_ (
    .A(_262_),
    .Y(_263_)
);

OAI21X1 _7267_ (
    .A(_243_),
    .B(_234_),
    .C(_172__bF$buf2),
    .Y(_264_)
);

OR2X2 _7268_ (
    .A(_264_),
    .B(_263_),
    .Y(_265_)
);

NOR2X1 _7269_ (
    .A(_243_),
    .B(_234_),
    .Y(_266_)
);

OAI21X1 _7270_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_266_),
    .C(_263_),
    .Y(_267_)
);

NAND3X1 _7271_ (
    .A(_255_),
    .B(_267_),
    .C(_265_),
    .Y(_268_)
);

NOR2X1 _7272_ (
    .A(_263_),
    .B(_264_),
    .Y(_269_)
);

AND2X2 _7273_ (
    .A(_264_),
    .B(_263_),
    .Y(_270_)
);

OAI21X1 _7274_ (
    .A(_269_),
    .B(_270_),
    .C(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_271_)
);

NAND2X1 _7275_ (
    .A(_271_),
    .B(_268_),
    .Y(_272_)
);

AOI21X1 _7276_ (
    .A(_254_),
    .B(_272_),
    .C(_160_),
    .Y(_273_)
);

OAI21X1 _7277_ (
    .A(_254_),
    .B(_272_),
    .C(_273_),
    .Y(_274_)
);

AOI22X1 _7278_ (
    .A(_105_),
    .B(_158__bF$buf0),
    .C(_274_),
    .D(_230_),
    .Y(_5_)
);

OAI21X1 _7279_ (
    .A(_272_),
    .B(_254_),
    .C(_271_),
    .Y(_275_)
);

INVX1 _7280_ (
    .A(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_276_)
);

NAND3X1 _7281_ (
    .A(_246_),
    .B(_263_),
    .C(_245_),
    .Y(_277_)
);

NAND2X1 _7282_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_278_)
);

INVX1 _7283_ (
    .A(_278_),
    .Y(_279_)
);

AOI21X1 _7284_ (
    .A(_237_),
    .B(_135__bF$buf3),
    .C(_279_),
    .Y(_280_)
);

NAND2X1 _7285_ (
    .A(_134__bF$buf4),
    .B(_191_),
    .Y(_281_)
);

OAI21X1 _7286_ (
    .A(_134__bF$buf3),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

NAND3X1 _7287_ (
    .A(_172__bF$buf1),
    .B(_282_),
    .C(_277_),
    .Y(_283_)
);

NOR3X1 _7288_ (
    .A(_243_),
    .B(_262_),
    .C(_234_),
    .Y(_284_)
);

INVX1 _7289_ (
    .A(_282_),
    .Y(_285_)
);

OAI21X1 _7290_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_284_),
    .C(_285_),
    .Y(_286_)
);

NAND3X1 _7291_ (
    .A(_276_),
    .B(_283_),
    .C(_286_),
    .Y(_287_)
);

AOI21X1 _7292_ (
    .A(_286_),
    .B(_283_),
    .C(_276_),
    .Y(_288_)
);

INVX1 _7293_ (
    .A(_288_),
    .Y(_289_)
);

NAND2X1 _7294_ (
    .A(_287_),
    .B(_289_),
    .Y(_290_)
);

AND2X2 _7295_ (
    .A(_275_),
    .B(_290_),
    .Y(_291_)
);

OAI21X1 _7296_ (
    .A(_290_),
    .B(_275_),
    .C(_227_),
    .Y(_292_)
);

OAI21X1 _7297_ (
    .A(_292_),
    .B(_291_),
    .C(_230_),
    .Y(_293_)
);

OAI21X1 _7298_ (
    .A(_113_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_293_),
    .Y(_6_)
);

INVX1 _7299_ (
    .A(\genblk1[0].u_ce.Ycalc [6]),
    .Y(_294_)
);

INVX1 _7300_ (
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_295_)
);

NAND3X1 _7301_ (
    .A(_263_),
    .B(_285_),
    .C(_266_),
    .Y(_296_)
);

AOI21X1 _7302_ (
    .A(_258_),
    .B(_135__bF$buf2),
    .C(_279_),
    .Y(_297_)
);

NAND2X1 _7303_ (
    .A(_134__bF$buf2),
    .B(_209_),
    .Y(_298_)
);

OAI21X1 _7304_ (
    .A(_134__bF$buf1),
    .B(_297_),
    .C(_298_),
    .Y(_299_)
);

NAND3X1 _7305_ (
    .A(_172__bF$buf0),
    .B(_299_),
    .C(_296_),
    .Y(_300_)
);

INVX1 _7306_ (
    .A(_299_),
    .Y(_301_)
);

OAI21X1 _7307_ (
    .A(_282_),
    .B(_277_),
    .C(_172__bF$buf5),
    .Y(_302_)
);

NAND2X1 _7308_ (
    .A(_301_),
    .B(_302_),
    .Y(_303_)
);

NAND3X1 _7309_ (
    .A(_295_),
    .B(_300_),
    .C(_303_),
    .Y(_304_)
);

NAND3X1 _7310_ (
    .A(_172__bF$buf4),
    .B(_301_),
    .C(_296_),
    .Y(_305_)
);

NAND2X1 _7311_ (
    .A(_299_),
    .B(_302_),
    .Y(_306_)
);

NAND3X1 _7312_ (
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .B(_305_),
    .C(_306_),
    .Y(_307_)
);

NAND2X1 _7313_ (
    .A(_304_),
    .B(_307_),
    .Y(_308_)
);

AOI21X1 _7314_ (
    .A(_265_),
    .B(_267_),
    .C(_255_),
    .Y(_309_)
);

NOR2X1 _7315_ (
    .A(_309_),
    .B(_288_),
    .Y(_310_)
);

OAI21X1 _7316_ (
    .A(_272_),
    .B(_254_),
    .C(_310_),
    .Y(_311_)
);

NAND2X1 _7317_ (
    .A(_287_),
    .B(_311_),
    .Y(_312_)
);

AOI21X1 _7318_ (
    .A(_312_),
    .B(_308_),
    .C(_160_),
    .Y(_313_)
);

OAI21X1 _7319_ (
    .A(_308_),
    .B(_312_),
    .C(_313_),
    .Y(_314_)
);

AOI22X1 _7320_ (
    .A(_294_),
    .B(_158__bF$buf4),
    .C(_314_),
    .D(_230_),
    .Y(_7_)
);

INVX1 _7321_ (
    .A(\genblk1[0].u_ce.Ycalc [7]),
    .Y(_315_)
);

AOI21X1 _7322_ (
    .A(_303_),
    .B(_300_),
    .C(_295_),
    .Y(_316_)
);

AND2X2 _7323_ (
    .A(_268_),
    .B(_271_),
    .Y(_317_)
);

NAND3X1 _7324_ (
    .A(_287_),
    .B(_289_),
    .C(_317_),
    .Y(_318_)
);

AOI21X1 _7325_ (
    .A(_309_),
    .B(_287_),
    .C(_288_),
    .Y(_319_)
);

OAI21X1 _7326_ (
    .A(_254_),
    .B(_318_),
    .C(_319_),
    .Y(_320_)
);

AOI21X1 _7327_ (
    .A(_320_),
    .B(_304_),
    .C(_316_),
    .Y(_321_)
);

INVX1 _7328_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_322_)
);

NAND3X1 _7329_ (
    .A(_285_),
    .B(_301_),
    .C(_284_),
    .Y(_323_)
);

INVX1 _7330_ (
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_324_)
);

NOR2X1 _7331_ (
    .A(_134__bF$buf0),
    .B(_324_),
    .Y(_325_)
);

INVX1 _7332_ (
    .A(_325_),
    .Y(_326_)
);

OAI21X1 _7333_ (
    .A(1'h0),
    .B(_239_),
    .C(_326_),
    .Y(_327_)
);

NAND3X1 _7334_ (
    .A(_172__bF$buf3),
    .B(_327_),
    .C(_323_),
    .Y(_328_)
);

INVX1 _7335_ (
    .A(_327_),
    .Y(_329_)
);

OAI21X1 _7336_ (
    .A(_299_),
    .B(_296_),
    .C(_172__bF$buf2),
    .Y(_330_)
);

NAND2X1 _7337_ (
    .A(_329_),
    .B(_330_),
    .Y(_331_)
);

NAND3X1 _7338_ (
    .A(_322_),
    .B(_328_),
    .C(_331_),
    .Y(_332_)
);

NAND3X1 _7339_ (
    .A(_172__bF$buf1),
    .B(_329_),
    .C(_323_),
    .Y(_333_)
);

NAND2X1 _7340_ (
    .A(_327_),
    .B(_330_),
    .Y(_334_)
);

NAND3X1 _7341_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(_333_),
    .C(_334_),
    .Y(_335_)
);

NAND2X1 _7342_ (
    .A(_332_),
    .B(_335_),
    .Y(_336_)
);

INVX1 _7343_ (
    .A(_336_),
    .Y(_337_)
);

NOR2X1 _7344_ (
    .A(_337_),
    .B(_321_),
    .Y(_338_)
);

OAI21X1 _7345_ (
    .A(_308_),
    .B(_312_),
    .C(_307_),
    .Y(_339_)
);

OAI21X1 _7346_ (
    .A(_336_),
    .B(_339_),
    .C(_227_),
    .Y(_340_)
);

OAI21X1 _7347_ (
    .A(_172__bF$buf0),
    .B(_227_),
    .C(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_341_)
);

INVX1 _7348_ (
    .A(_341_),
    .Y(_342_)
);

OAI21X1 _7349_ (
    .A(_340_),
    .B(_338_),
    .C(_342_),
    .Y(_343_)
);

OAI21X1 _7350_ (
    .A(_315_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_343_),
    .Y(_8_)
);

INVX1 _7351_ (
    .A(\genblk1[0].u_ce.Ycalc [8]),
    .Y(_344_)
);

OAI21X1 _7352_ (
    .A(_307_),
    .B(_336_),
    .C(_335_),
    .Y(_345_)
);

NOR2X1 _7353_ (
    .A(_308_),
    .B(_336_),
    .Y(_346_)
);

AOI21X1 _7354_ (
    .A(_346_),
    .B(_320_),
    .C(_345_),
    .Y(_347_)
);

INVX1 _7355_ (
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_348_)
);

OR2X2 _7356_ (
    .A(_323_),
    .B(_327_),
    .Y(_349_)
);

OAI21X1 _7357_ (
    .A(1'h0),
    .B(_260_),
    .C(_326_),
    .Y(_350_)
);

NAND3X1 _7358_ (
    .A(_172__bF$buf5),
    .B(_350_),
    .C(_349_),
    .Y(_351_)
);

NOR2X1 _7359_ (
    .A(_327_),
    .B(_323_),
    .Y(_352_)
);

INVX1 _7360_ (
    .A(_350_),
    .Y(_353_)
);

OAI21X1 _7361_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_352_),
    .C(_353_),
    .Y(_354_)
);

NAND3X1 _7362_ (
    .A(_348_),
    .B(_354_),
    .C(_351_),
    .Y(_355_)
);

NAND3X1 _7363_ (
    .A(_172__bF$buf4),
    .B(_353_),
    .C(_349_),
    .Y(_356_)
);

OAI21X1 _7364_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_352_),
    .C(_350_),
    .Y(_357_)
);

NAND3X1 _7365_ (
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .B(_357_),
    .C(_356_),
    .Y(_358_)
);

AND2X2 _7366_ (
    .A(_355_),
    .B(_358_),
    .Y(_359_)
);

INVX1 _7367_ (
    .A(_359_),
    .Y(_360_)
);

AOI21X1 _7368_ (
    .A(_347_),
    .B(_360_),
    .C(_160_),
    .Y(_361_)
);

OAI21X1 _7369_ (
    .A(_347_),
    .B(_360_),
    .C(_361_),
    .Y(_362_)
);

AOI22X1 _7370_ (
    .A(_344_),
    .B(_158__bF$buf3),
    .C(_362_),
    .D(_342_),
    .Y(_9_)
);

NAND2X1 _7371_ (
    .A(_316_),
    .B(_332_),
    .Y(_363_)
);

AND2X2 _7372_ (
    .A(_363_),
    .B(_335_),
    .Y(_364_)
);

AND2X2 _7373_ (
    .A(_304_),
    .B(_307_),
    .Y(_365_)
);

NAND3X1 _7374_ (
    .A(_332_),
    .B(_335_),
    .C(_365_),
    .Y(_366_)
);

OAI21X1 _7375_ (
    .A(_312_),
    .B(_366_),
    .C(_364_),
    .Y(_367_)
);

INVX1 _7376_ (
    .A(_358_),
    .Y(_368_)
);

AOI21X1 _7377_ (
    .A(_367_),
    .B(_355_),
    .C(_368_),
    .Y(_369_)
);

INVX1 _7378_ (
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_370_)
);

NOR3X1 _7379_ (
    .A(_327_),
    .B(_350_),
    .C(_323_),
    .Y(_371_)
);

INVX1 _7380_ (
    .A(_371_),
    .Y(_372_)
);

OAI21X1 _7381_ (
    .A(1'h0),
    .B(_280_),
    .C(_326_),
    .Y(_373_)
);

NAND3X1 _7382_ (
    .A(_172__bF$buf3),
    .B(_373_),
    .C(_372_),
    .Y(_374_)
);

INVX1 _7383_ (
    .A(_373_),
    .Y(_375_)
);

OAI21X1 _7384_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_371_),
    .C(_375_),
    .Y(_376_)
);

NAND3X1 _7385_ (
    .A(_370_),
    .B(_376_),
    .C(_374_),
    .Y(_377_)
);

NAND3X1 _7386_ (
    .A(_172__bF$buf2),
    .B(_375_),
    .C(_372_),
    .Y(_378_)
);

OAI21X1 _7387_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_371_),
    .C(_373_),
    .Y(_379_)
);

NAND3X1 _7388_ (
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .B(_379_),
    .C(_378_),
    .Y(_380_)
);

AND2X2 _7389_ (
    .A(_377_),
    .B(_380_),
    .Y(_381_)
);

AND2X2 _7390_ (
    .A(_369_),
    .B(_381_),
    .Y(_382_)
);

OAI21X1 _7391_ (
    .A(_381_),
    .B(_369_),
    .C(_227_),
    .Y(_383_)
);

OAI21X1 _7392_ (
    .A(_383_),
    .B(_382_),
    .C(_230_),
    .Y(_384_)
);

OAI21X1 _7393_ (
    .A(_110_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_384_),
    .Y(_10_)
);

INVX1 _7394_ (
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .Y(_385_)
);

OAI21X1 _7395_ (
    .A(1'h0),
    .B(_297_),
    .C(_326_),
    .Y(_386_)
);

INVX1 _7396_ (
    .A(_386_),
    .Y(_387_)
);

AOI21X1 _7397_ (
    .A(_371_),
    .B(_375_),
    .C(_387_),
    .Y(_388_)
);

NAND3X1 _7398_ (
    .A(_375_),
    .B(_387_),
    .C(_371_),
    .Y(_389_)
);

NAND2X1 _7399_ (
    .A(_172__bF$buf1),
    .B(_389_),
    .Y(_390_)
);

NAND2X1 _7400_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_386_),
    .Y(_391_)
);

OAI21X1 _7401_ (
    .A(_388_),
    .B(_390_),
    .C(_391_),
    .Y(_392_)
);

NAND2X1 _7402_ (
    .A(_385_),
    .B(_392_),
    .Y(_393_)
);

INVX1 _7403_ (
    .A(_388_),
    .Y(_394_)
);

AND2X2 _7404_ (
    .A(_389_),
    .B(_172__bF$buf0),
    .Y(_395_)
);

NAND2X1 _7405_ (
    .A(_394_),
    .B(_395_),
    .Y(_396_)
);

NAND3X1 _7406_ (
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .B(_391_),
    .C(_396_),
    .Y(_397_)
);

NAND2X1 _7407_ (
    .A(_393_),
    .B(_397_),
    .Y(_398_)
);

AOI21X1 _7408_ (
    .A(_374_),
    .B(_376_),
    .C(_370_),
    .Y(_399_)
);

AOI21X1 _7409_ (
    .A(_368_),
    .B(_377_),
    .C(_399_),
    .Y(_400_)
);

NAND3X1 _7410_ (
    .A(_359_),
    .B(_381_),
    .C(_367_),
    .Y(_401_)
);

AOI21X1 _7411_ (
    .A(_401_),
    .B(_400_),
    .C(_398_),
    .Y(_402_)
);

AND2X2 _7412_ (
    .A(_397_),
    .B(_393_),
    .Y(_403_)
);

NAND3X1 _7413_ (
    .A(_377_),
    .B(_380_),
    .C(_359_),
    .Y(_404_)
);

OAI21X1 _7414_ (
    .A(_404_),
    .B(_347_),
    .C(_400_),
    .Y(_405_)
);

OAI21X1 _7415_ (
    .A(_403_),
    .B(_405_),
    .C(_227_),
    .Y(_406_)
);

OR2X2 _7416_ (
    .A(_406_),
    .B(_402_),
    .Y(_407_)
);

AOI22X1 _7417_ (
    .A(_102_),
    .B(_158__bF$buf2),
    .C(_407_),
    .D(_230_),
    .Y(_11_)
);

NAND2X1 _7418_ (
    .A(\genblk1[0].u_ce.Ycalc [11]),
    .B(_158__bF$buf1),
    .Y(_408_)
);

INVX1 _7419_ (
    .A(_397_),
    .Y(_409_)
);

NAND2X1 _7420_ (
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .B(_324_),
    .Y(_410_)
);

INVX1 _7421_ (
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_411_)
);

NAND2X1 _7422_ (
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .B(_411_),
    .Y(_412_)
);

NAND2X1 _7423_ (
    .A(_410_),
    .B(_412_),
    .Y(_413_)
);

INVX1 _7424_ (
    .A(_413_),
    .Y(_414_)
);

NAND2X1 _7425_ (
    .A(_414_),
    .B(_390_),
    .Y(_415_)
);

NAND2X1 _7426_ (
    .A(_413_),
    .B(_395_),
    .Y(_416_)
);

NAND2X1 _7427_ (
    .A(_415_),
    .B(_416_),
    .Y(_417_)
);

INVX1 _7428_ (
    .A(_417_),
    .Y(_418_)
);

NOR3X1 _7429_ (
    .A(_409_),
    .B(_418_),
    .C(_402_),
    .Y(_419_)
);

AOI21X1 _7430_ (
    .A(_405_),
    .B(_403_),
    .C(_409_),
    .Y(_420_)
);

OAI21X1 _7431_ (
    .A(_417_),
    .B(_420_),
    .C(_227_),
    .Y(_421_)
);

OAI21X1 _7432_ (
    .A(_419_),
    .B(_421_),
    .C(_230_),
    .Y(_422_)
);

NAND2X1 _7433_ (
    .A(_408_),
    .B(_422_),
    .Y(_12_)
);

NAND2X1 _7434_ (
    .A(\genblk1[0].u_ce.Xcalc [0]),
    .B(_158__bF$buf0),
    .Y(_423_)
);

INVX1 _7435_ (
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_424_)
);

NAND2X1 _7436_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_425_)
);

OAI21X1 _7437_ (
    .A(1'h0),
    .B(_424_),
    .C(_425_),
    .Y(_426_)
);

NAND2X1 _7438_ (
    .A(1'h0),
    .B(_426_),
    .Y(_427_)
);

NOR2X1 _7439_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_428_)
);

NOR2X1 _7440_ (
    .A(1'h0),
    .B(_164_),
    .Y(_429_)
);

AOI22X1 _7441_ (
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .B(_428_),
    .C(_429_),
    .D(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_430_)
);

NAND3X1 _7442_ (
    .A(_134__bF$buf4),
    .B(_427_),
    .C(_430_),
    .Y(_431_)
);

NAND2X1 _7443_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_432_)
);

OAI21X1 _7444_ (
    .A(1'h0),
    .B(_295_),
    .C(_432_),
    .Y(_433_)
);

NAND2X1 _7445_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_434_)
);

OAI21X1 _7446_ (
    .A(1'h0),
    .B(_255_),
    .C(_434_),
    .Y(_435_)
);

MUX2X1 _7447_ (
    .A(_435_),
    .B(_433_),
    .S(_135__bF$buf1),
    .Y(_436_)
);

NAND2X1 _7448_ (
    .A(1'h0),
    .B(_436_),
    .Y(_437_)
);

AND2X2 _7449_ (
    .A(_431_),
    .B(_437_),
    .Y(_438_)
);

NOR2X1 _7450_ (
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .B(_438_),
    .Y(_439_)
);

NAND2X1 _7451_ (
    .A(_135__bF$buf0),
    .B(_435_),
    .Y(_440_)
);

NAND2X1 _7452_ (
    .A(1'h0),
    .B(_433_),
    .Y(_441_)
);

NAND2X1 _7453_ (
    .A(_440_),
    .B(_441_),
    .Y(_442_)
);

OAI21X1 _7454_ (
    .A(_134__bF$buf3),
    .B(_442_),
    .C(_431_),
    .Y(_443_)
);

OAI21X1 _7455_ (
    .A(_146_),
    .B(_443_),
    .C(_156_),
    .Y(_444_)
);

OAI21X1 _7456_ (
    .A(_444_),
    .B(_439_),
    .C(_423_),
    .Y(_13_)
);

NAND2X1 _7457_ (
    .A(\genblk1[0].u_ce.Xcalc [1]),
    .B(_158__bF$buf4),
    .Y(_445_)
);

NOR2X1 _7458_ (
    .A(_146_),
    .B(_443_),
    .Y(_446_)
);

NAND2X1 _7459_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_447_)
);

OAI21X1 _7460_ (
    .A(1'h0),
    .B(_233_),
    .C(_447_),
    .Y(_448_)
);

NAND2X1 _7461_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_449_)
);

OAI21X1 _7462_ (
    .A(1'h0),
    .B(_171_),
    .C(_449_),
    .Y(_450_)
);

MUX2X1 _7463_ (
    .A(_450_),
    .B(_448_),
    .S(_135__bF$buf4),
    .Y(_451_)
);

NAND2X1 _7464_ (
    .A(_134__bF$buf2),
    .B(_451_),
    .Y(_452_)
);

NAND2X1 _7465_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_453_)
);

OAI21X1 _7466_ (
    .A(1'h0),
    .B(_322_),
    .C(_453_),
    .Y(_454_)
);

INVX1 _7467_ (
    .A(_454_),
    .Y(_455_)
);

NAND2X1 _7468_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_456_)
);

OAI21X1 _7469_ (
    .A(1'h0),
    .B(_276_),
    .C(_456_),
    .Y(_457_)
);

NAND2X1 _7470_ (
    .A(_135__bF$buf3),
    .B(_457_),
    .Y(_458_)
);

OAI21X1 _7471_ (
    .A(_135__bF$buf2),
    .B(_455_),
    .C(_458_),
    .Y(_459_)
);

OAI21X1 _7472_ (
    .A(_134__bF$buf1),
    .B(_459_),
    .C(_452_),
    .Y(_460_)
);

NAND3X1 _7473_ (
    .A(_172__bF$buf5),
    .B(_460_),
    .C(_438_),
    .Y(_461_)
);

MUX2X1 _7474_ (
    .A(_457_),
    .B(_454_),
    .S(_135__bF$buf1),
    .Y(_462_)
);

MUX2X1 _7475_ (
    .A(_462_),
    .B(_451_),
    .S(1'h0),
    .Y(_463_)
);

OAI21X1 _7476_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_443_),
    .C(_463_),
    .Y(_464_)
);

AOI21X1 _7477_ (
    .A(_461_),
    .B(_464_),
    .C(_183_),
    .Y(_465_)
);

INVX1 _7478_ (
    .A(_465_),
    .Y(_466_)
);

NAND3X1 _7479_ (
    .A(_183_),
    .B(_464_),
    .C(_461_),
    .Y(_467_)
);

AND2X2 _7480_ (
    .A(_466_),
    .B(_467_),
    .Y(_468_)
);

NAND2X1 _7481_ (
    .A(_446_),
    .B(_468_),
    .Y(_469_)
);

OR2X2 _7482_ (
    .A(_468_),
    .B(_446_),
    .Y(_470_)
);

AOI21X1 _7483_ (
    .A(_470_),
    .B(_469_),
    .C(_160_),
    .Y(_471_)
);

OAI21X1 _7484_ (
    .A(_158__bF$buf3),
    .B(_471_),
    .C(_445_),
    .Y(_14_)
);

NAND2X1 _7485_ (
    .A(\genblk1[0].u_ce.Xcalc [2]),
    .B(_158__bF$buf2),
    .Y(_472_)
);

AOI21X1 _7486_ (
    .A(_446_),
    .B(_467_),
    .C(_465_),
    .Y(_473_)
);

NAND2X1 _7487_ (
    .A(_443_),
    .B(_460_),
    .Y(_474_)
);

NAND2X1 _7488_ (
    .A(1'h0),
    .B(_370_),
    .Y(_475_)
);

OAI21X1 _7489_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .C(_475_),
    .Y(_476_)
);

NAND2X1 _7490_ (
    .A(_135__bF$buf0),
    .B(_433_),
    .Y(_477_)
);

OAI21X1 _7491_ (
    .A(_135__bF$buf4),
    .B(_476_),
    .C(_477_),
    .Y(_478_)
);

NAND2X1 _7492_ (
    .A(_241_),
    .B(_426_),
    .Y(_479_)
);

NAND2X1 _7493_ (
    .A(_435_),
    .B(_240_),
    .Y(_480_)
);

NAND2X1 _7494_ (
    .A(_479_),
    .B(_480_),
    .Y(_481_)
);

AOI21X1 _7495_ (
    .A(_478_),
    .B(1'h0),
    .C(_481_),
    .Y(_482_)
);

INVX1 _7496_ (
    .A(_482_),
    .Y(_483_)
);

NAND3X1 _7497_ (
    .A(_172__bF$buf4),
    .B(_483_),
    .C(_474_),
    .Y(_484_)
);

AOI21X1 _7498_ (
    .A(_431_),
    .B(_437_),
    .C(_463_),
    .Y(_485_)
);

OAI21X1 _7499_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_485_),
    .C(_482_),
    .Y(_486_)
);

NAND3X1 _7500_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(_486_),
    .C(_484_),
    .Y(_487_)
);

INVX1 _7501_ (
    .A(_487_),
    .Y(_488_)
);

AOI21X1 _7502_ (
    .A(_484_),
    .B(_486_),
    .C(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_489_)
);

NOR2X1 _7503_ (
    .A(_489_),
    .B(_488_),
    .Y(_490_)
);

AND2X2 _7504_ (
    .A(_490_),
    .B(_473_),
    .Y(_491_)
);

NOR2X1 _7505_ (
    .A(_473_),
    .B(_490_),
    .Y(_492_)
);

OAI21X1 _7506_ (
    .A(_492_),
    .B(_491_),
    .C(_227_),
    .Y(_493_)
);

OAI21X1 _7507_ (
    .A(_158__bF$buf1),
    .B(_493_),
    .C(_472_),
    .Y(_15_)
);

OAI21X1 _7508_ (
    .A(_489_),
    .B(_473_),
    .C(_487_),
    .Y(_494_)
);

INVX1 _7509_ (
    .A(_494_),
    .Y(_495_)
);

NAND2X1 _7510_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [10]),
    .Y(_496_)
);

OAI21X1 _7511_ (
    .A(1'h0),
    .B(_370_),
    .C(_496_),
    .Y(_497_)
);

MUX2X1 _7512_ (
    .A(_497_),
    .B(_454_),
    .S(1'h0),
    .Y(_498_)
);

NOR2X1 _7513_ (
    .A(_134__bF$buf0),
    .B(_498_),
    .Y(_499_)
);

NAND2X1 _7514_ (
    .A(_241_),
    .B(_448_),
    .Y(_500_)
);

NAND2X1 _7515_ (
    .A(_457_),
    .B(_240_),
    .Y(_501_)
);

NAND2X1 _7516_ (
    .A(_500_),
    .B(_501_),
    .Y(_502_)
);

OR2X2 _7517_ (
    .A(_499_),
    .B(_502_),
    .Y(_503_)
);

OAI21X1 _7518_ (
    .A(_483_),
    .B(_474_),
    .C(_172__bF$buf3),
    .Y(_504_)
);

OR2X2 _7519_ (
    .A(_504_),
    .B(_503_),
    .Y(_505_)
);

OAI21X1 _7520_ (
    .A(_499_),
    .B(_502_),
    .C(_504_),
    .Y(_506_)
);

AOI21X1 _7521_ (
    .A(_505_),
    .B(_506_),
    .C(_180_),
    .Y(_507_)
);

INVX1 _7522_ (
    .A(_507_),
    .Y(_508_)
);

NAND3X1 _7523_ (
    .A(_180_),
    .B(_506_),
    .C(_505_),
    .Y(_509_)
);

NAND2X1 _7524_ (
    .A(_509_),
    .B(_508_),
    .Y(_510_)
);

OR2X2 _7525_ (
    .A(_510_),
    .B(_495_),
    .Y(_511_)
);

NAND2X1 _7526_ (
    .A(_495_),
    .B(_510_),
    .Y(_512_)
);

NAND2X1 _7527_ (
    .A(_512_),
    .B(_511_),
    .Y(_513_)
);

AOI22X1 _7528_ (
    .A(_126_),
    .B(_158__bF$buf0),
    .C(_513_),
    .D(_156_),
    .Y(_16_)
);

AOI21X1 _7529_ (
    .A(_494_),
    .B(_509_),
    .C(_507_),
    .Y(_514_)
);

NAND2X1 _7530_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_515_)
);

OAI21X1 _7531_ (
    .A(1'h0),
    .B(_385_),
    .C(_515_),
    .Y(_516_)
);

NAND2X1 _7532_ (
    .A(1'h0),
    .B(_516_),
    .Y(_517_)
);

OAI21X1 _7533_ (
    .A(1'h0),
    .B(_476_),
    .C(_517_),
    .Y(_518_)
);

NAND2X1 _7534_ (
    .A(1'h0),
    .B(_518_),
    .Y(_519_)
);

OAI21X1 _7535_ (
    .A(1'h0),
    .B(_436_),
    .C(_519_),
    .Y(_520_)
);

INVX1 _7536_ (
    .A(_520_),
    .Y(_521_)
);

NAND3X1 _7537_ (
    .A(_482_),
    .B(_443_),
    .C(_460_),
    .Y(_522_)
);

OAI21X1 _7538_ (
    .A(_503_),
    .B(_522_),
    .C(_172__bF$buf2),
    .Y(_523_)
);

OR2X2 _7539_ (
    .A(_523_),
    .B(_521_),
    .Y(_524_)
);

NOR2X1 _7540_ (
    .A(_503_),
    .B(_522_),
    .Y(_525_)
);

OAI21X1 _7541_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_525_),
    .C(_521_),
    .Y(_526_)
);

NAND3X1 _7542_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(_526_),
    .C(_524_),
    .Y(_527_)
);

OR2X2 _7543_ (
    .A(_523_),
    .B(_520_),
    .Y(_528_)
);

OAI21X1 _7544_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_525_),
    .C(_520_),
    .Y(_529_)
);

NAND3X1 _7545_ (
    .A(_139_),
    .B(_529_),
    .C(_528_),
    .Y(_530_)
);

NAND2X1 _7546_ (
    .A(_527_),
    .B(_530_),
    .Y(_531_)
);

OR2X2 _7547_ (
    .A(_514_),
    .B(_531_),
    .Y(_532_)
);

NAND2X1 _7548_ (
    .A(_531_),
    .B(_514_),
    .Y(_533_)
);

NAND2X1 _7549_ (
    .A(_533_),
    .B(_532_),
    .Y(_534_)
);

AOI22X1 _7550_ (
    .A(_121_),
    .B(_158__bF$buf4),
    .C(_534_),
    .D(_156_),
    .Y(_17_)
);

INVX1 _7551_ (
    .A(\genblk1[0].u_ce.Xcalc [5]),
    .Y(_535_)
);

OAI21X1 _7552_ (
    .A(_531_),
    .B(_514_),
    .C(_527_),
    .Y(_536_)
);

NAND2X1 _7553_ (
    .A(_521_),
    .B(_525_),
    .Y(_537_)
);

NOR2X1 _7554_ (
    .A(_135__bF$buf3),
    .B(_411_),
    .Y(_538_)
);

AOI21X1 _7555_ (
    .A(_135__bF$buf2),
    .B(_497_),
    .C(_538_),
    .Y(_539_)
);

NAND2X1 _7556_ (
    .A(_134__bF$buf4),
    .B(_459_),
    .Y(_540_)
);

OAI21X1 _7557_ (
    .A(_134__bF$buf3),
    .B(_539_),
    .C(_540_),
    .Y(_541_)
);

INVX1 _7558_ (
    .A(_541_),
    .Y(_542_)
);

NAND3X1 _7559_ (
    .A(_172__bF$buf1),
    .B(_542_),
    .C(_537_),
    .Y(_543_)
);

NOR2X1 _7560_ (
    .A(_502_),
    .B(_499_),
    .Y(_544_)
);

NAND3X1 _7561_ (
    .A(_482_),
    .B(_544_),
    .C(_485_),
    .Y(_545_)
);

OAI21X1 _7562_ (
    .A(_520_),
    .B(_545_),
    .C(_172__bF$buf0),
    .Y(_546_)
);

NAND2X1 _7563_ (
    .A(_541_),
    .B(_546_),
    .Y(_547_)
);

AOI21X1 _7564_ (
    .A(_543_),
    .B(_547_),
    .C(_176_),
    .Y(_548_)
);

INVX1 _7565_ (
    .A(_548_),
    .Y(_549_)
);

NAND3X1 _7566_ (
    .A(_176_),
    .B(_547_),
    .C(_543_),
    .Y(_550_)
);

NAND2X1 _7567_ (
    .A(_550_),
    .B(_549_),
    .Y(_551_)
);

NOR2X1 _7568_ (
    .A(_551_),
    .B(_536_),
    .Y(_552_)
);

AND2X2 _7569_ (
    .A(_536_),
    .B(_551_),
    .Y(_553_)
);

OAI21X1 _7570_ (
    .A(_552_),
    .B(_553_),
    .C(_156_),
    .Y(_554_)
);

OAI21X1 _7571_ (
    .A(_535_),
    .B(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .C(_554_),
    .Y(_18_)
);

INVX1 _7572_ (
    .A(\genblk1[0].u_ce.Xcalc [6]),
    .Y(_555_)
);

NAND3X1 _7573_ (
    .A(_521_),
    .B(_542_),
    .C(_525_),
    .Y(_556_)
);

AOI21X1 _7574_ (
    .A(_135__bF$buf1),
    .B(_516_),
    .C(_538_),
    .Y(_557_)
);

NAND2X1 _7575_ (
    .A(1'h0),
    .B(_557_),
    .Y(_558_)
);

OAI21X1 _7576_ (
    .A(1'h0),
    .B(_478_),
    .C(_558_),
    .Y(_559_)
);

NAND3X1 _7577_ (
    .A(_172__bF$buf5),
    .B(_559_),
    .C(_556_),
    .Y(_560_)
);

NOR3X1 _7578_ (
    .A(_520_),
    .B(_541_),
    .C(_545_),
    .Y(_561_)
);

INVX1 _7579_ (
    .A(_559_),
    .Y(_562_)
);

OAI21X1 _7580_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_561_),
    .C(_562_),
    .Y(_563_)
);

NAND2X1 _7581_ (
    .A(_560_),
    .B(_563_),
    .Y(_564_)
);

NAND2X1 _7582_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(_564_),
    .Y(_565_)
);

NAND3X1 _7583_ (
    .A(_136_),
    .B(_560_),
    .C(_563_),
    .Y(_566_)
);

NAND2X1 _7584_ (
    .A(_566_),
    .B(_565_),
    .Y(_567_)
);

AOI21X1 _7585_ (
    .A(_528_),
    .B(_529_),
    .C(_139_),
    .Y(_568_)
);

NOR2X1 _7586_ (
    .A(_568_),
    .B(_548_),
    .Y(_569_)
);

OAI21X1 _7587_ (
    .A(_531_),
    .B(_514_),
    .C(_569_),
    .Y(_570_)
);

NAND2X1 _7588_ (
    .A(_550_),
    .B(_570_),
    .Y(_571_)
);

NOR2X1 _7589_ (
    .A(_567_),
    .B(_571_),
    .Y(_572_)
);

AND2X2 _7590_ (
    .A(_565_),
    .B(_566_),
    .Y(_573_)
);

AND2X2 _7591_ (
    .A(_527_),
    .B(_530_),
    .Y(_574_)
);

NAND3X1 _7592_ (
    .A(_550_),
    .B(_574_),
    .C(_549_),
    .Y(_575_)
);

AOI21X1 _7593_ (
    .A(_568_),
    .B(_550_),
    .C(_548_),
    .Y(_576_)
);

OAI21X1 _7594_ (
    .A(_514_),
    .B(_575_),
    .C(_576_),
    .Y(_577_)
);

NOR2X1 _7595_ (
    .A(_573_),
    .B(_577_),
    .Y(_578_)
);

OAI21X1 _7596_ (
    .A(_578_),
    .B(_572_),
    .C(_227_),
    .Y(_579_)
);

NAND2X1 _7597_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_579_),
    .Y(_580_)
);

OAI21X1 _7598_ (
    .A(_555_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_580_),
    .Y(_19_)
);

INVX1 _7599_ (
    .A(\genblk1[0].u_ce.Xcalc [7]),
    .Y(_581_)
);

INVX1 _7600_ (
    .A(_565_),
    .Y(_582_)
);

NAND2X1 _7601_ (
    .A(_559_),
    .B(_561_),
    .Y(_583_)
);

NOR2X1 _7602_ (
    .A(_134__bF$buf2),
    .B(_411_),
    .Y(_584_)
);

INVX1 _7603_ (
    .A(_584_),
    .Y(_585_)
);

OAI21X1 _7604_ (
    .A(1'h0),
    .B(_498_),
    .C(_585_),
    .Y(_586_)
);

NAND3X1 _7605_ (
    .A(_172__bF$buf4),
    .B(_586_),
    .C(_583_),
    .Y(_587_)
);

INVX1 _7606_ (
    .A(_586_),
    .Y(_588_)
);

OAI21X1 _7607_ (
    .A(_562_),
    .B(_556_),
    .C(_172__bF$buf3),
    .Y(_589_)
);

NAND2X1 _7608_ (
    .A(_588_),
    .B(_589_),
    .Y(_590_)
);

NAND3X1 _7609_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(_587_),
    .C(_590_),
    .Y(_591_)
);

NAND3X1 _7610_ (
    .A(_172__bF$buf2),
    .B(_588_),
    .C(_583_),
    .Y(_592_)
);

NAND2X1 _7611_ (
    .A(_586_),
    .B(_589_),
    .Y(_593_)
);

NAND3X1 _7612_ (
    .A(_173_),
    .B(_592_),
    .C(_593_),
    .Y(_594_)
);

NAND2X1 _7613_ (
    .A(_591_),
    .B(_594_),
    .Y(_595_)
);

OAI21X1 _7614_ (
    .A(_582_),
    .B(_572_),
    .C(_595_),
    .Y(_596_)
);

NOR2X1 _7615_ (
    .A(_582_),
    .B(_572_),
    .Y(_597_)
);

INVX1 _7616_ (
    .A(_595_),
    .Y(_598_)
);

AOI21X1 _7617_ (
    .A(_597_),
    .B(_598_),
    .C(_155_),
    .Y(_599_)
);

AOI22X1 _7618_ (
    .A(_581_),
    .B(_158__bF$buf3),
    .C(_599_),
    .D(_596_),
    .Y(_20_)
);

OAI21X1 _7619_ (
    .A(_565_),
    .B(_595_),
    .C(_591_),
    .Y(_600_)
);

NOR2X1 _7620_ (
    .A(_567_),
    .B(_595_),
    .Y(_601_)
);

AOI21X1 _7621_ (
    .A(_601_),
    .B(_577_),
    .C(_600_),
    .Y(_602_)
);

INVX1 _7622_ (
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_603_)
);

NAND3X1 _7623_ (
    .A(_559_),
    .B(_588_),
    .C(_561_),
    .Y(_604_)
);

INVX1 _7624_ (
    .A(_518_),
    .Y(_605_)
);

OAI21X1 _7625_ (
    .A(1'h0),
    .B(_605_),
    .C(_585_),
    .Y(_606_)
);

INVX1 _7626_ (
    .A(_606_),
    .Y(_607_)
);

NAND3X1 _7627_ (
    .A(_172__bF$buf1),
    .B(_607_),
    .C(_604_),
    .Y(_608_)
);

OAI21X1 _7628_ (
    .A(_586_),
    .B(_583_),
    .C(_172__bF$buf0),
    .Y(_609_)
);

NAND2X1 _7629_ (
    .A(_606_),
    .B(_609_),
    .Y(_610_)
);

AOI21X1 _7630_ (
    .A(_610_),
    .B(_608_),
    .C(_603_),
    .Y(_611_)
);

NAND3X1 _7631_ (
    .A(_172__bF$buf5),
    .B(_606_),
    .C(_604_),
    .Y(_612_)
);

NAND2X1 _7632_ (
    .A(_607_),
    .B(_609_),
    .Y(_613_)
);

AOI21X1 _7633_ (
    .A(_613_),
    .B(_612_),
    .C(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_614_)
);

OAI21X1 _7634_ (
    .A(_611_),
    .B(_614_),
    .C(_602_),
    .Y(_615_)
);

INVX1 _7635_ (
    .A(_615_),
    .Y(_616_)
);

OR2X2 _7636_ (
    .A(_611_),
    .B(_614_),
    .Y(_617_)
);

OAI21X1 _7637_ (
    .A(_617_),
    .B(_602_),
    .C(_156_),
    .Y(_618_)
);

OAI22X1 _7638_ (
    .A(_118_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_618_),
    .D(_616_),
    .Y(_21_)
);

NAND2X1 _7639_ (
    .A(\genblk1[0].u_ce.Xcalc [9]),
    .B(_158__bF$buf2),
    .Y(_619_)
);

NOR2X1 _7640_ (
    .A(_617_),
    .B(_602_),
    .Y(_620_)
);

NOR2X1 _7641_ (
    .A(_611_),
    .B(_620_),
    .Y(_621_)
);

OAI21X1 _7642_ (
    .A(1'h0),
    .B(_539_),
    .C(_585_),
    .Y(_622_)
);

INVX1 _7643_ (
    .A(_622_),
    .Y(_623_)
);

OAI21X1 _7644_ (
    .A(_606_),
    .B(_604_),
    .C(_172__bF$buf4),
    .Y(_624_)
);

NAND2X1 _7645_ (
    .A(_623_),
    .B(_624_),
    .Y(_625_)
);

OR2X2 _7646_ (
    .A(_624_),
    .B(_623_),
    .Y(_626_)
);

NAND3X1 _7647_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(_625_),
    .C(_626_),
    .Y(_627_)
);

NAND2X1 _7648_ (
    .A(_625_),
    .B(_626_),
    .Y(_628_)
);

NAND2X1 _7649_ (
    .A(_235_),
    .B(_628_),
    .Y(_629_)
);

NAND2X1 _7650_ (
    .A(_627_),
    .B(_629_),
    .Y(_630_)
);

AND2X2 _7651_ (
    .A(_621_),
    .B(_630_),
    .Y(_631_)
);

OAI21X1 _7652_ (
    .A(_630_),
    .B(_621_),
    .C(_156_),
    .Y(_632_)
);

OAI21X1 _7653_ (
    .A(_632_),
    .B(_631_),
    .C(_619_),
    .Y(_22_)
);

INVX1 _7654_ (
    .A(\genblk1[0].u_ce.Xcalc [10]),
    .Y(_633_)
);

INVX1 _7655_ (
    .A(_627_),
    .Y(_634_)
);

AOI21X1 _7656_ (
    .A(_611_),
    .B(_629_),
    .C(_634_),
    .Y(_635_)
);

NOR2X1 _7657_ (
    .A(_611_),
    .B(_614_),
    .Y(_636_)
);

NAND3X1 _7658_ (
    .A(_627_),
    .B(_629_),
    .C(_636_),
    .Y(_637_)
);

OAI21X1 _7659_ (
    .A(_602_),
    .B(_637_),
    .C(_635_),
    .Y(_638_)
);

OAI21X1 _7660_ (
    .A(1'h0),
    .B(_557_),
    .C(_585_),
    .Y(_639_)
);

INVX1 _7661_ (
    .A(_639_),
    .Y(_640_)
);

OR2X2 _7662_ (
    .A(_604_),
    .B(_606_),
    .Y(_641_)
);

OAI21X1 _7663_ (
    .A(_622_),
    .B(_641_),
    .C(_172__bF$buf3),
    .Y(_642_)
);

NAND2X1 _7664_ (
    .A(_640_),
    .B(_642_),
    .Y(_643_)
);

OR2X2 _7665_ (
    .A(_642_),
    .B(_640_),
    .Y(_644_)
);

NAND3X1 _7666_ (
    .A(\genblk1[0].u_ce.Xin12b [10]),
    .B(_643_),
    .C(_644_),
    .Y(_645_)
);

AND2X2 _7667_ (
    .A(_642_),
    .B(_640_),
    .Y(_646_)
);

NOR2X1 _7668_ (
    .A(_640_),
    .B(_642_),
    .Y(_647_)
);

OAI21X1 _7669_ (
    .A(_647_),
    .B(_646_),
    .C(_256_),
    .Y(_648_)
);

NAND2X1 _7670_ (
    .A(_648_),
    .B(_645_),
    .Y(_649_)
);

AND2X2 _7671_ (
    .A(_638_),
    .B(_649_),
    .Y(_650_)
);

NOR2X1 _7672_ (
    .A(_649_),
    .B(_638_),
    .Y(_651_)
);

NOR2X1 _7673_ (
    .A(_650_),
    .B(_651_),
    .Y(_652_)
);

AOI22X1 _7674_ (
    .A(_633_),
    .B(_158__bF$buf1),
    .C(_652_),
    .D(_156_),
    .Y(_23_)
);

NAND2X1 _7675_ (
    .A(\genblk1[0].u_ce.Xcalc [11]),
    .B(_158__bF$buf0),
    .Y(_653_)
);

INVX1 _7676_ (
    .A(_645_),
    .Y(_654_)
);

AOI21X1 _7677_ (
    .A(_638_),
    .B(_648_),
    .C(_654_),
    .Y(_655_)
);

NAND2X1 _7678_ (
    .A(_172__bF$buf2),
    .B(_643_),
    .Y(_656_)
);

NOR2X1 _7679_ (
    .A(_413_),
    .B(_656_),
    .Y(_657_)
);

AOI21X1 _7680_ (
    .A(_643_),
    .B(_172__bF$buf1),
    .C(_414_),
    .Y(_658_)
);

NOR2X1 _7681_ (
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

AND2X2 _7682_ (
    .A(_655_),
    .B(_659_),
    .Y(_660_)
);

OAI21X1 _7683_ (
    .A(_659_),
    .B(_655_),
    .C(_156_),
    .Y(_661_)
);

OAI21X1 _7684_ (
    .A(_661_),
    .B(_660_),
    .C(_653_),
    .Y(_24_)
);

OAI21X1 _7685_ (
    .A(1'h0),
    .B(_135__bF$buf0),
    .C(_154_),
    .Y(_662_)
);

OAI21X1 _7686_ (
    .A(_429_),
    .B(_662_),
    .C(\genblk1[0].u_ce.Ain0 [0]),
    .Y(_663_)
);

INVX1 _7687_ (
    .A(\genblk1[0].u_ce.Ain0 [0]),
    .Y(_664_)
);

NOR2X1 _7688_ (
    .A(_429_),
    .B(_662_),
    .Y(_665_)
);

NAND2X1 _7689_ (
    .A(_664_),
    .B(_665_),
    .Y(_666_)
);

NAND2X1 _7690_ (
    .A(_663_),
    .B(_666_),
    .Y(_667_)
);

NAND2X1 _7691_ (
    .A(\genblk1[0].u_ce.Acalc [0]),
    .B(_158__bF$buf4),
    .Y(_668_)
);

OAI21X1 _7692_ (
    .A(_158__bF$buf3),
    .B(_667_),
    .C(_668_),
    .Y(_25_)
);

NAND2X1 _7693_ (
    .A(\genblk1[0].u_ce.Acalc [1]),
    .B(_158__bF$buf2),
    .Y(_669_)
);

INVX1 _7694_ (
    .A(_663_),
    .Y(_670_)
);

NOR2X1 _7695_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_671_)
);

AOI21X1 _7696_ (
    .A(_429_),
    .B(1'h0),
    .C(_671_),
    .Y(_672_)
);

NOR2X1 _7697_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_672_),
    .Y(_673_)
);

OAI21X1 _7698_ (
    .A(_429_),
    .B(_662_),
    .C(_172__bF$buf0),
    .Y(_674_)
);

AND2X2 _7699_ (
    .A(_674_),
    .B(_672_),
    .Y(_675_)
);

OR2X2 _7700_ (
    .A(_675_),
    .B(_673_),
    .Y(_676_)
);

OR2X2 _7701_ (
    .A(_676_),
    .B(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_677_)
);

OAI21X1 _7702_ (
    .A(_673_),
    .B(_675_),
    .C(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_678_)
);

NAND2X1 _7703_ (
    .A(_678_),
    .B(_677_),
    .Y(_679_)
);

NOR2X1 _7704_ (
    .A(_670_),
    .B(_679_),
    .Y(_680_)
);

NAND2X1 _7705_ (
    .A(_670_),
    .B(_679_),
    .Y(_681_)
);

NAND2X1 _7706_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .B(_681_),
    .Y(_682_)
);

OAI21X1 _7707_ (
    .A(_680_),
    .B(_682_),
    .C(_669_),
    .Y(_26_)
);

INVX1 _7708_ (
    .A(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_683_)
);

OAI21X1 _7709_ (
    .A(_683_),
    .B(_676_),
    .C(_681_),
    .Y(_684_)
);

OAI21X1 _7710_ (
    .A(_164_),
    .B(_135__bF$buf4),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_685_)
);

OAI21X1 _7711_ (
    .A(1'h0),
    .B(1'h0),
    .C(1'h0),
    .Y(_686_)
);

MUX2X1 _7712_ (
    .A(_686_),
    .B(1'h0),
    .S(_685_),
    .Y(_687_)
);

NAND2X1 _7713_ (
    .A(\genblk1[0].u_ce.Ain1 [0]),
    .B(_687_),
    .Y(_688_)
);

OR2X2 _7714_ (
    .A(_687_),
    .B(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_689_)
);

NAND2X1 _7715_ (
    .A(_688_),
    .B(_689_),
    .Y(_690_)
);

INVX1 _7716_ (
    .A(_690_),
    .Y(_691_)
);

NOR2X1 _7717_ (
    .A(_691_),
    .B(_684_),
    .Y(_692_)
);

NAND2X1 _7718_ (
    .A(_691_),
    .B(_684_),
    .Y(_693_)
);

NAND2X1 _7719_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_693_),
    .Y(_694_)
);

OAI22X1 _7720_ (
    .A(_80_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_692_),
    .D(_694_),
    .Y(_27_)
);

NOR2X1 _7721_ (
    .A(\genblk1[0].u_ce.Acalc [3]),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_695_)
);

NAND2X1 _7722_ (
    .A(_688_),
    .B(_693_),
    .Y(_696_)
);

INVX1 _7723_ (
    .A(_696_),
    .Y(_697_)
);

INVX1 _7724_ (
    .A(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_698_)
);

NOR2X1 _7725_ (
    .A(1'h0),
    .B(_135__bF$buf3),
    .Y(_699_)
);

OAI21X1 _7726_ (
    .A(_134__bF$buf1),
    .B(_699_),
    .C(_172__bF$buf5),
    .Y(_700_)
);

OAI21X1 _7727_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_701_)
);

OAI21X1 _7728_ (
    .A(_164_),
    .B(_701_),
    .C(_700_),
    .Y(_702_)
);

NOR2X1 _7729_ (
    .A(_698_),
    .B(_702_),
    .Y(_703_)
);

NAND2X1 _7730_ (
    .A(_698_),
    .B(_702_),
    .Y(_704_)
);

INVX1 _7731_ (
    .A(_704_),
    .Y(_705_)
);

NOR2X1 _7732_ (
    .A(_703_),
    .B(_705_),
    .Y(_706_)
);

OAI21X1 _7733_ (
    .A(_706_),
    .B(_697_),
    .C(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .Y(_707_)
);

AOI21X1 _7734_ (
    .A(_697_),
    .B(_706_),
    .C(_707_),
    .Y(_708_)
);

NOR2X1 _7735_ (
    .A(_695_),
    .B(_708_),
    .Y(_28_)
);

NAND2X1 _7736_ (
    .A(\genblk1[0].u_ce.Acalc [4]),
    .B(_158__bF$buf1),
    .Y(_709_)
);

INVX1 _7737_ (
    .A(\genblk1[0].u_ce.Ain12b [4]),
    .Y(_710_)
);

AOI21X1 _7738_ (
    .A(_429_),
    .B(1'h0),
    .C(_172__bF$buf4),
    .Y(_711_)
);

OAI21X1 _7739_ (
    .A(1'h0),
    .B(_429_),
    .C(_711_),
    .Y(_712_)
);

OAI21X1 _7740_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_672_),
    .C(_712_),
    .Y(_713_)
);

OR2X2 _7741_ (
    .A(_713_),
    .B(_710_),
    .Y(_714_)
);

NAND2X1 _7742_ (
    .A(_710_),
    .B(_713_),
    .Y(_715_)
);

NAND2X1 _7743_ (
    .A(_715_),
    .B(_714_),
    .Y(_716_)
);

AOI21X1 _7744_ (
    .A(_696_),
    .B(_704_),
    .C(_703_),
    .Y(_717_)
);

AND2X2 _7745_ (
    .A(_717_),
    .B(_716_),
    .Y(_718_)
);

OAI21X1 _7746_ (
    .A(_716_),
    .B(_717_),
    .C(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Y(_719_)
);

OAI21X1 _7747_ (
    .A(_719_),
    .B(_718_),
    .C(_709_),
    .Y(_29_)
);

OAI21X1 _7748_ (
    .A(_716_),
    .B(_717_),
    .C(_714_),
    .Y(_720_)
);

INVX1 _7749_ (
    .A(\genblk1[0].u_ce.Ain12b [5]),
    .Y(_721_)
);

OAI21X1 _7750_ (
    .A(_428_),
    .B(_241_),
    .C(_172__bF$buf3),
    .Y(_722_)
);

OAI21X1 _7751_ (
    .A(1'h0),
    .B(1'h0),
    .C(_154_),
    .Y(_723_)
);

OR2X2 _7752_ (
    .A(_723_),
    .B(_172__bF$buf2),
    .Y(_724_)
);

NAND2X1 _7753_ (
    .A(_722_),
    .B(_724_),
    .Y(_725_)
);

OR2X2 _7754_ (
    .A(_725_),
    .B(_721_),
    .Y(_726_)
);

NAND2X1 _7755_ (
    .A(_721_),
    .B(_725_),
    .Y(_727_)
);

NAND2X1 _7756_ (
    .A(_727_),
    .B(_726_),
    .Y(_728_)
);

INVX1 _7757_ (
    .A(_728_),
    .Y(_729_)
);

NOR2X1 _7758_ (
    .A(_729_),
    .B(_720_),
    .Y(_730_)
);

NAND2X1 _7759_ (
    .A(_729_),
    .B(_720_),
    .Y(_731_)
);

NAND2X1 _7760_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_731_),
    .Y(_732_)
);

OAI22X1 _7761_ (
    .A(_97_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_730_),
    .D(_732_),
    .Y(_30_)
);

NAND2X1 _7762_ (
    .A(\genblk1[0].u_ce.Acalc [6]),
    .B(_158__bF$buf0),
    .Y(_733_)
);

INVX1 _7763_ (
    .A(_716_),
    .Y(_734_)
);

NAND2X1 _7764_ (
    .A(_729_),
    .B(_734_),
    .Y(_735_)
);

OAI21X1 _7765_ (
    .A(_714_),
    .B(_728_),
    .C(_726_),
    .Y(_736_)
);

INVX1 _7766_ (
    .A(_736_),
    .Y(_737_)
);

OAI21X1 _7767_ (
    .A(_735_),
    .B(_717_),
    .C(_737_),
    .Y(_738_)
);

OAI21X1 _7768_ (
    .A(1'h0),
    .B(_164_),
    .C(_134__bF$buf0),
    .Y(_739_)
);

NOR2X1 _7769_ (
    .A(_739_),
    .B(_699_),
    .Y(_740_)
);

NAND2X1 _7770_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_740_),
    .Y(_741_)
);

OAI21X1 _7771_ (
    .A(_739_),
    .B(_699_),
    .C(_172__bF$buf1),
    .Y(_742_)
);

NAND2X1 _7772_ (
    .A(_742_),
    .B(_741_),
    .Y(_743_)
);

NAND2X1 _7773_ (
    .A(\genblk1[0].u_ce.Ain12b [6]),
    .B(_743_),
    .Y(_744_)
);

OR2X2 _7774_ (
    .A(_743_),
    .B(\genblk1[0].u_ce.Ain12b [6]),
    .Y(_745_)
);

NAND2X1 _7775_ (
    .A(_744_),
    .B(_745_),
    .Y(_746_)
);

INVX1 _7776_ (
    .A(_746_),
    .Y(_747_)
);

NOR2X1 _7777_ (
    .A(_747_),
    .B(_738_),
    .Y(_748_)
);

NAND2X1 _7778_ (
    .A(_747_),
    .B(_738_),
    .Y(_749_)
);

NAND2X1 _7779_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .B(_749_),
    .Y(_750_)
);

OAI21X1 _7780_ (
    .A(_748_),
    .B(_750_),
    .C(_733_),
    .Y(_31_)
);

INVX1 _7781_ (
    .A(\genblk1[0].u_ce.Acalc [7]),
    .Y(_751_)
);

NAND2X1 _7782_ (
    .A(_744_),
    .B(_749_),
    .Y(_752_)
);

INVX1 _7783_ (
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .Y(_753_)
);

NAND2X1 _7784_ (
    .A(_172__bF$buf0),
    .B(_671_),
    .Y(_754_)
);

OR2X2 _7785_ (
    .A(_671_),
    .B(_172__bF$buf5),
    .Y(_755_)
);

NAND2X1 _7786_ (
    .A(_754_),
    .B(_755_),
    .Y(_756_)
);

NOR2X1 _7787_ (
    .A(_753_),
    .B(_756_),
    .Y(_757_)
);

INVX1 _7788_ (
    .A(_757_),
    .Y(_758_)
);

NAND2X1 _7789_ (
    .A(_753_),
    .B(_756_),
    .Y(_759_)
);

NAND2X1 _7790_ (
    .A(_759_),
    .B(_758_),
    .Y(_760_)
);

OR2X2 _7791_ (
    .A(_752_),
    .B(_760_),
    .Y(_761_)
);

AOI21X1 _7792_ (
    .A(_752_),
    .B(_760_),
    .C(_158__bF$buf4),
    .Y(_762_)
);

AOI22X1 _7793_ (
    .A(_751_),
    .B(_158__bF$buf3),
    .C(_761_),
    .D(_762_),
    .Y(_32_)
);

NAND2X1 _7794_ (
    .A(\genblk1[0].u_ce.Acalc [8]),
    .B(_158__bF$buf2),
    .Y(_763_)
);

NOR2X1 _7795_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_154_),
    .Y(_764_)
);

INVX1 _7796_ (
    .A(_764_),
    .Y(_765_)
);

NAND3X1 _7797_ (
    .A(\genblk1[0].u_ce.Ain12b [8]),
    .B(_701_),
    .C(_765_),
    .Y(_766_)
);

INVX1 _7798_ (
    .A(_766_),
    .Y(_767_)
);

AOI21X1 _7799_ (
    .A(_765_),
    .B(_701_),
    .C(\genblk1[0].u_ce.Ain12b [8]),
    .Y(_768_)
);

NOR2X1 _7800_ (
    .A(_768_),
    .B(_767_),
    .Y(_769_)
);

OAI21X1 _7801_ (
    .A(_744_),
    .B(_760_),
    .C(_758_),
    .Y(_770_)
);

NOR2X1 _7802_ (
    .A(_760_),
    .B(_746_),
    .Y(_771_)
);

AOI21X1 _7803_ (
    .A(_771_),
    .B(_736_),
    .C(_770_),
    .Y(_772_)
);

NAND3X1 _7804_ (
    .A(_734_),
    .B(_729_),
    .C(_771_),
    .Y(_773_)
);

OAI21X1 _7805_ (
    .A(_773_),
    .B(_717_),
    .C(_772_),
    .Y(_774_)
);

NOR2X1 _7806_ (
    .A(_769_),
    .B(_774_),
    .Y(_775_)
);

NAND2X1 _7807_ (
    .A(_769_),
    .B(_774_),
    .Y(_776_)
);

NAND2X1 _7808_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .B(_776_),
    .Y(_777_)
);

OAI21X1 _7809_ (
    .A(_775_),
    .B(_777_),
    .C(_763_),
    .Y(_33_)
);

AOI21X1 _7810_ (
    .A(_774_),
    .B(_769_),
    .C(_767_),
    .Y(_778_)
);

OR2X2 _7811_ (
    .A(_172__bF$buf4),
    .B(\genblk1[0].u_ce.Ain12b [9]),
    .Y(_779_)
);

NAND2X1 _7812_ (
    .A(\genblk1[0].u_ce.Ain12b [9]),
    .B(_172__bF$buf3),
    .Y(_780_)
);

NAND2X1 _7813_ (
    .A(_780_),
    .B(_779_),
    .Y(_781_)
);

AND2X2 _7814_ (
    .A(_778_),
    .B(_781_),
    .Y(_782_)
);

OAI21X1 _7815_ (
    .A(_781_),
    .B(_778_),
    .C(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Y(_783_)
);

OAI22X1 _7816_ (
    .A(_94_),
    .B(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .C(_783_),
    .D(_782_),
    .Y(_34_)
);

NAND2X1 _7817_ (
    .A(\genblk1[0].u_ce.Acalc [10]),
    .B(_158__bF$buf1),
    .Y(_784_)
);

OAI21X1 _7818_ (
    .A(_781_),
    .B(_766_),
    .C(_780_),
    .Y(_785_)
);

NAND3X1 _7819_ (
    .A(_779_),
    .B(_780_),
    .C(_769_),
    .Y(_786_)
);

INVX1 _7820_ (
    .A(_786_),
    .Y(_787_)
);

AOI21X1 _7821_ (
    .A(_774_),
    .B(_787_),
    .C(_785_),
    .Y(_788_)
);

INVX1 _7822_ (
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .Y(_789_)
);

NAND2X1 _7823_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_789_),
    .Y(_790_)
);

NAND2X1 _7824_ (
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .B(_172__bF$buf2),
    .Y(_791_)
);

NAND2X1 _7825_ (
    .A(_790_),
    .B(_791_),
    .Y(_792_)
);

AND2X2 _7826_ (
    .A(_788_),
    .B(_792_),
    .Y(_793_)
);

OAI21X1 _7827_ (
    .A(_792_),
    .B(_788_),
    .C(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .Y(_794_)
);

OAI21X1 _7828_ (
    .A(_794_),
    .B(_793_),
    .C(_784_),
    .Y(_35_)
);

NAND2X1 _7829_ (
    .A(\genblk1[0].u_ce.Acalc [11]),
    .B(_158__bF$buf0),
    .Y(_795_)
);

OAI21X1 _7830_ (
    .A(_792_),
    .B(_788_),
    .C(_791_),
    .Y(_796_)
);

OAI21X1 _7831_ (
    .A(_158__bF$buf4),
    .B(_796_),
    .C(_795_),
    .Y(_36_)
);

NAND2X1 _7832_ (
    .A(\genblk1[0].u_ce.LoadCtl [5]),
    .B(_85_),
    .Y(_797_)
);

NAND2X1 _7833_ (
    .A(_86_),
    .B(_92_),
    .Y(_798_)
);

NOR2X1 _7834_ (
    .A(_797_),
    .B(_798_),
    .Y(_799_)
);

NAND2X1 _7835_ (
    .A(1'h0),
    .B(_799_),
    .Y(_800_)
);

OAI21X1 _7836_ (
    .A(_256_),
    .B(_799_),
    .C(_800_),
    .Y(_37_)
);

NAND2X1 _7837_ (
    .A(1'h0),
    .B(_799_),
    .Y(_801_)
);

OAI21X1 _7838_ (
    .A(_324_),
    .B(_799_),
    .C(_801_),
    .Y(_38_)
);

INVX1 _7839_ (
    .A(1'h0),
    .Y(_802_)
);

OR2X2 _7840_ (
    .A(_798_),
    .B(_85_),
    .Y(_803_)
);

OAI21X1 _7841_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_804_)
);

OAI21X1 _7842_ (
    .A(_802_),
    .B(_803_),
    .C(_804_),
    .Y(_39_)
);

INVX1 _7843_ (
    .A(1'h0),
    .Y(_805_)
);

OAI21X1 _7844_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Xin12b [9]),
    .Y(_806_)
);

OAI21X1 _7845_ (
    .A(_805_),
    .B(_803_),
    .C(_806_),
    .Y(_40_)
);

NAND2X1 _7846_ (
    .A(_92_),
    .B(_89_),
    .Y(_807_)
);

NAND2X1 _7847_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(_807_),
    .Y(_808_)
);

OAI21X1 _7848_ (
    .A(_802_),
    .B(_807_),
    .C(_808_),
    .Y(_41_)
);

NAND2X1 _7849_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(_807_),
    .Y(_809_)
);

OAI21X1 _7850_ (
    .A(_805_),
    .B(_807_),
    .C(_809_),
    .Y(_42_)
);

AND2X2 _7851_ (
    .A(_92_),
    .B(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_810_)
);

NAND2X1 _7852_ (
    .A(1'h0),
    .B(_810_),
    .Y(_811_)
);

OAI21X1 _7853_ (
    .A(_139_),
    .B(_810_),
    .C(_811_),
    .Y(_43_)
);

NAND2X1 _7854_ (
    .A(1'h0),
    .B(_810_),
    .Y(_812_)
);

OAI21X1 _7855_ (
    .A(_176_),
    .B(_810_),
    .C(_812_),
    .Y(_44_)
);

OAI21X1 _7856_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_813_)
);

OAI21X1 _7857_ (
    .A(_802_),
    .B(_83_),
    .C(_813_),
    .Y(_45_)
);

OAI21X1 _7858_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_814_)
);

OAI21X1 _7859_ (
    .A(_805_),
    .B(_83_),
    .C(_814_),
    .Y(_46_)
);

NAND2X1 _7860_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(1'h0),
    .Y(_815_)
);

OAI21X1 _7861_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_146_),
    .C(_815_),
    .Y(_47_)
);

NAND2X1 _7862_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(1'h0),
    .Y(_816_)
);

OAI21X1 _7863_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_183_),
    .C(_816_),
    .Y(_48_)
);

NAND2X1 _7864_ (
    .A(1'h0),
    .B(_799_),
    .Y(_817_)
);

OAI21X1 _7865_ (
    .A(_385_),
    .B(_799_),
    .C(_817_),
    .Y(_49_)
);

NAND2X1 _7866_ (
    .A(1'h0),
    .B(_799_),
    .Y(_818_)
);

OAI21X1 _7867_ (
    .A(_411_),
    .B(_799_),
    .C(_818_),
    .Y(_50_)
);

INVX1 _7868_ (
    .A(1'h0),
    .Y(_819_)
);

OAI21X1 _7869_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_820_)
);

OAI21X1 _7870_ (
    .A(_819_),
    .B(_803_),
    .C(_820_),
    .Y(_51_)
);

INVX1 _7871_ (
    .A(1'h0),
    .Y(_821_)
);

OAI21X1 _7872_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_822_)
);

OAI21X1 _7873_ (
    .A(_821_),
    .B(_803_),
    .C(_822_),
    .Y(_52_)
);

NAND2X1 _7874_ (
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .B(_807_),
    .Y(_823_)
);

OAI21X1 _7875_ (
    .A(_819_),
    .B(_807_),
    .C(_823_),
    .Y(_53_)
);

NAND2X1 _7876_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(_807_),
    .Y(_824_)
);

OAI21X1 _7877_ (
    .A(_821_),
    .B(_807_),
    .C(_824_),
    .Y(_54_)
);

NAND2X1 _7878_ (
    .A(1'h0),
    .B(_810_),
    .Y(_825_)
);

OAI21X1 _7879_ (
    .A(_255_),
    .B(_810_),
    .C(_825_),
    .Y(_55_)
);

NAND2X1 _7880_ (
    .A(1'h0),
    .B(_810_),
    .Y(_826_)
);

OAI21X1 _7881_ (
    .A(_276_),
    .B(_810_),
    .C(_826_),
    .Y(_56_)
);

OAI21X1 _7882_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_827_)
);

OAI21X1 _7883_ (
    .A(_819_),
    .B(_83_),
    .C(_827_),
    .Y(_57_)
);

OAI21X1 _7884_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_828_)
);

OAI21X1 _7885_ (
    .A(_821_),
    .B(_83_),
    .C(_828_),
    .Y(_58_)
);

NAND2X1 _7886_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(1'h0),
    .Y(_829_)
);

OAI21X1 _7887_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_133_),
    .C(_829_),
    .Y(_59_)
);

NAND2X1 _7888_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(1'h0),
    .Y(_830_)
);

OAI21X1 _7889_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_171_),
    .C(_830_),
    .Y(_60_)
);

NAND2X1 _7890_ (
    .A(\a[0] [0]),
    .B(_799_),
    .Y(_831_)
);

OAI21X1 _7891_ (
    .A(_789_),
    .B(_799_),
    .C(_831_),
    .Y(_61_)
);

NAND2X1 _7892_ (
    .A(\a[0] [1]),
    .B(_799_),
    .Y(_832_)
);

OAI21X1 _7893_ (
    .A(_172__bF$buf1),
    .B(_799_),
    .C(_832_),
    .Y(_62_)
);

INVX1 _7894_ (
    .A(\a[0] [0]),
    .Y(_833_)
);

OAI21X1 _7895_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Ain12b [8]),
    .Y(_834_)
);

OAI21X1 _7896_ (
    .A(_833_),
    .B(_803_),
    .C(_834_),
    .Y(_63_)
);

INVX1 _7897_ (
    .A(\a[0] [1]),
    .Y(_835_)
);

OAI21X1 _7898_ (
    .A(_85_),
    .B(_798_),
    .C(\genblk1[0].u_ce.Ain12b [9]),
    .Y(_836_)
);

OAI21X1 _7899_ (
    .A(_835_),
    .B(_803_),
    .C(_836_),
    .Y(_64_)
);

NAND2X1 _7900_ (
    .A(\genblk1[0].u_ce.Ain12b [6]),
    .B(_807_),
    .Y(_837_)
);

OAI21X1 _7901_ (
    .A(_833_),
    .B(_807_),
    .C(_837_),
    .Y(_65_)
);

NAND2X1 _7902_ (
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .B(_807_),
    .Y(_73_)
);

OAI21X1 _7903_ (
    .A(_835_),
    .B(_807_),
    .C(_73_),
    .Y(_66_)
);

NAND2X1 _7904_ (
    .A(\a[0] [0]),
    .B(_810_),
    .Y(_74_)
);

OAI21X1 _7905_ (
    .A(_710_),
    .B(_810_),
    .C(_74_),
    .Y(_67_)
);

NAND2X1 _7906_ (
    .A(\a[0] [1]),
    .B(_810_),
    .Y(_75_)
);

OAI21X1 _7907_ (
    .A(_721_),
    .B(_810_),
    .C(_75_),
    .Y(_68_)
);

OAI21X1 _7908_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_76_)
);

OAI21X1 _7909_ (
    .A(_833_),
    .B(_83_),
    .C(_76_),
    .Y(_69_)
);

OAI21X1 _7910_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_81_),
    .C(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_77_)
);

OAI21X1 _7911_ (
    .A(_835_),
    .B(_83_),
    .C(_77_),
    .Y(_70_)
);

NAND2X1 _7912_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[0] [0]),
    .Y(_78_)
);

OAI21X1 _7913_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_664_),
    .C(_78_),
    .Y(_71_)
);

NAND2X1 _7914_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[0] [1]),
    .Y(_79_)
);

OAI21X1 _7915_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_683_),
    .C(_79_),
    .Y(_72_)
);

DFFPOSX1 _7916_ (
    .CLK(clk_bF$buf7),
    .D(_0_),
    .Q(\genblk1[0].u_ce.Ycalc [0])
);

DFFPOSX1 _7917_ (
    .CLK(clk_bF$buf6),
    .D(_1_),
    .Q(\genblk1[0].u_ce.Ycalc [1])
);

DFFPOSX1 _7918_ (
    .CLK(clk_bF$buf5),
    .D(_2_),
    .Q(\genblk1[0].u_ce.ISout )
);

DFFPOSX1 _7919_ (
    .CLK(clk_bF$buf4),
    .D(_3_),
    .Q(\genblk1[0].u_ce.Ycalc [2])
);

DFFPOSX1 _7920_ (
    .CLK(clk_bF$buf3),
    .D(_4_),
    .Q(\genblk1[0].u_ce.Ycalc [3])
);

DFFPOSX1 _7921_ (
    .CLK(clk_bF$buf2),
    .D(_5_),
    .Q(\genblk1[0].u_ce.Ycalc [4])
);

DFFPOSX1 _7922_ (
    .CLK(clk_bF$buf1),
    .D(_6_),
    .Q(\genblk1[0].u_ce.Ycalc [5])
);

DFFPOSX1 _7923_ (
    .CLK(clk_bF$buf0),
    .D(_7_),
    .Q(\genblk1[0].u_ce.Ycalc [6])
);

DFFPOSX1 _7924_ (
    .CLK(clk_bF$buf78),
    .D(_8_),
    .Q(\genblk1[0].u_ce.Ycalc [7])
);

DFFPOSX1 _7925_ (
    .CLK(clk_bF$buf77),
    .D(_9_),
    .Q(\genblk1[0].u_ce.Ycalc [8])
);

DFFPOSX1 _7926_ (
    .CLK(clk_bF$buf76),
    .D(_10_),
    .Q(\genblk1[0].u_ce.Ycalc [9])
);

DFFPOSX1 _7927_ (
    .CLK(clk_bF$buf75),
    .D(_11_),
    .Q(\genblk1[0].u_ce.Ycalc [10])
);

DFFPOSX1 _7928_ (
    .CLK(clk_bF$buf74),
    .D(_12_),
    .Q(\genblk1[0].u_ce.Ycalc [11])
);

DFFPOSX1 _7929_ (
    .CLK(clk_bF$buf73),
    .D(_13_),
    .Q(\genblk1[0].u_ce.Xcalc [0])
);

DFFPOSX1 _7930_ (
    .CLK(clk_bF$buf72),
    .D(_14_),
    .Q(\genblk1[0].u_ce.Xcalc [1])
);

DFFPOSX1 _7931_ (
    .CLK(clk_bF$buf71),
    .D(_15_),
    .Q(\genblk1[0].u_ce.Xcalc [2])
);

DFFPOSX1 _7932_ (
    .CLK(clk_bF$buf70),
    .D(_16_),
    .Q(\genblk1[0].u_ce.Xcalc [3])
);

DFFPOSX1 _7933_ (
    .CLK(clk_bF$buf69),
    .D(_17_),
    .Q(\genblk1[0].u_ce.Xcalc [4])
);

DFFPOSX1 _7934_ (
    .CLK(clk_bF$buf68),
    .D(_18_),
    .Q(\genblk1[0].u_ce.Xcalc [5])
);

DFFPOSX1 _7935_ (
    .CLK(clk_bF$buf67),
    .D(_19_),
    .Q(\genblk1[0].u_ce.Xcalc [6])
);

DFFPOSX1 _7936_ (
    .CLK(clk_bF$buf66),
    .D(_20_),
    .Q(\genblk1[0].u_ce.Xcalc [7])
);

DFFPOSX1 _7937_ (
    .CLK(clk_bF$buf65),
    .D(_21_),
    .Q(\genblk1[0].u_ce.Xcalc [8])
);

DFFPOSX1 _7938_ (
    .CLK(clk_bF$buf64),
    .D(_22_),
    .Q(\genblk1[0].u_ce.Xcalc [9])
);

DFFPOSX1 _7939_ (
    .CLK(clk_bF$buf63),
    .D(_23_),
    .Q(\genblk1[0].u_ce.Xcalc [10])
);

DFFPOSX1 _7940_ (
    .CLK(clk_bF$buf62),
    .D(_24_),
    .Q(\genblk1[0].u_ce.Xcalc [11])
);

DFFPOSX1 _7941_ (
    .CLK(clk_bF$buf61),
    .D(_25_),
    .Q(\genblk1[0].u_ce.Acalc [0])
);

DFFPOSX1 _7942_ (
    .CLK(clk_bF$buf60),
    .D(_26_),
    .Q(\genblk1[0].u_ce.Acalc [1])
);

DFFPOSX1 _7943_ (
    .CLK(clk_bF$buf59),
    .D(_27_),
    .Q(\genblk1[0].u_ce.Acalc [2])
);

DFFPOSX1 _7944_ (
    .CLK(clk_bF$buf58),
    .D(_28_),
    .Q(\genblk1[0].u_ce.Acalc [3])
);

DFFPOSX1 _7945_ (
    .CLK(clk_bF$buf57),
    .D(_29_),
    .Q(\genblk1[0].u_ce.Acalc [4])
);

DFFPOSX1 _7946_ (
    .CLK(clk_bF$buf56),
    .D(_30_),
    .Q(\genblk1[0].u_ce.Acalc [5])
);

DFFPOSX1 _7947_ (
    .CLK(clk_bF$buf55),
    .D(_31_),
    .Q(\genblk1[0].u_ce.Acalc [6])
);

DFFPOSX1 _7948_ (
    .CLK(clk_bF$buf54),
    .D(_32_),
    .Q(\genblk1[0].u_ce.Acalc [7])
);

DFFPOSX1 _7949_ (
    .CLK(clk_bF$buf53),
    .D(_33_),
    .Q(\genblk1[0].u_ce.Acalc [8])
);

DFFPOSX1 _7950_ (
    .CLK(clk_bF$buf52),
    .D(_34_),
    .Q(\genblk1[0].u_ce.Acalc [9])
);

DFFPOSX1 _7951_ (
    .CLK(clk_bF$buf51),
    .D(_35_),
    .Q(\genblk1[0].u_ce.Acalc [10])
);

DFFPOSX1 _7952_ (
    .CLK(clk_bF$buf50),
    .D(_36_),
    .Q(\genblk1[0].u_ce.Acalc [11])
);

DFFPOSX1 _7953_ (
    .CLK(clk_bF$buf49),
    .D(_37_),
    .Q(\genblk1[0].u_ce.Xin12b [10])
);

DFFPOSX1 _7954_ (
    .CLK(clk_bF$buf48),
    .D(_38_),
    .Q(\genblk1[0].u_ce.Xin12b [11])
);

DFFPOSX1 _7955_ (
    .CLK(clk_bF$buf47),
    .D(_39_),
    .Q(\genblk1[0].u_ce.Xin12b [8])
);

DFFPOSX1 _7956_ (
    .CLK(clk_bF$buf46),
    .D(_40_),
    .Q(\genblk1[0].u_ce.Xin12b [9])
);

DFFPOSX1 _7957_ (
    .CLK(clk_bF$buf45),
    .D(_41_),
    .Q(\genblk1[0].u_ce.Xin12b [6])
);

DFFPOSX1 _7958_ (
    .CLK(clk_bF$buf44),
    .D(_42_),
    .Q(\genblk1[0].u_ce.Xin12b [7])
);

DFFPOSX1 _7959_ (
    .CLK(clk_bF$buf43),
    .D(_43_),
    .Q(\genblk1[0].u_ce.Xin12b [4])
);

DFFPOSX1 _7960_ (
    .CLK(clk_bF$buf42),
    .D(_44_),
    .Q(\genblk1[0].u_ce.Xin12b [5])
);

DFFPOSX1 _7961_ (
    .CLK(clk_bF$buf41),
    .D(_45_),
    .Q(\genblk1[0].u_ce.Xin1 [0])
);

DFFPOSX1 _7962_ (
    .CLK(clk_bF$buf40),
    .D(_46_),
    .Q(\genblk1[0].u_ce.Xin1 [1])
);

DFFPOSX1 _7963_ (
    .CLK(clk_bF$buf39),
    .D(_47_),
    .Q(\genblk1[0].u_ce.Xin0 [0])
);

DFFPOSX1 _7964_ (
    .CLK(clk_bF$buf38),
    .D(_48_),
    .Q(\genblk1[0].u_ce.Xin0 [1])
);

DFFPOSX1 _7965_ (
    .CLK(clk_bF$buf37),
    .D(_49_),
    .Q(\genblk1[0].u_ce.Yin12b [10])
);

DFFPOSX1 _7966_ (
    .CLK(clk_bF$buf36),
    .D(_50_),
    .Q(\genblk1[0].u_ce.Yin12b [11])
);

DFFPOSX1 _7967_ (
    .CLK(clk_bF$buf35),
    .D(_51_),
    .Q(\genblk1[0].u_ce.Yin12b [8])
);

DFFPOSX1 _7968_ (
    .CLK(clk_bF$buf34),
    .D(_52_),
    .Q(\genblk1[0].u_ce.Yin12b [9])
);

DFFPOSX1 _7969_ (
    .CLK(clk_bF$buf33),
    .D(_53_),
    .Q(\genblk1[0].u_ce.Yin12b [6])
);

DFFPOSX1 _7970_ (
    .CLK(clk_bF$buf32),
    .D(_54_),
    .Q(\genblk1[0].u_ce.Yin12b [7])
);

DFFPOSX1 _7971_ (
    .CLK(clk_bF$buf31),
    .D(_55_),
    .Q(\genblk1[0].u_ce.Yin12b [4])
);

DFFPOSX1 _7972_ (
    .CLK(clk_bF$buf30),
    .D(_56_),
    .Q(\genblk1[0].u_ce.Yin12b [5])
);

DFFPOSX1 _7973_ (
    .CLK(clk_bF$buf29),
    .D(_57_),
    .Q(\genblk1[0].u_ce.Yin1 [0])
);

DFFPOSX1 _7974_ (
    .CLK(clk_bF$buf28),
    .D(_58_),
    .Q(\genblk1[0].u_ce.Yin1 [1])
);

DFFPOSX1 _7975_ (
    .CLK(clk_bF$buf27),
    .D(_59_),
    .Q(\genblk1[0].u_ce.Yin0 [0])
);

DFFPOSX1 _7976_ (
    .CLK(clk_bF$buf26),
    .D(_60_),
    .Q(\genblk1[0].u_ce.Yin0 [1])
);

DFFPOSX1 _7977_ (
    .CLK(clk_bF$buf25),
    .D(_61_),
    .Q(\genblk1[0].u_ce.Ain12b [10])
);

DFFPOSX1 _7978_ (
    .CLK(clk_bF$buf24),
    .D(_62_),
    .Q(\genblk1[0].u_ce.Ain12b [11])
);

DFFPOSX1 _7979_ (
    .CLK(clk_bF$buf23),
    .D(_63_),
    .Q(\genblk1[0].u_ce.Ain12b [8])
);

DFFPOSX1 _7980_ (
    .CLK(clk_bF$buf22),
    .D(_64_),
    .Q(\genblk1[0].u_ce.Ain12b [9])
);

DFFPOSX1 _7981_ (
    .CLK(clk_bF$buf21),
    .D(_65_),
    .Q(\genblk1[0].u_ce.Ain12b [6])
);

DFFPOSX1 _7982_ (
    .CLK(clk_bF$buf20),
    .D(_66_),
    .Q(\genblk1[0].u_ce.Ain12b [7])
);

DFFPOSX1 _7983_ (
    .CLK(clk_bF$buf19),
    .D(_67_),
    .Q(\genblk1[0].u_ce.Ain12b [4])
);

DFFPOSX1 _7984_ (
    .CLK(clk_bF$buf18),
    .D(_68_),
    .Q(\genblk1[0].u_ce.Ain12b [5])
);

DFFPOSX1 _7985_ (
    .CLK(clk_bF$buf17),
    .D(_69_),
    .Q(\genblk1[0].u_ce.Ain1 [0])
);

DFFPOSX1 _7986_ (
    .CLK(clk_bF$buf16),
    .D(_70_),
    .Q(\genblk1[0].u_ce.Ain1 [1])
);

DFFPOSX1 _7987_ (
    .CLK(clk_bF$buf15),
    .D(_71_),
    .Q(\genblk1[0].u_ce.Ain0 [0])
);

DFFPOSX1 _7988_ (
    .CLK(clk_bF$buf14),
    .D(_72_),
    .Q(\genblk1[0].u_ce.Ain0 [1])
);

DFFPOSX1 _7989_ (
    .CLK(clk_bF$buf13),
    .D(\genblk1[0].u_ce.Rdy_bF$buf3 ),
    .Q(\genblk1[0].u_ce.LoadCtl [0])
);

DFFPOSX1 _7990_ (
    .CLK(clk_bF$buf12),
    .D(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[0].u_ce.LoadCtl [1])
);

DFFPOSX1 _7991_ (
    .CLK(clk_bF$buf11),
    .D(\genblk1[0].u_ce.LoadCtl [1]),
    .Q(\genblk1[0].u_ce.LoadCtl [2])
);

DFFPOSX1 _7992_ (
    .CLK(clk_bF$buf10),
    .D(\genblk1[0].u_ce.LoadCtl [2]),
    .Q(\genblk1[0].u_ce.LoadCtl [3])
);

DFFPOSX1 _7993_ (
    .CLK(clk_bF$buf9),
    .D(\genblk1[0].u_ce.LoadCtl [3]),
    .Q(\genblk1[0].u_ce.LoadCtl [4])
);

DFFPOSX1 _7994_ (
    .CLK(clk_bF$buf8),
    .D(\genblk1[0].u_ce.LoadCtl [4]),
    .Q(\genblk1[0].u_ce.LoadCtl [5])
);

DFFPOSX1 _7995_ (
    .CLK(clk_bF$buf7),
    .D(\genblk1[0].u_ce.LoadCtl [5]),
    .Q(\genblk1[0].u_ce.Vld )
);

INVX1 _7996_ (
    .A(\genblk1[1].u_ce.Acalc [2]),
    .Y(_918_)
);

INVX2 _7997_ (
    .A(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_919_)
);

NOR2X1 _7998_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_919_),
    .Y(_920_)
);

INVX2 _7999_ (
    .A(_920_),
    .Y(_921_)
);

NOR2X1 _8000_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [10]),
    .Y(_922_)
);

INVX4 _8001_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .Y(_923_)
);

NOR2X1 _8002_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.LoadCtl [3]),
    .Y(_924_)
);

OAI21X1 _8003_ (
    .A(_923_),
    .B(\genblk1[1].u_ce.Acalc [8]),
    .C(_924_),
    .Y(_925_)
);

INVX2 _8004_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_926_)
);

AND2X2 _8005_ (
    .A(_926_),
    .B(\genblk1[1].u_ce.LoadCtl [3]),
    .Y(_927_)
);

AOI22X1 _8006_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.Acalc [4]),
    .C(_927_),
    .D(\genblk1[1].u_ce.Acalc [6]),
    .Y(_928_)
);

OAI21X1 _8007_ (
    .A(_922_),
    .B(_925_),
    .C(_928_),
    .Y(_929_)
);

NOR2X1 _8008_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_930_)
);

AOI22X1 _8009_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.Acalc [0]),
    .C(_929_),
    .D(_930_),
    .Y(_931_)
);

OAI21X1 _8010_ (
    .A(_918_),
    .B(_921_),
    .C(_931_),
    .Y(\a[2] [0])
);

INVX1 _8011_ (
    .A(\genblk1[1].u_ce.Acalc [9]),
    .Y(_932_)
);

OAI21X1 _8012_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [11]),
    .C(_924_),
    .Y(_933_)
);

AOI21X1 _8013_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_932_),
    .C(_933_),
    .Y(_934_)
);

INVX1 _8014_ (
    .A(\genblk1[1].u_ce.Acalc [5]),
    .Y(_935_)
);

NAND2X1 _8015_ (
    .A(\genblk1[1].u_ce.Acalc [7]),
    .B(_927_),
    .Y(_936_)
);

OAI21X1 _8016_ (
    .A(_926_),
    .B(_935_),
    .C(_936_),
    .Y(_937_)
);

OAI21X1 _8017_ (
    .A(_934_),
    .B(_937_),
    .C(_930_),
    .Y(_938_)
);

AOI22X1 _8018_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Acalc [1]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Acalc [3]),
    .Y(_939_)
);

NAND2X1 _8019_ (
    .A(_939_),
    .B(_938_),
    .Y(\a[2] [1])
);

INVX1 _8020_ (
    .A(\genblk1[1].u_ce.Ycalc [10]),
    .Y(_940_)
);

OAI21X1 _8021_ (
    .A(_923_),
    .B(\genblk1[1].u_ce.Ycalc [8]),
    .C(_924_),
    .Y(_941_)
);

AOI21X1 _8022_ (
    .A(_923_),
    .B(_940_),
    .C(_941_),
    .Y(_942_)
);

INVX1 _8023_ (
    .A(\genblk1[1].u_ce.Ycalc [4]),
    .Y(_943_)
);

NAND2X1 _8024_ (
    .A(\genblk1[1].u_ce.Ycalc [6]),
    .B(_927_),
    .Y(_944_)
);

OAI21X1 _8025_ (
    .A(_926_),
    .B(_943_),
    .C(_944_),
    .Y(_945_)
);

OAI21X1 _8026_ (
    .A(_942_),
    .B(_945_),
    .C(_930_),
    .Y(_946_)
);

AOI22X1 _8027_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.Ycalc [0]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Ycalc [2]),
    .Y(_947_)
);

NAND2X1 _8028_ (
    .A(_947_),
    .B(_946_),
    .Y(\genblk1[1].u_ce.Y_ [0])
);

INVX1 _8029_ (
    .A(\genblk1[1].u_ce.Ycalc [9]),
    .Y(_948_)
);

OAI21X1 _8030_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Ycalc [11]),
    .C(_924_),
    .Y(_949_)
);

AOI21X1 _8031_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_948_),
    .C(_949_),
    .Y(_950_)
);

INVX1 _8032_ (
    .A(\genblk1[1].u_ce.Ycalc [5]),
    .Y(_951_)
);

NAND2X1 _8033_ (
    .A(\genblk1[1].u_ce.Ycalc [7]),
    .B(_927_),
    .Y(_952_)
);

OAI21X1 _8034_ (
    .A(_926_),
    .B(_951_),
    .C(_952_),
    .Y(_953_)
);

OAI21X1 _8035_ (
    .A(_950_),
    .B(_953_),
    .C(_930_),
    .Y(_954_)
);

AOI22X1 _8036_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[1].u_ce.Ycalc [1]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_955_)
);

NAND2X1 _8037_ (
    .A(_955_),
    .B(_954_),
    .Y(\genblk1[1].u_ce.Y_ [1])
);

INVX1 _8038_ (
    .A(\genblk1[1].u_ce.Xcalc [8]),
    .Y(_956_)
);

OAI21X1 _8039_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Xcalc [10]),
    .C(_924_),
    .Y(_957_)
);

AOI21X1 _8040_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_956_),
    .C(_957_),
    .Y(_958_)
);

INVX1 _8041_ (
    .A(\genblk1[1].u_ce.Xcalc [4]),
    .Y(_959_)
);

NAND2X1 _8042_ (
    .A(\genblk1[1].u_ce.Xcalc [6]),
    .B(_927_),
    .Y(_960_)
);

OAI21X1 _8043_ (
    .A(_926_),
    .B(_959_),
    .C(_960_),
    .Y(_961_)
);

OAI21X1 _8044_ (
    .A(_958_),
    .B(_961_),
    .C(_930_),
    .Y(_962_)
);

AOI22X1 _8045_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.Xcalc [0]),
    .C(_920_),
    .D(\genblk1[1].u_ce.Xcalc [2]),
    .Y(_963_)
);

NAND2X1 _8046_ (
    .A(_963_),
    .B(_962_),
    .Y(\genblk1[1].u_ce.X_ [0])
);

INVX1 _8047_ (
    .A(\genblk1[1].u_ce.Xcalc [3]),
    .Y(_964_)
);

NOR2X1 _8048_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Xcalc [11]),
    .Y(_965_)
);

OAI21X1 _8049_ (
    .A(_923_),
    .B(\genblk1[1].u_ce.Xcalc [9]),
    .C(_924_),
    .Y(_966_)
);

AOI22X1 _8050_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.Xcalc [5]),
    .C(_927_),
    .D(\genblk1[1].u_ce.Xcalc [7]),
    .Y(_967_)
);

OAI21X1 _8051_ (
    .A(_965_),
    .B(_966_),
    .C(_967_),
    .Y(_968_)
);

AOI22X1 _8052_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.Xcalc [1]),
    .C(_968_),
    .D(_930_),
    .Y(_969_)
);

OAI21X1 _8053_ (
    .A(_964_),
    .B(_921_),
    .C(_969_),
    .Y(\genblk1[1].u_ce.X_ [1])
);

INVX1 _8054_ (
    .A(\genblk1[1].u_ce.Ycalc [0]),
    .Y(_970_)
);

INVX1 _8055_ (
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .Y(_971_)
);

INVX8 _8056_ (
    .A(1'h0),
    .Y(_972_)
);

INVX8 _8057_ (
    .A(1'h0),
    .Y(_973_)
);

INVX1 _8058_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_974_)
);

NAND2X1 _8059_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_975_)
);

OAI21X1 _8060_ (
    .A(1'h1),
    .B(_974_),
    .C(_975_),
    .Y(_976_)
);

INVX1 _8061_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .Y(_977_)
);

NAND2X1 _8062_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_978_)
);

OAI21X1 _8063_ (
    .A(1'h1),
    .B(_977_),
    .C(_978_),
    .Y(_979_)
);

MUX2X1 _8064_ (
    .A(_979_),
    .B(_976_),
    .S(_973__bF$buf4),
    .Y(_980_)
);

INVX1 _8065_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_981_)
);

NAND2X1 _8066_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_982_)
);

OAI21X1 _8067_ (
    .A(1'h1),
    .B(_981_),
    .C(_982_),
    .Y(_983_)
);

INVX1 _8068_ (
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .Y(_984_)
);

NAND2X1 _8069_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_985_)
);

OAI21X1 _8070_ (
    .A(1'h1),
    .B(_984_),
    .C(_985_),
    .Y(_986_)
);

MUX2X1 _8071_ (
    .A(_986_),
    .B(_983_),
    .S(_973__bF$buf3),
    .Y(_987_)
);

MUX2X1 _8072_ (
    .A(_987_),
    .B(_980_),
    .S(_972__bF$buf4),
    .Y(_988_)
);

NOR2X1 _8073_ (
    .A(_971_),
    .B(_988_),
    .Y(_989_)
);

NAND2X1 _8074_ (
    .A(_971_),
    .B(_988_),
    .Y(_990_)
);

INVX1 _8075_ (
    .A(_990_),
    .Y(_991_)
);

NAND2X1 _8076_ (
    .A(_972__bF$buf3),
    .B(_973__bF$buf2),
    .Y(_992_)
);

OAI21X1 _8077_ (
    .A(1'h1),
    .B(_992_),
    .C(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .Y(_993_)
);

INVX2 _8078_ (
    .A(_993_),
    .Y(_994_)
);

OAI21X1 _8079_ (
    .A(_989_),
    .B(_991_),
    .C(_994_),
    .Y(_995_)
);

OAI21X1 _8080_ (
    .A(_970_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_995_),
    .Y(_838_)
);

INVX8 _8081_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_996_)
);

NAND2X1 _8082_ (
    .A(\genblk1[1].u_ce.Ycalc [1]),
    .B(_996__bF$buf4),
    .Y(_997_)
);

NOR2X1 _8083_ (
    .A(1'h1),
    .B(_992_),
    .Y(_998_)
);

MUX2X1 _8084_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(\genblk1[1].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_999_)
);

MUX2X1 _8085_ (
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .B(\genblk1[1].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_1000_)
);

MUX2X1 _8086_ (
    .A(_1000_),
    .B(_999_),
    .S(_973__bF$buf1),
    .Y(_1001_)
);

INVX2 _8087_ (
    .A(1'h1),
    .Y(_1002_)
);

NAND2X1 _8088_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(_1002_),
    .Y(_1003_)
);

AOI21X1 _8089_ (
    .A(_1003_),
    .B(_982_),
    .C(_973__bF$buf0),
    .Y(_1004_)
);

NAND3X1 _8090_ (
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .B(_1002_),
    .C(_973__bF$buf4),
    .Y(_1005_)
);

NAND3X1 _8091_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(1'h1),
    .C(_973__bF$buf3),
    .Y(_1006_)
);

NAND3X1 _8092_ (
    .A(_972__bF$buf2),
    .B(_1006_),
    .C(_1005_),
    .Y(_1007_)
);

OAI22X1 _8093_ (
    .A(_1004_),
    .B(_1007_),
    .C(_972__bF$buf1),
    .D(_1001_),
    .Y(_1008_)
);

INVX1 _8094_ (
    .A(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1009_)
);

INVX8 _8095_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1010_)
);

INVX1 _8096_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1011_)
);

NAND2X1 _8097_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1012_)
);

OAI21X1 _8098_ (
    .A(1'h1),
    .B(_1011_),
    .C(_1012_),
    .Y(_1013_)
);

INVX1 _8099_ (
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_1014_)
);

NAND2X1 _8100_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_1015_)
);

OAI21X1 _8101_ (
    .A(1'h1),
    .B(_1014_),
    .C(_1015_),
    .Y(_1016_)
);

MUX2X1 _8102_ (
    .A(_1016_),
    .B(_1013_),
    .S(_973__bF$buf2),
    .Y(_1017_)
);

INVX1 _8103_ (
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1018_)
);

NAND2X1 _8104_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [4]),
    .Y(_1019_)
);

OAI21X1 _8105_ (
    .A(1'h1),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_)
);

INVX1 _8106_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .Y(_1021_)
);

NAND2X1 _8107_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1022_)
);

OAI21X1 _8108_ (
    .A(1'h1),
    .B(_1021_),
    .C(_1022_),
    .Y(_1023_)
);

MUX2X1 _8109_ (
    .A(_1023_),
    .B(_1020_),
    .S(_973__bF$buf1),
    .Y(_1024_)
);

MUX2X1 _8110_ (
    .A(_1024_),
    .B(_1017_),
    .S(_972__bF$buf0),
    .Y(_1025_)
);

NAND3X1 _8111_ (
    .A(_1010__bF$buf5),
    .B(_988_),
    .C(_1025_),
    .Y(_1026_)
);

MUX2X1 _8112_ (
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_1027_)
);

MUX2X1 _8113_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_1028_)
);

MUX2X1 _8114_ (
    .A(_1028_),
    .B(_1027_),
    .S(_973__bF$buf0),
    .Y(_1029_)
);

MUX2X1 _8115_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_1030_)
);

MUX2X1 _8116_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(\genblk1[1].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_1031_)
);

MUX2X1 _8117_ (
    .A(_1031_),
    .B(_1030_),
    .S(_973__bF$buf4),
    .Y(_1032_)
);

MUX2X1 _8118_ (
    .A(_1032_),
    .B(_1029_),
    .S(_972__bF$buf4),
    .Y(_1033_)
);

OAI21X1 _8119_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1008_),
    .C(_1033_),
    .Y(_1034_)
);

AOI21X1 _8120_ (
    .A(_1034_),
    .B(_1026_),
    .C(_1009_),
    .Y(_1035_)
);

INVX1 _8121_ (
    .A(_1035_),
    .Y(_1036_)
);

NAND3X1 _8122_ (
    .A(_1009_),
    .B(_1026_),
    .C(_1034_),
    .Y(_1037_)
);

AND2X2 _8123_ (
    .A(_1036_),
    .B(_1037_),
    .Y(_1038_)
);

OAI21X1 _8124_ (
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .B(_1008_),
    .C(_1038_),
    .Y(_1039_)
);

OR2X2 _8125_ (
    .A(_1038_),
    .B(_990_),
    .Y(_1040_)
);

AOI21X1 _8126_ (
    .A(_1040_),
    .B(_1039_),
    .C(_998_),
    .Y(_1041_)
);

OAI21X1 _8127_ (
    .A(_996__bF$buf3),
    .B(_1041_),
    .C(_997_),
    .Y(_839_)
);

INVX1 _8128_ (
    .A(\genblk1[1].u_ce.ISout ),
    .Y(_1042_)
);

NAND2X1 _8129_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .B(\genblk1[0].u_ce.ISout ),
    .Y(_1043_)
);

OAI21X1 _8130_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .B(_1042_),
    .C(_1043_),
    .Y(_840_)
);

NAND2X1 _8131_ (
    .A(\genblk1[1].u_ce.Ycalc [2]),
    .B(_996__bF$buf2),
    .Y(_1044_)
);

AOI21X1 _8132_ (
    .A(_990_),
    .B(_1037_),
    .C(_1035_),
    .Y(_1045_)
);

MUX2X1 _8133_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(\genblk1[1].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_1046_)
);

MUX2X1 _8134_ (
    .A(_1046_),
    .B(_999_),
    .S(1'h0),
    .Y(_1047_)
);

MUX2X1 _8135_ (
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_1048_)
);

NAND2X1 _8136_ (
    .A(1'h0),
    .B(_972__bF$buf3),
    .Y(_1049_)
);

OAI22X1 _8137_ (
    .A(_1049_),
    .B(_1000_),
    .C(_1048_),
    .D(_992_),
    .Y(_1050_)
);

AOI21X1 _8138_ (
    .A(1'h0),
    .B(_1047_),
    .C(_1050_),
    .Y(_1051_)
);

AOI21X1 _8139_ (
    .A(_1033_),
    .B(_1008_),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_1052_)
);

NAND2X1 _8140_ (
    .A(_1051_),
    .B(_1052_),
    .Y(_1053_)
);

INVX1 _8141_ (
    .A(_1051_),
    .Y(_1054_)
);

OAI21X1 _8142_ (
    .A(_988_),
    .B(_1025_),
    .C(_1010__bF$buf4),
    .Y(_1055_)
);

NAND2X1 _8143_ (
    .A(_1054_),
    .B(_1055_),
    .Y(_1056_)
);

AOI21X1 _8144_ (
    .A(_1056_),
    .B(_1053_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1057_)
);

NAND3X1 _8145_ (
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .B(_1053_),
    .C(_1056_),
    .Y(_1058_)
);

INVX1 _8146_ (
    .A(_1058_),
    .Y(_1059_)
);

OR2X2 _8147_ (
    .A(_1059_),
    .B(_1057_),
    .Y(_1060_)
);

NOR2X1 _8148_ (
    .A(_1045_),
    .B(_1060_),
    .Y(_1061_)
);

INVX1 _8149_ (
    .A(_1061_),
    .Y(_1062_)
);

OAI21X1 _8150_ (
    .A(_1057_),
    .B(_1059_),
    .C(_1045_),
    .Y(_1063_)
);

AOI21X1 _8151_ (
    .A(_1062_),
    .B(_1063_),
    .C(_998_),
    .Y(_1064_)
);

INVX2 _8152_ (
    .A(_998_),
    .Y(_1065_)
);

OAI21X1 _8153_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1065_),
    .C(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .Y(_1066_)
);

OAI21X1 _8154_ (
    .A(_1066_),
    .B(_1064_),
    .C(_1044_),
    .Y(_841_)
);

INVX1 _8155_ (
    .A(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_1067_)
);

INVX2 _8156_ (
    .A(_1066_),
    .Y(_1068_)
);

OAI21X1 _8157_ (
    .A(_1057_),
    .B(_1045_),
    .C(_1058_),
    .Y(_1069_)
);

INVX1 _8158_ (
    .A(_1069_),
    .Y(_1070_)
);

INVX1 _8159_ (
    .A(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1071_)
);

NAND3X1 _8160_ (
    .A(_1008_),
    .B(_1033_),
    .C(_1051_),
    .Y(_1072_)
);

INVX1 _8161_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .Y(_1073_)
);

NAND2X1 _8162_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1074_)
);

OAI21X1 _8163_ (
    .A(1'h1),
    .B(_1073_),
    .C(_1074_),
    .Y(_1075_)
);

NAND2X1 _8164_ (
    .A(_973__bF$buf3),
    .B(_1027_),
    .Y(_1076_)
);

OAI21X1 _8165_ (
    .A(_973__bF$buf2),
    .B(_1075_),
    .C(_1076_),
    .Y(_1077_)
);

NOR2X1 _8166_ (
    .A(1'h0),
    .B(_973__bF$buf1),
    .Y(_1078_)
);

NOR2X1 _8167_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_1079_)
);

AOI22X1 _8168_ (
    .A(_1020_),
    .B(_1079_),
    .C(_1078_),
    .D(_1016_),
    .Y(_1080_)
);

OAI21X1 _8169_ (
    .A(_972__bF$buf2),
    .B(_1077_),
    .C(_1080_),
    .Y(_1081_)
);

NAND3X1 _8170_ (
    .A(_1010__bF$buf3),
    .B(_1081_),
    .C(_1072_),
    .Y(_1082_)
);

INVX1 _8171_ (
    .A(_1072_),
    .Y(_1083_)
);

INVX1 _8172_ (
    .A(_1081_),
    .Y(_1084_)
);

OAI21X1 _8173_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1083_),
    .C(_1084_),
    .Y(_1085_)
);

NAND3X1 _8174_ (
    .A(_1071_),
    .B(_1082_),
    .C(_1085_),
    .Y(_1086_)
);

AOI21X1 _8175_ (
    .A(_1085_),
    .B(_1082_),
    .C(_1071_),
    .Y(_1087_)
);

INVX1 _8176_ (
    .A(_1087_),
    .Y(_1088_)
);

NAND2X1 _8177_ (
    .A(_1086_),
    .B(_1088_),
    .Y(_1089_)
);

AOI21X1 _8178_ (
    .A(_1089_),
    .B(_1070_),
    .C(_998_),
    .Y(_1090_)
);

OAI21X1 _8179_ (
    .A(_1070_),
    .B(_1089_),
    .C(_1090_),
    .Y(_1091_)
);

AOI22X1 _8180_ (
    .A(_1067_),
    .B(_996__bF$buf1),
    .C(_1091_),
    .D(_1068_),
    .Y(_842_)
);

AOI21X1 _8181_ (
    .A(_1069_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1092_)
);

INVX1 _8182_ (
    .A(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1093_)
);

INVX1 _8183_ (
    .A(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1094_)
);

NAND2X1 _8184_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1095_)
);

OAI21X1 _8185_ (
    .A(1'h1),
    .B(_1094_),
    .C(_1095_),
    .Y(_1096_)
);

NAND2X1 _8186_ (
    .A(_973__bF$buf0),
    .B(_1046_),
    .Y(_1097_)
);

OAI21X1 _8187_ (
    .A(_973__bF$buf4),
    .B(_1096_),
    .C(_1097_),
    .Y(_1098_)
);

NAND2X1 _8188_ (
    .A(_972__bF$buf1),
    .B(_1001_),
    .Y(_1099_)
);

OAI21X1 _8189_ (
    .A(_972__bF$buf0),
    .B(_1098_),
    .C(_1099_),
    .Y(_1100_)
);

INVX2 _8190_ (
    .A(_1100_),
    .Y(_1101_)
);

OAI21X1 _8191_ (
    .A(_1081_),
    .B(_1072_),
    .C(_1010__bF$buf2),
    .Y(_1102_)
);

OR2X2 _8192_ (
    .A(_1102_),
    .B(_1101_),
    .Y(_1103_)
);

NOR2X1 _8193_ (
    .A(_1081_),
    .B(_1072_),
    .Y(_1104_)
);

OAI21X1 _8194_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1104_),
    .C(_1101_),
    .Y(_1105_)
);

NAND3X1 _8195_ (
    .A(_1093_),
    .B(_1105_),
    .C(_1103_),
    .Y(_1106_)
);

NOR2X1 _8196_ (
    .A(_1101_),
    .B(_1102_),
    .Y(_1107_)
);

AND2X2 _8197_ (
    .A(_1102_),
    .B(_1101_),
    .Y(_1108_)
);

OAI21X1 _8198_ (
    .A(_1107_),
    .B(_1108_),
    .C(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1109_)
);

NAND2X1 _8199_ (
    .A(_1109_),
    .B(_1106_),
    .Y(_1110_)
);

AOI21X1 _8200_ (
    .A(_1092_),
    .B(_1110_),
    .C(_998_),
    .Y(_1111_)
);

OAI21X1 _8201_ (
    .A(_1092_),
    .B(_1110_),
    .C(_1111_),
    .Y(_1112_)
);

AOI22X1 _8202_ (
    .A(_943_),
    .B(_996__bF$buf0),
    .C(_1112_),
    .D(_1068_),
    .Y(_843_)
);

OAI21X1 _8203_ (
    .A(_1110_),
    .B(_1092_),
    .C(_1109_),
    .Y(_1113_)
);

INVX1 _8204_ (
    .A(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1114_)
);

NAND3X1 _8205_ (
    .A(_1084_),
    .B(_1101_),
    .C(_1083_),
    .Y(_1115_)
);

NAND2X1 _8206_ (
    .A(1'h0),
    .B(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1116_)
);

INVX1 _8207_ (
    .A(_1116_),
    .Y(_1117_)
);

AOI21X1 _8208_ (
    .A(_1075_),
    .B(_973__bF$buf3),
    .C(_1117_),
    .Y(_1118_)
);

NAND2X1 _8209_ (
    .A(_972__bF$buf4),
    .B(_1029_),
    .Y(_1119_)
);

OAI21X1 _8210_ (
    .A(_972__bF$buf3),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_)
);

NAND3X1 _8211_ (
    .A(_1010__bF$buf1),
    .B(_1120_),
    .C(_1115_),
    .Y(_1121_)
);

NOR3X1 _8212_ (
    .A(_1081_),
    .B(_1100_),
    .C(_1072_),
    .Y(_1122_)
);

INVX1 _8213_ (
    .A(_1120_),
    .Y(_1123_)
);

OAI21X1 _8214_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1122_),
    .C(_1123_),
    .Y(_1124_)
);

NAND3X1 _8215_ (
    .A(_1114_),
    .B(_1121_),
    .C(_1124_),
    .Y(_1125_)
);

AOI21X1 _8216_ (
    .A(_1124_),
    .B(_1121_),
    .C(_1114_),
    .Y(_1126_)
);

INVX1 _8217_ (
    .A(_1126_),
    .Y(_1127_)
);

NAND2X1 _8218_ (
    .A(_1125_),
    .B(_1127_),
    .Y(_1128_)
);

AND2X2 _8219_ (
    .A(_1113_),
    .B(_1128_),
    .Y(_1129_)
);

OAI21X1 _8220_ (
    .A(_1128_),
    .B(_1113_),
    .C(_1065_),
    .Y(_1130_)
);

OAI21X1 _8221_ (
    .A(_1130_),
    .B(_1129_),
    .C(_1068_),
    .Y(_1131_)
);

OAI21X1 _8222_ (
    .A(_951_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_1131_),
    .Y(_844_)
);

INVX1 _8223_ (
    .A(\genblk1[1].u_ce.Ycalc [6]),
    .Y(_1132_)
);

INVX1 _8224_ (
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1133_)
);

NAND3X1 _8225_ (
    .A(_1101_),
    .B(_1123_),
    .C(_1104_),
    .Y(_1134_)
);

AOI21X1 _8226_ (
    .A(_1096_),
    .B(_973__bF$buf2),
    .C(_1117_),
    .Y(_1135_)
);

NAND2X1 _8227_ (
    .A(_972__bF$buf2),
    .B(_1047_),
    .Y(_1136_)
);

OAI21X1 _8228_ (
    .A(_972__bF$buf1),
    .B(_1135_),
    .C(_1136_),
    .Y(_1137_)
);

NAND3X1 _8229_ (
    .A(_1010__bF$buf0),
    .B(_1137_),
    .C(_1134_),
    .Y(_1138_)
);

INVX1 _8230_ (
    .A(_1137_),
    .Y(_1139_)
);

OAI21X1 _8231_ (
    .A(_1120_),
    .B(_1115_),
    .C(_1010__bF$buf5),
    .Y(_1140_)
);

NAND2X1 _8232_ (
    .A(_1139_),
    .B(_1140_),
    .Y(_1141_)
);

NAND3X1 _8233_ (
    .A(_1133_),
    .B(_1138_),
    .C(_1141_),
    .Y(_1142_)
);

NAND3X1 _8234_ (
    .A(_1010__bF$buf4),
    .B(_1139_),
    .C(_1134_),
    .Y(_1143_)
);

NAND2X1 _8235_ (
    .A(_1137_),
    .B(_1140_),
    .Y(_1144_)
);

NAND3X1 _8236_ (
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .B(_1143_),
    .C(_1144_),
    .Y(_1145_)
);

NAND2X1 _8237_ (
    .A(_1142_),
    .B(_1145_),
    .Y(_1146_)
);

AOI21X1 _8238_ (
    .A(_1103_),
    .B(_1105_),
    .C(_1093_),
    .Y(_1147_)
);

NOR2X1 _8239_ (
    .A(_1147_),
    .B(_1126_),
    .Y(_1148_)
);

OAI21X1 _8240_ (
    .A(_1110_),
    .B(_1092_),
    .C(_1148_),
    .Y(_1149_)
);

NAND2X1 _8241_ (
    .A(_1125_),
    .B(_1149_),
    .Y(_1150_)
);

AOI21X1 _8242_ (
    .A(_1150_),
    .B(_1146_),
    .C(_998_),
    .Y(_1151_)
);

OAI21X1 _8243_ (
    .A(_1146_),
    .B(_1150_),
    .C(_1151_),
    .Y(_1152_)
);

AOI22X1 _8244_ (
    .A(_1132_),
    .B(_996__bF$buf4),
    .C(_1152_),
    .D(_1068_),
    .Y(_845_)
);

INVX1 _8245_ (
    .A(\genblk1[1].u_ce.Ycalc [7]),
    .Y(_1153_)
);

AOI21X1 _8246_ (
    .A(_1141_),
    .B(_1138_),
    .C(_1133_),
    .Y(_1154_)
);

AND2X2 _8247_ (
    .A(_1106_),
    .B(_1109_),
    .Y(_1155_)
);

NAND3X1 _8248_ (
    .A(_1125_),
    .B(_1127_),
    .C(_1155_),
    .Y(_1156_)
);

AOI21X1 _8249_ (
    .A(_1147_),
    .B(_1125_),
    .C(_1126_),
    .Y(_1157_)
);

OAI21X1 _8250_ (
    .A(_1092_),
    .B(_1156_),
    .C(_1157_),
    .Y(_1158_)
);

AOI21X1 _8251_ (
    .A(_1158_),
    .B(_1142_),
    .C(_1154_),
    .Y(_1159_)
);

INVX1 _8252_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1160_)
);

NAND3X1 _8253_ (
    .A(_1123_),
    .B(_1139_),
    .C(_1122_),
    .Y(_1161_)
);

INVX1 _8254_ (
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1162_)
);

NOR2X1 _8255_ (
    .A(_972__bF$buf0),
    .B(_1162_),
    .Y(_1163_)
);

INVX1 _8256_ (
    .A(_1163_),
    .Y(_1164_)
);

OAI21X1 _8257_ (
    .A(1'h0),
    .B(_1077_),
    .C(_1164_),
    .Y(_1165_)
);

NAND3X1 _8258_ (
    .A(_1010__bF$buf3),
    .B(_1165_),
    .C(_1161_),
    .Y(_1166_)
);

INVX1 _8259_ (
    .A(_1165_),
    .Y(_1167_)
);

OAI21X1 _8260_ (
    .A(_1137_),
    .B(_1134_),
    .C(_1010__bF$buf2),
    .Y(_1168_)
);

NAND2X1 _8261_ (
    .A(_1167_),
    .B(_1168_),
    .Y(_1169_)
);

NAND3X1 _8262_ (
    .A(_1160_),
    .B(_1166_),
    .C(_1169_),
    .Y(_1170_)
);

NAND3X1 _8263_ (
    .A(_1010__bF$buf1),
    .B(_1167_),
    .C(_1161_),
    .Y(_1171_)
);

NAND2X1 _8264_ (
    .A(_1165_),
    .B(_1168_),
    .Y(_1172_)
);

NAND3X1 _8265_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(_1171_),
    .C(_1172_),
    .Y(_1173_)
);

NAND2X1 _8266_ (
    .A(_1170_),
    .B(_1173_),
    .Y(_1174_)
);

INVX1 _8267_ (
    .A(_1174_),
    .Y(_1175_)
);

NOR2X1 _8268_ (
    .A(_1175_),
    .B(_1159_),
    .Y(_1176_)
);

OAI21X1 _8269_ (
    .A(_1146_),
    .B(_1150_),
    .C(_1145_),
    .Y(_1177_)
);

OAI21X1 _8270_ (
    .A(_1174_),
    .B(_1177_),
    .C(_1065_),
    .Y(_1178_)
);

OAI21X1 _8271_ (
    .A(_1010__bF$buf0),
    .B(_1065_),
    .C(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_1179_)
);

INVX1 _8272_ (
    .A(_1179_),
    .Y(_1180_)
);

OAI21X1 _8273_ (
    .A(_1178_),
    .B(_1176_),
    .C(_1180_),
    .Y(_1181_)
);

OAI21X1 _8274_ (
    .A(_1153_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1181_),
    .Y(_846_)
);

INVX1 _8275_ (
    .A(\genblk1[1].u_ce.Ycalc [8]),
    .Y(_1182_)
);

OAI21X1 _8276_ (
    .A(_1145_),
    .B(_1174_),
    .C(_1173_),
    .Y(_1183_)
);

NOR2X1 _8277_ (
    .A(_1146_),
    .B(_1174_),
    .Y(_1184_)
);

AOI21X1 _8278_ (
    .A(_1184_),
    .B(_1158_),
    .C(_1183_),
    .Y(_1185_)
);

INVX1 _8279_ (
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1186_)
);

OR2X2 _8280_ (
    .A(_1161_),
    .B(_1165_),
    .Y(_1187_)
);

OAI21X1 _8281_ (
    .A(1'h0),
    .B(_1098_),
    .C(_1164_),
    .Y(_1188_)
);

NAND3X1 _8282_ (
    .A(_1010__bF$buf5),
    .B(_1188_),
    .C(_1187_),
    .Y(_1189_)
);

NOR2X1 _8283_ (
    .A(_1165_),
    .B(_1161_),
    .Y(_1190_)
);

INVX1 _8284_ (
    .A(_1188_),
    .Y(_1191_)
);

OAI21X1 _8285_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_)
);

NAND3X1 _8286_ (
    .A(_1186_),
    .B(_1192_),
    .C(_1189_),
    .Y(_1193_)
);

NAND3X1 _8287_ (
    .A(_1010__bF$buf4),
    .B(_1191_),
    .C(_1187_),
    .Y(_1194_)
);

OAI21X1 _8288_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1190_),
    .C(_1188_),
    .Y(_1195_)
);

NAND3X1 _8289_ (
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .B(_1195_),
    .C(_1194_),
    .Y(_1196_)
);

AND2X2 _8290_ (
    .A(_1193_),
    .B(_1196_),
    .Y(_1197_)
);

INVX1 _8291_ (
    .A(_1197_),
    .Y(_1198_)
);

AOI21X1 _8292_ (
    .A(_1185_),
    .B(_1198_),
    .C(_998_),
    .Y(_1199_)
);

OAI21X1 _8293_ (
    .A(_1185_),
    .B(_1198_),
    .C(_1199_),
    .Y(_1200_)
);

AOI22X1 _8294_ (
    .A(_1182_),
    .B(_996__bF$buf3),
    .C(_1200_),
    .D(_1180_),
    .Y(_847_)
);

NAND2X1 _8295_ (
    .A(_1154_),
    .B(_1170_),
    .Y(_1201_)
);

AND2X2 _8296_ (
    .A(_1201_),
    .B(_1173_),
    .Y(_1202_)
);

AND2X2 _8297_ (
    .A(_1142_),
    .B(_1145_),
    .Y(_1203_)
);

NAND3X1 _8298_ (
    .A(_1170_),
    .B(_1173_),
    .C(_1203_),
    .Y(_1204_)
);

OAI21X1 _8299_ (
    .A(_1150_),
    .B(_1204_),
    .C(_1202_),
    .Y(_1205_)
);

INVX1 _8300_ (
    .A(_1196_),
    .Y(_1206_)
);

AOI21X1 _8301_ (
    .A(_1205_),
    .B(_1193_),
    .C(_1206_),
    .Y(_1207_)
);

INVX1 _8302_ (
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1208_)
);

NOR3X1 _8303_ (
    .A(_1165_),
    .B(_1188_),
    .C(_1161_),
    .Y(_1209_)
);

INVX1 _8304_ (
    .A(_1209_),
    .Y(_1210_)
);

OAI21X1 _8305_ (
    .A(1'h0),
    .B(_1118_),
    .C(_1164_),
    .Y(_1211_)
);

NAND3X1 _8306_ (
    .A(_1010__bF$buf3),
    .B(_1211_),
    .C(_1210_),
    .Y(_1212_)
);

INVX1 _8307_ (
    .A(_1211_),
    .Y(_1213_)
);

OAI21X1 _8308_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1209_),
    .C(_1213_),
    .Y(_1214_)
);

NAND3X1 _8309_ (
    .A(_1208_),
    .B(_1214_),
    .C(_1212_),
    .Y(_1215_)
);

NAND3X1 _8310_ (
    .A(_1010__bF$buf2),
    .B(_1213_),
    .C(_1210_),
    .Y(_1216_)
);

OAI21X1 _8311_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1209_),
    .C(_1211_),
    .Y(_1217_)
);

NAND3X1 _8312_ (
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .B(_1217_),
    .C(_1216_),
    .Y(_1218_)
);

AND2X2 _8313_ (
    .A(_1215_),
    .B(_1218_),
    .Y(_1219_)
);

AND2X2 _8314_ (
    .A(_1207_),
    .B(_1219_),
    .Y(_1220_)
);

OAI21X1 _8315_ (
    .A(_1219_),
    .B(_1207_),
    .C(_1065_),
    .Y(_1221_)
);

OAI21X1 _8316_ (
    .A(_1221_),
    .B(_1220_),
    .C(_1068_),
    .Y(_1222_)
);

OAI21X1 _8317_ (
    .A(_948_),
    .B(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .C(_1222_),
    .Y(_848_)
);

INVX1 _8318_ (
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .Y(_1223_)
);

OAI21X1 _8319_ (
    .A(1'h0),
    .B(_1135_),
    .C(_1164_),
    .Y(_1224_)
);

INVX1 _8320_ (
    .A(_1224_),
    .Y(_1225_)
);

AOI21X1 _8321_ (
    .A(_1209_),
    .B(_1213_),
    .C(_1225_),
    .Y(_1226_)
);

NAND3X1 _8322_ (
    .A(_1213_),
    .B(_1225_),
    .C(_1209_),
    .Y(_1227_)
);

NAND2X1 _8323_ (
    .A(_1010__bF$buf1),
    .B(_1227_),
    .Y(_1228_)
);

NAND2X1 _8324_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1224_),
    .Y(_1229_)
);

OAI21X1 _8325_ (
    .A(_1226_),
    .B(_1228_),
    .C(_1229_),
    .Y(_1230_)
);

NAND2X1 _8326_ (
    .A(_1223_),
    .B(_1230_),
    .Y(_1231_)
);

INVX1 _8327_ (
    .A(_1226_),
    .Y(_1232_)
);

AND2X2 _8328_ (
    .A(_1227_),
    .B(_1010__bF$buf0),
    .Y(_1233_)
);

NAND2X1 _8329_ (
    .A(_1232_),
    .B(_1233_),
    .Y(_1234_)
);

NAND3X1 _8330_ (
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .B(_1229_),
    .C(_1234_),
    .Y(_1235_)
);

NAND2X1 _8331_ (
    .A(_1231_),
    .B(_1235_),
    .Y(_1236_)
);

AOI21X1 _8332_ (
    .A(_1212_),
    .B(_1214_),
    .C(_1208_),
    .Y(_1237_)
);

AOI21X1 _8333_ (
    .A(_1206_),
    .B(_1215_),
    .C(_1237_),
    .Y(_1238_)
);

NAND3X1 _8334_ (
    .A(_1197_),
    .B(_1219_),
    .C(_1205_),
    .Y(_1239_)
);

AOI21X1 _8335_ (
    .A(_1239_),
    .B(_1238_),
    .C(_1236_),
    .Y(_1240_)
);

AND2X2 _8336_ (
    .A(_1235_),
    .B(_1231_),
    .Y(_1241_)
);

NAND3X1 _8337_ (
    .A(_1215_),
    .B(_1218_),
    .C(_1197_),
    .Y(_1242_)
);

OAI21X1 _8338_ (
    .A(_1242_),
    .B(_1185_),
    .C(_1238_),
    .Y(_1243_)
);

OAI21X1 _8339_ (
    .A(_1241_),
    .B(_1243_),
    .C(_1065_),
    .Y(_1244_)
);

OR2X2 _8340_ (
    .A(_1244_),
    .B(_1240_),
    .Y(_1245_)
);

AOI22X1 _8341_ (
    .A(_940_),
    .B(_996__bF$buf2),
    .C(_1245_),
    .D(_1068_),
    .Y(_849_)
);

NAND2X1 _8342_ (
    .A(\genblk1[1].u_ce.Ycalc [11]),
    .B(_996__bF$buf1),
    .Y(_1246_)
);

INVX1 _8343_ (
    .A(_1235_),
    .Y(_1247_)
);

NAND2X1 _8344_ (
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .B(_1162_),
    .Y(_1248_)
);

INVX1 _8345_ (
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1249_)
);

NAND2X1 _8346_ (
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .B(_1249_),
    .Y(_1250_)
);

NAND2X1 _8347_ (
    .A(_1248_),
    .B(_1250_),
    .Y(_1251_)
);

INVX1 _8348_ (
    .A(_1251_),
    .Y(_1252_)
);

NAND2X1 _8349_ (
    .A(_1252_),
    .B(_1228_),
    .Y(_1253_)
);

NAND2X1 _8350_ (
    .A(_1251_),
    .B(_1233_),
    .Y(_1254_)
);

NAND2X1 _8351_ (
    .A(_1253_),
    .B(_1254_),
    .Y(_1255_)
);

INVX1 _8352_ (
    .A(_1255_),
    .Y(_1256_)
);

NOR3X1 _8353_ (
    .A(_1247_),
    .B(_1256_),
    .C(_1240_),
    .Y(_1257_)
);

AOI21X1 _8354_ (
    .A(_1243_),
    .B(_1241_),
    .C(_1247_),
    .Y(_1258_)
);

OAI21X1 _8355_ (
    .A(_1255_),
    .B(_1258_),
    .C(_1065_),
    .Y(_1259_)
);

OAI21X1 _8356_ (
    .A(_1257_),
    .B(_1259_),
    .C(_1068_),
    .Y(_1260_)
);

NAND2X1 _8357_ (
    .A(_1246_),
    .B(_1260_),
    .Y(_850_)
);

NAND2X1 _8358_ (
    .A(\genblk1[1].u_ce.Xcalc [0]),
    .B(_996__bF$buf0),
    .Y(_1261_)
);

INVX1 _8359_ (
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1262_)
);

NAND2X1 _8360_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1263_)
);

OAI21X1 _8361_ (
    .A(1'h1),
    .B(_1262_),
    .C(_1263_),
    .Y(_1264_)
);

NAND2X1 _8362_ (
    .A(1'h0),
    .B(_1264_),
    .Y(_1265_)
);

NOR2X1 _8363_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_1266_)
);

NOR2X1 _8364_ (
    .A(1'h0),
    .B(_1002_),
    .Y(_1267_)
);

AOI22X1 _8365_ (
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .B(_1266_),
    .C(_1267_),
    .D(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1268_)
);

NAND3X1 _8366_ (
    .A(_972__bF$buf4),
    .B(_1265_),
    .C(_1268_),
    .Y(_1269_)
);

NAND2X1 _8367_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1270_)
);

OAI21X1 _8368_ (
    .A(1'h1),
    .B(_1133_),
    .C(_1270_),
    .Y(_1271_)
);

NAND2X1 _8369_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1272_)
);

OAI21X1 _8370_ (
    .A(1'h1),
    .B(_1093_),
    .C(_1272_),
    .Y(_1273_)
);

MUX2X1 _8371_ (
    .A(_1273_),
    .B(_1271_),
    .S(_973__bF$buf1),
    .Y(_1274_)
);

NAND2X1 _8372_ (
    .A(1'h0),
    .B(_1274_),
    .Y(_1275_)
);

AND2X2 _8373_ (
    .A(_1269_),
    .B(_1275_),
    .Y(_1276_)
);

NOR2X1 _8374_ (
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .B(_1276_),
    .Y(_1277_)
);

NAND2X1 _8375_ (
    .A(_973__bF$buf0),
    .B(_1273_),
    .Y(_1278_)
);

NAND2X1 _8376_ (
    .A(1'h0),
    .B(_1271_),
    .Y(_1279_)
);

NAND2X1 _8377_ (
    .A(_1278_),
    .B(_1279_),
    .Y(_1280_)
);

OAI21X1 _8378_ (
    .A(_972__bF$buf3),
    .B(_1280_),
    .C(_1269_),
    .Y(_1281_)
);

OAI21X1 _8379_ (
    .A(_984_),
    .B(_1281_),
    .C(_994_),
    .Y(_1282_)
);

OAI21X1 _8380_ (
    .A(_1282_),
    .B(_1277_),
    .C(_1261_),
    .Y(_851_)
);

NAND2X1 _8381_ (
    .A(\genblk1[1].u_ce.Xcalc [1]),
    .B(_996__bF$buf4),
    .Y(_1283_)
);

NOR2X1 _8382_ (
    .A(_984_),
    .B(_1281_),
    .Y(_1284_)
);

NAND2X1 _8383_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1285_)
);

OAI21X1 _8384_ (
    .A(1'h1),
    .B(_1071_),
    .C(_1285_),
    .Y(_1286_)
);

NAND2X1 _8385_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1287_)
);

OAI21X1 _8386_ (
    .A(1'h1),
    .B(_1009_),
    .C(_1287_),
    .Y(_1288_)
);

MUX2X1 _8387_ (
    .A(_1288_),
    .B(_1286_),
    .S(_973__bF$buf4),
    .Y(_1289_)
);

NAND2X1 _8388_ (
    .A(_972__bF$buf2),
    .B(_1289_),
    .Y(_1290_)
);

NAND2X1 _8389_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1291_)
);

OAI21X1 _8390_ (
    .A(1'h1),
    .B(_1160_),
    .C(_1291_),
    .Y(_1292_)
);

INVX1 _8391_ (
    .A(_1292_),
    .Y(_1293_)
);

NAND2X1 _8392_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1294_)
);

OAI21X1 _8393_ (
    .A(1'h1),
    .B(_1114_),
    .C(_1294_),
    .Y(_1295_)
);

NAND2X1 _8394_ (
    .A(_973__bF$buf3),
    .B(_1295_),
    .Y(_1296_)
);

OAI21X1 _8395_ (
    .A(_973__bF$buf2),
    .B(_1293_),
    .C(_1296_),
    .Y(_1297_)
);

OAI21X1 _8396_ (
    .A(_972__bF$buf1),
    .B(_1297_),
    .C(_1290_),
    .Y(_1298_)
);

NAND3X1 _8397_ (
    .A(_1010__bF$buf5),
    .B(_1298_),
    .C(_1276_),
    .Y(_1299_)
);

MUX2X1 _8398_ (
    .A(_1295_),
    .B(_1292_),
    .S(_973__bF$buf1),
    .Y(_1300_)
);

MUX2X1 _8399_ (
    .A(_1300_),
    .B(_1289_),
    .S(1'h0),
    .Y(_1301_)
);

OAI21X1 _8400_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1281_),
    .C(_1301_),
    .Y(_1302_)
);

AOI21X1 _8401_ (
    .A(_1299_),
    .B(_1302_),
    .C(_1021_),
    .Y(_1303_)
);

INVX1 _8402_ (
    .A(_1303_),
    .Y(_1304_)
);

NAND3X1 _8403_ (
    .A(_1021_),
    .B(_1302_),
    .C(_1299_),
    .Y(_1305_)
);

AND2X2 _8404_ (
    .A(_1304_),
    .B(_1305_),
    .Y(_1306_)
);

NAND2X1 _8405_ (
    .A(_1284_),
    .B(_1306_),
    .Y(_1307_)
);

OR2X2 _8406_ (
    .A(_1306_),
    .B(_1284_),
    .Y(_1308_)
);

AOI21X1 _8407_ (
    .A(_1308_),
    .B(_1307_),
    .C(_998_),
    .Y(_1309_)
);

OAI21X1 _8408_ (
    .A(_996__bF$buf3),
    .B(_1309_),
    .C(_1283_),
    .Y(_852_)
);

NAND2X1 _8409_ (
    .A(\genblk1[1].u_ce.Xcalc [2]),
    .B(_996__bF$buf2),
    .Y(_1310_)
);

AOI21X1 _8410_ (
    .A(_1284_),
    .B(_1305_),
    .C(_1303_),
    .Y(_1311_)
);

NAND2X1 _8411_ (
    .A(_1281_),
    .B(_1298_),
    .Y(_1312_)
);

NAND2X1 _8412_ (
    .A(1'h1),
    .B(_1208_),
    .Y(_1313_)
);

OAI21X1 _8413_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .C(_1313_),
    .Y(_1314_)
);

NAND2X1 _8414_ (
    .A(_973__bF$buf0),
    .B(_1271_),
    .Y(_1315_)
);

OAI21X1 _8415_ (
    .A(_973__bF$buf4),
    .B(_1314_),
    .C(_1315_),
    .Y(_1316_)
);

NAND2X1 _8416_ (
    .A(_1079_),
    .B(_1264_),
    .Y(_1317_)
);

NAND2X1 _8417_ (
    .A(_1273_),
    .B(_1078_),
    .Y(_1318_)
);

NAND2X1 _8418_ (
    .A(_1317_),
    .B(_1318_),
    .Y(_1319_)
);

AOI21X1 _8419_ (
    .A(_1316_),
    .B(1'h0),
    .C(_1319_),
    .Y(_1320_)
);

INVX1 _8420_ (
    .A(_1320_),
    .Y(_1321_)
);

NAND3X1 _8421_ (
    .A(_1010__bF$buf4),
    .B(_1321_),
    .C(_1312_),
    .Y(_1322_)
);

AOI21X1 _8422_ (
    .A(_1269_),
    .B(_1275_),
    .C(_1301_),
    .Y(_1323_)
);

OAI21X1 _8423_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1323_),
    .C(_1320_),
    .Y(_1324_)
);

NAND3X1 _8424_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(_1324_),
    .C(_1322_),
    .Y(_1325_)
);

INVX1 _8425_ (
    .A(_1325_),
    .Y(_1326_)
);

AOI21X1 _8426_ (
    .A(_1322_),
    .B(_1324_),
    .C(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1327_)
);

NOR2X1 _8427_ (
    .A(_1327_),
    .B(_1326_),
    .Y(_1328_)
);

AND2X2 _8428_ (
    .A(_1328_),
    .B(_1311_),
    .Y(_1329_)
);

NOR2X1 _8429_ (
    .A(_1311_),
    .B(_1328_),
    .Y(_1330_)
);

OAI21X1 _8430_ (
    .A(_1330_),
    .B(_1329_),
    .C(_1065_),
    .Y(_1331_)
);

OAI21X1 _8431_ (
    .A(_996__bF$buf1),
    .B(_1331_),
    .C(_1310_),
    .Y(_853_)
);

OAI21X1 _8432_ (
    .A(_1327_),
    .B(_1311_),
    .C(_1325_),
    .Y(_1332_)
);

INVX1 _8433_ (
    .A(_1332_),
    .Y(_1333_)
);

NAND2X1 _8434_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [10]),
    .Y(_1334_)
);

OAI21X1 _8435_ (
    .A(1'h1),
    .B(_1208_),
    .C(_1334_),
    .Y(_1335_)
);

MUX2X1 _8436_ (
    .A(_1335_),
    .B(_1292_),
    .S(1'h0),
    .Y(_1336_)
);

NOR2X1 _8437_ (
    .A(_972__bF$buf0),
    .B(_1336_),
    .Y(_1337_)
);

NAND2X1 _8438_ (
    .A(_1079_),
    .B(_1286_),
    .Y(_1338_)
);

NAND2X1 _8439_ (
    .A(_1295_),
    .B(_1078_),
    .Y(_1339_)
);

NAND2X1 _8440_ (
    .A(_1338_),
    .B(_1339_),
    .Y(_1340_)
);

OR2X2 _8441_ (
    .A(_1337_),
    .B(_1340_),
    .Y(_1341_)
);

OAI21X1 _8442_ (
    .A(_1321_),
    .B(_1312_),
    .C(_1010__bF$buf3),
    .Y(_1342_)
);

OR2X2 _8443_ (
    .A(_1342_),
    .B(_1341_),
    .Y(_1343_)
);

OAI21X1 _8444_ (
    .A(_1337_),
    .B(_1340_),
    .C(_1342_),
    .Y(_1344_)
);

AOI21X1 _8445_ (
    .A(_1343_),
    .B(_1344_),
    .C(_1018_),
    .Y(_1345_)
);

INVX1 _8446_ (
    .A(_1345_),
    .Y(_1346_)
);

NAND3X1 _8447_ (
    .A(_1018_),
    .B(_1344_),
    .C(_1343_),
    .Y(_1347_)
);

NAND2X1 _8448_ (
    .A(_1347_),
    .B(_1346_),
    .Y(_1348_)
);

OR2X2 _8449_ (
    .A(_1348_),
    .B(_1333_),
    .Y(_1349_)
);

NAND2X1 _8450_ (
    .A(_1333_),
    .B(_1348_),
    .Y(_1350_)
);

NAND2X1 _8451_ (
    .A(_1350_),
    .B(_1349_),
    .Y(_1351_)
);

AOI22X1 _8452_ (
    .A(_964_),
    .B(_996__bF$buf0),
    .C(_1351_),
    .D(_994_),
    .Y(_854_)
);

AOI21X1 _8453_ (
    .A(_1332_),
    .B(_1347_),
    .C(_1345_),
    .Y(_1352_)
);

NAND2X1 _8454_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1353_)
);

OAI21X1 _8455_ (
    .A(1'h1),
    .B(_1223_),
    .C(_1353_),
    .Y(_1354_)
);

NAND2X1 _8456_ (
    .A(1'h0),
    .B(_1354_),
    .Y(_1355_)
);

OAI21X1 _8457_ (
    .A(1'h0),
    .B(_1314_),
    .C(_1355_),
    .Y(_1356_)
);

NAND2X1 _8458_ (
    .A(1'h0),
    .B(_1356_),
    .Y(_1357_)
);

OAI21X1 _8459_ (
    .A(1'h0),
    .B(_1274_),
    .C(_1357_),
    .Y(_1358_)
);

INVX1 _8460_ (
    .A(_1358_),
    .Y(_1359_)
);

NAND3X1 _8461_ (
    .A(_1320_),
    .B(_1281_),
    .C(_1298_),
    .Y(_1360_)
);

OAI21X1 _8462_ (
    .A(_1341_),
    .B(_1360_),
    .C(_1010__bF$buf2),
    .Y(_1361_)
);

OR2X2 _8463_ (
    .A(_1361_),
    .B(_1359_),
    .Y(_1362_)
);

NOR2X1 _8464_ (
    .A(_1341_),
    .B(_1360_),
    .Y(_1363_)
);

OAI21X1 _8465_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1363_),
    .C(_1359_),
    .Y(_1364_)
);

NAND3X1 _8466_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(_1364_),
    .C(_1362_),
    .Y(_1365_)
);

OR2X2 _8467_ (
    .A(_1361_),
    .B(_1358_),
    .Y(_1366_)
);

OAI21X1 _8468_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1363_),
    .C(_1358_),
    .Y(_1367_)
);

NAND3X1 _8469_ (
    .A(_977_),
    .B(_1367_),
    .C(_1366_),
    .Y(_1368_)
);

NAND2X1 _8470_ (
    .A(_1365_),
    .B(_1368_),
    .Y(_1369_)
);

OR2X2 _8471_ (
    .A(_1352_),
    .B(_1369_),
    .Y(_1370_)
);

NAND2X1 _8472_ (
    .A(_1369_),
    .B(_1352_),
    .Y(_1371_)
);

NAND2X1 _8473_ (
    .A(_1371_),
    .B(_1370_),
    .Y(_1372_)
);

AOI22X1 _8474_ (
    .A(_959_),
    .B(_996__bF$buf4),
    .C(_1372_),
    .D(_994_),
    .Y(_855_)
);

INVX1 _8475_ (
    .A(\genblk1[1].u_ce.Xcalc [5]),
    .Y(_1373_)
);

OAI21X1 _8476_ (
    .A(_1369_),
    .B(_1352_),
    .C(_1365_),
    .Y(_1374_)
);

NAND2X1 _8477_ (
    .A(_1359_),
    .B(_1363_),
    .Y(_1375_)
);

NOR2X1 _8478_ (
    .A(_973__bF$buf3),
    .B(_1249_),
    .Y(_1376_)
);

AOI21X1 _8479_ (
    .A(_973__bF$buf2),
    .B(_1335_),
    .C(_1376_),
    .Y(_1377_)
);

NAND2X1 _8480_ (
    .A(_972__bF$buf4),
    .B(_1297_),
    .Y(_1378_)
);

OAI21X1 _8481_ (
    .A(_972__bF$buf3),
    .B(_1377_),
    .C(_1378_),
    .Y(_1379_)
);

INVX1 _8482_ (
    .A(_1379_),
    .Y(_1380_)
);

NAND3X1 _8483_ (
    .A(_1010__bF$buf1),
    .B(_1380_),
    .C(_1375_),
    .Y(_1381_)
);

NOR2X1 _8484_ (
    .A(_1340_),
    .B(_1337_),
    .Y(_1382_)
);

NAND3X1 _8485_ (
    .A(_1320_),
    .B(_1382_),
    .C(_1323_),
    .Y(_1383_)
);

OAI21X1 _8486_ (
    .A(_1358_),
    .B(_1383_),
    .C(_1010__bF$buf0),
    .Y(_1384_)
);

NAND2X1 _8487_ (
    .A(_1379_),
    .B(_1384_),
    .Y(_1385_)
);

AOI21X1 _8488_ (
    .A(_1381_),
    .B(_1385_),
    .C(_1014_),
    .Y(_1386_)
);

INVX1 _8489_ (
    .A(_1386_),
    .Y(_1387_)
);

NAND3X1 _8490_ (
    .A(_1014_),
    .B(_1385_),
    .C(_1381_),
    .Y(_1388_)
);

NAND2X1 _8491_ (
    .A(_1388_),
    .B(_1387_),
    .Y(_1389_)
);

NOR2X1 _8492_ (
    .A(_1389_),
    .B(_1374_),
    .Y(_1390_)
);

AND2X2 _8493_ (
    .A(_1374_),
    .B(_1389_),
    .Y(_1391_)
);

OAI21X1 _8494_ (
    .A(_1390_),
    .B(_1391_),
    .C(_994_),
    .Y(_1392_)
);

OAI21X1 _8495_ (
    .A(_1373_),
    .B(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .C(_1392_),
    .Y(_856_)
);

INVX1 _8496_ (
    .A(\genblk1[1].u_ce.Xcalc [6]),
    .Y(_1393_)
);

NAND3X1 _8497_ (
    .A(_1359_),
    .B(_1380_),
    .C(_1363_),
    .Y(_1394_)
);

AOI21X1 _8498_ (
    .A(_973__bF$buf1),
    .B(_1354_),
    .C(_1376_),
    .Y(_1395_)
);

NAND2X1 _8499_ (
    .A(1'h0),
    .B(_1395_),
    .Y(_1396_)
);

OAI21X1 _8500_ (
    .A(1'h0),
    .B(_1316_),
    .C(_1396_),
    .Y(_1397_)
);

NAND3X1 _8501_ (
    .A(_1010__bF$buf5),
    .B(_1397_),
    .C(_1394_),
    .Y(_1398_)
);

NOR3X1 _8502_ (
    .A(_1358_),
    .B(_1379_),
    .C(_1383_),
    .Y(_1399_)
);

INVX1 _8503_ (
    .A(_1397_),
    .Y(_1400_)
);

OAI21X1 _8504_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1399_),
    .C(_1400_),
    .Y(_1401_)
);

NAND2X1 _8505_ (
    .A(_1398_),
    .B(_1401_),
    .Y(_1402_)
);

NAND2X1 _8506_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(_1402_),
    .Y(_1403_)
);

NAND3X1 _8507_ (
    .A(_974_),
    .B(_1398_),
    .C(_1401_),
    .Y(_1404_)
);

NAND2X1 _8508_ (
    .A(_1404_),
    .B(_1403_),
    .Y(_1405_)
);

AOI21X1 _8509_ (
    .A(_1366_),
    .B(_1367_),
    .C(_977_),
    .Y(_1406_)
);

NOR2X1 _8510_ (
    .A(_1406_),
    .B(_1386_),
    .Y(_1407_)
);

OAI21X1 _8511_ (
    .A(_1369_),
    .B(_1352_),
    .C(_1407_),
    .Y(_1408_)
);

NAND2X1 _8512_ (
    .A(_1388_),
    .B(_1408_),
    .Y(_1409_)
);

NOR2X1 _8513_ (
    .A(_1405_),
    .B(_1409_),
    .Y(_1410_)
);

AND2X2 _8514_ (
    .A(_1403_),
    .B(_1404_),
    .Y(_1411_)
);

AND2X2 _8515_ (
    .A(_1365_),
    .B(_1368_),
    .Y(_1412_)
);

NAND3X1 _8516_ (
    .A(_1388_),
    .B(_1412_),
    .C(_1387_),
    .Y(_1413_)
);

AOI21X1 _8517_ (
    .A(_1406_),
    .B(_1388_),
    .C(_1386_),
    .Y(_1414_)
);

OAI21X1 _8518_ (
    .A(_1352_),
    .B(_1413_),
    .C(_1414_),
    .Y(_1415_)
);

NOR2X1 _8519_ (
    .A(_1411_),
    .B(_1415_),
    .Y(_1416_)
);

OAI21X1 _8520_ (
    .A(_1416_),
    .B(_1410_),
    .C(_1065_),
    .Y(_1417_)
);

NAND2X1 _8521_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .B(_1417_),
    .Y(_1418_)
);

OAI21X1 _8522_ (
    .A(_1393_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1418_),
    .Y(_857_)
);

INVX1 _8523_ (
    .A(\genblk1[1].u_ce.Xcalc [7]),
    .Y(_1419_)
);

INVX1 _8524_ (
    .A(_1403_),
    .Y(_1420_)
);

NAND2X1 _8525_ (
    .A(_1397_),
    .B(_1399_),
    .Y(_1421_)
);

NOR2X1 _8526_ (
    .A(_972__bF$buf2),
    .B(_1249_),
    .Y(_1422_)
);

INVX1 _8527_ (
    .A(_1422_),
    .Y(_1423_)
);

OAI21X1 _8528_ (
    .A(1'h0),
    .B(_1336_),
    .C(_1423_),
    .Y(_1424_)
);

NAND3X1 _8529_ (
    .A(_1010__bF$buf4),
    .B(_1424_),
    .C(_1421_),
    .Y(_1425_)
);

INVX1 _8530_ (
    .A(_1424_),
    .Y(_1426_)
);

OAI21X1 _8531_ (
    .A(_1400_),
    .B(_1394_),
    .C(_1010__bF$buf3),
    .Y(_1427_)
);

NAND2X1 _8532_ (
    .A(_1426_),
    .B(_1427_),
    .Y(_1428_)
);

NAND3X1 _8533_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(_1425_),
    .C(_1428_),
    .Y(_1429_)
);

NAND3X1 _8534_ (
    .A(_1010__bF$buf2),
    .B(_1426_),
    .C(_1421_),
    .Y(_1430_)
);

NAND2X1 _8535_ (
    .A(_1424_),
    .B(_1427_),
    .Y(_1431_)
);

NAND3X1 _8536_ (
    .A(_1011_),
    .B(_1430_),
    .C(_1431_),
    .Y(_1432_)
);

NAND2X1 _8537_ (
    .A(_1429_),
    .B(_1432_),
    .Y(_1433_)
);

OAI21X1 _8538_ (
    .A(_1420_),
    .B(_1410_),
    .C(_1433_),
    .Y(_1434_)
);

NOR2X1 _8539_ (
    .A(_1420_),
    .B(_1410_),
    .Y(_1435_)
);

INVX1 _8540_ (
    .A(_1433_),
    .Y(_1436_)
);

AOI21X1 _8541_ (
    .A(_1435_),
    .B(_1436_),
    .C(_993_),
    .Y(_1437_)
);

AOI22X1 _8542_ (
    .A(_1419_),
    .B(_996__bF$buf3),
    .C(_1437_),
    .D(_1434_),
    .Y(_858_)
);

OAI21X1 _8543_ (
    .A(_1403_),
    .B(_1433_),
    .C(_1429_),
    .Y(_1438_)
);

NOR2X1 _8544_ (
    .A(_1405_),
    .B(_1433_),
    .Y(_1439_)
);

AOI21X1 _8545_ (
    .A(_1439_),
    .B(_1415_),
    .C(_1438_),
    .Y(_1440_)
);

INVX1 _8546_ (
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1441_)
);

NAND3X1 _8547_ (
    .A(_1397_),
    .B(_1426_),
    .C(_1399_),
    .Y(_1442_)
);

INVX1 _8548_ (
    .A(_1356_),
    .Y(_1443_)
);

OAI21X1 _8549_ (
    .A(1'h0),
    .B(_1443_),
    .C(_1423_),
    .Y(_1444_)
);

INVX1 _8550_ (
    .A(_1444_),
    .Y(_1445_)
);

NAND3X1 _8551_ (
    .A(_1010__bF$buf1),
    .B(_1445_),
    .C(_1442_),
    .Y(_1446_)
);

OAI21X1 _8552_ (
    .A(_1424_),
    .B(_1421_),
    .C(_1010__bF$buf0),
    .Y(_1447_)
);

NAND2X1 _8553_ (
    .A(_1444_),
    .B(_1447_),
    .Y(_1448_)
);

AOI21X1 _8554_ (
    .A(_1448_),
    .B(_1446_),
    .C(_1441_),
    .Y(_1449_)
);

NAND3X1 _8555_ (
    .A(_1010__bF$buf5),
    .B(_1444_),
    .C(_1442_),
    .Y(_1450_)
);

NAND2X1 _8556_ (
    .A(_1445_),
    .B(_1447_),
    .Y(_1451_)
);

AOI21X1 _8557_ (
    .A(_1451_),
    .B(_1450_),
    .C(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1452_)
);

OAI21X1 _8558_ (
    .A(_1449_),
    .B(_1452_),
    .C(_1440_),
    .Y(_1453_)
);

INVX1 _8559_ (
    .A(_1453_),
    .Y(_1454_)
);

OR2X2 _8560_ (
    .A(_1449_),
    .B(_1452_),
    .Y(_1455_)
);

OAI21X1 _8561_ (
    .A(_1455_),
    .B(_1440_),
    .C(_994_),
    .Y(_1456_)
);

OAI22X1 _8562_ (
    .A(_956_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1456_),
    .D(_1454_),
    .Y(_859_)
);

NAND2X1 _8563_ (
    .A(\genblk1[1].u_ce.Xcalc [9]),
    .B(_996__bF$buf2),
    .Y(_1457_)
);

NOR2X1 _8564_ (
    .A(_1455_),
    .B(_1440_),
    .Y(_1458_)
);

NOR2X1 _8565_ (
    .A(_1449_),
    .B(_1458_),
    .Y(_1459_)
);

OAI21X1 _8566_ (
    .A(1'h0),
    .B(_1377_),
    .C(_1423_),
    .Y(_1460_)
);

INVX1 _8567_ (
    .A(_1460_),
    .Y(_1461_)
);

OAI21X1 _8568_ (
    .A(_1444_),
    .B(_1442_),
    .C(_1010__bF$buf4),
    .Y(_1462_)
);

NAND2X1 _8569_ (
    .A(_1461_),
    .B(_1462_),
    .Y(_1463_)
);

OR2X2 _8570_ (
    .A(_1462_),
    .B(_1461_),
    .Y(_1464_)
);

NAND3X1 _8571_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(_1463_),
    .C(_1464_),
    .Y(_1465_)
);

NAND2X1 _8572_ (
    .A(_1463_),
    .B(_1464_),
    .Y(_1466_)
);

NAND2X1 _8573_ (
    .A(_1073_),
    .B(_1466_),
    .Y(_1467_)
);

NAND2X1 _8574_ (
    .A(_1465_),
    .B(_1467_),
    .Y(_1468_)
);

AND2X2 _8575_ (
    .A(_1459_),
    .B(_1468_),
    .Y(_1469_)
);

OAI21X1 _8576_ (
    .A(_1468_),
    .B(_1459_),
    .C(_994_),
    .Y(_1470_)
);

OAI21X1 _8577_ (
    .A(_1470_),
    .B(_1469_),
    .C(_1457_),
    .Y(_860_)
);

INVX1 _8578_ (
    .A(\genblk1[1].u_ce.Xcalc [10]),
    .Y(_1471_)
);

INVX1 _8579_ (
    .A(_1465_),
    .Y(_1472_)
);

AOI21X1 _8580_ (
    .A(_1449_),
    .B(_1467_),
    .C(_1472_),
    .Y(_1473_)
);

NOR2X1 _8581_ (
    .A(_1449_),
    .B(_1452_),
    .Y(_1474_)
);

NAND3X1 _8582_ (
    .A(_1465_),
    .B(_1467_),
    .C(_1474_),
    .Y(_1475_)
);

OAI21X1 _8583_ (
    .A(_1440_),
    .B(_1475_),
    .C(_1473_),
    .Y(_1476_)
);

OAI21X1 _8584_ (
    .A(1'h0),
    .B(_1395_),
    .C(_1423_),
    .Y(_1477_)
);

INVX1 _8585_ (
    .A(_1477_),
    .Y(_1478_)
);

OR2X2 _8586_ (
    .A(_1442_),
    .B(_1444_),
    .Y(_1479_)
);

OAI21X1 _8587_ (
    .A(_1460_),
    .B(_1479_),
    .C(_1010__bF$buf3),
    .Y(_1480_)
);

NAND2X1 _8588_ (
    .A(_1478_),
    .B(_1480_),
    .Y(_1481_)
);

OR2X2 _8589_ (
    .A(_1480_),
    .B(_1478_),
    .Y(_1482_)
);

NAND3X1 _8590_ (
    .A(\genblk1[1].u_ce.Xin12b [10]),
    .B(_1481_),
    .C(_1482_),
    .Y(_1483_)
);

AND2X2 _8591_ (
    .A(_1480_),
    .B(_1478_),
    .Y(_1484_)
);

NOR2X1 _8592_ (
    .A(_1478_),
    .B(_1480_),
    .Y(_1485_)
);

OAI21X1 _8593_ (
    .A(_1485_),
    .B(_1484_),
    .C(_1094_),
    .Y(_1486_)
);

NAND2X1 _8594_ (
    .A(_1486_),
    .B(_1483_),
    .Y(_1487_)
);

AND2X2 _8595_ (
    .A(_1476_),
    .B(_1487_),
    .Y(_1488_)
);

NOR2X1 _8596_ (
    .A(_1487_),
    .B(_1476_),
    .Y(_1489_)
);

NOR2X1 _8597_ (
    .A(_1488_),
    .B(_1489_),
    .Y(_1490_)
);

AOI22X1 _8598_ (
    .A(_1471_),
    .B(_996__bF$buf1),
    .C(_1490_),
    .D(_994_),
    .Y(_861_)
);

NAND2X1 _8599_ (
    .A(\genblk1[1].u_ce.Xcalc [11]),
    .B(_996__bF$buf0),
    .Y(_1491_)
);

INVX1 _8600_ (
    .A(_1483_),
    .Y(_1492_)
);

AOI21X1 _8601_ (
    .A(_1476_),
    .B(_1486_),
    .C(_1492_),
    .Y(_1493_)
);

NAND2X1 _8602_ (
    .A(_1010__bF$buf2),
    .B(_1481_),
    .Y(_1494_)
);

NOR2X1 _8603_ (
    .A(_1251_),
    .B(_1494_),
    .Y(_1495_)
);

AOI21X1 _8604_ (
    .A(_1481_),
    .B(_1010__bF$buf1),
    .C(_1252_),
    .Y(_1496_)
);

NOR2X1 _8605_ (
    .A(_1496_),
    .B(_1495_),
    .Y(_1497_)
);

AND2X2 _8606_ (
    .A(_1493_),
    .B(_1497_),
    .Y(_1498_)
);

OAI21X1 _8607_ (
    .A(_1497_),
    .B(_1493_),
    .C(_994_),
    .Y(_1499_)
);

OAI21X1 _8608_ (
    .A(_1499_),
    .B(_1498_),
    .C(_1491_),
    .Y(_862_)
);

OAI21X1 _8609_ (
    .A(1'h1),
    .B(_973__bF$buf0),
    .C(_992_),
    .Y(_1500_)
);

OAI21X1 _8610_ (
    .A(_1267_),
    .B(_1500_),
    .C(\genblk1[1].u_ce.Ain0 [0]),
    .Y(_1501_)
);

INVX1 _8611_ (
    .A(\genblk1[1].u_ce.Ain0 [0]),
    .Y(_1502_)
);

NOR2X1 _8612_ (
    .A(_1267_),
    .B(_1500_),
    .Y(_1503_)
);

NAND2X1 _8613_ (
    .A(_1502_),
    .B(_1503_),
    .Y(_1504_)
);

NAND2X1 _8614_ (
    .A(_1501_),
    .B(_1504_),
    .Y(_1505_)
);

NAND2X1 _8615_ (
    .A(\genblk1[1].u_ce.Acalc [0]),
    .B(_996__bF$buf4),
    .Y(_1506_)
);

OAI21X1 _8616_ (
    .A(_996__bF$buf3),
    .B(_1505_),
    .C(_1506_),
    .Y(_863_)
);

NAND2X1 _8617_ (
    .A(\genblk1[1].u_ce.Acalc [1]),
    .B(_996__bF$buf2),
    .Y(_1507_)
);

INVX1 _8618_ (
    .A(_1501_),
    .Y(_1508_)
);

NOR2X1 _8619_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_1509_)
);

AOI21X1 _8620_ (
    .A(_1267_),
    .B(1'h0),
    .C(_1509_),
    .Y(_1510_)
);

NOR2X1 _8621_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1510_),
    .Y(_1511_)
);

OAI21X1 _8622_ (
    .A(_1267_),
    .B(_1500_),
    .C(_1010__bF$buf0),
    .Y(_1512_)
);

AND2X2 _8623_ (
    .A(_1512_),
    .B(_1510_),
    .Y(_1513_)
);

OR2X2 _8624_ (
    .A(_1513_),
    .B(_1511_),
    .Y(_1514_)
);

OR2X2 _8625_ (
    .A(_1514_),
    .B(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1515_)
);

OAI21X1 _8626_ (
    .A(_1511_),
    .B(_1513_),
    .C(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1516_)
);

NAND2X1 _8627_ (
    .A(_1516_),
    .B(_1515_),
    .Y(_1517_)
);

NOR2X1 _8628_ (
    .A(_1508_),
    .B(_1517_),
    .Y(_1518_)
);

NAND2X1 _8629_ (
    .A(_1508_),
    .B(_1517_),
    .Y(_1519_)
);

NAND2X1 _8630_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .B(_1519_),
    .Y(_1520_)
);

OAI21X1 _8631_ (
    .A(_1518_),
    .B(_1520_),
    .C(_1507_),
    .Y(_864_)
);

INVX1 _8632_ (
    .A(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1521_)
);

OAI21X1 _8633_ (
    .A(_1521_),
    .B(_1514_),
    .C(_1519_),
    .Y(_1522_)
);

OAI21X1 _8634_ (
    .A(_1002_),
    .B(_973__bF$buf4),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_1523_)
);

OAI21X1 _8635_ (
    .A(1'h1),
    .B(1'h0),
    .C(1'h0),
    .Y(_1524_)
);

MUX2X1 _8636_ (
    .A(_1524_),
    .B(1'h0),
    .S(_1523_),
    .Y(_1525_)
);

NAND2X1 _8637_ (
    .A(\genblk1[1].u_ce.Ain1 [0]),
    .B(_1525_),
    .Y(_1526_)
);

OR2X2 _8638_ (
    .A(_1525_),
    .B(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_1527_)
);

NAND2X1 _8639_ (
    .A(_1526_),
    .B(_1527_),
    .Y(_1528_)
);

INVX1 _8640_ (
    .A(_1528_),
    .Y(_1529_)
);

NOR2X1 _8641_ (
    .A(_1529_),
    .B(_1522_),
    .Y(_1530_)
);

NAND2X1 _8642_ (
    .A(_1529_),
    .B(_1522_),
    .Y(_1531_)
);

NAND2X1 _8643_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1531_),
    .Y(_1532_)
);

OAI22X1 _8644_ (
    .A(_918_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_1530_),
    .D(_1532_),
    .Y(_865_)
);

NOR2X1 _8645_ (
    .A(\genblk1[1].u_ce.Acalc [3]),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_1533_)
);

NAND2X1 _8646_ (
    .A(_1526_),
    .B(_1531_),
    .Y(_1534_)
);

INVX1 _8647_ (
    .A(_1534_),
    .Y(_1535_)
);

INVX1 _8648_ (
    .A(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_1536_)
);

NOR2X1 _8649_ (
    .A(1'h1),
    .B(_973__bF$buf3),
    .Y(_1537_)
);

OAI21X1 _8650_ (
    .A(_972__bF$buf1),
    .B(_1537_),
    .C(_1010__bF$buf5),
    .Y(_1538_)
);

OAI21X1 _8651_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_1539_)
);

OAI21X1 _8652_ (
    .A(_1002_),
    .B(_1539_),
    .C(_1538_),
    .Y(_1540_)
);

NOR2X1 _8653_ (
    .A(_1536_),
    .B(_1540_),
    .Y(_1541_)
);

NAND2X1 _8654_ (
    .A(_1536_),
    .B(_1540_),
    .Y(_1542_)
);

INVX1 _8655_ (
    .A(_1542_),
    .Y(_1543_)
);

NOR2X1 _8656_ (
    .A(_1541_),
    .B(_1543_),
    .Y(_1544_)
);

OAI21X1 _8657_ (
    .A(_1544_),
    .B(_1535_),
    .C(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .Y(_1545_)
);

AOI21X1 _8658_ (
    .A(_1535_),
    .B(_1544_),
    .C(_1545_),
    .Y(_1546_)
);

NOR2X1 _8659_ (
    .A(_1533_),
    .B(_1546_),
    .Y(_866_)
);

NAND2X1 _8660_ (
    .A(\genblk1[1].u_ce.Acalc [4]),
    .B(_996__bF$buf1),
    .Y(_1547_)
);

INVX1 _8661_ (
    .A(\genblk1[1].u_ce.Ain12b [4]),
    .Y(_1548_)
);

AOI21X1 _8662_ (
    .A(_1267_),
    .B(1'h0),
    .C(_1010__bF$buf4),
    .Y(_1549_)
);

OAI21X1 _8663_ (
    .A(1'h0),
    .B(_1267_),
    .C(_1549_),
    .Y(_1550_)
);

OAI21X1 _8664_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1510_),
    .C(_1550_),
    .Y(_1551_)
);

OR2X2 _8665_ (
    .A(_1551_),
    .B(_1548_),
    .Y(_1552_)
);

NAND2X1 _8666_ (
    .A(_1548_),
    .B(_1551_),
    .Y(_1553_)
);

NAND2X1 _8667_ (
    .A(_1553_),
    .B(_1552_),
    .Y(_1554_)
);

AOI21X1 _8668_ (
    .A(_1534_),
    .B(_1542_),
    .C(_1541_),
    .Y(_1555_)
);

AND2X2 _8669_ (
    .A(_1555_),
    .B(_1554_),
    .Y(_1556_)
);

OAI21X1 _8670_ (
    .A(_1554_),
    .B(_1555_),
    .C(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_1557_)
);

OAI21X1 _8671_ (
    .A(_1557_),
    .B(_1556_),
    .C(_1547_),
    .Y(_867_)
);

OAI21X1 _8672_ (
    .A(_1554_),
    .B(_1555_),
    .C(_1552_),
    .Y(_1558_)
);

INVX1 _8673_ (
    .A(\genblk1[1].u_ce.Ain12b [5]),
    .Y(_1559_)
);

OAI21X1 _8674_ (
    .A(_1266_),
    .B(_1079_),
    .C(_1010__bF$buf3),
    .Y(_1560_)
);

OAI21X1 _8675_ (
    .A(1'h1),
    .B(1'h0),
    .C(_992_),
    .Y(_1561_)
);

OR2X2 _8676_ (
    .A(_1561_),
    .B(_1010__bF$buf2),
    .Y(_1562_)
);

NAND2X1 _8677_ (
    .A(_1560_),
    .B(_1562_),
    .Y(_1563_)
);

OR2X2 _8678_ (
    .A(_1563_),
    .B(_1559_),
    .Y(_1564_)
);

NAND2X1 _8679_ (
    .A(_1559_),
    .B(_1563_),
    .Y(_1565_)
);

NAND2X1 _8680_ (
    .A(_1565_),
    .B(_1564_),
    .Y(_1566_)
);

INVX1 _8681_ (
    .A(_1566_),
    .Y(_1567_)
);

NOR2X1 _8682_ (
    .A(_1567_),
    .B(_1558_),
    .Y(_1568_)
);

NAND2X1 _8683_ (
    .A(_1567_),
    .B(_1558_),
    .Y(_1569_)
);

NAND2X1 _8684_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1569_),
    .Y(_1570_)
);

OAI22X1 _8685_ (
    .A(_935_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_1568_),
    .D(_1570_),
    .Y(_868_)
);

NAND2X1 _8686_ (
    .A(\genblk1[1].u_ce.Acalc [6]),
    .B(_996__bF$buf0),
    .Y(_1571_)
);

INVX1 _8687_ (
    .A(_1554_),
    .Y(_1572_)
);

NAND2X1 _8688_ (
    .A(_1567_),
    .B(_1572_),
    .Y(_1573_)
);

OAI21X1 _8689_ (
    .A(_1552_),
    .B(_1566_),
    .C(_1564_),
    .Y(_1574_)
);

INVX1 _8690_ (
    .A(_1574_),
    .Y(_1575_)
);

OAI21X1 _8691_ (
    .A(_1573_),
    .B(_1555_),
    .C(_1575_),
    .Y(_1576_)
);

OAI21X1 _8692_ (
    .A(1'h0),
    .B(_1002_),
    .C(_972__bF$buf0),
    .Y(_1577_)
);

NOR2X1 _8693_ (
    .A(_1577_),
    .B(_1537_),
    .Y(_1578_)
);

NAND2X1 _8694_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1578_),
    .Y(_1579_)
);

OAI21X1 _8695_ (
    .A(_1577_),
    .B(_1537_),
    .C(_1010__bF$buf1),
    .Y(_1580_)
);

NAND2X1 _8696_ (
    .A(_1580_),
    .B(_1579_),
    .Y(_1581_)
);

NAND2X1 _8697_ (
    .A(\genblk1[1].u_ce.Ain12b [6]),
    .B(_1581_),
    .Y(_1582_)
);

OR2X2 _8698_ (
    .A(_1581_),
    .B(\genblk1[1].u_ce.Ain12b [6]),
    .Y(_1583_)
);

NAND2X1 _8699_ (
    .A(_1582_),
    .B(_1583_),
    .Y(_1584_)
);

INVX1 _8700_ (
    .A(_1584_),
    .Y(_1585_)
);

NOR2X1 _8701_ (
    .A(_1585_),
    .B(_1576_),
    .Y(_1586_)
);

NAND2X1 _8702_ (
    .A(_1585_),
    .B(_1576_),
    .Y(_1587_)
);

NAND2X1 _8703_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .B(_1587_),
    .Y(_1588_)
);

OAI21X1 _8704_ (
    .A(_1586_),
    .B(_1588_),
    .C(_1571_),
    .Y(_869_)
);

INVX1 _8705_ (
    .A(\genblk1[1].u_ce.Acalc [7]),
    .Y(_1589_)
);

NAND2X1 _8706_ (
    .A(_1582_),
    .B(_1587_),
    .Y(_1590_)
);

INVX1 _8707_ (
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .Y(_1591_)
);

NAND2X1 _8708_ (
    .A(_1010__bF$buf0),
    .B(_1509_),
    .Y(_1592_)
);

OR2X2 _8709_ (
    .A(_1509_),
    .B(_1010__bF$buf5),
    .Y(_1593_)
);

NAND2X1 _8710_ (
    .A(_1592_),
    .B(_1593_),
    .Y(_1594_)
);

NOR2X1 _8711_ (
    .A(_1591_),
    .B(_1594_),
    .Y(_1595_)
);

INVX1 _8712_ (
    .A(_1595_),
    .Y(_1596_)
);

NAND2X1 _8713_ (
    .A(_1591_),
    .B(_1594_),
    .Y(_1597_)
);

NAND2X1 _8714_ (
    .A(_1597_),
    .B(_1596_),
    .Y(_1598_)
);

OR2X2 _8715_ (
    .A(_1590_),
    .B(_1598_),
    .Y(_1599_)
);

AOI21X1 _8716_ (
    .A(_1590_),
    .B(_1598_),
    .C(_996__bF$buf4),
    .Y(_1600_)
);

AOI22X1 _8717_ (
    .A(_1589_),
    .B(_996__bF$buf3),
    .C(_1599_),
    .D(_1600_),
    .Y(_870_)
);

NAND2X1 _8718_ (
    .A(\genblk1[1].u_ce.Acalc [8]),
    .B(_996__bF$buf2),
    .Y(_1601_)
);

NOR2X1 _8719_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_992_),
    .Y(_1602_)
);

INVX1 _8720_ (
    .A(_1602_),
    .Y(_1603_)
);

NAND3X1 _8721_ (
    .A(\genblk1[1].u_ce.Ain12b [8]),
    .B(_1539_),
    .C(_1603_),
    .Y(_1604_)
);

INVX1 _8722_ (
    .A(_1604_),
    .Y(_1605_)
);

AOI21X1 _8723_ (
    .A(_1603_),
    .B(_1539_),
    .C(\genblk1[1].u_ce.Ain12b [8]),
    .Y(_1606_)
);

NOR2X1 _8724_ (
    .A(_1606_),
    .B(_1605_),
    .Y(_1607_)
);

OAI21X1 _8725_ (
    .A(_1582_),
    .B(_1598_),
    .C(_1596_),
    .Y(_1608_)
);

NOR2X1 _8726_ (
    .A(_1598_),
    .B(_1584_),
    .Y(_1609_)
);

AOI21X1 _8727_ (
    .A(_1609_),
    .B(_1574_),
    .C(_1608_),
    .Y(_1610_)
);

NAND3X1 _8728_ (
    .A(_1572_),
    .B(_1567_),
    .C(_1609_),
    .Y(_1611_)
);

OAI21X1 _8729_ (
    .A(_1611_),
    .B(_1555_),
    .C(_1610_),
    .Y(_1612_)
);

NOR2X1 _8730_ (
    .A(_1607_),
    .B(_1612_),
    .Y(_1613_)
);

NAND2X1 _8731_ (
    .A(_1607_),
    .B(_1612_),
    .Y(_1614_)
);

NAND2X1 _8732_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .B(_1614_),
    .Y(_1615_)
);

OAI21X1 _8733_ (
    .A(_1613_),
    .B(_1615_),
    .C(_1601_),
    .Y(_871_)
);

AOI21X1 _8734_ (
    .A(_1612_),
    .B(_1607_),
    .C(_1605_),
    .Y(_1616_)
);

OR2X2 _8735_ (
    .A(_1010__bF$buf4),
    .B(\genblk1[1].u_ce.Ain12b [9]),
    .Y(_1617_)
);

NAND2X1 _8736_ (
    .A(\genblk1[1].u_ce.Ain12b [9]),
    .B(_1010__bF$buf3),
    .Y(_1618_)
);

NAND2X1 _8737_ (
    .A(_1618_),
    .B(_1617_),
    .Y(_1619_)
);

AND2X2 _8738_ (
    .A(_1616_),
    .B(_1619_),
    .Y(_1620_)
);

OAI21X1 _8739_ (
    .A(_1619_),
    .B(_1616_),
    .C(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_1621_)
);

OAI22X1 _8740_ (
    .A(_932_),
    .B(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .C(_1621_),
    .D(_1620_),
    .Y(_872_)
);

NAND2X1 _8741_ (
    .A(\genblk1[1].u_ce.Acalc [10]),
    .B(_996__bF$buf1),
    .Y(_1622_)
);

OAI21X1 _8742_ (
    .A(_1619_),
    .B(_1604_),
    .C(_1618_),
    .Y(_1623_)
);

NAND3X1 _8743_ (
    .A(_1617_),
    .B(_1618_),
    .C(_1607_),
    .Y(_1624_)
);

INVX1 _8744_ (
    .A(_1624_),
    .Y(_1625_)
);

AOI21X1 _8745_ (
    .A(_1612_),
    .B(_1625_),
    .C(_1623_),
    .Y(_1626_)
);

INVX1 _8746_ (
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .Y(_1627_)
);

NAND2X1 _8747_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1627_),
    .Y(_1628_)
);

NAND2X1 _8748_ (
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .B(_1010__bF$buf2),
    .Y(_1629_)
);

NAND2X1 _8749_ (
    .A(_1628_),
    .B(_1629_),
    .Y(_1630_)
);

AND2X2 _8750_ (
    .A(_1626_),
    .B(_1630_),
    .Y(_1631_)
);

OAI21X1 _8751_ (
    .A(_1630_),
    .B(_1626_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1632_)
);

OAI21X1 _8752_ (
    .A(_1632_),
    .B(_1631_),
    .C(_1622_),
    .Y(_873_)
);

NAND2X1 _8753_ (
    .A(\genblk1[1].u_ce.Acalc [11]),
    .B(_996__bF$buf0),
    .Y(_1633_)
);

OAI21X1 _8754_ (
    .A(_1630_),
    .B(_1626_),
    .C(_1629_),
    .Y(_1634_)
);

OAI21X1 _8755_ (
    .A(_996__bF$buf4),
    .B(_1634_),
    .C(_1633_),
    .Y(_874_)
);

NAND2X1 _8756_ (
    .A(\genblk1[1].u_ce.LoadCtl [5]),
    .B(_923_),
    .Y(_1635_)
);

NAND2X1 _8757_ (
    .A(_924_),
    .B(_930_),
    .Y(_1636_)
);

NOR2X1 _8758_ (
    .A(_1635_),
    .B(_1636_),
    .Y(_1637_)
);

NAND2X1 _8759_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1637_),
    .Y(_1638_)
);

OAI21X1 _8760_ (
    .A(_1094_),
    .B(_1637_),
    .C(_1638_),
    .Y(_875_)
);

NAND2X1 _8761_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1637_),
    .Y(_1639_)
);

OAI21X1 _8762_ (
    .A(_1162_),
    .B(_1637_),
    .C(_1639_),
    .Y(_876_)
);

INVX1 _8763_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .Y(_1640_)
);

OR2X2 _8764_ (
    .A(_1636_),
    .B(_923_),
    .Y(_1641_)
);

OAI21X1 _8765_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1642_)
);

OAI21X1 _8766_ (
    .A(_1640_),
    .B(_1641_),
    .C(_1642_),
    .Y(_877_)
);

INVX1 _8767_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .Y(_1643_)
);

OAI21X1 _8768_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Xin12b [9]),
    .Y(_1644_)
);

OAI21X1 _8769_ (
    .A(_1643_),
    .B(_1641_),
    .C(_1644_),
    .Y(_878_)
);

NAND2X1 _8770_ (
    .A(_930_),
    .B(_927_),
    .Y(_1645_)
);

NAND2X1 _8771_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(_1645_),
    .Y(_1646_)
);

OAI21X1 _8772_ (
    .A(_1640_),
    .B(_1645_),
    .C(_1646_),
    .Y(_879_)
);

NAND2X1 _8773_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(_1645_),
    .Y(_1647_)
);

OAI21X1 _8774_ (
    .A(_1643_),
    .B(_1645_),
    .C(_1647_),
    .Y(_880_)
);

AND2X2 _8775_ (
    .A(_930_),
    .B(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_1648_)
);

NAND2X1 _8776_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1648_),
    .Y(_1649_)
);

OAI21X1 _8777_ (
    .A(_977_),
    .B(_1648_),
    .C(_1649_),
    .Y(_881_)
);

NAND2X1 _8778_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1648_),
    .Y(_1650_)
);

OAI21X1 _8779_ (
    .A(_1014_),
    .B(_1648_),
    .C(_1650_),
    .Y(_882_)
);

OAI21X1 _8780_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1651_)
);

OAI21X1 _8781_ (
    .A(_1640_),
    .B(_921_),
    .C(_1651_),
    .Y(_883_)
);

OAI21X1 _8782_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1652_)
);

OAI21X1 _8783_ (
    .A(_1643_),
    .B(_921_),
    .C(_1652_),
    .Y(_884_)
);

NAND2X1 _8784_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.X_ [0]),
    .Y(_1653_)
);

OAI21X1 _8785_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_984_),
    .C(_1653_),
    .Y(_885_)
);

NAND2X1 _8786_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.X_ [1]),
    .Y(_1654_)
);

OAI21X1 _8787_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1021_),
    .C(_1654_),
    .Y(_886_)
);

NAND2X1 _8788_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1637_),
    .Y(_1655_)
);

OAI21X1 _8789_ (
    .A(_1223_),
    .B(_1637_),
    .C(_1655_),
    .Y(_887_)
);

NAND2X1 _8790_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1637_),
    .Y(_1656_)
);

OAI21X1 _8791_ (
    .A(_1249_),
    .B(_1637_),
    .C(_1656_),
    .Y(_888_)
);

INVX1 _8792_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .Y(_1657_)
);

OAI21X1 _8793_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1658_)
);

OAI21X1 _8794_ (
    .A(_1657_),
    .B(_1641_),
    .C(_1658_),
    .Y(_889_)
);

INVX1 _8795_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .Y(_1659_)
);

OAI21X1 _8796_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1660_)
);

OAI21X1 _8797_ (
    .A(_1659_),
    .B(_1641_),
    .C(_1660_),
    .Y(_890_)
);

NAND2X1 _8798_ (
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .B(_1645_),
    .Y(_1661_)
);

OAI21X1 _8799_ (
    .A(_1657_),
    .B(_1645_),
    .C(_1661_),
    .Y(_891_)
);

NAND2X1 _8800_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(_1645_),
    .Y(_1662_)
);

OAI21X1 _8801_ (
    .A(_1659_),
    .B(_1645_),
    .C(_1662_),
    .Y(_892_)
);

NAND2X1 _8802_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1648_),
    .Y(_1663_)
);

OAI21X1 _8803_ (
    .A(_1093_),
    .B(_1648_),
    .C(_1663_),
    .Y(_893_)
);

NAND2X1 _8804_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1648_),
    .Y(_1664_)
);

OAI21X1 _8805_ (
    .A(_1114_),
    .B(_1648_),
    .C(_1664_),
    .Y(_894_)
);

OAI21X1 _8806_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1665_)
);

OAI21X1 _8807_ (
    .A(_1657_),
    .B(_921_),
    .C(_1665_),
    .Y(_895_)
);

OAI21X1 _8808_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1666_)
);

OAI21X1 _8809_ (
    .A(_1659_),
    .B(_921_),
    .C(_1666_),
    .Y(_896_)
);

NAND2X1 _8810_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.Y_ [0]),
    .Y(_1667_)
);

OAI21X1 _8811_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_971_),
    .C(_1667_),
    .Y(_897_)
);

NAND2X1 _8812_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.Y_ [1]),
    .Y(_1668_)
);

OAI21X1 _8813_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1009_),
    .C(_1668_),
    .Y(_898_)
);

NAND2X1 _8814_ (
    .A(\a[1] [0]),
    .B(_1637_),
    .Y(_1669_)
);

OAI21X1 _8815_ (
    .A(_1627_),
    .B(_1637_),
    .C(_1669_),
    .Y(_899_)
);

NAND2X1 _8816_ (
    .A(\a[1] [1]),
    .B(_1637_),
    .Y(_1670_)
);

OAI21X1 _8817_ (
    .A(_1010__bF$buf1),
    .B(_1637_),
    .C(_1670_),
    .Y(_900_)
);

INVX1 _8818_ (
    .A(\a[1] [0]),
    .Y(_1671_)
);

OAI21X1 _8819_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Ain12b [8]),
    .Y(_1672_)
);

OAI21X1 _8820_ (
    .A(_1671_),
    .B(_1641_),
    .C(_1672_),
    .Y(_901_)
);

INVX1 _8821_ (
    .A(\a[1] [1]),
    .Y(_1673_)
);

OAI21X1 _8822_ (
    .A(_923_),
    .B(_1636_),
    .C(\genblk1[1].u_ce.Ain12b [9]),
    .Y(_1674_)
);

OAI21X1 _8823_ (
    .A(_1673_),
    .B(_1641_),
    .C(_1674_),
    .Y(_902_)
);

NAND2X1 _8824_ (
    .A(\genblk1[1].u_ce.Ain12b [6]),
    .B(_1645_),
    .Y(_1675_)
);

OAI21X1 _8825_ (
    .A(_1671_),
    .B(_1645_),
    .C(_1675_),
    .Y(_903_)
);

NAND2X1 _8826_ (
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .B(_1645_),
    .Y(_911_)
);

OAI21X1 _8827_ (
    .A(_1673_),
    .B(_1645_),
    .C(_911_),
    .Y(_904_)
);

NAND2X1 _8828_ (
    .A(\a[1] [0]),
    .B(_1648_),
    .Y(_912_)
);

OAI21X1 _8829_ (
    .A(_1548_),
    .B(_1648_),
    .C(_912_),
    .Y(_905_)
);

NAND2X1 _8830_ (
    .A(\a[1] [1]),
    .B(_1648_),
    .Y(_913_)
);

OAI21X1 _8831_ (
    .A(_1559_),
    .B(_1648_),
    .C(_913_),
    .Y(_906_)
);

OAI21X1 _8832_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_914_)
);

OAI21X1 _8833_ (
    .A(_1671_),
    .B(_921_),
    .C(_914_),
    .Y(_907_)
);

OAI21X1 _8834_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_919_),
    .C(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_915_)
);

OAI21X1 _8835_ (
    .A(_1673_),
    .B(_921_),
    .C(_915_),
    .Y(_908_)
);

NAND2X1 _8836_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[1] [0]),
    .Y(_916_)
);

OAI21X1 _8837_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1502_),
    .C(_916_),
    .Y(_909_)
);

NAND2X1 _8838_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[1] [1]),
    .Y(_917_)
);

OAI21X1 _8839_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1521_),
    .C(_917_),
    .Y(_910_)
);

DFFPOSX1 _8840_ (
    .CLK(clk_bF$buf6),
    .D(_838_),
    .Q(\genblk1[1].u_ce.Ycalc [0])
);

DFFPOSX1 _8841_ (
    .CLK(clk_bF$buf5),
    .D(_839_),
    .Q(\genblk1[1].u_ce.Ycalc [1])
);

DFFPOSX1 _8842_ (
    .CLK(clk_bF$buf4),
    .D(_840_),
    .Q(\genblk1[1].u_ce.ISout )
);

DFFPOSX1 _8843_ (
    .CLK(clk_bF$buf3),
    .D(_841_),
    .Q(\genblk1[1].u_ce.Ycalc [2])
);

DFFPOSX1 _8844_ (
    .CLK(clk_bF$buf2),
    .D(_842_),
    .Q(\genblk1[1].u_ce.Ycalc [3])
);

DFFPOSX1 _8845_ (
    .CLK(clk_bF$buf1),
    .D(_843_),
    .Q(\genblk1[1].u_ce.Ycalc [4])
);

DFFPOSX1 _8846_ (
    .CLK(clk_bF$buf0),
    .D(_844_),
    .Q(\genblk1[1].u_ce.Ycalc [5])
);

DFFPOSX1 _8847_ (
    .CLK(clk_bF$buf78),
    .D(_845_),
    .Q(\genblk1[1].u_ce.Ycalc [6])
);

DFFPOSX1 _8848_ (
    .CLK(clk_bF$buf77),
    .D(_846_),
    .Q(\genblk1[1].u_ce.Ycalc [7])
);

DFFPOSX1 _8849_ (
    .CLK(clk_bF$buf76),
    .D(_847_),
    .Q(\genblk1[1].u_ce.Ycalc [8])
);

DFFPOSX1 _8850_ (
    .CLK(clk_bF$buf75),
    .D(_848_),
    .Q(\genblk1[1].u_ce.Ycalc [9])
);

DFFPOSX1 _8851_ (
    .CLK(clk_bF$buf74),
    .D(_849_),
    .Q(\genblk1[1].u_ce.Ycalc [10])
);

DFFPOSX1 _8852_ (
    .CLK(clk_bF$buf73),
    .D(_850_),
    .Q(\genblk1[1].u_ce.Ycalc [11])
);

DFFPOSX1 _8853_ (
    .CLK(clk_bF$buf72),
    .D(_851_),
    .Q(\genblk1[1].u_ce.Xcalc [0])
);

DFFPOSX1 _8854_ (
    .CLK(clk_bF$buf71),
    .D(_852_),
    .Q(\genblk1[1].u_ce.Xcalc [1])
);

DFFPOSX1 _8855_ (
    .CLK(clk_bF$buf70),
    .D(_853_),
    .Q(\genblk1[1].u_ce.Xcalc [2])
);

DFFPOSX1 _8856_ (
    .CLK(clk_bF$buf69),
    .D(_854_),
    .Q(\genblk1[1].u_ce.Xcalc [3])
);

DFFPOSX1 _8857_ (
    .CLK(clk_bF$buf68),
    .D(_855_),
    .Q(\genblk1[1].u_ce.Xcalc [4])
);

DFFPOSX1 _8858_ (
    .CLK(clk_bF$buf67),
    .D(_856_),
    .Q(\genblk1[1].u_ce.Xcalc [5])
);

DFFPOSX1 _8859_ (
    .CLK(clk_bF$buf66),
    .D(_857_),
    .Q(\genblk1[1].u_ce.Xcalc [6])
);

DFFPOSX1 _8860_ (
    .CLK(clk_bF$buf65),
    .D(_858_),
    .Q(\genblk1[1].u_ce.Xcalc [7])
);

DFFPOSX1 _8861_ (
    .CLK(clk_bF$buf64),
    .D(_859_),
    .Q(\genblk1[1].u_ce.Xcalc [8])
);

DFFPOSX1 _8862_ (
    .CLK(clk_bF$buf63),
    .D(_860_),
    .Q(\genblk1[1].u_ce.Xcalc [9])
);

DFFPOSX1 _8863_ (
    .CLK(clk_bF$buf62),
    .D(_861_),
    .Q(\genblk1[1].u_ce.Xcalc [10])
);

DFFPOSX1 _8864_ (
    .CLK(clk_bF$buf61),
    .D(_862_),
    .Q(\genblk1[1].u_ce.Xcalc [11])
);

DFFPOSX1 _8865_ (
    .CLK(clk_bF$buf60),
    .D(_863_),
    .Q(\genblk1[1].u_ce.Acalc [0])
);

DFFPOSX1 _8866_ (
    .CLK(clk_bF$buf59),
    .D(_864_),
    .Q(\genblk1[1].u_ce.Acalc [1])
);

DFFPOSX1 _8867_ (
    .CLK(clk_bF$buf58),
    .D(_865_),
    .Q(\genblk1[1].u_ce.Acalc [2])
);

DFFPOSX1 _8868_ (
    .CLK(clk_bF$buf57),
    .D(_866_),
    .Q(\genblk1[1].u_ce.Acalc [3])
);

DFFPOSX1 _8869_ (
    .CLK(clk_bF$buf56),
    .D(_867_),
    .Q(\genblk1[1].u_ce.Acalc [4])
);

DFFPOSX1 _8870_ (
    .CLK(clk_bF$buf55),
    .D(_868_),
    .Q(\genblk1[1].u_ce.Acalc [5])
);

DFFPOSX1 _8871_ (
    .CLK(clk_bF$buf54),
    .D(_869_),
    .Q(\genblk1[1].u_ce.Acalc [6])
);

DFFPOSX1 _8872_ (
    .CLK(clk_bF$buf53),
    .D(_870_),
    .Q(\genblk1[1].u_ce.Acalc [7])
);

DFFPOSX1 _8873_ (
    .CLK(clk_bF$buf52),
    .D(_871_),
    .Q(\genblk1[1].u_ce.Acalc [8])
);

DFFPOSX1 _8874_ (
    .CLK(clk_bF$buf51),
    .D(_872_),
    .Q(\genblk1[1].u_ce.Acalc [9])
);

DFFPOSX1 _8875_ (
    .CLK(clk_bF$buf50),
    .D(_873_),
    .Q(\genblk1[1].u_ce.Acalc [10])
);

DFFPOSX1 _8876_ (
    .CLK(clk_bF$buf49),
    .D(_874_),
    .Q(\genblk1[1].u_ce.Acalc [11])
);

DFFPOSX1 _8877_ (
    .CLK(clk_bF$buf48),
    .D(_875_),
    .Q(\genblk1[1].u_ce.Xin12b [10])
);

DFFPOSX1 _8878_ (
    .CLK(clk_bF$buf47),
    .D(_876_),
    .Q(\genblk1[1].u_ce.Xin12b [11])
);

DFFPOSX1 _8879_ (
    .CLK(clk_bF$buf46),
    .D(_877_),
    .Q(\genblk1[1].u_ce.Xin12b [8])
);

DFFPOSX1 _8880_ (
    .CLK(clk_bF$buf45),
    .D(_878_),
    .Q(\genblk1[1].u_ce.Xin12b [9])
);

DFFPOSX1 _8881_ (
    .CLK(clk_bF$buf44),
    .D(_879_),
    .Q(\genblk1[1].u_ce.Xin12b [6])
);

DFFPOSX1 _8882_ (
    .CLK(clk_bF$buf43),
    .D(_880_),
    .Q(\genblk1[1].u_ce.Xin12b [7])
);

DFFPOSX1 _8883_ (
    .CLK(clk_bF$buf42),
    .D(_881_),
    .Q(\genblk1[1].u_ce.Xin12b [4])
);

DFFPOSX1 _8884_ (
    .CLK(clk_bF$buf41),
    .D(_882_),
    .Q(\genblk1[1].u_ce.Xin12b [5])
);

DFFPOSX1 _8885_ (
    .CLK(clk_bF$buf40),
    .D(_883_),
    .Q(\genblk1[1].u_ce.Xin1 [0])
);

DFFPOSX1 _8886_ (
    .CLK(clk_bF$buf39),
    .D(_884_),
    .Q(\genblk1[1].u_ce.Xin1 [1])
);

DFFPOSX1 _8887_ (
    .CLK(clk_bF$buf38),
    .D(_885_),
    .Q(\genblk1[1].u_ce.Xin0 [0])
);

DFFPOSX1 _8888_ (
    .CLK(clk_bF$buf37),
    .D(_886_),
    .Q(\genblk1[1].u_ce.Xin0 [1])
);

DFFPOSX1 _8889_ (
    .CLK(clk_bF$buf36),
    .D(_887_),
    .Q(\genblk1[1].u_ce.Yin12b [10])
);

DFFPOSX1 _8890_ (
    .CLK(clk_bF$buf35),
    .D(_888_),
    .Q(\genblk1[1].u_ce.Yin12b [11])
);

DFFPOSX1 _8891_ (
    .CLK(clk_bF$buf34),
    .D(_889_),
    .Q(\genblk1[1].u_ce.Yin12b [8])
);

DFFPOSX1 _8892_ (
    .CLK(clk_bF$buf33),
    .D(_890_),
    .Q(\genblk1[1].u_ce.Yin12b [9])
);

DFFPOSX1 _8893_ (
    .CLK(clk_bF$buf32),
    .D(_891_),
    .Q(\genblk1[1].u_ce.Yin12b [6])
);

DFFPOSX1 _8894_ (
    .CLK(clk_bF$buf31),
    .D(_892_),
    .Q(\genblk1[1].u_ce.Yin12b [7])
);

DFFPOSX1 _8895_ (
    .CLK(clk_bF$buf30),
    .D(_893_),
    .Q(\genblk1[1].u_ce.Yin12b [4])
);

DFFPOSX1 _8896_ (
    .CLK(clk_bF$buf29),
    .D(_894_),
    .Q(\genblk1[1].u_ce.Yin12b [5])
);

DFFPOSX1 _8897_ (
    .CLK(clk_bF$buf28),
    .D(_895_),
    .Q(\genblk1[1].u_ce.Yin1 [0])
);

DFFPOSX1 _8898_ (
    .CLK(clk_bF$buf27),
    .D(_896_),
    .Q(\genblk1[1].u_ce.Yin1 [1])
);

DFFPOSX1 _8899_ (
    .CLK(clk_bF$buf26),
    .D(_897_),
    .Q(\genblk1[1].u_ce.Yin0 [0])
);

DFFPOSX1 _8900_ (
    .CLK(clk_bF$buf25),
    .D(_898_),
    .Q(\genblk1[1].u_ce.Yin0 [1])
);

DFFPOSX1 _8901_ (
    .CLK(clk_bF$buf24),
    .D(_899_),
    .Q(\genblk1[1].u_ce.Ain12b [10])
);

DFFPOSX1 _8902_ (
    .CLK(clk_bF$buf23),
    .D(_900_),
    .Q(\genblk1[1].u_ce.Ain12b [11])
);

DFFPOSX1 _8903_ (
    .CLK(clk_bF$buf22),
    .D(_901_),
    .Q(\genblk1[1].u_ce.Ain12b [8])
);

DFFPOSX1 _8904_ (
    .CLK(clk_bF$buf21),
    .D(_902_),
    .Q(\genblk1[1].u_ce.Ain12b [9])
);

DFFPOSX1 _8905_ (
    .CLK(clk_bF$buf20),
    .D(_903_),
    .Q(\genblk1[1].u_ce.Ain12b [6])
);

DFFPOSX1 _8906_ (
    .CLK(clk_bF$buf19),
    .D(_904_),
    .Q(\genblk1[1].u_ce.Ain12b [7])
);

DFFPOSX1 _8907_ (
    .CLK(clk_bF$buf18),
    .D(_905_),
    .Q(\genblk1[1].u_ce.Ain12b [4])
);

DFFPOSX1 _8908_ (
    .CLK(clk_bF$buf17),
    .D(_906_),
    .Q(\genblk1[1].u_ce.Ain12b [5])
);

DFFPOSX1 _8909_ (
    .CLK(clk_bF$buf16),
    .D(_907_),
    .Q(\genblk1[1].u_ce.Ain1 [0])
);

DFFPOSX1 _8910_ (
    .CLK(clk_bF$buf15),
    .D(_908_),
    .Q(\genblk1[1].u_ce.Ain1 [1])
);

DFFPOSX1 _8911_ (
    .CLK(clk_bF$buf14),
    .D(_909_),
    .Q(\genblk1[1].u_ce.Ain0 [0])
);

DFFPOSX1 _8912_ (
    .CLK(clk_bF$buf13),
    .D(_910_),
    .Q(\genblk1[1].u_ce.Ain0 [1])
);

DFFPOSX1 _8913_ (
    .CLK(clk_bF$buf12),
    .D(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[1].u_ce.LoadCtl [0])
);

DFFPOSX1 _8914_ (
    .CLK(clk_bF$buf11),
    .D(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[1].u_ce.LoadCtl [1])
);

DFFPOSX1 _8915_ (
    .CLK(clk_bF$buf10),
    .D(\genblk1[1].u_ce.LoadCtl [1]),
    .Q(\genblk1[1].u_ce.LoadCtl [2])
);

DFFPOSX1 _8916_ (
    .CLK(clk_bF$buf9),
    .D(\genblk1[1].u_ce.LoadCtl [2]),
    .Q(\genblk1[1].u_ce.LoadCtl [3])
);

DFFPOSX1 _8917_ (
    .CLK(clk_bF$buf8),
    .D(\genblk1[1].u_ce.LoadCtl [3]),
    .Q(\genblk1[1].u_ce.LoadCtl [4])
);

DFFPOSX1 _8918_ (
    .CLK(clk_bF$buf7),
    .D(\genblk1[1].u_ce.LoadCtl [4]),
    .Q(\genblk1[1].u_ce.LoadCtl [5])
);

DFFPOSX1 _8919_ (
    .CLK(clk_bF$buf6),
    .D(\genblk1[1].u_ce.LoadCtl [5]),
    .Q(\genblk1[1].u_ce.Vld )
);

INVX1 _8920_ (
    .A(\genblk1[2].u_ce.Acalc [2]),
    .Y(_1756_)
);

INVX2 _8921_ (
    .A(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1757_)
);

NOR2X1 _8922_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1757_),
    .Y(_1758_)
);

INVX2 _8923_ (
    .A(_1758_),
    .Y(_1759_)
);

NOR2X1 _8924_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [10]),
    .Y(_1760_)
);

INVX4 _8925_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .Y(_1761_)
);

NOR2X1 _8926_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.LoadCtl [3]),
    .Y(_1762_)
);

OAI21X1 _8927_ (
    .A(_1761_),
    .B(\genblk1[2].u_ce.Acalc [8]),
    .C(_1762_),
    .Y(_1763_)
);

INVX2 _8928_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_1764_)
);

AND2X2 _8929_ (
    .A(_1764_),
    .B(\genblk1[2].u_ce.LoadCtl [3]),
    .Y(_1765_)
);

AOI22X1 _8930_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.Acalc [4]),
    .C(_1765_),
    .D(\genblk1[2].u_ce.Acalc [6]),
    .Y(_1766_)
);

OAI21X1 _8931_ (
    .A(_1760_),
    .B(_1763_),
    .C(_1766_),
    .Y(_1767_)
);

NOR2X1 _8932_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1768_)
);

AOI22X1 _8933_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Acalc [0]),
    .C(_1767_),
    .D(_1768_),
    .Y(_1769_)
);

OAI21X1 _8934_ (
    .A(_1756_),
    .B(_1759_),
    .C(_1769_),
    .Y(\a[3] [0])
);

INVX1 _8935_ (
    .A(\genblk1[2].u_ce.Acalc [9]),
    .Y(_1770_)
);

OAI21X1 _8936_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [11]),
    .C(_1762_),
    .Y(_1771_)
);

AOI21X1 _8937_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1770_),
    .C(_1771_),
    .Y(_1772_)
);

INVX1 _8938_ (
    .A(\genblk1[2].u_ce.Acalc [5]),
    .Y(_1773_)
);

NAND2X1 _8939_ (
    .A(\genblk1[2].u_ce.Acalc [7]),
    .B(_1765_),
    .Y(_1774_)
);

OAI21X1 _8940_ (
    .A(_1764_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1775_)
);

OAI21X1 _8941_ (
    .A(_1772_),
    .B(_1775_),
    .C(_1768_),
    .Y(_1776_)
);

AOI22X1 _8942_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[2].u_ce.Acalc [1]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Acalc [3]),
    .Y(_1777_)
);

NAND2X1 _8943_ (
    .A(_1777_),
    .B(_1776_),
    .Y(\a[3] [1])
);

INVX1 _8944_ (
    .A(\genblk1[2].u_ce.Ycalc [10]),
    .Y(_1778_)
);

OAI21X1 _8945_ (
    .A(_1761_),
    .B(\genblk1[2].u_ce.Ycalc [8]),
    .C(_1762_),
    .Y(_1779_)
);

AOI21X1 _8946_ (
    .A(_1761_),
    .B(_1778_),
    .C(_1779_),
    .Y(_1780_)
);

INVX1 _8947_ (
    .A(\genblk1[2].u_ce.Ycalc [4]),
    .Y(_1781_)
);

NAND2X1 _8948_ (
    .A(\genblk1[2].u_ce.Ycalc [6]),
    .B(_1765_),
    .Y(_1782_)
);

OAI21X1 _8949_ (
    .A(_1764_),
    .B(_1781_),
    .C(_1782_),
    .Y(_1783_)
);

OAI21X1 _8950_ (
    .A(_1780_),
    .B(_1783_),
    .C(_1768_),
    .Y(_1784_)
);

AOI22X1 _8951_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.Ycalc [0]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Ycalc [2]),
    .Y(_1785_)
);

NAND2X1 _8952_ (
    .A(_1785_),
    .B(_1784_),
    .Y(\genblk1[2].u_ce.Y_ [0])
);

INVX1 _8953_ (
    .A(\genblk1[2].u_ce.Ycalc [9]),
    .Y(_1786_)
);

OAI21X1 _8954_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Ycalc [11]),
    .C(_1762_),
    .Y(_1787_)
);

AOI21X1 _8955_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1786_),
    .C(_1787_),
    .Y(_1788_)
);

INVX1 _8956_ (
    .A(\genblk1[2].u_ce.Ycalc [5]),
    .Y(_1789_)
);

NAND2X1 _8957_ (
    .A(\genblk1[2].u_ce.Ycalc [7]),
    .B(_1765_),
    .Y(_1790_)
);

OAI21X1 _8958_ (
    .A(_1764_),
    .B(_1789_),
    .C(_1790_),
    .Y(_1791_)
);

OAI21X1 _8959_ (
    .A(_1788_),
    .B(_1791_),
    .C(_1768_),
    .Y(_1792_)
);

AOI22X1 _8960_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[2].u_ce.Ycalc [1]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1793_)
);

NAND2X1 _8961_ (
    .A(_1793_),
    .B(_1792_),
    .Y(\genblk1[2].u_ce.Y_ [1])
);

INVX1 _8962_ (
    .A(\genblk1[2].u_ce.Xcalc [8]),
    .Y(_1794_)
);

OAI21X1 _8963_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Xcalc [10]),
    .C(_1762_),
    .Y(_1795_)
);

AOI21X1 _8964_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1794_),
    .C(_1795_),
    .Y(_1796_)
);

INVX1 _8965_ (
    .A(\genblk1[2].u_ce.Xcalc [4]),
    .Y(_1797_)
);

NAND2X1 _8966_ (
    .A(\genblk1[2].u_ce.Xcalc [6]),
    .B(_1765_),
    .Y(_1798_)
);

OAI21X1 _8967_ (
    .A(_1764_),
    .B(_1797_),
    .C(_1798_),
    .Y(_1799_)
);

OAI21X1 _8968_ (
    .A(_1796_),
    .B(_1799_),
    .C(_1768_),
    .Y(_1800_)
);

AOI22X1 _8969_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[2].u_ce.Xcalc [0]),
    .C(_1758_),
    .D(\genblk1[2].u_ce.Xcalc [2]),
    .Y(_1801_)
);

NAND2X1 _8970_ (
    .A(_1801_),
    .B(_1800_),
    .Y(\genblk1[2].u_ce.X_ [0])
);

INVX1 _8971_ (
    .A(\genblk1[2].u_ce.Xcalc [3]),
    .Y(_1802_)
);

NOR2X1 _8972_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Xcalc [11]),
    .Y(_1803_)
);

OAI21X1 _8973_ (
    .A(_1761_),
    .B(\genblk1[2].u_ce.Xcalc [9]),
    .C(_1762_),
    .Y(_1804_)
);

AOI22X1 _8974_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.Xcalc [5]),
    .C(_1765_),
    .D(\genblk1[2].u_ce.Xcalc [7]),
    .Y(_1805_)
);

OAI21X1 _8975_ (
    .A(_1803_),
    .B(_1804_),
    .C(_1805_),
    .Y(_1806_)
);

AOI22X1 _8976_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Xcalc [1]),
    .C(_1806_),
    .D(_1768_),
    .Y(_1807_)
);

OAI21X1 _8977_ (
    .A(_1802_),
    .B(_1759_),
    .C(_1807_),
    .Y(\genblk1[2].u_ce.X_ [1])
);

INVX1 _8978_ (
    .A(\genblk1[2].u_ce.Ycalc [0]),
    .Y(_1808_)
);

INVX1 _8979_ (
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .Y(_1809_)
);

INVX8 _8980_ (
    .A(1'h0),
    .Y(_1810_)
);

INVX8 _8981_ (
    .A(1'h1),
    .Y(_1811_)
);

INVX1 _8982_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_1812_)
);

NAND2X1 _8983_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1813_)
);

OAI21X1 _8984_ (
    .A(1'h0),
    .B(_1812_),
    .C(_1813_),
    .Y(_1814_)
);

INVX1 _8985_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .Y(_1815_)
);

NAND2X1 _8986_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1816_)
);

OAI21X1 _8987_ (
    .A(1'h0),
    .B(_1815_),
    .C(_1816_),
    .Y(_1817_)
);

MUX2X1 _8988_ (
    .A(_1817_),
    .B(_1814_),
    .S(_1811__bF$buf4),
    .Y(_1818_)
);

INVX1 _8989_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1819_)
);

NAND2X1 _8990_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1820_)
);

OAI21X1 _8991_ (
    .A(1'h0),
    .B(_1819_),
    .C(_1820_),
    .Y(_1821_)
);

INVX1 _8992_ (
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .Y(_1822_)
);

NAND2X1 _8993_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_1823_)
);

OAI21X1 _8994_ (
    .A(1'h0),
    .B(_1822_),
    .C(_1823_),
    .Y(_1824_)
);

MUX2X1 _8995_ (
    .A(_1824_),
    .B(_1821_),
    .S(_1811__bF$buf3),
    .Y(_1825_)
);

MUX2X1 _8996_ (
    .A(_1825_),
    .B(_1818_),
    .S(_1810__bF$buf4),
    .Y(_1826_)
);

NOR2X1 _8997_ (
    .A(_1809_),
    .B(_1826_),
    .Y(_1827_)
);

NAND2X1 _8998_ (
    .A(_1809_),
    .B(_1826_),
    .Y(_1828_)
);

INVX1 _8999_ (
    .A(_1828_),
    .Y(_1829_)
);

NAND2X1 _9000_ (
    .A(_1810__bF$buf3),
    .B(_1811__bF$buf2),
    .Y(_1830_)
);

OAI21X1 _9001_ (
    .A(1'h0),
    .B(_1830_),
    .C(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .Y(_1831_)
);

INVX2 _9002_ (
    .A(_1831_),
    .Y(_1832_)
);

OAI21X1 _9003_ (
    .A(_1827_),
    .B(_1829_),
    .C(_1832_),
    .Y(_1833_)
);

OAI21X1 _9004_ (
    .A(_1808_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_1833_),
    .Y(_1676_)
);

INVX8 _9005_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_1834_)
);

NAND2X1 _9006_ (
    .A(\genblk1[2].u_ce.Ycalc [1]),
    .B(_1834__bF$buf4),
    .Y(_1835_)
);

NOR2X1 _9007_ (
    .A(1'h0),
    .B(_1830_),
    .Y(_1836_)
);

MUX2X1 _9008_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(\genblk1[2].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_1837_)
);

MUX2X1 _9009_ (
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .B(\genblk1[2].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_1838_)
);

MUX2X1 _9010_ (
    .A(_1838_),
    .B(_1837_),
    .S(_1811__bF$buf1),
    .Y(_1839_)
);

INVX2 _9011_ (
    .A(1'h0),
    .Y(_1840_)
);

NAND2X1 _9012_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(_1840_),
    .Y(_1841_)
);

AOI21X1 _9013_ (
    .A(_1841_),
    .B(_1820_),
    .C(_1811__bF$buf0),
    .Y(_1842_)
);

NAND3X1 _9014_ (
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .B(_1840_),
    .C(_1811__bF$buf4),
    .Y(_1843_)
);

NAND3X1 _9015_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(1'h0),
    .C(_1811__bF$buf3),
    .Y(_1844_)
);

NAND3X1 _9016_ (
    .A(_1810__bF$buf2),
    .B(_1844_),
    .C(_1843_),
    .Y(_1845_)
);

OAI22X1 _9017_ (
    .A(_1842_),
    .B(_1845_),
    .C(_1810__bF$buf1),
    .D(_1839_),
    .Y(_1846_)
);

INVX1 _9018_ (
    .A(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_1847_)
);

INVX8 _9019_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1848_)
);

INVX1 _9020_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1849_)
);

NAND2X1 _9021_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_1850_)
);

OAI21X1 _9022_ (
    .A(1'h0),
    .B(_1849_),
    .C(_1850_),
    .Y(_1851_)
);

INVX1 _9023_ (
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1852_)
);

NAND2X1 _9024_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_1853_)
);

OAI21X1 _9025_ (
    .A(1'h0),
    .B(_1852_),
    .C(_1853_),
    .Y(_1854_)
);

MUX2X1 _9026_ (
    .A(_1854_),
    .B(_1851_),
    .S(_1811__bF$buf2),
    .Y(_1855_)
);

INVX1 _9027_ (
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1856_)
);

NAND2X1 _9028_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [4]),
    .Y(_1857_)
);

OAI21X1 _9029_ (
    .A(1'h0),
    .B(_1856_),
    .C(_1857_),
    .Y(_1858_)
);

INVX1 _9030_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .Y(_1859_)
);

NAND2X1 _9031_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1860_)
);

OAI21X1 _9032_ (
    .A(1'h0),
    .B(_1859_),
    .C(_1860_),
    .Y(_1861_)
);

MUX2X1 _9033_ (
    .A(_1861_),
    .B(_1858_),
    .S(_1811__bF$buf1),
    .Y(_1862_)
);

MUX2X1 _9034_ (
    .A(_1862_),
    .B(_1855_),
    .S(_1810__bF$buf0),
    .Y(_1863_)
);

NAND3X1 _9035_ (
    .A(_1848__bF$buf5),
    .B(_1826_),
    .C(_1863_),
    .Y(_1864_)
);

MUX2X1 _9036_ (
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_1865_)
);

MUX2X1 _9037_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_1866_)
);

MUX2X1 _9038_ (
    .A(_1866_),
    .B(_1865_),
    .S(_1811__bF$buf0),
    .Y(_1867_)
);

MUX2X1 _9039_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_1868_)
);

MUX2X1 _9040_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(\genblk1[2].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_1869_)
);

MUX2X1 _9041_ (
    .A(_1869_),
    .B(_1868_),
    .S(_1811__bF$buf4),
    .Y(_1870_)
);

MUX2X1 _9042_ (
    .A(_1870_),
    .B(_1867_),
    .S(_1810__bF$buf4),
    .Y(_1871_)
);

OAI21X1 _9043_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1846_),
    .C(_1871_),
    .Y(_1872_)
);

AOI21X1 _9044_ (
    .A(_1872_),
    .B(_1864_),
    .C(_1847_),
    .Y(_1873_)
);

INVX1 _9045_ (
    .A(_1873_),
    .Y(_1874_)
);

NAND3X1 _9046_ (
    .A(_1847_),
    .B(_1864_),
    .C(_1872_),
    .Y(_1875_)
);

AND2X2 _9047_ (
    .A(_1874_),
    .B(_1875_),
    .Y(_1876_)
);

OAI21X1 _9048_ (
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .B(_1846_),
    .C(_1876_),
    .Y(_1877_)
);

OR2X2 _9049_ (
    .A(_1876_),
    .B(_1828_),
    .Y(_1878_)
);

AOI21X1 _9050_ (
    .A(_1878_),
    .B(_1877_),
    .C(_1836_),
    .Y(_1879_)
);

OAI21X1 _9051_ (
    .A(_1834__bF$buf3),
    .B(_1879_),
    .C(_1835_),
    .Y(_1677_)
);

INVX1 _9052_ (
    .A(\genblk1[2].u_ce.ISout ),
    .Y(_1880_)
);

NAND2X1 _9053_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .B(\genblk1[1].u_ce.ISout ),
    .Y(_1881_)
);

OAI21X1 _9054_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_1880_),
    .C(_1881_),
    .Y(_1678_)
);

NAND2X1 _9055_ (
    .A(\genblk1[2].u_ce.Ycalc [2]),
    .B(_1834__bF$buf2),
    .Y(_1882_)
);

AOI21X1 _9056_ (
    .A(_1828_),
    .B(_1875_),
    .C(_1873_),
    .Y(_1883_)
);

MUX2X1 _9057_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(\genblk1[2].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_1884_)
);

MUX2X1 _9058_ (
    .A(_1884_),
    .B(_1837_),
    .S(1'h1),
    .Y(_1885_)
);

MUX2X1 _9059_ (
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_1886_)
);

NAND2X1 _9060_ (
    .A(1'h1),
    .B(_1810__bF$buf3),
    .Y(_1887_)
);

OAI22X1 _9061_ (
    .A(_1887_),
    .B(_1838_),
    .C(_1886_),
    .D(_1830_),
    .Y(_1888_)
);

AOI21X1 _9062_ (
    .A(1'h0),
    .B(_1885_),
    .C(_1888_),
    .Y(_1889_)
);

AOI21X1 _9063_ (
    .A(_1871_),
    .B(_1846_),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_1890_)
);

NAND2X1 _9064_ (
    .A(_1889_),
    .B(_1890_),
    .Y(_1891_)
);

INVX1 _9065_ (
    .A(_1889_),
    .Y(_1892_)
);

OAI21X1 _9066_ (
    .A(_1826_),
    .B(_1863_),
    .C(_1848__bF$buf4),
    .Y(_1893_)
);

NAND2X1 _9067_ (
    .A(_1892_),
    .B(_1893_),
    .Y(_1894_)
);

AOI21X1 _9068_ (
    .A(_1894_),
    .B(_1891_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_1895_)
);

NAND3X1 _9069_ (
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .B(_1891_),
    .C(_1894_),
    .Y(_1896_)
);

INVX1 _9070_ (
    .A(_1896_),
    .Y(_1897_)
);

OR2X2 _9071_ (
    .A(_1897_),
    .B(_1895_),
    .Y(_1898_)
);

NOR2X1 _9072_ (
    .A(_1883_),
    .B(_1898_),
    .Y(_1899_)
);

INVX1 _9073_ (
    .A(_1899_),
    .Y(_1900_)
);

OAI21X1 _9074_ (
    .A(_1895_),
    .B(_1897_),
    .C(_1883_),
    .Y(_1901_)
);

AOI21X1 _9075_ (
    .A(_1900_),
    .B(_1901_),
    .C(_1836_),
    .Y(_1902_)
);

INVX2 _9076_ (
    .A(_1836_),
    .Y(_1903_)
);

OAI21X1 _9077_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1903_),
    .C(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .Y(_1904_)
);

OAI21X1 _9078_ (
    .A(_1904_),
    .B(_1902_),
    .C(_1882_),
    .Y(_1679_)
);

INVX1 _9079_ (
    .A(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1905_)
);

INVX2 _9080_ (
    .A(_1904_),
    .Y(_1906_)
);

OAI21X1 _9081_ (
    .A(_1895_),
    .B(_1883_),
    .C(_1896_),
    .Y(_1907_)
);

INVX1 _9082_ (
    .A(_1907_),
    .Y(_1908_)
);

INVX1 _9083_ (
    .A(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_1909_)
);

NAND3X1 _9084_ (
    .A(_1846_),
    .B(_1871_),
    .C(_1889_),
    .Y(_1910_)
);

INVX1 _9085_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .Y(_1911_)
);

NAND2X1 _9086_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_1912_)
);

OAI21X1 _9087_ (
    .A(1'h0),
    .B(_1911_),
    .C(_1912_),
    .Y(_1913_)
);

NAND2X1 _9088_ (
    .A(_1811__bF$buf3),
    .B(_1865_),
    .Y(_1914_)
);

OAI21X1 _9089_ (
    .A(_1811__bF$buf2),
    .B(_1913_),
    .C(_1914_),
    .Y(_1915_)
);

NOR2X1 _9090_ (
    .A(1'h0),
    .B(_1811__bF$buf1),
    .Y(_1916_)
);

NOR2X1 _9091_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_1917_)
);

AOI22X1 _9092_ (
    .A(_1858_),
    .B(_1917_),
    .C(_1916_),
    .D(_1854_),
    .Y(_1918_)
);

OAI21X1 _9093_ (
    .A(_1810__bF$buf2),
    .B(_1915_),
    .C(_1918_),
    .Y(_1919_)
);

NAND3X1 _9094_ (
    .A(_1848__bF$buf3),
    .B(_1919_),
    .C(_1910_),
    .Y(_1920_)
);

INVX1 _9095_ (
    .A(_1910_),
    .Y(_1921_)
);

INVX1 _9096_ (
    .A(_1919_),
    .Y(_1922_)
);

OAI21X1 _9097_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1921_),
    .C(_1922_),
    .Y(_1923_)
);

NAND3X1 _9098_ (
    .A(_1909_),
    .B(_1920_),
    .C(_1923_),
    .Y(_1924_)
);

AOI21X1 _9099_ (
    .A(_1923_),
    .B(_1920_),
    .C(_1909_),
    .Y(_1925_)
);

INVX1 _9100_ (
    .A(_1925_),
    .Y(_1926_)
);

NAND2X1 _9101_ (
    .A(_1924_),
    .B(_1926_),
    .Y(_1927_)
);

AOI21X1 _9102_ (
    .A(_1927_),
    .B(_1908_),
    .C(_1836_),
    .Y(_1928_)
);

OAI21X1 _9103_ (
    .A(_1908_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_)
);

AOI22X1 _9104_ (
    .A(_1905_),
    .B(_1834__bF$buf1),
    .C(_1929_),
    .D(_1906_),
    .Y(_1680_)
);

AOI21X1 _9105_ (
    .A(_1907_),
    .B(_1924_),
    .C(_1925_),
    .Y(_1930_)
);

INVX1 _9106_ (
    .A(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_1931_)
);

INVX1 _9107_ (
    .A(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_1932_)
);

NAND2X1 _9108_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_1933_)
);

OAI21X1 _9109_ (
    .A(1'h0),
    .B(_1932_),
    .C(_1933_),
    .Y(_1934_)
);

NAND2X1 _9110_ (
    .A(_1811__bF$buf0),
    .B(_1884_),
    .Y(_1935_)
);

OAI21X1 _9111_ (
    .A(_1811__bF$buf4),
    .B(_1934_),
    .C(_1935_),
    .Y(_1936_)
);

NAND2X1 _9112_ (
    .A(_1810__bF$buf1),
    .B(_1839_),
    .Y(_1937_)
);

OAI21X1 _9113_ (
    .A(_1810__bF$buf0),
    .B(_1936_),
    .C(_1937_),
    .Y(_1938_)
);

INVX2 _9114_ (
    .A(_1938_),
    .Y(_1939_)
);

OAI21X1 _9115_ (
    .A(_1919_),
    .B(_1910_),
    .C(_1848__bF$buf2),
    .Y(_1940_)
);

OR2X2 _9116_ (
    .A(_1940_),
    .B(_1939_),
    .Y(_1941_)
);

NOR2X1 _9117_ (
    .A(_1919_),
    .B(_1910_),
    .Y(_1942_)
);

OAI21X1 _9118_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1942_),
    .C(_1939_),
    .Y(_1943_)
);

NAND3X1 _9119_ (
    .A(_1931_),
    .B(_1943_),
    .C(_1941_),
    .Y(_1944_)
);

NOR2X1 _9120_ (
    .A(_1939_),
    .B(_1940_),
    .Y(_1945_)
);

AND2X2 _9121_ (
    .A(_1940_),
    .B(_1939_),
    .Y(_1946_)
);

OAI21X1 _9122_ (
    .A(_1945_),
    .B(_1946_),
    .C(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_1947_)
);

NAND2X1 _9123_ (
    .A(_1947_),
    .B(_1944_),
    .Y(_1948_)
);

AOI21X1 _9124_ (
    .A(_1930_),
    .B(_1948_),
    .C(_1836_),
    .Y(_1949_)
);

OAI21X1 _9125_ (
    .A(_1930_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1950_)
);

AOI22X1 _9126_ (
    .A(_1781_),
    .B(_1834__bF$buf0),
    .C(_1950_),
    .D(_1906_),
    .Y(_1681_)
);

OAI21X1 _9127_ (
    .A(_1948_),
    .B(_1930_),
    .C(_1947_),
    .Y(_1951_)
);

INVX1 _9128_ (
    .A(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_1952_)
);

NAND3X1 _9129_ (
    .A(_1922_),
    .B(_1939_),
    .C(_1921_),
    .Y(_1953_)
);

NAND2X1 _9130_ (
    .A(1'h1),
    .B(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_1954_)
);

INVX1 _9131_ (
    .A(_1954_),
    .Y(_1955_)
);

AOI21X1 _9132_ (
    .A(_1913_),
    .B(_1811__bF$buf3),
    .C(_1955_),
    .Y(_1956_)
);

NAND2X1 _9133_ (
    .A(_1810__bF$buf4),
    .B(_1867_),
    .Y(_1957_)
);

OAI21X1 _9134_ (
    .A(_1810__bF$buf3),
    .B(_1956_),
    .C(_1957_),
    .Y(_1958_)
);

NAND3X1 _9135_ (
    .A(_1848__bF$buf1),
    .B(_1958_),
    .C(_1953_),
    .Y(_1959_)
);

NOR3X1 _9136_ (
    .A(_1919_),
    .B(_1938_),
    .C(_1910_),
    .Y(_1960_)
);

INVX1 _9137_ (
    .A(_1958_),
    .Y(_1961_)
);

OAI21X1 _9138_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1960_),
    .C(_1961_),
    .Y(_1962_)
);

NAND3X1 _9139_ (
    .A(_1952_),
    .B(_1959_),
    .C(_1962_),
    .Y(_1963_)
);

AOI21X1 _9140_ (
    .A(_1962_),
    .B(_1959_),
    .C(_1952_),
    .Y(_1964_)
);

INVX1 _9141_ (
    .A(_1964_),
    .Y(_1965_)
);

NAND2X1 _9142_ (
    .A(_1963_),
    .B(_1965_),
    .Y(_1966_)
);

AND2X2 _9143_ (
    .A(_1951_),
    .B(_1966_),
    .Y(_1967_)
);

OAI21X1 _9144_ (
    .A(_1966_),
    .B(_1951_),
    .C(_1903_),
    .Y(_1968_)
);

OAI21X1 _9145_ (
    .A(_1968_),
    .B(_1967_),
    .C(_1906_),
    .Y(_1969_)
);

OAI21X1 _9146_ (
    .A(_1789_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_1969_),
    .Y(_1682_)
);

INVX1 _9147_ (
    .A(\genblk1[2].u_ce.Ycalc [6]),
    .Y(_1970_)
);

INVX1 _9148_ (
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_1971_)
);

NAND3X1 _9149_ (
    .A(_1939_),
    .B(_1961_),
    .C(_1942_),
    .Y(_1972_)
);

AOI21X1 _9150_ (
    .A(_1934_),
    .B(_1811__bF$buf2),
    .C(_1955_),
    .Y(_1973_)
);

NAND2X1 _9151_ (
    .A(_1810__bF$buf2),
    .B(_1885_),
    .Y(_1974_)
);

OAI21X1 _9152_ (
    .A(_1810__bF$buf1),
    .B(_1973_),
    .C(_1974_),
    .Y(_1975_)
);

NAND3X1 _9153_ (
    .A(_1848__bF$buf0),
    .B(_1975_),
    .C(_1972_),
    .Y(_1976_)
);

INVX1 _9154_ (
    .A(_1975_),
    .Y(_1977_)
);

OAI21X1 _9155_ (
    .A(_1958_),
    .B(_1953_),
    .C(_1848__bF$buf5),
    .Y(_1978_)
);

NAND2X1 _9156_ (
    .A(_1977_),
    .B(_1978_),
    .Y(_1979_)
);

NAND3X1 _9157_ (
    .A(_1971_),
    .B(_1976_),
    .C(_1979_),
    .Y(_1980_)
);

NAND3X1 _9158_ (
    .A(_1848__bF$buf4),
    .B(_1977_),
    .C(_1972_),
    .Y(_1981_)
);

NAND2X1 _9159_ (
    .A(_1975_),
    .B(_1978_),
    .Y(_1982_)
);

NAND3X1 _9160_ (
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .B(_1981_),
    .C(_1982_),
    .Y(_1983_)
);

NAND2X1 _9161_ (
    .A(_1980_),
    .B(_1983_),
    .Y(_1984_)
);

AOI21X1 _9162_ (
    .A(_1941_),
    .B(_1943_),
    .C(_1931_),
    .Y(_1985_)
);

NOR2X1 _9163_ (
    .A(_1985_),
    .B(_1964_),
    .Y(_1986_)
);

OAI21X1 _9164_ (
    .A(_1948_),
    .B(_1930_),
    .C(_1986_),
    .Y(_1987_)
);

NAND2X1 _9165_ (
    .A(_1963_),
    .B(_1987_),
    .Y(_1988_)
);

AOI21X1 _9166_ (
    .A(_1988_),
    .B(_1984_),
    .C(_1836_),
    .Y(_1989_)
);

OAI21X1 _9167_ (
    .A(_1984_),
    .B(_1988_),
    .C(_1989_),
    .Y(_1990_)
);

AOI22X1 _9168_ (
    .A(_1970_),
    .B(_1834__bF$buf4),
    .C(_1990_),
    .D(_1906_),
    .Y(_1683_)
);

INVX1 _9169_ (
    .A(\genblk1[2].u_ce.Ycalc [7]),
    .Y(_1991_)
);

AOI21X1 _9170_ (
    .A(_1979_),
    .B(_1976_),
    .C(_1971_),
    .Y(_1992_)
);

AND2X2 _9171_ (
    .A(_1944_),
    .B(_1947_),
    .Y(_1993_)
);

NAND3X1 _9172_ (
    .A(_1963_),
    .B(_1965_),
    .C(_1993_),
    .Y(_1994_)
);

AOI21X1 _9173_ (
    .A(_1985_),
    .B(_1963_),
    .C(_1964_),
    .Y(_1995_)
);

OAI21X1 _9174_ (
    .A(_1930_),
    .B(_1994_),
    .C(_1995_),
    .Y(_1996_)
);

AOI21X1 _9175_ (
    .A(_1996_),
    .B(_1980_),
    .C(_1992_),
    .Y(_1997_)
);

INVX1 _9176_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_1998_)
);

NAND3X1 _9177_ (
    .A(_1961_),
    .B(_1977_),
    .C(_1960_),
    .Y(_1999_)
);

INVX1 _9178_ (
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_2000_)
);

NOR2X1 _9179_ (
    .A(_1810__bF$buf0),
    .B(_2000_),
    .Y(_2001_)
);

INVX1 _9180_ (
    .A(_2001_),
    .Y(_2002_)
);

OAI21X1 _9181_ (
    .A(1'h0),
    .B(_1915_),
    .C(_2002_),
    .Y(_2003_)
);

NAND3X1 _9182_ (
    .A(_1848__bF$buf3),
    .B(_2003_),
    .C(_1999_),
    .Y(_2004_)
);

INVX1 _9183_ (
    .A(_2003_),
    .Y(_2005_)
);

OAI21X1 _9184_ (
    .A(_1975_),
    .B(_1972_),
    .C(_1848__bF$buf2),
    .Y(_2006_)
);

NAND2X1 _9185_ (
    .A(_2005_),
    .B(_2006_),
    .Y(_2007_)
);

NAND3X1 _9186_ (
    .A(_1998_),
    .B(_2004_),
    .C(_2007_),
    .Y(_2008_)
);

NAND3X1 _9187_ (
    .A(_1848__bF$buf1),
    .B(_2005_),
    .C(_1999_),
    .Y(_2009_)
);

NAND2X1 _9188_ (
    .A(_2003_),
    .B(_2006_),
    .Y(_2010_)
);

NAND3X1 _9189_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(_2009_),
    .C(_2010_),
    .Y(_2011_)
);

NAND2X1 _9190_ (
    .A(_2008_),
    .B(_2011_),
    .Y(_2012_)
);

INVX1 _9191_ (
    .A(_2012_),
    .Y(_2013_)
);

NOR2X1 _9192_ (
    .A(_2013_),
    .B(_1997_),
    .Y(_2014_)
);

OAI21X1 _9193_ (
    .A(_1984_),
    .B(_1988_),
    .C(_1983_),
    .Y(_2015_)
);

OAI21X1 _9194_ (
    .A(_2012_),
    .B(_2015_),
    .C(_1903_),
    .Y(_2016_)
);

OAI21X1 _9195_ (
    .A(_1848__bF$buf0),
    .B(_1903_),
    .C(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2017_)
);

INVX1 _9196_ (
    .A(_2017_),
    .Y(_2018_)
);

OAI21X1 _9197_ (
    .A(_2016_),
    .B(_2014_),
    .C(_2018_),
    .Y(_2019_)
);

OAI21X1 _9198_ (
    .A(_1991_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2019_),
    .Y(_1684_)
);

INVX1 _9199_ (
    .A(\genblk1[2].u_ce.Ycalc [8]),
    .Y(_2020_)
);

OAI21X1 _9200_ (
    .A(_1983_),
    .B(_2012_),
    .C(_2011_),
    .Y(_2021_)
);

NOR2X1 _9201_ (
    .A(_1984_),
    .B(_2012_),
    .Y(_2022_)
);

AOI21X1 _9202_ (
    .A(_2022_),
    .B(_1996_),
    .C(_2021_),
    .Y(_2023_)
);

INVX1 _9203_ (
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2024_)
);

OR2X2 _9204_ (
    .A(_1999_),
    .B(_2003_),
    .Y(_2025_)
);

OAI21X1 _9205_ (
    .A(1'h0),
    .B(_1936_),
    .C(_2002_),
    .Y(_2026_)
);

NAND3X1 _9206_ (
    .A(_1848__bF$buf5),
    .B(_2026_),
    .C(_2025_),
    .Y(_2027_)
);

NOR2X1 _9207_ (
    .A(_2003_),
    .B(_1999_),
    .Y(_2028_)
);

INVX1 _9208_ (
    .A(_2026_),
    .Y(_2029_)
);

OAI21X1 _9209_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2028_),
    .C(_2029_),
    .Y(_2030_)
);

NAND3X1 _9210_ (
    .A(_2024_),
    .B(_2030_),
    .C(_2027_),
    .Y(_2031_)
);

NAND3X1 _9211_ (
    .A(_1848__bF$buf4),
    .B(_2029_),
    .C(_2025_),
    .Y(_2032_)
);

OAI21X1 _9212_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2028_),
    .C(_2026_),
    .Y(_2033_)
);

NAND3X1 _9213_ (
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .B(_2033_),
    .C(_2032_),
    .Y(_2034_)
);

AND2X2 _9214_ (
    .A(_2031_),
    .B(_2034_),
    .Y(_2035_)
);

INVX1 _9215_ (
    .A(_2035_),
    .Y(_2036_)
);

AOI21X1 _9216_ (
    .A(_2023_),
    .B(_2036_),
    .C(_1836_),
    .Y(_2037_)
);

OAI21X1 _9217_ (
    .A(_2023_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_)
);

AOI22X1 _9218_ (
    .A(_2020_),
    .B(_1834__bF$buf3),
    .C(_2038_),
    .D(_2018_),
    .Y(_1685_)
);

NAND2X1 _9219_ (
    .A(_1992_),
    .B(_2008_),
    .Y(_2039_)
);

AND2X2 _9220_ (
    .A(_2039_),
    .B(_2011_),
    .Y(_2040_)
);

AND2X2 _9221_ (
    .A(_1980_),
    .B(_1983_),
    .Y(_2041_)
);

NAND3X1 _9222_ (
    .A(_2008_),
    .B(_2011_),
    .C(_2041_),
    .Y(_2042_)
);

OAI21X1 _9223_ (
    .A(_1988_),
    .B(_2042_),
    .C(_2040_),
    .Y(_2043_)
);

INVX1 _9224_ (
    .A(_2034_),
    .Y(_2044_)
);

AOI21X1 _9225_ (
    .A(_2043_),
    .B(_2031_),
    .C(_2044_),
    .Y(_2045_)
);

INVX1 _9226_ (
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2046_)
);

NOR3X1 _9227_ (
    .A(_2003_),
    .B(_2026_),
    .C(_1999_),
    .Y(_2047_)
);

INVX1 _9228_ (
    .A(_2047_),
    .Y(_2048_)
);

OAI21X1 _9229_ (
    .A(1'h0),
    .B(_1956_),
    .C(_2002_),
    .Y(_2049_)
);

NAND3X1 _9230_ (
    .A(_1848__bF$buf3),
    .B(_2049_),
    .C(_2048_),
    .Y(_2050_)
);

INVX1 _9231_ (
    .A(_2049_),
    .Y(_2051_)
);

OAI21X1 _9232_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2047_),
    .C(_2051_),
    .Y(_2052_)
);

NAND3X1 _9233_ (
    .A(_2046_),
    .B(_2052_),
    .C(_2050_),
    .Y(_2053_)
);

NAND3X1 _9234_ (
    .A(_1848__bF$buf2),
    .B(_2051_),
    .C(_2048_),
    .Y(_2054_)
);

OAI21X1 _9235_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2047_),
    .C(_2049_),
    .Y(_2055_)
);

NAND3X1 _9236_ (
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .B(_2055_),
    .C(_2054_),
    .Y(_2056_)
);

AND2X2 _9237_ (
    .A(_2053_),
    .B(_2056_),
    .Y(_2057_)
);

AND2X2 _9238_ (
    .A(_2045_),
    .B(_2057_),
    .Y(_2058_)
);

OAI21X1 _9239_ (
    .A(_2057_),
    .B(_2045_),
    .C(_1903_),
    .Y(_2059_)
);

OAI21X1 _9240_ (
    .A(_2059_),
    .B(_2058_),
    .C(_1906_),
    .Y(_2060_)
);

OAI21X1 _9241_ (
    .A(_1786_),
    .B(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .C(_2060_),
    .Y(_1686_)
);

INVX1 _9242_ (
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .Y(_2061_)
);

OAI21X1 _9243_ (
    .A(1'h0),
    .B(_1973_),
    .C(_2002_),
    .Y(_2062_)
);

INVX1 _9244_ (
    .A(_2062_),
    .Y(_2063_)
);

AOI21X1 _9245_ (
    .A(_2047_),
    .B(_2051_),
    .C(_2063_),
    .Y(_2064_)
);

NAND3X1 _9246_ (
    .A(_2051_),
    .B(_2063_),
    .C(_2047_),
    .Y(_2065_)
);

NAND2X1 _9247_ (
    .A(_1848__bF$buf1),
    .B(_2065_),
    .Y(_2066_)
);

NAND2X1 _9248_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2062_),
    .Y(_2067_)
);

OAI21X1 _9249_ (
    .A(_2064_),
    .B(_2066_),
    .C(_2067_),
    .Y(_2068_)
);

NAND2X1 _9250_ (
    .A(_2061_),
    .B(_2068_),
    .Y(_2069_)
);

INVX1 _9251_ (
    .A(_2064_),
    .Y(_2070_)
);

AND2X2 _9252_ (
    .A(_2065_),
    .B(_1848__bF$buf0),
    .Y(_2071_)
);

NAND2X1 _9253_ (
    .A(_2070_),
    .B(_2071_),
    .Y(_2072_)
);

NAND3X1 _9254_ (
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .B(_2067_),
    .C(_2072_),
    .Y(_2073_)
);

NAND2X1 _9255_ (
    .A(_2069_),
    .B(_2073_),
    .Y(_2074_)
);

AOI21X1 _9256_ (
    .A(_2050_),
    .B(_2052_),
    .C(_2046_),
    .Y(_2075_)
);

AOI21X1 _9257_ (
    .A(_2044_),
    .B(_2053_),
    .C(_2075_),
    .Y(_2076_)
);

NAND3X1 _9258_ (
    .A(_2035_),
    .B(_2057_),
    .C(_2043_),
    .Y(_2077_)
);

AOI21X1 _9259_ (
    .A(_2077_),
    .B(_2076_),
    .C(_2074_),
    .Y(_2078_)
);

AND2X2 _9260_ (
    .A(_2073_),
    .B(_2069_),
    .Y(_2079_)
);

NAND3X1 _9261_ (
    .A(_2053_),
    .B(_2056_),
    .C(_2035_),
    .Y(_2080_)
);

OAI21X1 _9262_ (
    .A(_2080_),
    .B(_2023_),
    .C(_2076_),
    .Y(_2081_)
);

OAI21X1 _9263_ (
    .A(_2079_),
    .B(_2081_),
    .C(_1903_),
    .Y(_2082_)
);

OR2X2 _9264_ (
    .A(_2082_),
    .B(_2078_),
    .Y(_2083_)
);

AOI22X1 _9265_ (
    .A(_1778_),
    .B(_1834__bF$buf2),
    .C(_2083_),
    .D(_1906_),
    .Y(_1687_)
);

NAND2X1 _9266_ (
    .A(\genblk1[2].u_ce.Ycalc [11]),
    .B(_1834__bF$buf1),
    .Y(_2084_)
);

INVX1 _9267_ (
    .A(_2073_),
    .Y(_2085_)
);

NAND2X1 _9268_ (
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .B(_2000_),
    .Y(_2086_)
);

INVX1 _9269_ (
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2087_)
);

NAND2X1 _9270_ (
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .B(_2087_),
    .Y(_2088_)
);

NAND2X1 _9271_ (
    .A(_2086_),
    .B(_2088_),
    .Y(_2089_)
);

INVX1 _9272_ (
    .A(_2089_),
    .Y(_2090_)
);

NAND2X1 _9273_ (
    .A(_2090_),
    .B(_2066_),
    .Y(_2091_)
);

NAND2X1 _9274_ (
    .A(_2089_),
    .B(_2071_),
    .Y(_2092_)
);

NAND2X1 _9275_ (
    .A(_2091_),
    .B(_2092_),
    .Y(_2093_)
);

INVX1 _9276_ (
    .A(_2093_),
    .Y(_2094_)
);

NOR3X1 _9277_ (
    .A(_2085_),
    .B(_2094_),
    .C(_2078_),
    .Y(_2095_)
);

AOI21X1 _9278_ (
    .A(_2081_),
    .B(_2079_),
    .C(_2085_),
    .Y(_2096_)
);

OAI21X1 _9279_ (
    .A(_2093_),
    .B(_2096_),
    .C(_1903_),
    .Y(_2097_)
);

OAI21X1 _9280_ (
    .A(_2095_),
    .B(_2097_),
    .C(_1906_),
    .Y(_2098_)
);

NAND2X1 _9281_ (
    .A(_2084_),
    .B(_2098_),
    .Y(_1688_)
);

NAND2X1 _9282_ (
    .A(\genblk1[2].u_ce.Xcalc [0]),
    .B(_1834__bF$buf0),
    .Y(_2099_)
);

INVX1 _9283_ (
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2100_)
);

NAND2X1 _9284_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2101_)
);

OAI21X1 _9285_ (
    .A(1'h0),
    .B(_2100_),
    .C(_2101_),
    .Y(_2102_)
);

NAND2X1 _9286_ (
    .A(1'h1),
    .B(_2102_),
    .Y(_2103_)
);

NOR2X1 _9287_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_2104_)
);

NOR2X1 _9288_ (
    .A(1'h1),
    .B(_1840_),
    .Y(_2105_)
);

AOI22X1 _9289_ (
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .B(_2104_),
    .C(_2105_),
    .D(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_2106_)
);

NAND3X1 _9290_ (
    .A(_1810__bF$buf4),
    .B(_2103_),
    .C(_2106_),
    .Y(_2107_)
);

NAND2X1 _9291_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_2108_)
);

OAI21X1 _9292_ (
    .A(1'h0),
    .B(_1971_),
    .C(_2108_),
    .Y(_2109_)
);

NAND2X1 _9293_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_2110_)
);

OAI21X1 _9294_ (
    .A(1'h0),
    .B(_1931_),
    .C(_2110_),
    .Y(_2111_)
);

MUX2X1 _9295_ (
    .A(_2111_),
    .B(_2109_),
    .S(_1811__bF$buf1),
    .Y(_2112_)
);

NAND2X1 _9296_ (
    .A(1'h0),
    .B(_2112_),
    .Y(_2113_)
);

AND2X2 _9297_ (
    .A(_2107_),
    .B(_2113_),
    .Y(_2114_)
);

NOR2X1 _9298_ (
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .B(_2114_),
    .Y(_2115_)
);

NAND2X1 _9299_ (
    .A(_1811__bF$buf0),
    .B(_2111_),
    .Y(_2116_)
);

NAND2X1 _9300_ (
    .A(1'h1),
    .B(_2109_),
    .Y(_2117_)
);

NAND2X1 _9301_ (
    .A(_2116_),
    .B(_2117_),
    .Y(_2118_)
);

OAI21X1 _9302_ (
    .A(_1810__bF$buf3),
    .B(_2118_),
    .C(_2107_),
    .Y(_2119_)
);

OAI21X1 _9303_ (
    .A(_1822_),
    .B(_2119_),
    .C(_1832_),
    .Y(_2120_)
);

OAI21X1 _9304_ (
    .A(_2120_),
    .B(_2115_),
    .C(_2099_),
    .Y(_1689_)
);

NAND2X1 _9305_ (
    .A(\genblk1[2].u_ce.Xcalc [1]),
    .B(_1834__bF$buf4),
    .Y(_2121_)
);

NOR2X1 _9306_ (
    .A(_1822_),
    .B(_2119_),
    .Y(_2122_)
);

NAND2X1 _9307_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_2123_)
);

OAI21X1 _9308_ (
    .A(1'h0),
    .B(_1909_),
    .C(_2123_),
    .Y(_2124_)
);

NAND2X1 _9309_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2125_)
);

OAI21X1 _9310_ (
    .A(1'h0),
    .B(_1847_),
    .C(_2125_),
    .Y(_2126_)
);

MUX2X1 _9311_ (
    .A(_2126_),
    .B(_2124_),
    .S(_1811__bF$buf4),
    .Y(_2127_)
);

NAND2X1 _9312_ (
    .A(_1810__bF$buf2),
    .B(_2127_),
    .Y(_2128_)
);

NAND2X1 _9313_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2129_)
);

OAI21X1 _9314_ (
    .A(1'h0),
    .B(_1998_),
    .C(_2129_),
    .Y(_2130_)
);

INVX1 _9315_ (
    .A(_2130_),
    .Y(_2131_)
);

NAND2X1 _9316_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_2132_)
);

OAI21X1 _9317_ (
    .A(1'h0),
    .B(_1952_),
    .C(_2132_),
    .Y(_2133_)
);

NAND2X1 _9318_ (
    .A(_1811__bF$buf3),
    .B(_2133_),
    .Y(_2134_)
);

OAI21X1 _9319_ (
    .A(_1811__bF$buf2),
    .B(_2131_),
    .C(_2134_),
    .Y(_2135_)
);

OAI21X1 _9320_ (
    .A(_1810__bF$buf1),
    .B(_2135_),
    .C(_2128_),
    .Y(_2136_)
);

NAND3X1 _9321_ (
    .A(_1848__bF$buf5),
    .B(_2136_),
    .C(_2114_),
    .Y(_2137_)
);

MUX2X1 _9322_ (
    .A(_2133_),
    .B(_2130_),
    .S(_1811__bF$buf1),
    .Y(_2138_)
);

MUX2X1 _9323_ (
    .A(_2138_),
    .B(_2127_),
    .S(1'h0),
    .Y(_2139_)
);

OAI21X1 _9324_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2119_),
    .C(_2139_),
    .Y(_2140_)
);

AOI21X1 _9325_ (
    .A(_2137_),
    .B(_2140_),
    .C(_1859_),
    .Y(_2141_)
);

INVX1 _9326_ (
    .A(_2141_),
    .Y(_2142_)
);

NAND3X1 _9327_ (
    .A(_1859_),
    .B(_2140_),
    .C(_2137_),
    .Y(_2143_)
);

AND2X2 _9328_ (
    .A(_2142_),
    .B(_2143_),
    .Y(_2144_)
);

NAND2X1 _9329_ (
    .A(_2122_),
    .B(_2144_),
    .Y(_2145_)
);

OR2X2 _9330_ (
    .A(_2144_),
    .B(_2122_),
    .Y(_2146_)
);

AOI21X1 _9331_ (
    .A(_2146_),
    .B(_2145_),
    .C(_1836_),
    .Y(_2147_)
);

OAI21X1 _9332_ (
    .A(_1834__bF$buf3),
    .B(_2147_),
    .C(_2121_),
    .Y(_1690_)
);

NAND2X1 _9333_ (
    .A(\genblk1[2].u_ce.Xcalc [2]),
    .B(_1834__bF$buf2),
    .Y(_2148_)
);

AOI21X1 _9334_ (
    .A(_2122_),
    .B(_2143_),
    .C(_2141_),
    .Y(_2149_)
);

NAND2X1 _9335_ (
    .A(_2119_),
    .B(_2136_),
    .Y(_2150_)
);

NAND2X1 _9336_ (
    .A(1'h0),
    .B(_2046_),
    .Y(_2151_)
);

OAI21X1 _9337_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .C(_2151_),
    .Y(_2152_)
);

NAND2X1 _9338_ (
    .A(_1811__bF$buf0),
    .B(_2109_),
    .Y(_2153_)
);

OAI21X1 _9339_ (
    .A(_1811__bF$buf4),
    .B(_2152_),
    .C(_2153_),
    .Y(_2154_)
);

NAND2X1 _9340_ (
    .A(_1917_),
    .B(_2102_),
    .Y(_2155_)
);

NAND2X1 _9341_ (
    .A(_2111_),
    .B(_1916_),
    .Y(_2156_)
);

NAND2X1 _9342_ (
    .A(_2155_),
    .B(_2156_),
    .Y(_2157_)
);

AOI21X1 _9343_ (
    .A(_2154_),
    .B(1'h0),
    .C(_2157_),
    .Y(_2158_)
);

INVX1 _9344_ (
    .A(_2158_),
    .Y(_2159_)
);

NAND3X1 _9345_ (
    .A(_1848__bF$buf4),
    .B(_2159_),
    .C(_2150_),
    .Y(_2160_)
);

AOI21X1 _9346_ (
    .A(_2107_),
    .B(_2113_),
    .C(_2139_),
    .Y(_2161_)
);

OAI21X1 _9347_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2161_),
    .C(_2158_),
    .Y(_2162_)
);

NAND3X1 _9348_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(_2162_),
    .C(_2160_),
    .Y(_2163_)
);

INVX1 _9349_ (
    .A(_2163_),
    .Y(_2164_)
);

AOI21X1 _9350_ (
    .A(_2160_),
    .B(_2162_),
    .C(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_2165_)
);

NOR2X1 _9351_ (
    .A(_2165_),
    .B(_2164_),
    .Y(_2166_)
);

AND2X2 _9352_ (
    .A(_2166_),
    .B(_2149_),
    .Y(_2167_)
);

NOR2X1 _9353_ (
    .A(_2149_),
    .B(_2166_),
    .Y(_2168_)
);

OAI21X1 _9354_ (
    .A(_2168_),
    .B(_2167_),
    .C(_1903_),
    .Y(_2169_)
);

OAI21X1 _9355_ (
    .A(_1834__bF$buf1),
    .B(_2169_),
    .C(_2148_),
    .Y(_1691_)
);

OAI21X1 _9356_ (
    .A(_2165_),
    .B(_2149_),
    .C(_2163_),
    .Y(_2170_)
);

INVX1 _9357_ (
    .A(_2170_),
    .Y(_2171_)
);

NAND2X1 _9358_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [10]),
    .Y(_2172_)
);

OAI21X1 _9359_ (
    .A(1'h0),
    .B(_2046_),
    .C(_2172_),
    .Y(_2173_)
);

MUX2X1 _9360_ (
    .A(_2173_),
    .B(_2130_),
    .S(1'h1),
    .Y(_2174_)
);

NOR2X1 _9361_ (
    .A(_1810__bF$buf0),
    .B(_2174_),
    .Y(_2175_)
);

NAND2X1 _9362_ (
    .A(_1917_),
    .B(_2124_),
    .Y(_2176_)
);

NAND2X1 _9363_ (
    .A(_2133_),
    .B(_1916_),
    .Y(_2177_)
);

NAND2X1 _9364_ (
    .A(_2176_),
    .B(_2177_),
    .Y(_2178_)
);

OR2X2 _9365_ (
    .A(_2175_),
    .B(_2178_),
    .Y(_2179_)
);

OAI21X1 _9366_ (
    .A(_2159_),
    .B(_2150_),
    .C(_1848__bF$buf3),
    .Y(_2180_)
);

OR2X2 _9367_ (
    .A(_2180_),
    .B(_2179_),
    .Y(_2181_)
);

OAI21X1 _9368_ (
    .A(_2175_),
    .B(_2178_),
    .C(_2180_),
    .Y(_2182_)
);

AOI21X1 _9369_ (
    .A(_2181_),
    .B(_2182_),
    .C(_1856_),
    .Y(_2183_)
);

INVX1 _9370_ (
    .A(_2183_),
    .Y(_2184_)
);

NAND3X1 _9371_ (
    .A(_1856_),
    .B(_2182_),
    .C(_2181_),
    .Y(_2185_)
);

NAND2X1 _9372_ (
    .A(_2185_),
    .B(_2184_),
    .Y(_2186_)
);

OR2X2 _9373_ (
    .A(_2186_),
    .B(_2171_),
    .Y(_2187_)
);

NAND2X1 _9374_ (
    .A(_2171_),
    .B(_2186_),
    .Y(_2188_)
);

NAND2X1 _9375_ (
    .A(_2188_),
    .B(_2187_),
    .Y(_2189_)
);

AOI22X1 _9376_ (
    .A(_1802_),
    .B(_1834__bF$buf0),
    .C(_2189_),
    .D(_1832_),
    .Y(_1692_)
);

AOI21X1 _9377_ (
    .A(_2170_),
    .B(_2185_),
    .C(_2183_),
    .Y(_2190_)
);

NAND2X1 _9378_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2191_)
);

OAI21X1 _9379_ (
    .A(1'h0),
    .B(_2061_),
    .C(_2191_),
    .Y(_2192_)
);

NAND2X1 _9380_ (
    .A(1'h1),
    .B(_2192_),
    .Y(_2193_)
);

OAI21X1 _9381_ (
    .A(1'h1),
    .B(_2152_),
    .C(_2193_),
    .Y(_2194_)
);

NAND2X1 _9382_ (
    .A(1'h0),
    .B(_2194_),
    .Y(_2195_)
);

OAI21X1 _9383_ (
    .A(1'h0),
    .B(_2112_),
    .C(_2195_),
    .Y(_2196_)
);

INVX1 _9384_ (
    .A(_2196_),
    .Y(_2197_)
);

NAND3X1 _9385_ (
    .A(_2158_),
    .B(_2119_),
    .C(_2136_),
    .Y(_2198_)
);

OAI21X1 _9386_ (
    .A(_2179_),
    .B(_2198_),
    .C(_1848__bF$buf2),
    .Y(_2199_)
);

OR2X2 _9387_ (
    .A(_2199_),
    .B(_2197_),
    .Y(_2200_)
);

NOR2X1 _9388_ (
    .A(_2179_),
    .B(_2198_),
    .Y(_2201_)
);

OAI21X1 _9389_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2201_),
    .C(_2197_),
    .Y(_2202_)
);

NAND3X1 _9390_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(_2202_),
    .C(_2200_),
    .Y(_2203_)
);

OR2X2 _9391_ (
    .A(_2199_),
    .B(_2196_),
    .Y(_2204_)
);

OAI21X1 _9392_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2201_),
    .C(_2196_),
    .Y(_2205_)
);

NAND3X1 _9393_ (
    .A(_1815_),
    .B(_2205_),
    .C(_2204_),
    .Y(_2206_)
);

NAND2X1 _9394_ (
    .A(_2203_),
    .B(_2206_),
    .Y(_2207_)
);

OR2X2 _9395_ (
    .A(_2190_),
    .B(_2207_),
    .Y(_2208_)
);

NAND2X1 _9396_ (
    .A(_2207_),
    .B(_2190_),
    .Y(_2209_)
);

NAND2X1 _9397_ (
    .A(_2209_),
    .B(_2208_),
    .Y(_2210_)
);

AOI22X1 _9398_ (
    .A(_1797_),
    .B(_1834__bF$buf4),
    .C(_2210_),
    .D(_1832_),
    .Y(_1693_)
);

INVX1 _9399_ (
    .A(\genblk1[2].u_ce.Xcalc [5]),
    .Y(_2211_)
);

OAI21X1 _9400_ (
    .A(_2207_),
    .B(_2190_),
    .C(_2203_),
    .Y(_2212_)
);

NAND2X1 _9401_ (
    .A(_2197_),
    .B(_2201_),
    .Y(_2213_)
);

NOR2X1 _9402_ (
    .A(_1811__bF$buf3),
    .B(_2087_),
    .Y(_2214_)
);

AOI21X1 _9403_ (
    .A(_1811__bF$buf2),
    .B(_2173_),
    .C(_2214_),
    .Y(_2215_)
);

NAND2X1 _9404_ (
    .A(_1810__bF$buf4),
    .B(_2135_),
    .Y(_2216_)
);

OAI21X1 _9405_ (
    .A(_1810__bF$buf3),
    .B(_2215_),
    .C(_2216_),
    .Y(_2217_)
);

INVX1 _9406_ (
    .A(_2217_),
    .Y(_2218_)
);

NAND3X1 _9407_ (
    .A(_1848__bF$buf1),
    .B(_2218_),
    .C(_2213_),
    .Y(_2219_)
);

NOR2X1 _9408_ (
    .A(_2178_),
    .B(_2175_),
    .Y(_2220_)
);

NAND3X1 _9409_ (
    .A(_2158_),
    .B(_2220_),
    .C(_2161_),
    .Y(_2221_)
);

OAI21X1 _9410_ (
    .A(_2196_),
    .B(_2221_),
    .C(_1848__bF$buf0),
    .Y(_2222_)
);

NAND2X1 _9411_ (
    .A(_2217_),
    .B(_2222_),
    .Y(_2223_)
);

AOI21X1 _9412_ (
    .A(_2219_),
    .B(_2223_),
    .C(_1852_),
    .Y(_2224_)
);

INVX1 _9413_ (
    .A(_2224_),
    .Y(_2225_)
);

NAND3X1 _9414_ (
    .A(_1852_),
    .B(_2223_),
    .C(_2219_),
    .Y(_2226_)
);

NAND2X1 _9415_ (
    .A(_2226_),
    .B(_2225_),
    .Y(_2227_)
);

NOR2X1 _9416_ (
    .A(_2227_),
    .B(_2212_),
    .Y(_2228_)
);

AND2X2 _9417_ (
    .A(_2212_),
    .B(_2227_),
    .Y(_2229_)
);

OAI21X1 _9418_ (
    .A(_2228_),
    .B(_2229_),
    .C(_1832_),
    .Y(_2230_)
);

OAI21X1 _9419_ (
    .A(_2211_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2230_),
    .Y(_1694_)
);

INVX1 _9420_ (
    .A(\genblk1[2].u_ce.Xcalc [6]),
    .Y(_2231_)
);

NAND3X1 _9421_ (
    .A(_2197_),
    .B(_2218_),
    .C(_2201_),
    .Y(_2232_)
);

AOI21X1 _9422_ (
    .A(_1811__bF$buf1),
    .B(_2192_),
    .C(_2214_),
    .Y(_2233_)
);

NAND2X1 _9423_ (
    .A(1'h0),
    .B(_2233_),
    .Y(_2234_)
);

OAI21X1 _9424_ (
    .A(1'h0),
    .B(_2154_),
    .C(_2234_),
    .Y(_2235_)
);

NAND3X1 _9425_ (
    .A(_1848__bF$buf5),
    .B(_2235_),
    .C(_2232_),
    .Y(_2236_)
);

NOR3X1 _9426_ (
    .A(_2196_),
    .B(_2217_),
    .C(_2221_),
    .Y(_2237_)
);

INVX1 _9427_ (
    .A(_2235_),
    .Y(_2238_)
);

OAI21X1 _9428_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2237_),
    .C(_2238_),
    .Y(_2239_)
);

NAND2X1 _9429_ (
    .A(_2236_),
    .B(_2239_),
    .Y(_2240_)
);

NAND2X1 _9430_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(_2240_),
    .Y(_2241_)
);

NAND3X1 _9431_ (
    .A(_1812_),
    .B(_2236_),
    .C(_2239_),
    .Y(_2242_)
);

NAND2X1 _9432_ (
    .A(_2242_),
    .B(_2241_),
    .Y(_2243_)
);

AOI21X1 _9433_ (
    .A(_2204_),
    .B(_2205_),
    .C(_1815_),
    .Y(_2244_)
);

NOR2X1 _9434_ (
    .A(_2244_),
    .B(_2224_),
    .Y(_2245_)
);

OAI21X1 _9435_ (
    .A(_2207_),
    .B(_2190_),
    .C(_2245_),
    .Y(_2246_)
);

NAND2X1 _9436_ (
    .A(_2226_),
    .B(_2246_),
    .Y(_2247_)
);

NOR2X1 _9437_ (
    .A(_2243_),
    .B(_2247_),
    .Y(_2248_)
);

AND2X2 _9438_ (
    .A(_2241_),
    .B(_2242_),
    .Y(_2249_)
);

AND2X2 _9439_ (
    .A(_2203_),
    .B(_2206_),
    .Y(_2250_)
);

NAND3X1 _9440_ (
    .A(_2226_),
    .B(_2250_),
    .C(_2225_),
    .Y(_2251_)
);

AOI21X1 _9441_ (
    .A(_2244_),
    .B(_2226_),
    .C(_2224_),
    .Y(_2252_)
);

OAI21X1 _9442_ (
    .A(_2190_),
    .B(_2251_),
    .C(_2252_),
    .Y(_2253_)
);

NOR2X1 _9443_ (
    .A(_2249_),
    .B(_2253_),
    .Y(_2254_)
);

OAI21X1 _9444_ (
    .A(_2254_),
    .B(_2248_),
    .C(_1903_),
    .Y(_2255_)
);

NAND2X1 _9445_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .B(_2255_),
    .Y(_2256_)
);

OAI21X1 _9446_ (
    .A(_2231_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_2256_),
    .Y(_1695_)
);

INVX1 _9447_ (
    .A(\genblk1[2].u_ce.Xcalc [7]),
    .Y(_2257_)
);

INVX1 _9448_ (
    .A(_2241_),
    .Y(_2258_)
);

NAND2X1 _9449_ (
    .A(_2235_),
    .B(_2237_),
    .Y(_2259_)
);

NOR2X1 _9450_ (
    .A(_1810__bF$buf2),
    .B(_2087_),
    .Y(_2260_)
);

INVX1 _9451_ (
    .A(_2260_),
    .Y(_2261_)
);

OAI21X1 _9452_ (
    .A(1'h0),
    .B(_2174_),
    .C(_2261_),
    .Y(_2262_)
);

NAND3X1 _9453_ (
    .A(_1848__bF$buf4),
    .B(_2262_),
    .C(_2259_),
    .Y(_2263_)
);

INVX1 _9454_ (
    .A(_2262_),
    .Y(_2264_)
);

OAI21X1 _9455_ (
    .A(_2238_),
    .B(_2232_),
    .C(_1848__bF$buf3),
    .Y(_2265_)
);

NAND2X1 _9456_ (
    .A(_2264_),
    .B(_2265_),
    .Y(_2266_)
);

NAND3X1 _9457_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(_2263_),
    .C(_2266_),
    .Y(_2267_)
);

NAND3X1 _9458_ (
    .A(_1848__bF$buf2),
    .B(_2264_),
    .C(_2259_),
    .Y(_2268_)
);

NAND2X1 _9459_ (
    .A(_2262_),
    .B(_2265_),
    .Y(_2269_)
);

NAND3X1 _9460_ (
    .A(_1849_),
    .B(_2268_),
    .C(_2269_),
    .Y(_2270_)
);

NAND2X1 _9461_ (
    .A(_2267_),
    .B(_2270_),
    .Y(_2271_)
);

OAI21X1 _9462_ (
    .A(_2258_),
    .B(_2248_),
    .C(_2271_),
    .Y(_2272_)
);

NOR2X1 _9463_ (
    .A(_2258_),
    .B(_2248_),
    .Y(_2273_)
);

INVX1 _9464_ (
    .A(_2271_),
    .Y(_2274_)
);

AOI21X1 _9465_ (
    .A(_2273_),
    .B(_2274_),
    .C(_1831_),
    .Y(_2275_)
);

AOI22X1 _9466_ (
    .A(_2257_),
    .B(_1834__bF$buf3),
    .C(_2275_),
    .D(_2272_),
    .Y(_1696_)
);

OAI21X1 _9467_ (
    .A(_2241_),
    .B(_2271_),
    .C(_2267_),
    .Y(_2276_)
);

NOR2X1 _9468_ (
    .A(_2243_),
    .B(_2271_),
    .Y(_2277_)
);

AOI21X1 _9469_ (
    .A(_2277_),
    .B(_2253_),
    .C(_2276_),
    .Y(_2278_)
);

INVX1 _9470_ (
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2279_)
);

NAND3X1 _9471_ (
    .A(_2235_),
    .B(_2264_),
    .C(_2237_),
    .Y(_2280_)
);

INVX1 _9472_ (
    .A(_2194_),
    .Y(_2281_)
);

OAI21X1 _9473_ (
    .A(1'h0),
    .B(_2281_),
    .C(_2261_),
    .Y(_2282_)
);

INVX1 _9474_ (
    .A(_2282_),
    .Y(_2283_)
);

NAND3X1 _9475_ (
    .A(_1848__bF$buf1),
    .B(_2283_),
    .C(_2280_),
    .Y(_2284_)
);

OAI21X1 _9476_ (
    .A(_2262_),
    .B(_2259_),
    .C(_1848__bF$buf0),
    .Y(_2285_)
);

NAND2X1 _9477_ (
    .A(_2282_),
    .B(_2285_),
    .Y(_2286_)
);

AOI21X1 _9478_ (
    .A(_2286_),
    .B(_2284_),
    .C(_2279_),
    .Y(_2287_)
);

NAND3X1 _9479_ (
    .A(_1848__bF$buf5),
    .B(_2282_),
    .C(_2280_),
    .Y(_2288_)
);

NAND2X1 _9480_ (
    .A(_2283_),
    .B(_2285_),
    .Y(_2289_)
);

AOI21X1 _9481_ (
    .A(_2289_),
    .B(_2288_),
    .C(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2290_)
);

OAI21X1 _9482_ (
    .A(_2287_),
    .B(_2290_),
    .C(_2278_),
    .Y(_2291_)
);

INVX1 _9483_ (
    .A(_2291_),
    .Y(_2292_)
);

OR2X2 _9484_ (
    .A(_2287_),
    .B(_2290_),
    .Y(_2293_)
);

OAI21X1 _9485_ (
    .A(_2293_),
    .B(_2278_),
    .C(_1832_),
    .Y(_2294_)
);

OAI22X1 _9486_ (
    .A(_1794_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2294_),
    .D(_2292_),
    .Y(_1697_)
);

NAND2X1 _9487_ (
    .A(\genblk1[2].u_ce.Xcalc [9]),
    .B(_1834__bF$buf2),
    .Y(_2295_)
);

NOR2X1 _9488_ (
    .A(_2293_),
    .B(_2278_),
    .Y(_2296_)
);

NOR2X1 _9489_ (
    .A(_2287_),
    .B(_2296_),
    .Y(_2297_)
);

OAI21X1 _9490_ (
    .A(1'h0),
    .B(_2215_),
    .C(_2261_),
    .Y(_2298_)
);

INVX1 _9491_ (
    .A(_2298_),
    .Y(_2299_)
);

OAI21X1 _9492_ (
    .A(_2282_),
    .B(_2280_),
    .C(_1848__bF$buf4),
    .Y(_2300_)
);

NAND2X1 _9493_ (
    .A(_2299_),
    .B(_2300_),
    .Y(_2301_)
);

OR2X2 _9494_ (
    .A(_2300_),
    .B(_2299_),
    .Y(_2302_)
);

NAND3X1 _9495_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(_2301_),
    .C(_2302_),
    .Y(_2303_)
);

NAND2X1 _9496_ (
    .A(_2301_),
    .B(_2302_),
    .Y(_2304_)
);

NAND2X1 _9497_ (
    .A(_1911_),
    .B(_2304_),
    .Y(_2305_)
);

NAND2X1 _9498_ (
    .A(_2303_),
    .B(_2305_),
    .Y(_2306_)
);

AND2X2 _9499_ (
    .A(_2297_),
    .B(_2306_),
    .Y(_2307_)
);

OAI21X1 _9500_ (
    .A(_2306_),
    .B(_2297_),
    .C(_1832_),
    .Y(_2308_)
);

OAI21X1 _9501_ (
    .A(_2308_),
    .B(_2307_),
    .C(_2295_),
    .Y(_1698_)
);

INVX1 _9502_ (
    .A(\genblk1[2].u_ce.Xcalc [10]),
    .Y(_2309_)
);

INVX1 _9503_ (
    .A(_2303_),
    .Y(_2310_)
);

AOI21X1 _9504_ (
    .A(_2287_),
    .B(_2305_),
    .C(_2310_),
    .Y(_2311_)
);

NOR2X1 _9505_ (
    .A(_2287_),
    .B(_2290_),
    .Y(_2312_)
);

NAND3X1 _9506_ (
    .A(_2303_),
    .B(_2305_),
    .C(_2312_),
    .Y(_2313_)
);

OAI21X1 _9507_ (
    .A(_2278_),
    .B(_2313_),
    .C(_2311_),
    .Y(_2314_)
);

OAI21X1 _9508_ (
    .A(1'h0),
    .B(_2233_),
    .C(_2261_),
    .Y(_2315_)
);

INVX1 _9509_ (
    .A(_2315_),
    .Y(_2316_)
);

OR2X2 _9510_ (
    .A(_2280_),
    .B(_2282_),
    .Y(_2317_)
);

OAI21X1 _9511_ (
    .A(_2298_),
    .B(_2317_),
    .C(_1848__bF$buf3),
    .Y(_2318_)
);

NAND2X1 _9512_ (
    .A(_2316_),
    .B(_2318_),
    .Y(_2319_)
);

OR2X2 _9513_ (
    .A(_2318_),
    .B(_2316_),
    .Y(_2320_)
);

NAND3X1 _9514_ (
    .A(\genblk1[2].u_ce.Xin12b [10]),
    .B(_2319_),
    .C(_2320_),
    .Y(_2321_)
);

AND2X2 _9515_ (
    .A(_2318_),
    .B(_2316_),
    .Y(_2322_)
);

NOR2X1 _9516_ (
    .A(_2316_),
    .B(_2318_),
    .Y(_2323_)
);

OAI21X1 _9517_ (
    .A(_2323_),
    .B(_2322_),
    .C(_1932_),
    .Y(_2324_)
);

NAND2X1 _9518_ (
    .A(_2324_),
    .B(_2321_),
    .Y(_2325_)
);

AND2X2 _9519_ (
    .A(_2314_),
    .B(_2325_),
    .Y(_2326_)
);

NOR2X1 _9520_ (
    .A(_2325_),
    .B(_2314_),
    .Y(_2327_)
);

NOR2X1 _9521_ (
    .A(_2326_),
    .B(_2327_),
    .Y(_2328_)
);

AOI22X1 _9522_ (
    .A(_2309_),
    .B(_1834__bF$buf1),
    .C(_2328_),
    .D(_1832_),
    .Y(_1699_)
);

NAND2X1 _9523_ (
    .A(\genblk1[2].u_ce.Xcalc [11]),
    .B(_1834__bF$buf0),
    .Y(_2329_)
);

INVX1 _9524_ (
    .A(_2321_),
    .Y(_2330_)
);

AOI21X1 _9525_ (
    .A(_2314_),
    .B(_2324_),
    .C(_2330_),
    .Y(_2331_)
);

NAND2X1 _9526_ (
    .A(_1848__bF$buf2),
    .B(_2319_),
    .Y(_2332_)
);

NOR2X1 _9527_ (
    .A(_2089_),
    .B(_2332_),
    .Y(_2333_)
);

AOI21X1 _9528_ (
    .A(_2319_),
    .B(_1848__bF$buf1),
    .C(_2090_),
    .Y(_2334_)
);

NOR2X1 _9529_ (
    .A(_2334_),
    .B(_2333_),
    .Y(_2335_)
);

AND2X2 _9530_ (
    .A(_2331_),
    .B(_2335_),
    .Y(_2336_)
);

OAI21X1 _9531_ (
    .A(_2335_),
    .B(_2331_),
    .C(_1832_),
    .Y(_2337_)
);

OAI21X1 _9532_ (
    .A(_2337_),
    .B(_2336_),
    .C(_2329_),
    .Y(_1700_)
);

OAI21X1 _9533_ (
    .A(1'h0),
    .B(_1811__bF$buf0),
    .C(_1830_),
    .Y(_2338_)
);

OAI21X1 _9534_ (
    .A(_2105_),
    .B(_2338_),
    .C(\genblk1[2].u_ce.Ain0 [0]),
    .Y(_2339_)
);

INVX1 _9535_ (
    .A(\genblk1[2].u_ce.Ain0 [0]),
    .Y(_2340_)
);

NOR2X1 _9536_ (
    .A(_2105_),
    .B(_2338_),
    .Y(_2341_)
);

NAND2X1 _9537_ (
    .A(_2340_),
    .B(_2341_),
    .Y(_2342_)
);

NAND2X1 _9538_ (
    .A(_2339_),
    .B(_2342_),
    .Y(_2343_)
);

NAND2X1 _9539_ (
    .A(\genblk1[2].u_ce.Acalc [0]),
    .B(_1834__bF$buf4),
    .Y(_2344_)
);

OAI21X1 _9540_ (
    .A(_1834__bF$buf3),
    .B(_2343_),
    .C(_2344_),
    .Y(_1701_)
);

NAND2X1 _9541_ (
    .A(\genblk1[2].u_ce.Acalc [1]),
    .B(_1834__bF$buf2),
    .Y(_2345_)
);

INVX1 _9542_ (
    .A(_2339_),
    .Y(_2346_)
);

NOR2X1 _9543_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_2347_)
);

AOI21X1 _9544_ (
    .A(_2105_),
    .B(1'h0),
    .C(_2347_),
    .Y(_2348_)
);

NOR2X1 _9545_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2348_),
    .Y(_2349_)
);

OAI21X1 _9546_ (
    .A(_2105_),
    .B(_2338_),
    .C(_1848__bF$buf0),
    .Y(_2350_)
);

AND2X2 _9547_ (
    .A(_2350_),
    .B(_2348_),
    .Y(_2351_)
);

OR2X2 _9548_ (
    .A(_2351_),
    .B(_2349_),
    .Y(_2352_)
);

OR2X2 _9549_ (
    .A(_2352_),
    .B(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2353_)
);

OAI21X1 _9550_ (
    .A(_2349_),
    .B(_2351_),
    .C(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2354_)
);

NAND2X1 _9551_ (
    .A(_2354_),
    .B(_2353_),
    .Y(_2355_)
);

NOR2X1 _9552_ (
    .A(_2346_),
    .B(_2355_),
    .Y(_2356_)
);

NAND2X1 _9553_ (
    .A(_2346_),
    .B(_2355_),
    .Y(_2357_)
);

NAND2X1 _9554_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_2357_),
    .Y(_2358_)
);

OAI21X1 _9555_ (
    .A(_2356_),
    .B(_2358_),
    .C(_2345_),
    .Y(_1702_)
);

INVX1 _9556_ (
    .A(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2359_)
);

OAI21X1 _9557_ (
    .A(_2359_),
    .B(_2352_),
    .C(_2357_),
    .Y(_2360_)
);

OAI21X1 _9558_ (
    .A(_1840_),
    .B(_1811__bF$buf4),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_2361_)
);

OAI21X1 _9559_ (
    .A(1'h0),
    .B(1'h1),
    .C(1'h0),
    .Y(_2362_)
);

MUX2X1 _9560_ (
    .A(_2362_),
    .B(1'h0),
    .S(_2361_),
    .Y(_2363_)
);

NAND2X1 _9561_ (
    .A(\genblk1[2].u_ce.Ain1 [0]),
    .B(_2363_),
    .Y(_2364_)
);

OR2X2 _9562_ (
    .A(_2363_),
    .B(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_2365_)
);

NAND2X1 _9563_ (
    .A(_2364_),
    .B(_2365_),
    .Y(_2366_)
);

INVX1 _9564_ (
    .A(_2366_),
    .Y(_2367_)
);

NOR2X1 _9565_ (
    .A(_2367_),
    .B(_2360_),
    .Y(_2368_)
);

NAND2X1 _9566_ (
    .A(_2367_),
    .B(_2360_),
    .Y(_2369_)
);

NAND2X1 _9567_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2369_),
    .Y(_2370_)
);

OAI22X1 _9568_ (
    .A(_1756_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_2368_),
    .D(_2370_),
    .Y(_1703_)
);

NOR2X1 _9569_ (
    .A(\genblk1[2].u_ce.Acalc [3]),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2371_)
);

NAND2X1 _9570_ (
    .A(_2364_),
    .B(_2369_),
    .Y(_2372_)
);

INVX1 _9571_ (
    .A(_2372_),
    .Y(_2373_)
);

INVX1 _9572_ (
    .A(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_2374_)
);

NOR2X1 _9573_ (
    .A(1'h0),
    .B(_1811__bF$buf3),
    .Y(_2375_)
);

OAI21X1 _9574_ (
    .A(_1810__bF$buf1),
    .B(_2375_),
    .C(_1848__bF$buf5),
    .Y(_2376_)
);

OAI21X1 _9575_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_2377_)
);

OAI21X1 _9576_ (
    .A(_1840_),
    .B(_2377_),
    .C(_2376_),
    .Y(_2378_)
);

NOR2X1 _9577_ (
    .A(_2374_),
    .B(_2378_),
    .Y(_2379_)
);

NAND2X1 _9578_ (
    .A(_2374_),
    .B(_2378_),
    .Y(_2380_)
);

INVX1 _9579_ (
    .A(_2380_),
    .Y(_2381_)
);

NOR2X1 _9580_ (
    .A(_2379_),
    .B(_2381_),
    .Y(_2382_)
);

OAI21X1 _9581_ (
    .A(_2382_),
    .B(_2373_),
    .C(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .Y(_2383_)
);

AOI21X1 _9582_ (
    .A(_2373_),
    .B(_2382_),
    .C(_2383_),
    .Y(_2384_)
);

NOR2X1 _9583_ (
    .A(_2371_),
    .B(_2384_),
    .Y(_1704_)
);

NAND2X1 _9584_ (
    .A(\genblk1[2].u_ce.Acalc [4]),
    .B(_1834__bF$buf1),
    .Y(_2385_)
);

INVX1 _9585_ (
    .A(\genblk1[2].u_ce.Ain12b [4]),
    .Y(_2386_)
);

AOI21X1 _9586_ (
    .A(_2105_),
    .B(1'h0),
    .C(_1848__bF$buf4),
    .Y(_2387_)
);

OAI21X1 _9587_ (
    .A(1'h0),
    .B(_2105_),
    .C(_2387_),
    .Y(_2388_)
);

OAI21X1 _9588_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2348_),
    .C(_2388_),
    .Y(_2389_)
);

OR2X2 _9589_ (
    .A(_2389_),
    .B(_2386_),
    .Y(_2390_)
);

NAND2X1 _9590_ (
    .A(_2386_),
    .B(_2389_),
    .Y(_2391_)
);

NAND2X1 _9591_ (
    .A(_2391_),
    .B(_2390_),
    .Y(_2392_)
);

AOI21X1 _9592_ (
    .A(_2372_),
    .B(_2380_),
    .C(_2379_),
    .Y(_2393_)
);

AND2X2 _9593_ (
    .A(_2393_),
    .B(_2392_),
    .Y(_2394_)
);

OAI21X1 _9594_ (
    .A(_2392_),
    .B(_2393_),
    .C(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .Y(_2395_)
);

OAI21X1 _9595_ (
    .A(_2395_),
    .B(_2394_),
    .C(_2385_),
    .Y(_1705_)
);

OAI21X1 _9596_ (
    .A(_2392_),
    .B(_2393_),
    .C(_2390_),
    .Y(_2396_)
);

INVX1 _9597_ (
    .A(\genblk1[2].u_ce.Ain12b [5]),
    .Y(_2397_)
);

OAI21X1 _9598_ (
    .A(_2104_),
    .B(_1917_),
    .C(_1848__bF$buf3),
    .Y(_2398_)
);

OAI21X1 _9599_ (
    .A(1'h0),
    .B(1'h1),
    .C(_1830_),
    .Y(_2399_)
);

OR2X2 _9600_ (
    .A(_2399_),
    .B(_1848__bF$buf2),
    .Y(_2400_)
);

NAND2X1 _9601_ (
    .A(_2398_),
    .B(_2400_),
    .Y(_2401_)
);

OR2X2 _9602_ (
    .A(_2401_),
    .B(_2397_),
    .Y(_2402_)
);

NAND2X1 _9603_ (
    .A(_2397_),
    .B(_2401_),
    .Y(_2403_)
);

NAND2X1 _9604_ (
    .A(_2403_),
    .B(_2402_),
    .Y(_2404_)
);

INVX1 _9605_ (
    .A(_2404_),
    .Y(_2405_)
);

NOR2X1 _9606_ (
    .A(_2405_),
    .B(_2396_),
    .Y(_2406_)
);

NAND2X1 _9607_ (
    .A(_2405_),
    .B(_2396_),
    .Y(_2407_)
);

NAND2X1 _9608_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2407_),
    .Y(_2408_)
);

OAI22X1 _9609_ (
    .A(_1773_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_2406_),
    .D(_2408_),
    .Y(_1706_)
);

NAND2X1 _9610_ (
    .A(\genblk1[2].u_ce.Acalc [6]),
    .B(_1834__bF$buf0),
    .Y(_2409_)
);

INVX1 _9611_ (
    .A(_2392_),
    .Y(_2410_)
);

NAND2X1 _9612_ (
    .A(_2405_),
    .B(_2410_),
    .Y(_2411_)
);

OAI21X1 _9613_ (
    .A(_2390_),
    .B(_2404_),
    .C(_2402_),
    .Y(_2412_)
);

INVX1 _9614_ (
    .A(_2412_),
    .Y(_2413_)
);

OAI21X1 _9615_ (
    .A(_2411_),
    .B(_2393_),
    .C(_2413_),
    .Y(_2414_)
);

OAI21X1 _9616_ (
    .A(1'h1),
    .B(_1840_),
    .C(_1810__bF$buf0),
    .Y(_2415_)
);

NOR2X1 _9617_ (
    .A(_2415_),
    .B(_2375_),
    .Y(_2416_)
);

NAND2X1 _9618_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2416_),
    .Y(_2417_)
);

OAI21X1 _9619_ (
    .A(_2415_),
    .B(_2375_),
    .C(_1848__bF$buf1),
    .Y(_2418_)
);

NAND2X1 _9620_ (
    .A(_2418_),
    .B(_2417_),
    .Y(_2419_)
);

NAND2X1 _9621_ (
    .A(\genblk1[2].u_ce.Ain12b [6]),
    .B(_2419_),
    .Y(_2420_)
);

OR2X2 _9622_ (
    .A(_2419_),
    .B(\genblk1[2].u_ce.Ain12b [6]),
    .Y(_2421_)
);

NAND2X1 _9623_ (
    .A(_2420_),
    .B(_2421_),
    .Y(_2422_)
);

INVX1 _9624_ (
    .A(_2422_),
    .Y(_2423_)
);

NOR2X1 _9625_ (
    .A(_2423_),
    .B(_2414_),
    .Y(_2424_)
);

NAND2X1 _9626_ (
    .A(_2423_),
    .B(_2414_),
    .Y(_2425_)
);

NAND2X1 _9627_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .B(_2425_),
    .Y(_2426_)
);

OAI21X1 _9628_ (
    .A(_2424_),
    .B(_2426_),
    .C(_2409_),
    .Y(_1707_)
);

INVX1 _9629_ (
    .A(\genblk1[2].u_ce.Acalc [7]),
    .Y(_2427_)
);

NAND2X1 _9630_ (
    .A(_2420_),
    .B(_2425_),
    .Y(_2428_)
);

INVX1 _9631_ (
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .Y(_2429_)
);

NAND2X1 _9632_ (
    .A(_1848__bF$buf0),
    .B(_2347_),
    .Y(_2430_)
);

OR2X2 _9633_ (
    .A(_2347_),
    .B(_1848__bF$buf5),
    .Y(_2431_)
);

NAND2X1 _9634_ (
    .A(_2430_),
    .B(_2431_),
    .Y(_2432_)
);

NOR2X1 _9635_ (
    .A(_2429_),
    .B(_2432_),
    .Y(_2433_)
);

INVX1 _9636_ (
    .A(_2433_),
    .Y(_2434_)
);

NAND2X1 _9637_ (
    .A(_2429_),
    .B(_2432_),
    .Y(_2435_)
);

NAND2X1 _9638_ (
    .A(_2435_),
    .B(_2434_),
    .Y(_2436_)
);

OR2X2 _9639_ (
    .A(_2428_),
    .B(_2436_),
    .Y(_2437_)
);

AOI21X1 _9640_ (
    .A(_2428_),
    .B(_2436_),
    .C(_1834__bF$buf4),
    .Y(_2438_)
);

AOI22X1 _9641_ (
    .A(_2427_),
    .B(_1834__bF$buf3),
    .C(_2437_),
    .D(_2438_),
    .Y(_1708_)
);

NAND2X1 _9642_ (
    .A(\genblk1[2].u_ce.Acalc [8]),
    .B(_1834__bF$buf2),
    .Y(_2439_)
);

NOR2X1 _9643_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1830_),
    .Y(_2440_)
);

INVX1 _9644_ (
    .A(_2440_),
    .Y(_2441_)
);

NAND3X1 _9645_ (
    .A(\genblk1[2].u_ce.Ain12b [8]),
    .B(_2377_),
    .C(_2441_),
    .Y(_2442_)
);

INVX1 _9646_ (
    .A(_2442_),
    .Y(_2443_)
);

AOI21X1 _9647_ (
    .A(_2441_),
    .B(_2377_),
    .C(\genblk1[2].u_ce.Ain12b [8]),
    .Y(_2444_)
);

NOR2X1 _9648_ (
    .A(_2444_),
    .B(_2443_),
    .Y(_2445_)
);

OAI21X1 _9649_ (
    .A(_2420_),
    .B(_2436_),
    .C(_2434_),
    .Y(_2446_)
);

NOR2X1 _9650_ (
    .A(_2436_),
    .B(_2422_),
    .Y(_2447_)
);

AOI21X1 _9651_ (
    .A(_2447_),
    .B(_2412_),
    .C(_2446_),
    .Y(_2448_)
);

NAND3X1 _9652_ (
    .A(_2410_),
    .B(_2405_),
    .C(_2447_),
    .Y(_2449_)
);

OAI21X1 _9653_ (
    .A(_2449_),
    .B(_2393_),
    .C(_2448_),
    .Y(_2450_)
);

NOR2X1 _9654_ (
    .A(_2445_),
    .B(_2450_),
    .Y(_2451_)
);

NAND2X1 _9655_ (
    .A(_2445_),
    .B(_2450_),
    .Y(_2452_)
);

NAND2X1 _9656_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .B(_2452_),
    .Y(_2453_)
);

OAI21X1 _9657_ (
    .A(_2451_),
    .B(_2453_),
    .C(_2439_),
    .Y(_1709_)
);

AOI21X1 _9658_ (
    .A(_2450_),
    .B(_2445_),
    .C(_2443_),
    .Y(_2454_)
);

OR2X2 _9659_ (
    .A(_1848__bF$buf4),
    .B(\genblk1[2].u_ce.Ain12b [9]),
    .Y(_2455_)
);

NAND2X1 _9660_ (
    .A(\genblk1[2].u_ce.Ain12b [9]),
    .B(_1848__bF$buf3),
    .Y(_2456_)
);

NAND2X1 _9661_ (
    .A(_2456_),
    .B(_2455_),
    .Y(_2457_)
);

AND2X2 _9662_ (
    .A(_2454_),
    .B(_2457_),
    .Y(_2458_)
);

OAI21X1 _9663_ (
    .A(_2457_),
    .B(_2454_),
    .C(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .Y(_2459_)
);

OAI22X1 _9664_ (
    .A(_1770_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2459_),
    .D(_2458_),
    .Y(_1710_)
);

NAND2X1 _9665_ (
    .A(\genblk1[2].u_ce.Acalc [10]),
    .B(_1834__bF$buf1),
    .Y(_2460_)
);

OAI21X1 _9666_ (
    .A(_2457_),
    .B(_2442_),
    .C(_2456_),
    .Y(_2461_)
);

NAND3X1 _9667_ (
    .A(_2455_),
    .B(_2456_),
    .C(_2445_),
    .Y(_2462_)
);

INVX1 _9668_ (
    .A(_2462_),
    .Y(_2463_)
);

AOI21X1 _9669_ (
    .A(_2450_),
    .B(_2463_),
    .C(_2461_),
    .Y(_2464_)
);

INVX1 _9670_ (
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .Y(_2465_)
);

NAND2X1 _9671_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2465_),
    .Y(_2466_)
);

NAND2X1 _9672_ (
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .B(_1848__bF$buf2),
    .Y(_2467_)
);

NAND2X1 _9673_ (
    .A(_2466_),
    .B(_2467_),
    .Y(_2468_)
);

AND2X2 _9674_ (
    .A(_2464_),
    .B(_2468_),
    .Y(_2469_)
);

OAI21X1 _9675_ (
    .A(_2468_),
    .B(_2464_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2470_)
);

OAI21X1 _9676_ (
    .A(_2470_),
    .B(_2469_),
    .C(_2460_),
    .Y(_1711_)
);

NAND2X1 _9677_ (
    .A(\genblk1[2].u_ce.Acalc [11]),
    .B(_1834__bF$buf0),
    .Y(_2471_)
);

OAI21X1 _9678_ (
    .A(_2468_),
    .B(_2464_),
    .C(_2467_),
    .Y(_2472_)
);

OAI21X1 _9679_ (
    .A(_1834__bF$buf4),
    .B(_2472_),
    .C(_2471_),
    .Y(_1712_)
);

NAND2X1 _9680_ (
    .A(\genblk1[2].u_ce.LoadCtl [5]),
    .B(_1761_),
    .Y(_2473_)
);

NAND2X1 _9681_ (
    .A(_1762_),
    .B(_1768_),
    .Y(_2474_)
);

NOR2X1 _9682_ (
    .A(_2473_),
    .B(_2474_),
    .Y(_2475_)
);

NAND2X1 _9683_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2475_),
    .Y(_2476_)
);

OAI21X1 _9684_ (
    .A(_1932_),
    .B(_2475_),
    .C(_2476_),
    .Y(_1713_)
);

NAND2X1 _9685_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2475_),
    .Y(_2477_)
);

OAI21X1 _9686_ (
    .A(_2000_),
    .B(_2475_),
    .C(_2477_),
    .Y(_1714_)
);

INVX1 _9687_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .Y(_2478_)
);

OR2X2 _9688_ (
    .A(_2474_),
    .B(_1761_),
    .Y(_2479_)
);

OAI21X1 _9689_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2480_)
);

OAI21X1 _9690_ (
    .A(_2478_),
    .B(_2479_),
    .C(_2480_),
    .Y(_1715_)
);

INVX1 _9691_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .Y(_2481_)
);

OAI21X1 _9692_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Xin12b [9]),
    .Y(_2482_)
);

OAI21X1 _9693_ (
    .A(_2481_),
    .B(_2479_),
    .C(_2482_),
    .Y(_1716_)
);

NAND2X1 _9694_ (
    .A(_1768_),
    .B(_1765_),
    .Y(_2483_)
);

NAND2X1 _9695_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(_2483_),
    .Y(_2484_)
);

OAI21X1 _9696_ (
    .A(_2478_),
    .B(_2483_),
    .C(_2484_),
    .Y(_1717_)
);

NAND2X1 _9697_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(_2483_),
    .Y(_2485_)
);

OAI21X1 _9698_ (
    .A(_2481_),
    .B(_2483_),
    .C(_2485_),
    .Y(_1718_)
);

AND2X2 _9699_ (
    .A(_1768_),
    .B(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_2486_)
);

NAND2X1 _9700_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2486_),
    .Y(_2487_)
);

OAI21X1 _9701_ (
    .A(_1815_),
    .B(_2486_),
    .C(_2487_),
    .Y(_1719_)
);

NAND2X1 _9702_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2486_),
    .Y(_2488_)
);

OAI21X1 _9703_ (
    .A(_1852_),
    .B(_2486_),
    .C(_2488_),
    .Y(_1720_)
);

OAI21X1 _9704_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_2489_)
);

OAI21X1 _9705_ (
    .A(_2478_),
    .B(_1759_),
    .C(_2489_),
    .Y(_1721_)
);

OAI21X1 _9706_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_2490_)
);

OAI21X1 _9707_ (
    .A(_2481_),
    .B(_1759_),
    .C(_2490_),
    .Y(_1722_)
);

NAND2X1 _9708_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[1].u_ce.X_ [0]),
    .Y(_2491_)
);

OAI21X1 _9709_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1822_),
    .C(_2491_),
    .Y(_1723_)
);

NAND2X1 _9710_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.X_ [1]),
    .Y(_2492_)
);

OAI21X1 _9711_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1859_),
    .C(_2492_),
    .Y(_1724_)
);

NAND2X1 _9712_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2475_),
    .Y(_2493_)
);

OAI21X1 _9713_ (
    .A(_2061_),
    .B(_2475_),
    .C(_2493_),
    .Y(_1725_)
);

NAND2X1 _9714_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2475_),
    .Y(_2494_)
);

OAI21X1 _9715_ (
    .A(_2087_),
    .B(_2475_),
    .C(_2494_),
    .Y(_1726_)
);

INVX1 _9716_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .Y(_2495_)
);

OAI21X1 _9717_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2496_)
);

OAI21X1 _9718_ (
    .A(_2495_),
    .B(_2479_),
    .C(_2496_),
    .Y(_1727_)
);

INVX1 _9719_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .Y(_2497_)
);

OAI21X1 _9720_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2498_)
);

OAI21X1 _9721_ (
    .A(_2497_),
    .B(_2479_),
    .C(_2498_),
    .Y(_1728_)
);

NAND2X1 _9722_ (
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .B(_2483_),
    .Y(_2499_)
);

OAI21X1 _9723_ (
    .A(_2495_),
    .B(_2483_),
    .C(_2499_),
    .Y(_1729_)
);

NAND2X1 _9724_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(_2483_),
    .Y(_2500_)
);

OAI21X1 _9725_ (
    .A(_2497_),
    .B(_2483_),
    .C(_2500_),
    .Y(_1730_)
);

NAND2X1 _9726_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2486_),
    .Y(_2501_)
);

OAI21X1 _9727_ (
    .A(_1931_),
    .B(_2486_),
    .C(_2501_),
    .Y(_1731_)
);

NAND2X1 _9728_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2486_),
    .Y(_2502_)
);

OAI21X1 _9729_ (
    .A(_1952_),
    .B(_2486_),
    .C(_2502_),
    .Y(_1732_)
);

OAI21X1 _9730_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2503_)
);

OAI21X1 _9731_ (
    .A(_2495_),
    .B(_1759_),
    .C(_2503_),
    .Y(_1733_)
);

OAI21X1 _9732_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2504_)
);

OAI21X1 _9733_ (
    .A(_2497_),
    .B(_1759_),
    .C(_2504_),
    .Y(_1734_)
);

NAND2X1 _9734_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.Y_ [0]),
    .Y(_2505_)
);

OAI21X1 _9735_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_1809_),
    .C(_2505_),
    .Y(_1735_)
);

NAND2X1 _9736_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Y_ [1]),
    .Y(_2506_)
);

OAI21X1 _9737_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1847_),
    .C(_2506_),
    .Y(_1736_)
);

NAND2X1 _9738_ (
    .A(\a[2] [0]),
    .B(_2475_),
    .Y(_2507_)
);

OAI21X1 _9739_ (
    .A(_2465_),
    .B(_2475_),
    .C(_2507_),
    .Y(_1737_)
);

NAND2X1 _9740_ (
    .A(\a[2] [1]),
    .B(_2475_),
    .Y(_2508_)
);

OAI21X1 _9741_ (
    .A(_1848__bF$buf1),
    .B(_2475_),
    .C(_2508_),
    .Y(_1738_)
);

INVX1 _9742_ (
    .A(\a[2] [0]),
    .Y(_2509_)
);

OAI21X1 _9743_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Ain12b [8]),
    .Y(_2510_)
);

OAI21X1 _9744_ (
    .A(_2509_),
    .B(_2479_),
    .C(_2510_),
    .Y(_1739_)
);

INVX1 _9745_ (
    .A(\a[2] [1]),
    .Y(_2511_)
);

OAI21X1 _9746_ (
    .A(_1761_),
    .B(_2474_),
    .C(\genblk1[2].u_ce.Ain12b [9]),
    .Y(_2512_)
);

OAI21X1 _9747_ (
    .A(_2511_),
    .B(_2479_),
    .C(_2512_),
    .Y(_1740_)
);

NAND2X1 _9748_ (
    .A(\genblk1[2].u_ce.Ain12b [6]),
    .B(_2483_),
    .Y(_2513_)
);

OAI21X1 _9749_ (
    .A(_2509_),
    .B(_2483_),
    .C(_2513_),
    .Y(_1741_)
);

NAND2X1 _9750_ (
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .B(_2483_),
    .Y(_1749_)
);

OAI21X1 _9751_ (
    .A(_2511_),
    .B(_2483_),
    .C(_1749_),
    .Y(_1742_)
);

NAND2X1 _9752_ (
    .A(\a[2] [0]),
    .B(_2486_),
    .Y(_1750_)
);

OAI21X1 _9753_ (
    .A(_2386_),
    .B(_2486_),
    .C(_1750_),
    .Y(_1743_)
);

NAND2X1 _9754_ (
    .A(\a[2] [1]),
    .B(_2486_),
    .Y(_1751_)
);

OAI21X1 _9755_ (
    .A(_2397_),
    .B(_2486_),
    .C(_1751_),
    .Y(_1744_)
);

OAI21X1 _9756_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_1752_)
);

OAI21X1 _9757_ (
    .A(_2509_),
    .B(_1759_),
    .C(_1752_),
    .Y(_1745_)
);

OAI21X1 _9758_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1757_),
    .C(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_1753_)
);

OAI21X1 _9759_ (
    .A(_2511_),
    .B(_1759_),
    .C(_1753_),
    .Y(_1746_)
);

NAND2X1 _9760_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[2] [0]),
    .Y(_1754_)
);

OAI21X1 _9761_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2340_),
    .C(_1754_),
    .Y(_1747_)
);

NAND2X1 _9762_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[2] [1]),
    .Y(_1755_)
);

OAI21X1 _9763_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2359_),
    .C(_1755_),
    .Y(_1748_)
);

DFFPOSX1 _9764_ (
    .CLK(clk_bF$buf5),
    .D(_1676_),
    .Q(\genblk1[2].u_ce.Ycalc [0])
);

DFFPOSX1 _9765_ (
    .CLK(clk_bF$buf4),
    .D(_1677_),
    .Q(\genblk1[2].u_ce.Ycalc [1])
);

DFFPOSX1 _9766_ (
    .CLK(clk_bF$buf3),
    .D(_1678_),
    .Q(\genblk1[2].u_ce.ISout )
);

DFFPOSX1 _9767_ (
    .CLK(clk_bF$buf2),
    .D(_1679_),
    .Q(\genblk1[2].u_ce.Ycalc [2])
);

DFFPOSX1 _9768_ (
    .CLK(clk_bF$buf1),
    .D(_1680_),
    .Q(\genblk1[2].u_ce.Ycalc [3])
);

DFFPOSX1 _9769_ (
    .CLK(clk_bF$buf0),
    .D(_1681_),
    .Q(\genblk1[2].u_ce.Ycalc [4])
);

DFFPOSX1 _9770_ (
    .CLK(clk_bF$buf78),
    .D(_1682_),
    .Q(\genblk1[2].u_ce.Ycalc [5])
);

DFFPOSX1 _9771_ (
    .CLK(clk_bF$buf77),
    .D(_1683_),
    .Q(\genblk1[2].u_ce.Ycalc [6])
);

DFFPOSX1 _9772_ (
    .CLK(clk_bF$buf76),
    .D(_1684_),
    .Q(\genblk1[2].u_ce.Ycalc [7])
);

DFFPOSX1 _9773_ (
    .CLK(clk_bF$buf75),
    .D(_1685_),
    .Q(\genblk1[2].u_ce.Ycalc [8])
);

DFFPOSX1 _9774_ (
    .CLK(clk_bF$buf74),
    .D(_1686_),
    .Q(\genblk1[2].u_ce.Ycalc [9])
);

DFFPOSX1 _9775_ (
    .CLK(clk_bF$buf73),
    .D(_1687_),
    .Q(\genblk1[2].u_ce.Ycalc [10])
);

DFFPOSX1 _9776_ (
    .CLK(clk_bF$buf72),
    .D(_1688_),
    .Q(\genblk1[2].u_ce.Ycalc [11])
);

DFFPOSX1 _9777_ (
    .CLK(clk_bF$buf71),
    .D(_1689_),
    .Q(\genblk1[2].u_ce.Xcalc [0])
);

DFFPOSX1 _9778_ (
    .CLK(clk_bF$buf70),
    .D(_1690_),
    .Q(\genblk1[2].u_ce.Xcalc [1])
);

DFFPOSX1 _9779_ (
    .CLK(clk_bF$buf69),
    .D(_1691_),
    .Q(\genblk1[2].u_ce.Xcalc [2])
);

DFFPOSX1 _9780_ (
    .CLK(clk_bF$buf68),
    .D(_1692_),
    .Q(\genblk1[2].u_ce.Xcalc [3])
);

DFFPOSX1 _9781_ (
    .CLK(clk_bF$buf67),
    .D(_1693_),
    .Q(\genblk1[2].u_ce.Xcalc [4])
);

DFFPOSX1 _9782_ (
    .CLK(clk_bF$buf66),
    .D(_1694_),
    .Q(\genblk1[2].u_ce.Xcalc [5])
);

DFFPOSX1 _9783_ (
    .CLK(clk_bF$buf65),
    .D(_1695_),
    .Q(\genblk1[2].u_ce.Xcalc [6])
);

DFFPOSX1 _9784_ (
    .CLK(clk_bF$buf64),
    .D(_1696_),
    .Q(\genblk1[2].u_ce.Xcalc [7])
);

DFFPOSX1 _9785_ (
    .CLK(clk_bF$buf63),
    .D(_1697_),
    .Q(\genblk1[2].u_ce.Xcalc [8])
);

DFFPOSX1 _9786_ (
    .CLK(clk_bF$buf62),
    .D(_1698_),
    .Q(\genblk1[2].u_ce.Xcalc [9])
);

DFFPOSX1 _9787_ (
    .CLK(clk_bF$buf61),
    .D(_1699_),
    .Q(\genblk1[2].u_ce.Xcalc [10])
);

DFFPOSX1 _9788_ (
    .CLK(clk_bF$buf60),
    .D(_1700_),
    .Q(\genblk1[2].u_ce.Xcalc [11])
);

DFFPOSX1 _9789_ (
    .CLK(clk_bF$buf59),
    .D(_1701_),
    .Q(\genblk1[2].u_ce.Acalc [0])
);

DFFPOSX1 _9790_ (
    .CLK(clk_bF$buf58),
    .D(_1702_),
    .Q(\genblk1[2].u_ce.Acalc [1])
);

DFFPOSX1 _9791_ (
    .CLK(clk_bF$buf57),
    .D(_1703_),
    .Q(\genblk1[2].u_ce.Acalc [2])
);

DFFPOSX1 _9792_ (
    .CLK(clk_bF$buf56),
    .D(_1704_),
    .Q(\genblk1[2].u_ce.Acalc [3])
);

DFFPOSX1 _9793_ (
    .CLK(clk_bF$buf55),
    .D(_1705_),
    .Q(\genblk1[2].u_ce.Acalc [4])
);

DFFPOSX1 _9794_ (
    .CLK(clk_bF$buf54),
    .D(_1706_),
    .Q(\genblk1[2].u_ce.Acalc [5])
);

DFFPOSX1 _9795_ (
    .CLK(clk_bF$buf53),
    .D(_1707_),
    .Q(\genblk1[2].u_ce.Acalc [6])
);

DFFPOSX1 _9796_ (
    .CLK(clk_bF$buf52),
    .D(_1708_),
    .Q(\genblk1[2].u_ce.Acalc [7])
);

DFFPOSX1 _9797_ (
    .CLK(clk_bF$buf51),
    .D(_1709_),
    .Q(\genblk1[2].u_ce.Acalc [8])
);

DFFPOSX1 _9798_ (
    .CLK(clk_bF$buf50),
    .D(_1710_),
    .Q(\genblk1[2].u_ce.Acalc [9])
);

DFFPOSX1 _9799_ (
    .CLK(clk_bF$buf49),
    .D(_1711_),
    .Q(\genblk1[2].u_ce.Acalc [10])
);

DFFPOSX1 _9800_ (
    .CLK(clk_bF$buf48),
    .D(_1712_),
    .Q(\genblk1[2].u_ce.Acalc [11])
);

DFFPOSX1 _9801_ (
    .CLK(clk_bF$buf47),
    .D(_1713_),
    .Q(\genblk1[2].u_ce.Xin12b [10])
);

DFFPOSX1 _9802_ (
    .CLK(clk_bF$buf46),
    .D(_1714_),
    .Q(\genblk1[2].u_ce.Xin12b [11])
);

DFFPOSX1 _9803_ (
    .CLK(clk_bF$buf45),
    .D(_1715_),
    .Q(\genblk1[2].u_ce.Xin12b [8])
);

DFFPOSX1 _9804_ (
    .CLK(clk_bF$buf44),
    .D(_1716_),
    .Q(\genblk1[2].u_ce.Xin12b [9])
);

DFFPOSX1 _9805_ (
    .CLK(clk_bF$buf43),
    .D(_1717_),
    .Q(\genblk1[2].u_ce.Xin12b [6])
);

DFFPOSX1 _9806_ (
    .CLK(clk_bF$buf42),
    .D(_1718_),
    .Q(\genblk1[2].u_ce.Xin12b [7])
);

DFFPOSX1 _9807_ (
    .CLK(clk_bF$buf41),
    .D(_1719_),
    .Q(\genblk1[2].u_ce.Xin12b [4])
);

DFFPOSX1 _9808_ (
    .CLK(clk_bF$buf40),
    .D(_1720_),
    .Q(\genblk1[2].u_ce.Xin12b [5])
);

DFFPOSX1 _9809_ (
    .CLK(clk_bF$buf39),
    .D(_1721_),
    .Q(\genblk1[2].u_ce.Xin1 [0])
);

DFFPOSX1 _9810_ (
    .CLK(clk_bF$buf38),
    .D(_1722_),
    .Q(\genblk1[2].u_ce.Xin1 [1])
);

DFFPOSX1 _9811_ (
    .CLK(clk_bF$buf37),
    .D(_1723_),
    .Q(\genblk1[2].u_ce.Xin0 [0])
);

DFFPOSX1 _9812_ (
    .CLK(clk_bF$buf36),
    .D(_1724_),
    .Q(\genblk1[2].u_ce.Xin0 [1])
);

DFFPOSX1 _9813_ (
    .CLK(clk_bF$buf35),
    .D(_1725_),
    .Q(\genblk1[2].u_ce.Yin12b [10])
);

DFFPOSX1 _9814_ (
    .CLK(clk_bF$buf34),
    .D(_1726_),
    .Q(\genblk1[2].u_ce.Yin12b [11])
);

DFFPOSX1 _9815_ (
    .CLK(clk_bF$buf33),
    .D(_1727_),
    .Q(\genblk1[2].u_ce.Yin12b [8])
);

DFFPOSX1 _9816_ (
    .CLK(clk_bF$buf32),
    .D(_1728_),
    .Q(\genblk1[2].u_ce.Yin12b [9])
);

DFFPOSX1 _9817_ (
    .CLK(clk_bF$buf31),
    .D(_1729_),
    .Q(\genblk1[2].u_ce.Yin12b [6])
);

DFFPOSX1 _9818_ (
    .CLK(clk_bF$buf30),
    .D(_1730_),
    .Q(\genblk1[2].u_ce.Yin12b [7])
);

DFFPOSX1 _9819_ (
    .CLK(clk_bF$buf29),
    .D(_1731_),
    .Q(\genblk1[2].u_ce.Yin12b [4])
);

DFFPOSX1 _9820_ (
    .CLK(clk_bF$buf28),
    .D(_1732_),
    .Q(\genblk1[2].u_ce.Yin12b [5])
);

DFFPOSX1 _9821_ (
    .CLK(clk_bF$buf27),
    .D(_1733_),
    .Q(\genblk1[2].u_ce.Yin1 [0])
);

DFFPOSX1 _9822_ (
    .CLK(clk_bF$buf26),
    .D(_1734_),
    .Q(\genblk1[2].u_ce.Yin1 [1])
);

DFFPOSX1 _9823_ (
    .CLK(clk_bF$buf25),
    .D(_1735_),
    .Q(\genblk1[2].u_ce.Yin0 [0])
);

DFFPOSX1 _9824_ (
    .CLK(clk_bF$buf24),
    .D(_1736_),
    .Q(\genblk1[2].u_ce.Yin0 [1])
);

DFFPOSX1 _9825_ (
    .CLK(clk_bF$buf23),
    .D(_1737_),
    .Q(\genblk1[2].u_ce.Ain12b [10])
);

DFFPOSX1 _9826_ (
    .CLK(clk_bF$buf22),
    .D(_1738_),
    .Q(\genblk1[2].u_ce.Ain12b [11])
);

DFFPOSX1 _9827_ (
    .CLK(clk_bF$buf21),
    .D(_1739_),
    .Q(\genblk1[2].u_ce.Ain12b [8])
);

DFFPOSX1 _9828_ (
    .CLK(clk_bF$buf20),
    .D(_1740_),
    .Q(\genblk1[2].u_ce.Ain12b [9])
);

DFFPOSX1 _9829_ (
    .CLK(clk_bF$buf19),
    .D(_1741_),
    .Q(\genblk1[2].u_ce.Ain12b [6])
);

DFFPOSX1 _9830_ (
    .CLK(clk_bF$buf18),
    .D(_1742_),
    .Q(\genblk1[2].u_ce.Ain12b [7])
);

DFFPOSX1 _9831_ (
    .CLK(clk_bF$buf17),
    .D(_1743_),
    .Q(\genblk1[2].u_ce.Ain12b [4])
);

DFFPOSX1 _9832_ (
    .CLK(clk_bF$buf16),
    .D(_1744_),
    .Q(\genblk1[2].u_ce.Ain12b [5])
);

DFFPOSX1 _9833_ (
    .CLK(clk_bF$buf15),
    .D(_1745_),
    .Q(\genblk1[2].u_ce.Ain1 [0])
);

DFFPOSX1 _9834_ (
    .CLK(clk_bF$buf14),
    .D(_1746_),
    .Q(\genblk1[2].u_ce.Ain1 [1])
);

DFFPOSX1 _9835_ (
    .CLK(clk_bF$buf13),
    .D(_1747_),
    .Q(\genblk1[2].u_ce.Ain0 [0])
);

DFFPOSX1 _9836_ (
    .CLK(clk_bF$buf12),
    .D(_1748_),
    .Q(\genblk1[2].u_ce.Ain0 [1])
);

DFFPOSX1 _9837_ (
    .CLK(clk_bF$buf11),
    .D(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[2].u_ce.LoadCtl [0])
);

DFFPOSX1 _9838_ (
    .CLK(clk_bF$buf10),
    .D(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[2].u_ce.LoadCtl [1])
);

DFFPOSX1 _9839_ (
    .CLK(clk_bF$buf9),
    .D(\genblk1[2].u_ce.LoadCtl [1]),
    .Q(\genblk1[2].u_ce.LoadCtl [2])
);

DFFPOSX1 _9840_ (
    .CLK(clk_bF$buf8),
    .D(\genblk1[2].u_ce.LoadCtl [2]),
    .Q(\genblk1[2].u_ce.LoadCtl [3])
);

DFFPOSX1 _9841_ (
    .CLK(clk_bF$buf7),
    .D(\genblk1[2].u_ce.LoadCtl [3]),
    .Q(\genblk1[2].u_ce.LoadCtl [4])
);

DFFPOSX1 _9842_ (
    .CLK(clk_bF$buf6),
    .D(\genblk1[2].u_ce.LoadCtl [4]),
    .Q(\genblk1[2].u_ce.LoadCtl [5])
);

DFFPOSX1 _9843_ (
    .CLK(clk_bF$buf5),
    .D(\genblk1[2].u_ce.LoadCtl [5]),
    .Q(\genblk1[2].u_ce.Vld )
);

INVX1 _9844_ (
    .A(\genblk1[3].u_ce.Acalc [2]),
    .Y(_2594_)
);

INVX2 _9845_ (
    .A(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2595_)
);

NOR2X1 _9846_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_2595_),
    .Y(_2596_)
);

INVX2 _9847_ (
    .A(_2596_),
    .Y(_2597_)
);

NOR2X1 _9848_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [10]),
    .Y(_2598_)
);

INVX4 _9849_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .Y(_2599_)
);

NOR2X1 _9850_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.LoadCtl [3]),
    .Y(_2600_)
);

OAI21X1 _9851_ (
    .A(_2599_),
    .B(\genblk1[3].u_ce.Acalc [8]),
    .C(_2600_),
    .Y(_2601_)
);

INVX2 _9852_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_2602_)
);

AND2X2 _9853_ (
    .A(_2602_),
    .B(\genblk1[3].u_ce.LoadCtl [3]),
    .Y(_2603_)
);

AOI22X1 _9854_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.Acalc [4]),
    .C(_2603_),
    .D(\genblk1[3].u_ce.Acalc [6]),
    .Y(_2604_)
);

OAI21X1 _9855_ (
    .A(_2598_),
    .B(_2601_),
    .C(_2604_),
    .Y(_2605_)
);

NOR2X1 _9856_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2606_)
);

AOI22X1 _9857_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.Acalc [0]),
    .C(_2605_),
    .D(_2606_),
    .Y(_2607_)
);

OAI21X1 _9858_ (
    .A(_2594_),
    .B(_2597_),
    .C(_2607_),
    .Y(\a[4] [0])
);

INVX1 _9859_ (
    .A(\genblk1[3].u_ce.Acalc [9]),
    .Y(_2608_)
);

OAI21X1 _9860_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [11]),
    .C(_2600_),
    .Y(_2609_)
);

AOI21X1 _9861_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2608_),
    .C(_2609_),
    .Y(_2610_)
);

INVX1 _9862_ (
    .A(\genblk1[3].u_ce.Acalc [5]),
    .Y(_2611_)
);

NAND2X1 _9863_ (
    .A(\genblk1[3].u_ce.Acalc [7]),
    .B(_2603_),
    .Y(_2612_)
);

OAI21X1 _9864_ (
    .A(_2602_),
    .B(_2611_),
    .C(_2612_),
    .Y(_2613_)
);

OAI21X1 _9865_ (
    .A(_2610_),
    .B(_2613_),
    .C(_2606_),
    .Y(_2614_)
);

AOI22X1 _9866_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Acalc [1]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Acalc [3]),
    .Y(_2615_)
);

NAND2X1 _9867_ (
    .A(_2615_),
    .B(_2614_),
    .Y(\a[4] [1])
);

INVX1 _9868_ (
    .A(\genblk1[3].u_ce.Ycalc [10]),
    .Y(_2616_)
);

OAI21X1 _9869_ (
    .A(_2599_),
    .B(\genblk1[3].u_ce.Ycalc [8]),
    .C(_2600_),
    .Y(_2617_)
);

AOI21X1 _9870_ (
    .A(_2599_),
    .B(_2616_),
    .C(_2617_),
    .Y(_2618_)
);

INVX1 _9871_ (
    .A(\genblk1[3].u_ce.Ycalc [4]),
    .Y(_2619_)
);

NAND2X1 _9872_ (
    .A(\genblk1[3].u_ce.Ycalc [6]),
    .B(_2603_),
    .Y(_2620_)
);

OAI21X1 _9873_ (
    .A(_2602_),
    .B(_2619_),
    .C(_2620_),
    .Y(_2621_)
);

OAI21X1 _9874_ (
    .A(_2618_),
    .B(_2621_),
    .C(_2606_),
    .Y(_2622_)
);

AOI22X1 _9875_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.Ycalc [0]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Ycalc [2]),
    .Y(_2623_)
);

NAND2X1 _9876_ (
    .A(_2623_),
    .B(_2622_),
    .Y(\genblk1[3].u_ce.Y_ [0])
);

INVX1 _9877_ (
    .A(\genblk1[3].u_ce.Ycalc [9]),
    .Y(_2624_)
);

OAI21X1 _9878_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Ycalc [11]),
    .C(_2600_),
    .Y(_2625_)
);

AOI21X1 _9879_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2624_),
    .C(_2625_),
    .Y(_2626_)
);

INVX1 _9880_ (
    .A(\genblk1[3].u_ce.Ycalc [5]),
    .Y(_2627_)
);

NAND2X1 _9881_ (
    .A(\genblk1[3].u_ce.Ycalc [7]),
    .B(_2603_),
    .Y(_2628_)
);

OAI21X1 _9882_ (
    .A(_2602_),
    .B(_2627_),
    .C(_2628_),
    .Y(_2629_)
);

OAI21X1 _9883_ (
    .A(_2626_),
    .B(_2629_),
    .C(_2606_),
    .Y(_2630_)
);

AOI22X1 _9884_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[3].u_ce.Ycalc [1]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2631_)
);

NAND2X1 _9885_ (
    .A(_2631_),
    .B(_2630_),
    .Y(\genblk1[3].u_ce.Y_ [1])
);

INVX1 _9886_ (
    .A(\genblk1[3].u_ce.Xcalc [8]),
    .Y(_2632_)
);

OAI21X1 _9887_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Xcalc [10]),
    .C(_2600_),
    .Y(_2633_)
);

AOI21X1 _9888_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2632_),
    .C(_2633_),
    .Y(_2634_)
);

INVX1 _9889_ (
    .A(\genblk1[3].u_ce.Xcalc [4]),
    .Y(_2635_)
);

NAND2X1 _9890_ (
    .A(\genblk1[3].u_ce.Xcalc [6]),
    .B(_2603_),
    .Y(_2636_)
);

OAI21X1 _9891_ (
    .A(_2602_),
    .B(_2635_),
    .C(_2636_),
    .Y(_2637_)
);

OAI21X1 _9892_ (
    .A(_2634_),
    .B(_2637_),
    .C(_2606_),
    .Y(_2638_)
);

AOI22X1 _9893_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.Xcalc [0]),
    .C(_2596_),
    .D(\genblk1[3].u_ce.Xcalc [2]),
    .Y(_2639_)
);

NAND2X1 _9894_ (
    .A(_2639_),
    .B(_2638_),
    .Y(\genblk1[3].u_ce.X_ [0])
);

INVX1 _9895_ (
    .A(\genblk1[3].u_ce.Xcalc [3]),
    .Y(_2640_)
);

NOR2X1 _9896_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Xcalc [11]),
    .Y(_2641_)
);

OAI21X1 _9897_ (
    .A(_2599_),
    .B(\genblk1[3].u_ce.Xcalc [9]),
    .C(_2600_),
    .Y(_2642_)
);

AOI22X1 _9898_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.Xcalc [5]),
    .C(_2603_),
    .D(\genblk1[3].u_ce.Xcalc [7]),
    .Y(_2643_)
);

OAI21X1 _9899_ (
    .A(_2641_),
    .B(_2642_),
    .C(_2643_),
    .Y(_2644_)
);

AOI22X1 _9900_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.Xcalc [1]),
    .C(_2644_),
    .D(_2606_),
    .Y(_2645_)
);

OAI21X1 _9901_ (
    .A(_2640_),
    .B(_2597_),
    .C(_2645_),
    .Y(\genblk1[3].u_ce.X_ [1])
);

INVX1 _9902_ (
    .A(\genblk1[3].u_ce.Ycalc [0]),
    .Y(_2646_)
);

INVX1 _9903_ (
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .Y(_2647_)
);

INVX8 _9904_ (
    .A(1'h0),
    .Y(_2648_)
);

INVX8 _9905_ (
    .A(1'h1),
    .Y(_2649_)
);

INVX1 _9906_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_2650_)
);

NAND2X1 _9907_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2651_)
);

OAI21X1 _9908_ (
    .A(1'h1),
    .B(_2650_),
    .C(_2651_),
    .Y(_2652_)
);

INVX1 _9909_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .Y(_2653_)
);

NAND2X1 _9910_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2654_)
);

OAI21X1 _9911_ (
    .A(1'h1),
    .B(_2653_),
    .C(_2654_),
    .Y(_2655_)
);

MUX2X1 _9912_ (
    .A(_2655_),
    .B(_2652_),
    .S(_2649__bF$buf3),
    .Y(_2656_)
);

INVX1 _9913_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2657_)
);

NAND2X1 _9914_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2658_)
);

OAI21X1 _9915_ (
    .A(1'h1),
    .B(_2657_),
    .C(_2658_),
    .Y(_2659_)
);

INVX1 _9916_ (
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .Y(_2660_)
);

NAND2X1 _9917_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_2661_)
);

OAI21X1 _9918_ (
    .A(1'h1),
    .B(_2660_),
    .C(_2661_),
    .Y(_2662_)
);

MUX2X1 _9919_ (
    .A(_2662_),
    .B(_2659_),
    .S(_2649__bF$buf2),
    .Y(_2663_)
);

MUX2X1 _9920_ (
    .A(_2663_),
    .B(_2656_),
    .S(_2648__bF$buf1),
    .Y(_2664_)
);

NOR2X1 _9921_ (
    .A(_2647_),
    .B(_2664_),
    .Y(_2665_)
);

NAND2X1 _9922_ (
    .A(_2647_),
    .B(_2664_),
    .Y(_2666_)
);

INVX1 _9923_ (
    .A(_2666_),
    .Y(_2667_)
);

NAND2X1 _9924_ (
    .A(_2648__bF$buf0),
    .B(_2649__bF$buf1),
    .Y(_2668_)
);

OAI21X1 _9925_ (
    .A(1'h1),
    .B(_2668_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_2669_)
);

INVX2 _9926_ (
    .A(_2669_),
    .Y(_2670_)
);

OAI21X1 _9927_ (
    .A(_2665_),
    .B(_2667_),
    .C(_2670_),
    .Y(_2671_)
);

OAI21X1 _9928_ (
    .A(_2646_),
    .B(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .C(_2671_),
    .Y(_2514_)
);

INVX8 _9929_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_2672_)
);

NAND2X1 _9930_ (
    .A(\genblk1[3].u_ce.Ycalc [1]),
    .B(_2672__bF$buf1),
    .Y(_2673_)
);

NOR2X1 _9931_ (
    .A(1'h1),
    .B(_2668_),
    .Y(_2674_)
);

MUX2X1 _9932_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(\genblk1[3].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_2675_)
);

MUX2X1 _9933_ (
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .B(\genblk1[3].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_2676_)
);

MUX2X1 _9934_ (
    .A(_2676_),
    .B(_2675_),
    .S(_2649__bF$buf0),
    .Y(_2677_)
);

INVX2 _9935_ (
    .A(1'h1),
    .Y(_2678_)
);

NAND2X1 _9936_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(_2678_),
    .Y(_2679_)
);

AOI21X1 _9937_ (
    .A(_2679_),
    .B(_2658_),
    .C(_2649__bF$buf4),
    .Y(_2680_)
);

NAND3X1 _9938_ (
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .B(_2678_),
    .C(_2649__bF$buf3),
    .Y(_2681_)
);

NAND3X1 _9939_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(1'h1),
    .C(_2649__bF$buf2),
    .Y(_2682_)
);

NAND3X1 _9940_ (
    .A(_2648__bF$buf4),
    .B(_2682_),
    .C(_2681_),
    .Y(_2683_)
);

OAI22X1 _9941_ (
    .A(_2680_),
    .B(_2683_),
    .C(_2648__bF$buf3),
    .D(_2677_),
    .Y(_2684_)
);

INVX1 _9942_ (
    .A(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2685_)
);

INVX8 _9943_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_2686_)
);

INVX1 _9944_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2687_)
);

NAND2X1 _9945_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_2688_)
);

OAI21X1 _9946_ (
    .A(1'h1),
    .B(_2687_),
    .C(_2688_),
    .Y(_2689_)
);

INVX1 _9947_ (
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2690_)
);

NAND2X1 _9948_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_2691_)
);

OAI21X1 _9949_ (
    .A(1'h1),
    .B(_2690_),
    .C(_2691_),
    .Y(_2692_)
);

MUX2X1 _9950_ (
    .A(_2692_),
    .B(_2689_),
    .S(_2649__bF$buf1),
    .Y(_2693_)
);

INVX1 _9951_ (
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2694_)
);

NAND2X1 _9952_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [4]),
    .Y(_2695_)
);

OAI21X1 _9953_ (
    .A(1'h1),
    .B(_2694_),
    .C(_2695_),
    .Y(_2696_)
);

INVX1 _9954_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .Y(_2697_)
);

NAND2X1 _9955_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2698_)
);

OAI21X1 _9956_ (
    .A(1'h1),
    .B(_2697_),
    .C(_2698_),
    .Y(_2699_)
);

MUX2X1 _9957_ (
    .A(_2699_),
    .B(_2696_),
    .S(_2649__bF$buf0),
    .Y(_2700_)
);

MUX2X1 _9958_ (
    .A(_2700_),
    .B(_2693_),
    .S(_2648__bF$buf2),
    .Y(_2701_)
);

NAND3X1 _9959_ (
    .A(_2686__bF$buf2),
    .B(_2664_),
    .C(_2701_),
    .Y(_2702_)
);

MUX2X1 _9960_ (
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_2703_)
);

MUX2X1 _9961_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_2704_)
);

MUX2X1 _9962_ (
    .A(_2704_),
    .B(_2703_),
    .S(_2649__bF$buf4),
    .Y(_2705_)
);

MUX2X1 _9963_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_2706_)
);

MUX2X1 _9964_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(\genblk1[3].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_2707_)
);

MUX2X1 _9965_ (
    .A(_2707_),
    .B(_2706_),
    .S(_2649__bF$buf3),
    .Y(_2708_)
);

MUX2X1 _9966_ (
    .A(_2708_),
    .B(_2705_),
    .S(_2648__bF$buf1),
    .Y(_2709_)
);

OAI21X1 _9967_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2684_),
    .C(_2709_),
    .Y(_2710_)
);

AOI21X1 _9968_ (
    .A(_2710_),
    .B(_2702_),
    .C(_2685_),
    .Y(_2711_)
);

INVX1 _9969_ (
    .A(_2711_),
    .Y(_2712_)
);

NAND3X1 _9970_ (
    .A(_2685_),
    .B(_2702_),
    .C(_2710_),
    .Y(_2713_)
);

AND2X2 _9971_ (
    .A(_2712_),
    .B(_2713_),
    .Y(_2714_)
);

OAI21X1 _9972_ (
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .B(_2684_),
    .C(_2714_),
    .Y(_2715_)
);

OR2X2 _9973_ (
    .A(_2714_),
    .B(_2666_),
    .Y(_2716_)
);

AOI21X1 _9974_ (
    .A(_2716_),
    .B(_2715_),
    .C(_2674_),
    .Y(_2717_)
);

OAI21X1 _9975_ (
    .A(_2672__bF$buf0),
    .B(_2717_),
    .C(_2673_),
    .Y(_2515_)
);

INVX1 _9976_ (
    .A(\genblk1[3].u_ce.ISout ),
    .Y(_2718_)
);

NAND2X1 _9977_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .B(\genblk1[2].u_ce.ISout ),
    .Y(_2719_)
);

OAI21X1 _9978_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .B(_2718_),
    .C(_2719_),
    .Y(_2516_)
);

NAND2X1 _9979_ (
    .A(\genblk1[3].u_ce.Ycalc [2]),
    .B(_2672__bF$buf4),
    .Y(_2720_)
);

AOI21X1 _9980_ (
    .A(_2666_),
    .B(_2713_),
    .C(_2711_),
    .Y(_2721_)
);

MUX2X1 _9981_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(\genblk1[3].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_2722_)
);

MUX2X1 _9982_ (
    .A(_2722_),
    .B(_2675_),
    .S(1'h1),
    .Y(_2723_)
);

MUX2X1 _9983_ (
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_2724_)
);

NAND2X1 _9984_ (
    .A(1'h1),
    .B(_2648__bF$buf0),
    .Y(_2725_)
);

OAI22X1 _9985_ (
    .A(_2725_),
    .B(_2676_),
    .C(_2724_),
    .D(_2668_),
    .Y(_2726_)
);

AOI21X1 _9986_ (
    .A(1'h0),
    .B(_2723_),
    .C(_2726_),
    .Y(_2727_)
);

AOI21X1 _9987_ (
    .A(_2709_),
    .B(_2684_),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_2728_)
);

NAND2X1 _9988_ (
    .A(_2727_),
    .B(_2728_),
    .Y(_2729_)
);

INVX1 _9989_ (
    .A(_2727_),
    .Y(_2730_)
);

OAI21X1 _9990_ (
    .A(_2664_),
    .B(_2701_),
    .C(_2686__bF$buf1),
    .Y(_2731_)
);

NAND2X1 _9991_ (
    .A(_2730_),
    .B(_2731_),
    .Y(_2732_)
);

AOI21X1 _9992_ (
    .A(_2732_),
    .B(_2729_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2733_)
);

NAND3X1 _9993_ (
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .B(_2729_),
    .C(_2732_),
    .Y(_2734_)
);

INVX1 _9994_ (
    .A(_2734_),
    .Y(_2735_)
);

OR2X2 _9995_ (
    .A(_2735_),
    .B(_2733_),
    .Y(_2736_)
);

NOR2X1 _9996_ (
    .A(_2721_),
    .B(_2736_),
    .Y(_2737_)
);

INVX1 _9997_ (
    .A(_2737_),
    .Y(_2738_)
);

OAI21X1 _9998_ (
    .A(_2733_),
    .B(_2735_),
    .C(_2721_),
    .Y(_2739_)
);

AOI21X1 _9999_ (
    .A(_2738_),
    .B(_2739_),
    .C(_2674_),
    .Y(_2740_)
);

endmodule
