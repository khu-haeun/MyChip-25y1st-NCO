magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect -122 -162 306 734
<< ntransistor >>
rect 103 480 113 604
<< ptransistor >>
rect 43 0 53 124
rect 103 0 113 124
<< ndiffusion >>
rect 60 562 103 604
rect 60 550 72 562
rect 84 550 103 562
rect 60 506 103 550
rect 60 494 72 506
rect 84 494 103 506
rect 60 480 103 494
rect 113 562 156 604
rect 113 550 132 562
rect 144 550 156 562
rect 113 506 156 550
rect 113 494 132 506
rect 144 494 156 506
rect 113 480 156 494
<< ndcontact >>
rect 72 550 84 562
rect 72 494 84 506
rect 132 550 144 562
rect 132 494 144 506
<< psubstratepdiff >>
rect 0 110 43 124
rect 0 98 12 110
rect 24 98 43 110
rect 0 54 43 98
rect 0 42 12 54
rect 24 42 43 54
rect 0 0 43 42
rect 53 110 103 124
rect 53 98 72 110
rect 84 98 103 110
rect 53 54 103 98
rect 53 42 72 54
rect 84 42 103 54
rect 53 0 103 42
rect 113 110 156 124
rect 113 98 132 110
rect 144 98 156 110
rect 113 54 156 98
rect 113 42 132 54
rect 144 42 156 54
rect 113 0 156 42
<< psubstratepcontact >>
rect 12 98 24 110
rect 12 42 24 54
rect 72 98 84 110
rect 72 42 84 54
rect 132 98 144 110
rect 132 42 144 54
<< polysilicon >>
rect 103 604 113 614
rect 103 456 113 480
rect 43 124 53 148
rect 103 124 113 148
rect 43 -10 53 0
rect 103 -10 113 0
<< genericcontact >>
rect 72 550 84 562
rect 132 550 144 562
rect 72 494 84 506
rect 132 494 144 506
rect 12 98 24 110
rect 72 98 84 110
rect 132 98 144 110
rect 12 42 24 54
rect 72 42 84 54
rect 132 42 144 54
<< metal1 >>
rect 58 562 100 606
rect 58 550 72 562
rect 84 550 100 562
rect 58 506 100 550
rect 58 494 72 506
rect 84 494 100 506
rect 58 478 100 494
rect 116 562 158 606
rect 116 550 132 562
rect 144 550 158 562
rect 116 506 158 550
rect 116 494 132 506
rect 144 494 158 506
rect 116 478 158 494
rect 30 418 126 462
rect 2 146 126 186
rect -2 110 40 126
rect -2 98 12 110
rect 24 98 40 110
rect -2 54 40 98
rect -2 42 12 54
rect 24 42 40 54
rect -2 -18 40 42
rect 56 110 100 126
rect 56 98 72 110
rect 84 98 100 110
rect 56 54 100 98
rect 56 42 72 54
rect 84 42 100 54
rect 56 -2 100 42
rect 116 110 158 126
rect 116 98 132 110
rect 144 98 158 110
rect 116 54 158 98
rect 116 42 132 54
rect 144 42 158 54
rect 116 -18 158 42
rect -2 -42 158 -18
<< metal2 >>
rect 58 478 98 606
rect 118 526 158 606
rect 118 478 186 526
rect 30 418 126 458
rect 78 186 106 418
rect 2 146 126 186
rect 146 126 186 478
rect 58 -2 98 126
rect 118 78 186 126
rect 118 -2 158 78
<< metal3 >>
rect 58 478 98 606
rect 58 -2 98 126
rect 118 -2 158 126
use CONT$4  CONT$4_0
timestamp 1569543463
transform -1 0 18 0 -1 76
box -6 -6 6 6
use CONT$4  CONT$4_1
timestamp 1569543463
transform -1 0 18 0 -1 20
box -6 -6 6 6
use poly1cont_CDNS_704676826053$2  poly1cont_CDNS_704676826053$2_0
timestamp 1569543463
transform 1 0 90 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053$2  poly1cont_CDNS_704676826053$2_1
timestamp 1569543463
transform -1 0 126 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053$2  poly1cont_CDNS_704676826053$2_2
timestamp 1569543463
transform 1 0 30 0 1 146
box 0 0 36 36
use VIA1$4  VIA1$4_0
timestamp 1569543463
transform -1 0 138 0 -1 76
box -8 -8 8 8
use VIA1$4  VIA1$4_1
timestamp 1569543463
transform 1 0 78 0 1 528
box -8 -8 8 8
use VIA1$4  VIA1$4_2
timestamp 1569543463
transform 1 0 78 0 1 584
box -8 -8 8 8
use VIA1$4  VIA1$4_3
timestamp 1569543463
transform 1 0 138 0 1 528
box -8 -8 8 8
use VIA1$4  VIA1$4_4
timestamp 1569543463
transform -1 0 138 0 -1 20
box -8 -8 8 8
use VIA1$4  VIA1$4_5
timestamp 1569543463
transform 1 0 50 0 1 438
box -8 -8 8 8
use VIA1$4  VIA1$4_6
timestamp 1569543463
transform 1 0 22 0 1 166
box -8 -8 8 8
use VIA1$4  VIA1$4_7
timestamp 1569543463
transform -1 0 78 0 -1 76
box -8 -8 8 8
use VIA1$4  VIA1$4_8
timestamp 1569543463
transform 1 0 138 0 1 584
box -8 -8 8 8
use VIA1$4  VIA1$4_9
timestamp 1569543463
transform 1 0 78 0 1 166
box -8 -8 8 8
use VIA1$4  VIA1$4_10
timestamp 1569543463
transform 1 0 82 0 1 438
box -8 -8 8 8
use VIA1$4  VIA1$4_11
timestamp 1569543463
transform -1 0 78 0 -1 20
box -8 -8 8 8
use VIA2$4  VIA2$4_0
timestamp 1569543463
transform 1 0 78 0 1 500
box -8 -8 8 8
use VIA2$4  VIA2$4_1
timestamp 1569543463
transform -1 0 78 0 -1 48
box -8 -8 8 8
use VIA2$4  VIA2$4_2
timestamp 1569543463
transform 1 0 78 0 1 556
box -8 -8 8 8
use VIA2$4  VIA2$4_3
timestamp 1569543463
transform -1 0 78 0 -1 104
box -8 -8 8 8
<< end >>
