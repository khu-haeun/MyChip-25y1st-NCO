magic
tech scmos
magscale 1 30
timestamp 1740931377
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 58700 143400 140900 144900
rect 139800 139100 140900 143400
rect 48300 132600 50500 138400
rect 73700 46700 119700 47100
rect 60200 45900 120500 46300
<< m2contact >>
rect 50300 143400 58700 144900
rect 45400 132600 48300 138400
rect 73300 46700 73700 47100
rect 119700 46700 120100 47100
rect 59800 45900 60200 46300
rect 120500 45900 120900 46300
<< metal2 >>
rect 50300 144900 58700 145900
rect 62400 140400 62900 145900
rect 75900 142300 76400 145900
rect 89400 142500 89900 145900
rect 102900 141400 103400 145900
rect 102900 140900 126800 141400
rect 62400 139900 117585 140400
rect 126300 140000 126800 140900
rect 131700 140000 132200 142000
rect 44000 132600 45400 138400
rect 144200 129900 145900 130400
rect 44100 116300 45100 116800
rect 143200 116400 145900 116900
rect 44100 102800 46100 103300
rect 47100 89800 47600 112000
rect 44100 89300 47600 89800
rect 48100 76300 48600 111300
rect 143300 102900 145900 103400
rect 144300 89400 145900 89900
rect 44100 75800 48600 76300
rect 44100 48700 46900 49400
rect 75800 48300 76200 48900
rect 76600 47500 77000 48900
rect 59800 44100 60200 45900
rect 73300 44100 73700 46700
rect 78600 46700 79000 48900
rect 80300 45900 80700 48900
rect 81100 44900 81500 48900
rect 119700 47100 120100 48900
rect 81100 44500 87200 44900
rect 86800 44100 87200 44500
rect 100300 44100 100700 45500
rect 113700 44100 114100 46300
rect 120500 46300 120900 48900
rect 127300 44100 127700 47100
rect 140800 44100 141200 47900
<< m3contact >>
rect 75900 140800 76400 142300
rect 89400 142000 89900 142500
rect 131700 142000 132200 142500
rect 142700 129900 144200 130400
rect 45100 115300 45600 116800
rect 141700 116400 143200 116900
rect 47100 112000 47600 113500
rect 46100 102800 46600 104300
rect 48100 111300 48600 112800
rect 141800 102900 143300 103400
rect 142800 89400 144300 89900
rect 46900 48700 49000 49400
rect 75800 47900 76200 48300
rect 76600 47100 77000 47500
rect 78600 46300 79000 46700
rect 80300 45500 80700 45900
rect 113700 46300 114100 46700
rect 100300 45500 100700 45900
rect 140800 47900 141200 48300
rect 127300 47100 127700 47500
<< metal3 >>
rect 89900 142000 131700 142500
rect 76400 140800 86700 141300
rect 86200 139500 86700 140800
rect 140300 137900 143200 138400
rect 48700 137100 50400 137600
rect 48700 131300 49100 137100
rect 140300 137000 142200 137500
rect 46100 130800 49100 131300
rect 45100 98000 45600 115300
rect 46100 104300 46600 130800
rect 141700 116900 142200 137000
rect 142700 130400 143200 137900
rect 47600 113100 50500 113500
rect 48600 112400 50500 112800
rect 45100 97500 50400 98000
rect 141800 83600 142300 102900
rect 140200 83100 142300 83600
rect 142800 80200 143300 89400
rect 140200 79700 143300 80200
rect 48300 68900 50400 69600
rect 48300 49400 49000 68900
rect 76200 47900 140800 48300
rect 77000 47100 127300 47500
rect 79000 46300 113700 46700
rect 80700 45500 100300 45900
<< end >>
