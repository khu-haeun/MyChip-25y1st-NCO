//      // verilator_coverage annotation
        /* Verilog module written by vlog2Verilog (qflow) */
        
        module cordic_element(
 037078     input [1:0] Ain,
 037853     output [1:0] Aout,
 001963     input ISin,
 001956     output ISout,
 039624     input Rdy,
 381100     input [2:0] Stg,
 114044     output Vld,
 051639     input [1:0] Xin,
 057160     output [1:0] Xout,
 049025     input [1:0] Yin,
 054951     output [1:0] Yout,
 362248     input clk
        );
        /* verilator coverage_off */
        wire vdd = 1'b1;
        wire gnd = 1'b0;
        /* verilator coverage_on */
        
        wire _588_ ;
        wire _168_ ;
        wire _800_ ;
        wire _60_ ;
        wire _397_ ;
        wire _703_ ;
        wire _19_ ;
        wire _512_ ;
 114044 wire [6:0] LoadCtl ;
        wire _741_ ;
        wire _321_ ;
        wire _57_ ;
        wire _550_ ;
        wire _130_ ;
        wire _606_ ;
        wire _835_ ;
        wire _415_ ;
        wire _95_ ;
        wire _644_ ;
        wire _224_ ;
        wire _453_ ;
        wire _509_ ;
        wire _682_ ;
        wire _262_ ;
        wire _738_ ;
        wire _318_ ;
        wire _491_ ;
        wire _547_ ;
        wire _127_ ;
        wire _776_ ;
        wire _356_ ;
        wire _585_ ;
        wire _165_ ;
        wire _394_ ;
        wire _679_ ;
        wire _259_ ;
        wire _488_ ;
        wire _700_ ;
        wire _297_ ;
        wire _16_ ;
        wire _54_ ;
        wire _603_ ;
        wire _832_ ;
        wire _412_ ;
        wire _92_ ;
        wire _641_ ;
        wire _221_ ;
        wire _450_ ;
        //wire ISin ;
        wire _506_ ;
 005205 wire [11:0] Acalc ;
        wire _735_ ;
        wire _315_ ;
        wire _544_ ;
        wire _124_ ;
        wire _773_ ;
        wire _353_ ;
        wire _829_ ;
        wire _409_ ;
        wire _89_ ;
        wire _582_ ;
        wire _162_ ;
        wire _638_ ;
        wire _218_ ;
        wire _391_ ;
        wire _447_ ;
        wire _676_ ;
        wire _256_ ;
        wire _485_ ;
        wire _294_ ;
        wire _13_ ;
        wire _579_ ;
        wire _159_ ;
        wire _51_ ;
        wire _388_ ;
        wire _600_ ;
        //wire Rdy ;
        wire _197_ ;
        wire _7_ ;
        wire _503_ ;
        wire _732_ ;
        wire _312_ ;
        wire _48_ ;
        wire _541_ ;
        wire _121_ ;
        //wire ISout ;
        wire _770_ ;
        wire _350_ ;
        wire _826_ ;
        wire _406_ ;
        wire _86_ ;
        wire _635_ ;
        wire _215_ ;
        wire _444_ ;
        wire _673_ ;
        wire _253_ ;
        wire _729_ ;
        wire _309_ ;
        wire _482_ ;
        wire _538_ ;
        wire _118_ ;
        wire _291_ ;
        wire _10_ ;
        wire _767_ ;
        wire _347_ ;
        wire _576_ ;
        wire _156_ ;
        wire _385_ ;
        wire _194_ ;
        wire _479_ ;
        wire _288_ ;
        wire _4_ ;
        wire _500_ ;
        wire _45_ ;
        wire _823_ ;
        wire _403_ ;
        wire _83_ ;
        wire _632_ ;
        wire _212_ ;
        wire [1:0] _861_ ;
        wire _441_ ;
        wire _670_ ;
        wire _250_ ;
        wire _726_ ;
        wire _306_ ;
        wire _535_ ;
        wire _115_ ;
        wire _764_ ;
        wire _344_ ;
        wire _573_ ;
        wire _153_ ;
        wire _629_ ;
        wire _209_ ;
        wire _382_ ;
        wire _858_ ;
        wire _438_ ;
        wire _191_ ;
        wire _667_ ;
        wire _247_ ;
        wire _476_ ;
 362248 wire clk_bF$buf0 ;
 362248 wire clk_bF$buf1 ;
 362248 wire clk_bF$buf2 ;
 362248 wire clk_bF$buf3 ;
 362248 wire clk_bF$buf4 ;
 362248 wire clk_bF$buf5 ;
 362248 wire clk_bF$buf6 ;
 362248 wire clk_bF$buf7 ;
        wire _285_ ;
        wire _1_ ;
        //wire [2:0] Stg ;
        wire _42_ ;
        wire _799_ ;
        wire _379_ ;
        wire _188_ ;
        wire _820_ ;
        wire _400_ ;
        wire _80_ ;
        wire _723_ ;
        wire _303_ ;
        wire _39_ ;
        wire _532_ ;
        wire _112_ ;
        wire _761_ ;
        wire _341_ ;
        //wire clk ;
        wire _817_ ;
        wire _77_ ;
        wire _570_ ;
        wire _150_ ;
        wire _626_ ;
        wire _206_ ;
        wire _855_ ;
        wire _435_ ;
        wire _664_ ;
        wire _244_ ;
        wire _473_ ;
        wire _529_ ;
        wire _109_ ;
        wire _282_ ;
        wire _758_ ;
        wire _338_ ;
        wire _567_ ;
        wire _147_ ;
        wire _796_ ;
        wire _376_ ;
        wire _185_ ;
        wire _699_ ;
        wire _279_ ;
        wire _720_ ;
        wire _300_ ;
        wire _36_ ;
        wire _814_ ;
        wire _74_ ;
        wire _623_ ;
        wire _203_ ;
        wire _852_ ;
        wire _432_ ;
        wire _661_ ;
        wire _241_ ;
        wire _717_ ;
        wire _470_ ;
        wire _526_ ;
        wire _106_ ;
        wire _755_ ;
        wire _335_ ;
        wire _564_ ;
        wire _144_ ;
        wire _793_ ;
        wire _373_ ;
        wire _849_ ;
        wire _429_ ;
        wire _182_ ;
 039616 wire LoadCtl_0_bF$buf0 ;
 039616 wire LoadCtl_0_bF$buf1 ;
 039616 wire LoadCtl_0_bF$buf2 ;
 039616 wire LoadCtl_0_bF$buf3 ;
        wire _658_ ;
        wire _238_ ;
        wire _467_ ;
        wire _696_ ;
        wire _276_ ;
 381100 wire Stg_0_bF$buf0 ;
 381100 wire Stg_0_bF$buf1 ;
 381100 wire Stg_0_bF$buf2 ;
 381100 wire Stg_0_bF$buf3 ;
 381100 wire Stg_0_bF$buf4 ;
 381100 wire Stg_0_bF$buf5 ;
 381100 wire Stg_0_bF$buf6 ;
        wire _33_ ;
        wire _599_ ;
        wire _179_ ;
        wire _811_ ;
        wire _71_ ;
        wire _620_ ;
        wire _200_ ;
 003598 wire [11:0] Ycalc ;
        wire _714_ ;
        wire _523_ ;
        wire _103_ ;
        wire _752_ ;
        wire _332_ ;
        wire _808_ ;
        wire _68_ ;
        wire _561_ ;
        wire _141_ ;
        wire _617_ ;
        wire _790_ ;
        wire _370_ ;
        wire _846_ ;
        wire _426_ ;
        wire _655_ ;
        wire _235_ ;
        wire _464_ ;
        wire _693_ ;
        wire _273_ ;
        wire _749_ ;
        wire _329_ ;
        wire _558_ ;
        wire _138_ ;
        wire _30_ ;
        wire _787_ ;
        wire _367_ ;
        wire _596_ ;
        wire _176_ ;
        wire _499_ ;
        wire _711_ ;
        wire _27_ ;
        wire _520_ ;
        wire _100_ ;
        wire _805_ ;
        wire _65_ ;
        wire _614_ ;
        wire _843_ ;
        wire _423_ ;
        wire _652_ ;
        wire _232_ ;
        wire _708_ ;
        wire _461_ ;
        wire _517_ ;
        wire _690_ ;
        wire _270_ ;
        wire _746_ ;
        wire _326_ ;
        wire _555_ ;
        wire _135_ ;
        wire _784_ ;
        wire _364_ ;
        wire _593_ ;
        wire _173_ ;
        wire _649_ ;
        wire _229_ ;
        wire _458_ ;
        wire _687_ ;
        wire _267_ ;
        wire _496_ ;
        wire _24_ ;
        wire _802_ ;
        wire _62_ ;
        wire _399_ ;
        wire _611_ ;
        wire _840_ ;
        wire _420_ ;
        wire _705_ ;
        wire _514_ ;
        wire _743_ ;
        wire _323_ ;
        wire _59_ ;
        wire _552_ ;
        wire _132_ ;
        wire _608_ ;
        wire _781_ ;
        wire _361_ ;
        wire _837_ ;
        wire _417_ ;
        wire _97_ ;
        wire _590_ ;
        wire _170_ ;
        wire _646_ ;
        wire _226_ ;
        wire _188__bF$buf0 ;
        wire _188__bF$buf1 ;
        wire _188__bF$buf2 ;
        wire _188__bF$buf3 ;
        wire _188__bF$buf4 ;
        wire _455_ ;
        wire _684_ ;
        wire _264_ ;
        wire _493_ ;
        wire _549_ ;
        wire _129_ ;
        wire _21_ ;
        wire _778_ ;
        wire _358_ ;
        wire _587_ ;
        wire _167_ ;
        wire _396_ ;
        wire _702_ ;
        wire _299_ ;
        wire _18_ ;
        wire _511_ ;
        wire _740_ ;
        wire _320_ ;
        wire _56_ ;
        wire _605_ ;
        wire _834_ ;
        wire _414_ ;
        wire _94_ ;
        wire _643_ ;
        wire _223_ ;
        wire _452_ ;
        wire _508_ ;
        wire _681_ ;
        wire _261_ ;
        wire _737_ ;
        wire _317_ ;
        wire _490_ ;
        wire _546_ ;
        wire _126_ ;
        wire _775_ ;
        wire _355_ ;
        wire _584_ ;
        wire _164_ ;
        wire _393_ ;
        wire _449_ ;
        wire _678_ ;
        wire _258_ ;
        wire _487_ ;
        wire _296_ ;
        wire _15_ ;
 014431 wire [1:0] Ain0 ;
 025480 wire [1:0] Ain1 ;
        wire _53_ ;
        wire _602_ ;
        wire _199_ ;
        wire _831_ ;
        wire _411_ ;
        wire _91_ ;
        wire _640_ ;
        wire _220_ ;
        wire _9_ ;
        wire _505_ ;
        wire _734_ ;
        wire _314_ ;
        wire _543_ ;
        wire _123_ ;
        wire _772_ ;
        wire _352_ ;
        wire _828_ ;
        wire _408_ ;
        wire _88_ ;
 381100 wire Stg_2_bF$buf0 ;
 381100 wire Stg_2_bF$buf1 ;
 381100 wire Stg_2_bF$buf2 ;
 381100 wire Stg_2_bF$buf3 ;
 381100 wire Stg_2_bF$buf4 ;
        wire _581_ ;
        wire _161_ ;
        wire _637_ ;
        wire _217_ ;
        wire _390_ ;
        wire _446_ ;
~002595 wire [11:0] Xin12b ;
        //wire [1:0] Yin ;
        wire _675_ ;
        wire _255_ ;
        wire _484_ ;
        wire _293_ ;
        wire _12_ ;
        wire _769_ ;
        wire _349_ ;
        wire _578_ ;
        wire _158_ ;
        wire _50_ ;
        wire _387_ ;
        wire _196_ ;
        wire _6_ ;
        wire _502_ ;
        wire _731_ ;
        wire _311_ ;
        wire _47_ ;
        wire _540_ ;
        wire _120_ ;
        wire _825_ ;
        wire _405_ ;
        wire _85_ ;
 003184 wire [11:0] Xcalc ;
 003724 wire [1:0] Yin0 ;
 004258 wire [1:0] Yin1 ;
        wire _634_ ;
        wire _214_ ;
        wire _443_ ;
        wire _672_ ;
        wire _252_ ;
        wire _728_ ;
        wire _308_ ;
        wire _481_ ;
        wire _537_ ;
        wire _117_ ;
        wire _290_ ;
        wire _766_ ;
        wire _346_ ;
        wire _575_ ;
        wire _155_ ;
        wire _384_ ;
        //wire [1:0] Aout ;
        wire _193_ ;
        wire _669_ ;
        wire _249_ ;
        wire _478_ ;
        wire _287_ ;
        wire _3_ ;
        wire _44_ ;
        wire _201__bF$buf0 ;
        wire _201__bF$buf1 ;
        wire _201__bF$buf2 ;
        wire _201__bF$buf3 ;
        wire _201__bF$buf4 ;
        wire _201__bF$buf5 ;
        wire _201__bF$buf6 ;
        wire _822_ ;
        wire _402_ ;
        wire _82_ ;
        wire _631_ ;
        wire _211_ ;
        wire _860_ ;
        wire _440_ ;
        wire _725_ ;
        wire _305_ ;
 004705 wire [1:0] Xin0 ;
 002300 wire [1:0] Xin1 ;
        wire _534_ ;
        wire _114_ ;
 003012 wire Ain12b_11_bF$buf0 ;
 003012 wire Ain12b_11_bF$buf1 ;
 003012 wire Ain12b_11_bF$buf2 ;
 003012 wire Ain12b_11_bF$buf3 ;
 003012 wire Ain12b_11_bF$buf4 ;
        wire _763_ ;
        wire _343_ ;
        wire _819_ ;
        wire _79_ ;
        wire _572_ ;
        wire _152_ ;
        wire _628_ ;
        wire _208_ ;
        wire _381_ ;
        wire _857_ ;
        wire _437_ ;
        wire _190_ ;
        wire _666_ ;
        wire _246_ ;
        wire _475_ ;
        wire _284_ ;
        wire _0_ ;
        wire _569_ ;
        wire _149_ ;
        wire _41_ ;
        wire _798_ ;
        wire _378_ ;
        wire _187_ ;
        //wire [1:0] Yout ;
        wire _722_ ;
        wire _302_ ;
        wire _38_ ;
        wire _531_ ;
        wire _111_ ;
        wire _760_ ;
        wire _340_ ;
        wire _816_ ;
        wire _76_ ;
        //wire [1:0] Ain ;
        wire _625_ ;
        wire _205_ ;
        wire _854_ ;
        wire _434_ ;
        wire _663_ ;
        wire _243_ ;
        wire _719_ ;
        wire _472_ ;
        wire _528_ ;
        wire _108_ ;
        wire _281_ ;
        wire _757_ ;
        wire _337_ ;
        wire _566_ ;
        wire _146_ ;
        wire _795_ ;
        wire _375_ ;
        wire _184_ ;
        wire _469_ ;
        wire _698_ ;
        wire _278_ ;
        wire _35_ ;
        //wire [1:0] Xout ;
        wire _813_ ;
        wire _73_ ;
        wire _622_ ;
        wire _202_ ;
        wire _851_ ;
        wire _431_ ;
        wire _660_ ;
        wire _240_ ;
        wire _716_ ;
        wire _525_ ;
        wire _105_ ;
        wire _754_ ;
        wire _334_ ;
        wire _563_ ;
        wire _143_ ;
        wire _619_ ;
        wire _792_ ;
        wire _372_ ;
        wire _848_ ;
        wire _428_ ;
        wire _181_ ;
        wire _657_ ;
        wire _237_ ;
        wire _466_ ;
~012931 wire [11:0] Ain12b ;
        wire _695_ ;
        wire _275_ ;
        wire _32_ ;
        wire _789_ ;
        wire _369_ ;
        wire _598_ ;
        wire _178_ ;
        wire _810_ ;
        wire _70_ ;
        wire _713_ ;
        wire _29_ ;
        wire _522_ ;
        wire _102_ ;
        wire _751_ ;
        wire _331_ ;
        wire _807_ ;
        wire _67_ ;
        wire _560_ ;
        wire _140_ ;
        wire _616_ ;
        wire _845_ ;
        wire _425_ ;
        wire _654_ ;
        wire _234_ ;
        wire _463_ ;
        wire _519_ ;
        wire _692_ ;
        wire _272_ ;
        wire _748_ ;
        wire _328_ ;
        wire _557_ ;
        wire _137_ ;
        wire _786_ ;
        wire _366_ ;
        wire _595_ ;
        wire _175_ ;
        wire _689_ ;
        wire _269_ ;
        wire _498_ ;
        wire _710_ ;
        wire _26_ ;
        wire _804_ ;
        wire _64_ ;
        wire _613_ ;
        wire _842_ ;
        wire _422_ ;
        wire _651_ ;
        wire _231_ ;
        wire _707_ ;
        wire _460_ ;
        wire _516_ ;
        wire _745_ ;
        wire _325_ ;
        wire _554_ ;
        wire _134_ ;
        wire _783_ ;
        wire _363_ ;
        wire _839_ ;
        wire _419_ ;
        wire _99_ ;
        wire _592_ ;
        wire _172_ ;
        //wire Vld ;
        wire _648_ ;
        wire _228_ ;
        wire _457_ ;
        wire _686_ ;
        wire _266_ ;
        wire _495_ ;
        wire _23_ ;
        wire _589_ ;
        wire _169_ ;
        wire _801_ ;
        wire _61_ ;
        wire _398_ ;
        wire _610_ ;
        wire _704_ ;
        wire _513_ ;
        wire _742_ ;
        wire _322_ ;
        wire _58_ ;
        wire _551_ ;
        wire _131_ ;
        wire _607_ ;
        wire _780_ ;
        wire _360_ ;
        wire _836_ ;
        wire _416_ ;
        wire _96_ ;
        wire _645_ ;
        wire _225_ ;
        wire _454_ ;
        wire _683_ ;
        wire _263_ ;
        wire _739_ ;
        wire _319_ ;
        wire _492_ ;
        wire _548_ ;
        wire _128_ ;
        wire _20_ ;
        wire _777_ ;
        wire _357_ ;
        wire _586_ ;
        wire _166_ ;
        wire _395_ ;
        wire _164__bF$buf0 ;
        wire _164__bF$buf1 ;
        wire _164__bF$buf2 ;
        wire _164__bF$buf3 ;
        wire _164__bF$buf4 ;
        wire _489_ ;
        wire _701_ ;
        wire _298_ ;
        wire _17_ ;
        wire _510_ ;
        wire _55_ ;
        wire _604_ ;
        wire _183__bF$buf0 ;
        wire _183__bF$buf1 ;
        wire _183__bF$buf2 ;
        wire _183__bF$buf3 ;
        wire _833_ ;
        wire _413_ ;
        wire _93_ ;
        wire _642_ ;
        wire _222_ ;
        wire _451_ ;
        wire _507_ ;
        wire _680_ ;
        wire _260_ ;
        wire _736_ ;
        wire _316_ ;
        wire _545_ ;
        wire _125_ ;
        wire _774_ ;
        wire _354_ ;
        wire _583_ ;
        wire _163_ ;
        wire _639_ ;
        wire _219_ ;
        wire _392_ ;
        wire _448_ ;
        wire _677_ ;
        wire _257_ ;
        wire _486_ ;
        wire _295_ ;
        wire _14_ ;
        wire _52_ ;
        wire _389_ ;
        wire _601_ ;
        wire _198_ ;
        wire _830_ ;
        wire _410_ ;
        wire _90_ ;
        wire _8_ ;
        wire _504_ ;
        wire _733_ ;
        wire _313_ ;
        wire _49_ ;
        wire _542_ ;
        wire _122_ ;
        wire _771_ ;
        wire _351_ ;
        wire _827_ ;
        wire _407_ ;
        wire _87_ ;
        wire _580_ ;
        wire _160_ ;
        wire _636_ ;
        wire _216_ ;
        wire _445_ ;
        wire _674_ ;
        wire _254_ ;
        wire _483_ ;
 114044 wire LoadCtl_6_bF$buf0 ;
 114044 wire LoadCtl_6_bF$buf1 ;
 114044 wire LoadCtl_6_bF$buf2 ;
 114044 wire LoadCtl_6_bF$buf3 ;
 114044 wire LoadCtl_6_bF$buf4 ;
        wire _539_ ;
        wire _119_ ;
        wire _292_ ;
        wire _11_ ;
        wire _768_ ;
        wire _348_ ;
~002879 wire [11:0] Yin12b ;
        wire _577_ ;
        wire _157_ ;
        wire _386_ ;
        wire _195_ ;
        wire _289_ ;
        wire _5_ ;
        wire _501_ ;
        wire _730_ ;
        wire _310_ ;
        wire _46_ ;
        wire _824_ ;
        wire _404_ ;
        wire _84_ ;
        wire _633_ ;
        wire _213_ ;
        wire [1:0] _862_ ;
        wire _442_ ;
        wire _671_ ;
        wire _251_ ;
        wire _727_ ;
        wire _307_ ;
        wire _480_ ;
        wire _536_ ;
        wire _116_ ;
        wire _765_ ;
        wire _345_ ;
        wire _574_ ;
        wire _154_ ;
        wire _383_ ;
        wire [1:0] _859_ ;
        wire _439_ ;
        wire _192_ ;
        wire _668_ ;
        wire _248_ ;
        wire _477_ ;
        wire _286_ ;
        wire _2_ ;
        wire _43_ ;
        wire _189_ ;
        wire _821_ ;
        wire _401_ ;
        wire _81_ ;
        wire _630_ ;
        wire _210_ ;
 381100 wire Stg_1_bF$buf0 ;
 381100 wire Stg_1_bF$buf1 ;
 381100 wire Stg_1_bF$buf2 ;
 381100 wire Stg_1_bF$buf3 ;
        wire _724_ ;
        wire _304_ ;
        wire _533_ ;
        wire _113_ ;
        wire _762_ ;
        wire _342_ ;
        wire _818_ ;
        wire _78_ ;
        wire _571_ ;
        wire _151_ ;
        wire _627_ ;
        wire _207_ ;
        wire _380_ ;
        wire _856_ ;
        wire _436_ ;
        //wire [1:0] Xin ;
        wire _665_ ;
        wire _245_ ;
        wire _474_ ;
        wire _283_ ;
        wire _759_ ;
        wire _339_ ;
        wire _568_ ;
        wire _148_ ;
        wire _40_ ;
        wire _797_ ;
        wire _377_ ;
        wire _186_ ;
        wire _721_ ;
        wire _301_ ;
        wire _37_ ;
        wire _530_ ;
        wire _110_ ;
        wire _815_ ;
        wire _75_ ;
        wire _624_ ;
        wire _204_ ;
        wire _853_ ;
        wire _433_ ;
        wire _662_ ;
        wire _242_ ;
        wire _718_ ;
        wire _471_ ;
        wire _527_ ;
        wire _107_ ;
        wire _280_ ;
        wire _756_ ;
        wire _336_ ;
        wire _565_ ;
        wire _145_ ;
        wire _794_ ;
        wire _374_ ;
        wire _183_ ;
        wire _659_ ;
        wire _239_ ;
        wire _468_ ;
        wire _697_ ;
        wire _277_ ;
        wire _34_ ;
        wire _812_ ;
        wire _72_ ;
        wire _621_ ;
        wire _201_ ;
        wire _850_ ;
        wire _430_ ;
        wire _715_ ;
        wire _524_ ;
        wire _104_ ;
        wire _753_ ;
        wire _333_ ;
        wire _809_ ;
        wire _69_ ;
        wire _562_ ;
        wire _142_ ;
        wire _618_ ;
        wire _791_ ;
        wire _371_ ;
        wire _847_ ;
        wire _427_ ;
        wire _180_ ;
        wire _656_ ;
        wire _236_ ;
        wire _465_ ;
        wire _694_ ;
        wire _274_ ;
        wire _559_ ;
        wire _139_ ;
        wire _31_ ;
        wire _788_ ;
        wire _368_ ;
        wire _597_ ;
        wire _177_ ;
        wire _712_ ;
        wire _28_ ;
        wire _521_ ;
        wire _101_ ;
        wire _750_ ;
        wire _330_ ;
        wire _806_ ;
        wire _66_ ;
        wire _615_ ;
        wire _844_ ;
        wire _424_ ;
        wire _653_ ;
        wire _233_ ;
        wire _709_ ;
        wire _462_ ;
        wire _518_ ;
        wire _691_ ;
        wire _271_ ;
        wire _747_ ;
        wire _327_ ;
        wire _556_ ;
        wire _136_ ;
        wire _785_ ;
        wire _365_ ;
        wire _594_ ;
        wire _174_ ;
        wire _459_ ;
        wire _688_ ;
        wire _268_ ;
        wire _497_ ;
        wire _25_ ;
        wire _803_ ;
        wire _63_ ;
        wire _612_ ;
        wire _841_ ;
        wire _421_ ;
        wire _650_ ;
        wire _230_ ;
        wire _706_ ;
        wire _515_ ;
        wire _744_ ;
        wire _324_ ;
        wire _553_ ;
        wire _133_ ;
        wire _609_ ;
        wire _782_ ;
        wire _362_ ;
        wire _838_ ;
        wire _418_ ;
        wire _98_ ;
        wire _591_ ;
        wire _171_ ;
        wire _647_ ;
        wire _227_ ;
        wire _456_ ;
        wire _685_ ;
        wire _265_ ;
        wire _494_ ;
        wire _22_ ;
        wire _779_ ;
        wire _359_ ;
        
        BUFX2 BUFX2_insert58 (
            .A(_201_),
            .Y(_201__bF$buf0)
        );
        
        BUFX2 BUFX2_insert57 (
            .A(_201_),
            .Y(_201__bF$buf1)
        );
        
        BUFX2 BUFX2_insert56 (
            .A(_201_),
            .Y(_201__bF$buf2)
        );
        
        BUFX2 BUFX2_insert55 (
            .A(_201_),
            .Y(_201__bF$buf3)
        );
        
        BUFX2 BUFX2_insert54 (
            .A(_201_),
            .Y(_201__bF$buf4)
        );
        
        BUFX2 BUFX2_insert53 (
            .A(_201_),
            .Y(_201__bF$buf5)
        );
        
        BUFX2 BUFX2_insert52 (
            .A(_201_),
            .Y(_201__bF$buf6)
        );
        
        BUFX2 BUFX2_insert51 (
            .A(Ain12b[11]),
            .Y(Ain12b_11_bF$buf0)
        );
        
        BUFX2 BUFX2_insert50 (
            .A(Ain12b[11]),
            .Y(Ain12b_11_bF$buf1)
        );
        
        BUFX2 BUFX2_insert49 (
            .A(Ain12b[11]),
            .Y(Ain12b_11_bF$buf2)
        );
        
        BUFX2 BUFX2_insert48 (
            .A(Ain12b[11]),
            .Y(Ain12b_11_bF$buf3)
        );
        
        BUFX2 BUFX2_insert47 (
            .A(Ain12b[11]),
            .Y(Ain12b_11_bF$buf4)
        );
        
        BUFX2 BUFX2_insert46 (
            .A(_183_),
            .Y(_183__bF$buf0)
        );
        
        BUFX2 BUFX2_insert45 (
            .A(_183_),
            .Y(_183__bF$buf1)
        );
        
        BUFX2 BUFX2_insert44 (
            .A(_183_),
            .Y(_183__bF$buf2)
        );
        
        BUFX2 BUFX2_insert43 (
            .A(_183_),
            .Y(_183__bF$buf3)
        );
        
        BUFX2 BUFX2_insert42 (
            .A(Stg[1]),
            .Y(Stg_1_bF$buf0)
        );
        
        BUFX2 BUFX2_insert41 (
            .A(Stg[1]),
            .Y(Stg_1_bF$buf1)
        );
        
        BUFX2 BUFX2_insert40 (
            .A(Stg[1]),
            .Y(Stg_1_bF$buf2)
        );
        
        BUFX2 BUFX2_insert39 (
            .A(Stg[1]),
            .Y(Stg_1_bF$buf3)
        );
        
        BUFX2 BUFX2_insert38 (
            .A(LoadCtl[0]),
            .Y(LoadCtl_0_bF$buf0)
        );
        
        BUFX2 BUFX2_insert37 (
            .A(LoadCtl[0]),
            .Y(LoadCtl_0_bF$buf1)
        );
        
        BUFX2 BUFX2_insert36 (
            .A(LoadCtl[0]),
            .Y(LoadCtl_0_bF$buf2)
        );
        
        BUFX2 BUFX2_insert35 (
            .A(LoadCtl[0]),
            .Y(LoadCtl_0_bF$buf3)
        );
        
        BUFX2 BUFX2_insert34 (
            .A(Stg[2]),
            .Y(Stg_2_bF$buf0)
        );
        
        BUFX2 BUFX2_insert33 (
            .A(Stg[2]),
            .Y(Stg_2_bF$buf1)
        );
        
        BUFX2 BUFX2_insert32 (
            .A(Stg[2]),
            .Y(Stg_2_bF$buf2)
        );
        
        BUFX2 BUFX2_insert31 (
            .A(Stg[2]),
            .Y(Stg_2_bF$buf3)
        );
        
        BUFX2 BUFX2_insert30 (
            .A(Stg[2]),
            .Y(Stg_2_bF$buf4)
        );
        
        BUFX2 BUFX2_insert29 (
            .A(LoadCtl[6]),
            .Y(LoadCtl_6_bF$buf0)
        );
        
        BUFX2 BUFX2_insert28 (
            .A(LoadCtl[6]),
            .Y(LoadCtl_6_bF$buf1)
        );
        
        BUFX2 BUFX2_insert27 (
            .A(LoadCtl[6]),
            .Y(LoadCtl_6_bF$buf2)
        );
        
        BUFX2 BUFX2_insert26 (
            .A(LoadCtl[6]),
            .Y(LoadCtl_6_bF$buf3)
        );
        
        BUFX2 BUFX2_insert25 (
            .A(LoadCtl[6]),
            .Y(LoadCtl_6_bF$buf4)
        );
        
        BUFX2 BUFX2_insert24 (
            .A(_164_),
            .Y(_164__bF$buf0)
        );
        
        BUFX2 BUFX2_insert23 (
            .A(_164_),
            .Y(_164__bF$buf1)
        );
        
        BUFX2 BUFX2_insert22 (
            .A(_164_),
            .Y(_164__bF$buf2)
        );
        
        BUFX2 BUFX2_insert21 (
            .A(_164_),
            .Y(_164__bF$buf3)
        );
        
        BUFX2 BUFX2_insert20 (
            .A(_164_),
            .Y(_164__bF$buf4)
        );
        
        CLKBUF1 CLKBUF1_insert19 (
            .A(clk),
            .Y(clk_bF$buf0)
        );
        
        CLKBUF1 CLKBUF1_insert18 (
            .A(clk),
            .Y(clk_bF$buf1)
        );
        
        CLKBUF1 CLKBUF1_insert17 (
            .A(clk),
            .Y(clk_bF$buf2)
        );
        
        CLKBUF1 CLKBUF1_insert16 (
            .A(clk),
            .Y(clk_bF$buf3)
        );
        
        CLKBUF1 CLKBUF1_insert15 (
            .A(clk),
            .Y(clk_bF$buf4)
        );
        
        CLKBUF1 CLKBUF1_insert14 (
            .A(clk),
            .Y(clk_bF$buf5)
        );
        
        CLKBUF1 CLKBUF1_insert13 (
            .A(clk),
            .Y(clk_bF$buf6)
        );
        
        CLKBUF1 CLKBUF1_insert12 (
            .A(clk),
            .Y(clk_bF$buf7)
        );
        
        BUFX2 BUFX2_insert11 (
            .A(_188_),
            .Y(_188__bF$buf0)
        );
        
        BUFX2 BUFX2_insert10 (
            .A(_188_),
            .Y(_188__bF$buf1)
        );
        
        BUFX2 BUFX2_insert9 (
            .A(_188_),
            .Y(_188__bF$buf2)
        );
        
        BUFX2 BUFX2_insert8 (
            .A(_188_),
            .Y(_188__bF$buf3)
        );
        
        BUFX2 BUFX2_insert7 (
            .A(_188_),
            .Y(_188__bF$buf4)
        );
        
        BUFX2 BUFX2_insert6 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf0)
        );
        
        BUFX2 BUFX2_insert5 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf1)
        );
        
        BUFX2 BUFX2_insert4 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf2)
        );
        
        BUFX2 BUFX2_insert3 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf3)
        );
        
        BUFX2 BUFX2_insert2 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf4)
        );
        
        BUFX2 BUFX2_insert1 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf5)
        );
        
        BUFX2 BUFX2_insert0 (
            .A(Stg[0]),
            .Y(Stg_0_bF$buf6)
        );
        
        NAND2X1 _1000_ (
            .A(Stg_0_bF$buf6),
            .B(Yin1[1]),
            .Y(_235_)
        );
        
        OAI21X1 _1001_ (
            .A(Stg_0_bF$buf5),
            .B(_234_),
            .C(_235_),
            .Y(_236_)
        );
        
        NAND2X1 _1002_ (
            .A(Stg_0_bF$buf4),
            .B(Yin0[1]),
            .Y(_237_)
        );
        
        OAI21X1 _1003_ (
            .A(Stg_0_bF$buf3),
            .B(_163_),
            .C(_237_),
            .Y(_238_)
        );
        
        MUX2X1 _1004_ (
            .A(_238_),
            .B(_236_),
            .S(_164__bF$buf4),
            .Y(_239_)
        );
        
        NAND2X1 _1005_ (
            .A(_183__bF$buf3),
            .B(_239_),
            .Y(_240_)
        );
        
        INVX1 _1006_ (
            .A(Yin12b[6]),
            .Y(_241_)
        );
        
        NAND2X1 _1007_ (
            .A(Stg_0_bF$buf2),
            .B(Yin12b[7]),
            .Y(_242_)
        );
        
        OAI21X1 _1008_ (
            .A(Stg_0_bF$buf1),
            .B(_241_),
            .C(_242_),
            .Y(_243_)
        );
        
        INVX1 _1009_ (
            .A(Yin12b[4]),
            .Y(_244_)
        );
        
        NAND2X1 _1010_ (
            .A(Stg_0_bF$buf0),
            .B(Yin12b[5]),
            .Y(_245_)
        );
        
        OAI21X1 _1011_ (
            .A(Stg_0_bF$buf6),
            .B(_244_),
            .C(_245_),
            .Y(_246_)
        );
        
        MUX2X1 _1012_ (
            .A(_246_),
            .B(_243_),
            .S(_164__bF$buf3),
            .Y(_247_)
        );
        
        NAND2X1 _1013_ (
            .A(Stg_2_bF$buf4),
            .B(_247_),
            .Y(_248_)
        );
        
        AND2X2 _1014_ (
            .A(_240_),
            .B(_248_),
            .Y(_249_)
        );
        
        NOR2X1 _1015_ (
            .A(Xin0[0]),
            .B(_249_),
            .Y(_250_)
        );
        
        INVX1 _1016_ (
            .A(_247_),
            .Y(_251_)
        );
        
        OAI21X1 _1017_ (
            .A(_183__bF$buf2),
            .B(_251_),
            .C(_240_),
            .Y(_252_)
        );
        
        OAI21X1 _1018_ (
            .A(_168_),
            .B(_252_),
            .C(_186_),
            .Y(_253_)
        );
        
        OAI21X1 _1019_ (
            .A(_253_),
            .B(_250_),
            .C(_233_),
            .Y(_2_)
        );
        
        NAND2X1 _1020_ (
            .A(Xcalc[1]),
            .B(_188__bF$buf4),
            .Y(_254_)
        );
        
        NOR2X1 _1021_ (
            .A(_168_),
            .B(_252_),
            .Y(_255_)
        );
        
        INVX1 _1022_ (
            .A(Yin1[1]),
            .Y(_256_)
        );
        
        NAND2X1 _1023_ (
            .A(Stg_0_bF$buf5),
            .B(Yin12b[4]),
            .Y(_257_)
        );
        
        OAI21X1 _1024_ (
            .A(Stg_0_bF$buf4),
            .B(_256_),
            .C(_257_),
            .Y(_258_)
        );
        
        NAND2X1 _1025_ (
            .A(Stg_0_bF$buf3),
            .B(Yin1[0]),
            .Y(_259_)
        );
        
        OAI21X1 _1026_ (
            .A(Stg_0_bF$buf2),
            .B(_200_),
            .C(_259_),
            .Y(_260_)
        );
        
        MUX2X1 _1027_ (
            .A(_260_),
            .B(_258_),
            .S(_164__bF$buf2),
            .Y(_261_)
        );
        
        INVX1 _1028_ (
            .A(Yin12b[7]),
            .Y(_262_)
        );
        
        NAND2X1 _1029_ (
            .A(Stg_0_bF$buf1),
            .B(Yin12b[8]),
            .Y(_263_)
        );
        
        OAI21X1 _1030_ (
            .A(Stg_0_bF$buf0),
            .B(_262_),
            .C(_263_),
            .Y(_264_)
        );
        
        INVX1 _1031_ (
            .A(Yin12b[5]),
            .Y(_265_)
        );
        
        NAND2X1 _1032_ (
            .A(Stg_0_bF$buf6),
            .B(Yin12b[6]),
            .Y(_266_)
        );
        
        OAI21X1 _1033_ (
            .A(Stg_0_bF$buf5),
            .B(_265_),
            .C(_266_),
            .Y(_267_)
        );
        
        MUX2X1 _1034_ (
            .A(_267_),
            .B(_264_),
            .S(_164__bF$buf1),
            .Y(_268_)
        );
        
        MUX2X1 _1035_ (
            .A(_268_),
            .B(_261_),
            .S(Stg_2_bF$buf3),
            .Y(_269_)
        );
        
        OAI21X1 _1036_ (
            .A(Ain12b_11_bF$buf4),
            .B(_252_),
            .C(_269_),
            .Y(_270_)
        );
        
        INVX1 _1037_ (
            .A(_269_),
            .Y(_271_)
        );
        
        NAND3X1 _1038_ (
            .A(_201__bF$buf6),
            .B(_271_),
            .C(_249_),
            .Y(_272_)
        );
        
        AOI21X1 _1039_ (
            .A(_270_),
            .B(_272_),
            .C(_205_),
            .Y(_273_)
        );
        
        INVX1 _1040_ (
            .A(_273_),
            .Y(_274_)
        );
        
        NAND3X1 _1041_ (
            .A(_205_),
            .B(_272_),
            .C(_270_),
            .Y(_275_)
        );
        
        NAND3X1 _1042_ (
            .A(_255_),
            .B(_275_),
            .C(_274_),
            .Y(_276_)
        );
        
        INVX1 _1043_ (
            .A(_255_),
            .Y(_277_)
        );
        
        INVX1 _1044_ (
            .A(_275_),
            .Y(_278_)
        );
        
        OAI21X1 _1045_ (
            .A(_273_),
            .B(_278_),
            .C(_277_),
            .Y(_279_)
        );
        
        AOI21X1 _1046_ (
            .A(_279_),
            .B(_276_),
            .C(_192_),
            .Y(_280_)
        );
        
        OAI21X1 _1047_ (
            .A(_188__bF$buf3),
            .B(_280_),
            .C(_254_),
            .Y(_3_)
        );
        
        NAND2X1 _1048_ (
            .A(Xcalc[2]),
            .B(_188__bF$buf2),
            .Y(_281_)
        );
        
        AOI21X1 _1049_ (
            .A(_255_),
            .B(_275_),
            .C(_273_),
            .Y(_282_)
        );
        
        INVX1 _1050_ (
            .A(_282_),
            .Y(_283_)
        );
        
        INVX1 _1051_ (
            .A(Yin12b[9]),
            .Y(_284_)
        );
        
        NAND2X1 _1052_ (
            .A(Stg_0_bF$buf4),
            .B(_284_),
            .Y(_285_)
        );
        
        OAI21X1 _1053_ (
            .A(Stg_0_bF$buf3),
            .B(Yin12b[8]),
            .C(_285_),
            .Y(_286_)
        );
        
        NAND2X1 _1054_ (
            .A(_164__bF$buf0),
            .B(_243_),
            .Y(_287_)
        );
        
        OAI21X1 _1055_ (
            .A(_164__bF$buf4),
            .B(_286_),
            .C(_287_),
            .Y(_288_)
        );
        
        NAND2X1 _1056_ (
            .A(Stg_1_bF$buf3),
            .B(_183__bF$buf1),
            .Y(_289_)
        );
        
        INVX1 _1057_ (
            .A(_289_),
            .Y(_290_)
        );
        
        NAND2X1 _1058_ (
            .A(_246_),
            .B(_290_),
            .Y(_291_)
        );
        
        INVX1 _1059_ (
            .A(_184_),
            .Y(_292_)
        );
        
        NAND2X1 _1060_ (
            .A(_236_),
            .B(_292_),
            .Y(_293_)
        );
        
        NAND2X1 _1061_ (
            .A(_291_),
            .B(_293_),
            .Y(_294_)
        );
        
        AOI21X1 _1062_ (
            .A(_288_),
            .B(Stg_2_bF$buf2),
            .C(_294_),
            .Y(_295_)
        );
        
        OAI21X1 _1063_ (
            .A(_269_),
            .B(_249_),
            .C(_201__bF$buf5),
            .Y(_296_)
        );
        
        OR2X2 _1064_ (
            .A(_296_),
            .B(_295_),
            .Y(_297_)
        );
        
        AOI21X1 _1065_ (
            .A(_240_),
            .B(_248_),
            .C(_269_),
            .Y(_298_)
        );
        
        OAI21X1 _1066_ (
            .A(Ain12b_11_bF$buf3),
            .B(_298_),
            .C(_295_),
            .Y(_299_)
        );
        
        NAND3X1 _1067_ (
            .A(Xin1[0]),
            .B(_299_),
            .C(_297_),
            .Y(_300_)
        );
        
        INVX1 _1068_ (
            .A(_300_),
            .Y(_301_)
        );
        
        AOI21X1 _1069_ (
            .A(_297_),
            .B(_299_),
            .C(Xin1[0]),
            .Y(_302_)
        );
        
        NOR2X1 _1070_ (
            .A(_302_),
            .B(_301_),
            .Y(_303_)
        );
        
        NOR2X1 _1071_ (
            .A(_283_),
            .B(_303_),
            .Y(_304_)
        );
        
        INVX1 _1072_ (
            .A(_303_),
            .Y(_305_)
        );
        
        OAI21X1 _1073_ (
            .A(_282_),
            .B(_305_),
            .C(_186_),
            .Y(_306_)
        );
        
        OAI21X1 _1074_ (
            .A(_304_),
            .B(_306_),
            .C(_281_),
            .Y(_4_)
        );
        
        NAND2X1 _1075_ (
            .A(Xcalc[3]),
            .B(_188__bF$buf1),
            .Y(_307_)
        );
        
        OAI21X1 _1076_ (
            .A(_282_),
            .B(_302_),
            .C(_300_),
            .Y(_308_)
        );
        
        INVX1 _1077_ (
            .A(_308_),
            .Y(_309_)
        );
        
        NAND2X1 _1078_ (
            .A(_295_),
            .B(_298_),
            .Y(_310_)
        );
        
        INVX1 _1079_ (
            .A(Yin12b[10]),
            .Y(_311_)
        );
        
        NAND2X1 _1080_ (
            .A(Stg_0_bF$buf2),
            .B(_311_),
            .Y(_312_)
        );
        
        OAI21X1 _1081_ (
            .A(Stg_0_bF$buf1),
            .B(Yin12b[9]),
            .C(_312_),
            .Y(_313_)
        );
        
        NAND2X1 _1082_ (
            .A(_164__bF$buf3),
            .B(_264_),
            .Y(_314_)
        );
        
        OAI21X1 _1083_ (
            .A(_164__bF$buf2),
            .B(_313_),
            .C(_314_),
            .Y(_315_)
        );
        
        NAND2X1 _1084_ (
            .A(_267_),
            .B(_290_),
            .Y(_316_)
        );
        
        NAND2X1 _1085_ (
            .A(_258_),
            .B(_292_),
            .Y(_317_)
        );
        
        NAND2X1 _1086_ (
            .A(_316_),
            .B(_317_),
            .Y(_318_)
        );
        
        AOI21X1 _1087_ (
            .A(_315_),
            .B(Stg_2_bF$buf1),
            .C(_318_),
            .Y(_319_)
        );
        
        NAND3X1 _1088_ (
            .A(_201__bF$buf4),
            .B(_319_),
            .C(_310_),
            .Y(_320_)
        );
        
        INVX1 _1089_ (
            .A(_310_),
            .Y(_321_)
        );
        
        INVX1 _1090_ (
            .A(_319_),
            .Y(_322_)
        );
        
        OAI21X1 _1091_ (
            .A(Ain12b_11_bF$buf2),
            .B(_321_),
            .C(_322_),
            .Y(_323_)
        );
        
        AOI21X1 _1092_ (
            .A(_323_),
            .B(_320_),
            .C(_202_),
            .Y(_324_)
        );
        
        INVX1 _1093_ (
            .A(_324_),
            .Y(_325_)
        );
        
        NAND3X1 _1094_ (
            .A(_202_),
            .B(_320_),
            .C(_323_),
            .Y(_326_)
        );
        
        NAND2X1 _1095_ (
            .A(_326_),
            .B(_325_),
            .Y(_327_)
        );
        
        OR2X2 _1096_ (
            .A(_327_),
            .B(_309_),
            .Y(_328_)
        );
        
        NAND2X1 _1097_ (
            .A(_309_),
            .B(_327_),
            .Y(_329_)
        );
        
        AOI21X1 _1098_ (
            .A(_328_),
            .B(_329_),
            .C(_192_),
            .Y(_330_)
        );
        
        OAI21X1 _1099_ (
            .A(_188__bF$buf0),
            .B(_330_),
            .C(_307_),
            .Y(_5_)
        );
        
        AOI21X1 _1100_ (
            .A(_308_),
            .B(_326_),
            .C(_324_),
            .Y(_331_)
        );
        
        NAND3X1 _1101_ (
            .A(_295_),
            .B(_319_),
            .C(_298_),
            .Y(_332_)
        );
        
        NAND2X1 _1102_ (
            .A(Stg_0_bF$buf0),
            .B(Yin12b[11]),
            .Y(_333_)
        );
        
        OAI21X1 _1103_ (
            .A(Stg_0_bF$buf6),
            .B(_311_),
            .C(_333_),
            .Y(_334_)
        );
        
        NAND2X1 _1104_ (
            .A(Stg_1_bF$buf2),
            .B(_334_),
            .Y(_335_)
        );
        
        OAI21X1 _1105_ (
            .A(Stg_1_bF$buf1),
            .B(_286_),
            .C(_335_),
            .Y(_336_)
        );
        
        NAND2X1 _1106_ (
            .A(Stg_2_bF$buf0),
            .B(_336_),
            .Y(_337_)
        );
        
        OAI21X1 _1107_ (
            .A(Stg_2_bF$buf4),
            .B(_247_),
            .C(_337_),
            .Y(_338_)
        );
        
        INVX1 _1108_ (
            .A(_338_),
            .Y(_339_)
        );
        
        NAND3X1 _1109_ (
            .A(_201__bF$buf3),
            .B(_339_),
            .C(_332_),
            .Y(_340_)
        );
        
        INVX1 _1110_ (
            .A(_340_),
            .Y(_341_)
        );
        
        AOI21X1 _1111_ (
            .A(_332_),
            .B(_201__bF$buf2),
            .C(_339_),
            .Y(_342_)
        );
        
        OAI21X1 _1112_ (
            .A(_342_),
            .B(_341_),
            .C(Xin12b[4]),
            .Y(_343_)
        );
        
        OAI21X1 _1113_ (
            .A(_322_),
            .B(_310_),
            .C(_201__bF$buf1),
            .Y(_344_)
        );
        
        NAND2X1 _1114_ (
            .A(_338_),
            .B(_344_),
            .Y(_345_)
        );
        
        NAND3X1 _1115_ (
            .A(_175_),
            .B(_340_),
            .C(_345_),
            .Y(_346_)
        );
        
        AND2X2 _1116_ (
            .A(_343_),
            .B(_346_),
            .Y(_347_)
        );
        
        INVX1 _1117_ (
            .A(_347_),
            .Y(_348_)
        );
        
        OR2X2 _1118_ (
            .A(_331_),
            .B(_348_),
            .Y(_349_)
        );
        
        NAND2X1 _1119_ (
            .A(_348_),
            .B(_331_),
            .Y(_350_)
        );
        
        NAND2X1 _1120_ (
            .A(_350_),
            .B(_349_),
            .Y(_351_)
        );
        
        AOI22X1 _1121_ (
            .A(_150_),
            .B(_188__bF$buf4),
            .C(_351_),
            .D(_186_),
            .Y(_6_)
        );
        
        OAI21X1 _1122_ (
            .A(_348_),
            .B(_331_),
            .C(_343_),
            .Y(_352_)
        );
        
        NOR2X1 _1123_ (
            .A(_338_),
            .B(_332_),
            .Y(_353_)
        );
        
        INVX1 _1124_ (
            .A(_353_),
            .Y(_354_)
        );
        
        NOR2X1 _1125_ (
            .A(Stg_1_bF$buf0),
            .B(_313_),
            .Y(_355_)
        );
        
        INVX1 _1126_ (
            .A(Yin12b[11]),
            .Y(_356_)
        );
        
        NOR2X1 _1127_ (
            .A(_164__bF$buf1),
            .B(_356_),
            .Y(_357_)
        );
        
        OAI21X1 _1128_ (
            .A(_357_),
            .B(_355_),
            .C(Stg_2_bF$buf3),
            .Y(_358_)
        );
        
        OAI21X1 _1129_ (
            .A(Stg_2_bF$buf2),
            .B(_268_),
            .C(_358_),
            .Y(_359_)
        );
        
        NAND3X1 _1130_ (
            .A(_201__bF$buf0),
            .B(_359_),
            .C(_354_),
            .Y(_360_)
        );
        
        INVX1 _1131_ (
            .A(_359_),
            .Y(_361_)
        );
        
        OAI21X1 _1132_ (
            .A(Ain12b_11_bF$buf1),
            .B(_353_),
            .C(_361_),
            .Y(_362_)
        );
        
        NAND3X1 _1133_ (
            .A(Xin12b[5]),
            .B(_362_),
            .C(_360_),
            .Y(_363_)
        );
        
        NAND3X1 _1134_ (
            .A(_201__bF$buf6),
            .B(_361_),
            .C(_354_),
            .Y(_364_)
        );
        
        OAI21X1 _1135_ (
            .A(Ain12b_11_bF$buf0),
            .B(_353_),
            .C(_359_),
            .Y(_365_)
        );
        
        NAND3X1 _1136_ (
            .A(_212_),
            .B(_365_),
            .C(_364_),
            .Y(_366_)
        );
        
        NAND2X1 _1137_ (
            .A(_363_),
            .B(_366_),
            .Y(_367_)
        );
        
        INVX1 _1138_ (
            .A(_367_),
            .Y(_368_)
        );
        
        AND2X2 _1139_ (
            .A(_352_),
            .B(_368_),
            .Y(_369_)
        );
        
        OAI21X1 _1140_ (
            .A(_368_),
            .B(_352_),
            .C(_186_),
            .Y(_370_)
        );
        
        OAI22X1 _1141_ (
            .A(_158_),
            .B(LoadCtl_6_bF$buf4),
            .C(_370_),
            .D(_369_),
            .Y(_7_)
        );
        
        NOR3X1 _1142_ (
            .A(_338_),
            .B(_359_),
            .C(_332_),
            .Y(_371_)
        );
        
        INVX1 _1143_ (
            .A(_371_),
            .Y(_372_)
        );
        
        AOI21X1 _1144_ (
            .A(_164__bF$buf0),
            .B(_334_),
            .C(_357_),
            .Y(_373_)
        );
        
        NAND2X1 _1145_ (
            .A(_183__bF$buf0),
            .B(_288_),
            .Y(_374_)
        );
        
        OAI21X1 _1146_ (
            .A(_183__bF$buf3),
            .B(_373_),
            .C(_374_),
            .Y(_375_)
        );
        
        INVX1 _1147_ (
            .A(_375_),
            .Y(_376_)
        );
        
        NAND3X1 _1148_ (
            .A(_201__bF$buf5),
            .B(_376_),
            .C(_372_),
            .Y(_377_)
        );
        
        OAI21X1 _1149_ (
            .A(Ain12b_11_bF$buf4),
            .B(_371_),
            .C(_375_),
            .Y(_378_)
        );
        
        NAND2X1 _1150_ (
            .A(_378_),
            .B(_377_),
            .Y(_379_)
        );
        
        NAND2X1 _1151_ (
            .A(Xin12b[6]),
            .B(_379_),
            .Y(_380_)
        );
        
        NAND3X1 _1152_ (
            .A(_172_),
            .B(_378_),
            .C(_377_),
            .Y(_381_)
        );
        
        AND2X2 _1153_ (
            .A(_380_),
            .B(_381_),
            .Y(_382_)
        );
        
        NAND3X1 _1154_ (
            .A(_363_),
            .B(_366_),
            .C(_347_),
            .Y(_383_)
        );
        
        INVX1 _1155_ (
            .A(_343_),
            .Y(_384_)
        );
        
        AOI21X1 _1156_ (
            .A(_364_),
            .B(_365_),
            .C(_212_),
            .Y(_385_)
        );
        
        AOI21X1 _1157_ (
            .A(_384_),
            .B(_366_),
            .C(_385_),
            .Y(_386_)
        );
        
        OAI21X1 _1158_ (
            .A(_331_),
            .B(_383_),
            .C(_386_),
            .Y(_387_)
        );
        
        AND2X2 _1159_ (
            .A(_387_),
            .B(_382_),
            .Y(_388_)
        );
        
        NOR2X1 _1160_ (
            .A(_382_),
            .B(_387_),
            .Y(_389_)
        );
        
        OAI21X1 _1161_ (
            .A(_389_),
            .B(_388_),
            .C(_191_),
            .Y(_390_)
        );
        
        NAND2X1 _1162_ (
            .A(LoadCtl_6_bF$buf3),
            .B(_390_),
            .Y(_391_)
        );
        
        OAI21X1 _1163_ (
            .A(_149_),
            .B(LoadCtl_6_bF$buf2),
            .C(_391_),
            .Y(_8_)
        );
        
        AOI21X1 _1164_ (
            .A(_377_),
            .B(_378_),
            .C(_172_),
            .Y(_392_)
        );
        
        NOR2X1 _1165_ (
            .A(_392_),
            .B(_388_),
            .Y(_393_)
        );
        
        NAND3X1 _1166_ (
            .A(_361_),
            .B(_376_),
            .C(_353_),
            .Y(_394_)
        );
        
        NOR2X1 _1167_ (
            .A(_183__bF$buf2),
            .B(_356_),
            .Y(_395_)
        );
        
        AOI21X1 _1168_ (
            .A(_315_),
            .B(_183__bF$buf1),
            .C(_395_),
            .Y(_396_)
        );
        
        NAND3X1 _1169_ (
            .A(_201__bF$buf4),
            .B(_396_),
            .C(_394_),
            .Y(_397_)
        );
        
        INVX1 _1170_ (
            .A(_397_),
            .Y(_398_)
        );
        
        AOI21X1 _1171_ (
            .A(_394_),
            .B(_201__bF$buf3),
            .C(_396_),
            .Y(_399_)
        );
        
        OAI21X1 _1172_ (
            .A(_399_),
            .B(_398_),
            .C(Xin12b[7]),
            .Y(_400_)
        );
        
        INVX1 _1173_ (
            .A(_396_),
            .Y(_401_)
        );
        
        NAND2X1 _1174_ (
            .A(_201__bF$buf2),
            .B(_394_),
            .Y(_402_)
        );
        
        NAND2X1 _1175_ (
            .A(_401_),
            .B(_402_),
            .Y(_403_)
        );
        
        NAND3X1 _1176_ (
            .A(_209_),
            .B(_397_),
            .C(_403_),
            .Y(_404_)
        );
        
        AND2X2 _1177_ (
            .A(_400_),
            .B(_404_),
            .Y(_405_)
        );
        
        OR2X2 _1178_ (
            .A(_393_),
            .B(_405_),
            .Y(_406_)
        );
        
        AOI21X1 _1179_ (
            .A(_393_),
            .B(_405_),
            .C(_185_),
            .Y(_407_)
        );
        
        AOI22X1 _1180_ (
            .A(_157_),
            .B(_188__bF$buf3),
            .C(_406_),
            .D(_407_),
            .Y(_9_)
        );
        
        NAND2X1 _1181_ (
            .A(Xcalc[8]),
            .B(_188__bF$buf2),
            .Y(_408_)
        );
        
        NAND2X1 _1182_ (
            .A(_392_),
            .B(_404_),
            .Y(_409_)
        );
        
        AND2X2 _1183_ (
            .A(_409_),
            .B(_400_),
            .Y(_410_)
        );
        
        NAND3X1 _1184_ (
            .A(_382_),
            .B(_387_),
            .C(_405_),
            .Y(_411_)
        );
        
        NAND2X1 _1185_ (
            .A(_410_),
            .B(_411_),
            .Y(_412_)
        );
        
        NAND3X1 _1186_ (
            .A(_376_),
            .B(_396_),
            .C(_371_),
            .Y(_413_)
        );
        
        INVX1 _1187_ (
            .A(_336_),
            .Y(_414_)
        );
        
        INVX1 _1188_ (
            .A(_395_),
            .Y(_415_)
        );
        
        OAI21X1 _1189_ (
            .A(Stg_2_bF$buf1),
            .B(_414_),
            .C(_415_),
            .Y(_416_)
        );
        
        NAND3X1 _1190_ (
            .A(_201__bF$buf1),
            .B(_416_),
            .C(_413_),
            .Y(_417_)
        );
        
        INVX1 _1191_ (
            .A(_416_),
            .Y(_418_)
        );
        
        OAI21X1 _1192_ (
            .A(_401_),
            .B(_394_),
            .C(_201__bF$buf0),
            .Y(_419_)
        );
        
        NAND2X1 _1193_ (
            .A(_418_),
            .B(_419_),
            .Y(_420_)
        );
        
        NAND3X1 _1194_ (
            .A(Xin12b[8]),
            .B(_417_),
            .C(_420_),
            .Y(_421_)
        );
        
        INVX1 _1195_ (
            .A(Xin12b[8]),
            .Y(_422_)
        );
        
        NAND3X1 _1196_ (
            .A(_201__bF$buf6),
            .B(_418_),
            .C(_413_),
            .Y(_423_)
        );
        
        NAND2X1 _1197_ (
            .A(_416_),
            .B(_419_),
            .Y(_424_)
        );
        
        NAND3X1 _1198_ (
            .A(_422_),
            .B(_423_),
            .C(_424_),
            .Y(_425_)
        );
        
        AND2X2 _1199_ (
            .A(_421_),
            .B(_425_),
            .Y(_426_)
        );
        
        OR2X2 _1200_ (
            .A(_412_),
            .B(_426_),
            .Y(_427_)
        );
        
        INVX1 _1201_ (
            .A(_427_),
            .Y(_428_)
        );
        
        INVX1 _1202_ (
            .A(_426_),
            .Y(_429_)
        );
        
        AOI21X1 _1203_ (
            .A(_411_),
            .B(_410_),
            .C(_429_),
            .Y(_430_)
        );
        
        INVX1 _1204_ (
            .A(_430_),
            .Y(_431_)
        );
        
        NAND2X1 _1205_ (
            .A(_186_),
            .B(_431_),
            .Y(_432_)
        );
        
        OAI21X1 _1206_ (
            .A(_432_),
            .B(_428_),
            .C(_408_),
            .Y(_10_)
        );
        
        INVX1 _1207_ (
            .A(Xcalc[9]),
            .Y(_433_)
        );
        
        INVX1 _1208_ (
            .A(_421_),
            .Y(_434_)
        );
        
        OR2X2 _1209_ (
            .A(_355_),
            .B(_357_),
            .Y(_435_)
        );
        
        AOI21X1 _1210_ (
            .A(_435_),
            .B(_183__bF$buf0),
            .C(_395_),
            .Y(_436_)
        );
        
        OAI21X1 _1211_ (
            .A(_416_),
            .B(_413_),
            .C(_201__bF$buf5),
            .Y(_437_)
        );
        
        NAND2X1 _1212_ (
            .A(_436_),
            .B(_437_),
            .Y(_438_)
        );
        
        OR2X2 _1213_ (
            .A(_437_),
            .B(_436_),
            .Y(_439_)
        );
        
        NAND3X1 _1214_ (
            .A(Xin12b[9]),
            .B(_438_),
            .C(_439_),
            .Y(_440_)
        );
        
        INVX1 _1215_ (
            .A(Xin12b[9]),
            .Y(_441_)
        );
        
        AND2X2 _1216_ (
            .A(_437_),
            .B(_436_),
            .Y(_442_)
        );
        
        NOR2X1 _1217_ (
            .A(_436_),
            .B(_437_),
            .Y(_443_)
        );
        
        OAI21X1 _1218_ (
            .A(_443_),
            .B(_442_),
            .C(_441_),
            .Y(_444_)
        );
        
        NAND2X1 _1219_ (
            .A(_444_),
            .B(_440_),
            .Y(_445_)
        );
        
        NOR3X1 _1220_ (
            .A(_434_),
            .B(_445_),
            .C(_430_),
            .Y(_446_)
        );
        
        AOI22X1 _1221_ (
            .A(_440_),
            .B(_444_),
            .C(_431_),
            .D(_421_),
            .Y(_447_)
        );
        
        OAI21X1 _1222_ (
            .A(_446_),
            .B(_447_),
            .C(_186_),
            .Y(_448_)
        );
        
        OAI21X1 _1223_ (
            .A(_433_),
            .B(LoadCtl_6_bF$buf1),
            .C(_448_),
            .Y(_11_)
        );
        
        OAI21X1 _1224_ (
            .A(Stg_2_bF$buf0),
            .B(_373_),
            .C(_415_),
            .Y(_449_)
        );
        
        OR2X2 _1225_ (
            .A(_413_),
            .B(_416_),
            .Y(_450_)
        );
        
        INVX1 _1226_ (
            .A(_436_),
            .Y(_451_)
        );
        
        OAI21X1 _1227_ (
            .A(_451_),
            .B(_450_),
            .C(_201__bF$buf4),
            .Y(_452_)
        );
        
        NOR2X1 _1228_ (
            .A(_449_),
            .B(_452_),
            .Y(_453_)
        );
        
        INVX1 _1229_ (
            .A(_449_),
            .Y(_454_)
        );
        
        OAI21X1 _1230_ (
            .A(Ain12b_11_bF$buf3),
            .B(_436_),
            .C(_437_),
            .Y(_455_)
        );
        
        NOR2X1 _1231_ (
            .A(_454_),
            .B(_455_),
            .Y(_456_)
        );
        
        OAI21X1 _1232_ (
            .A(_456_),
            .B(_453_),
            .C(Xin12b[10]),
            .Y(_457_)
        );
        
        INVX1 _1233_ (
            .A(Xin12b[10]),
            .Y(_458_)
        );
        
        NOR2X1 _1234_ (
            .A(_449_),
            .B(_455_),
            .Y(_459_)
        );
        
        NOR2X1 _1235_ (
            .A(_454_),
            .B(_452_),
            .Y(_460_)
        );
        
        OAI21X1 _1236_ (
            .A(_459_),
            .B(_460_),
            .C(_458_),
            .Y(_461_)
        );
        
        AND2X2 _1237_ (
            .A(_457_),
            .B(_461_),
            .Y(_462_)
        );
        
        OAI21X1 _1238_ (
            .A(_421_),
            .B(_445_),
            .C(_440_),
            .Y(_463_)
        );
        
        NAND3X1 _1239_ (
            .A(_440_),
            .B(_444_),
            .C(_426_),
            .Y(_464_)
        );
        
        AOI21X1 _1240_ (
            .A(_410_),
            .B(_411_),
            .C(_464_),
            .Y(_465_)
        );
        
        OAI21X1 _1241_ (
            .A(_463_),
            .B(_465_),
            .C(_462_),
            .Y(_466_)
        );
        
        INVX1 _1242_ (
            .A(_462_),
            .Y(_467_)
        );
        
        NOR2X1 _1243_ (
            .A(_463_),
            .B(_465_),
            .Y(_468_)
        );
        
        NAND2X1 _1244_ (
            .A(_467_),
            .B(_468_),
            .Y(_469_)
        );
        
        NAND2X1 _1245_ (
            .A(_466_),
            .B(_469_),
            .Y(_470_)
        );
        
        AOI22X1 _1246_ (
            .A(_146_),
            .B(_188__bF$buf1),
            .C(_470_),
            .D(_186_),
            .Y(_12_)
        );
        
        INVX1 _1247_ (
            .A(Xin12b[11]),
            .Y(_471_)
        );
        
        NAND2X1 _1248_ (
            .A(Yin12b[11]),
            .B(_471_),
            .Y(_472_)
        );
        
        NAND2X1 _1249_ (
            .A(Xin12b[11]),
            .B(_356_),
            .Y(_473_)
        );
        
        NAND2X1 _1250_ (
            .A(_472_),
            .B(_473_),
            .Y(_474_)
        );
        
        INVX1 _1251_ (
            .A(_474_),
            .Y(_475_)
        );
        
        OAI21X1 _1252_ (
            .A(Ain12b_11_bF$buf2),
            .B(_459_),
            .C(_475_),
            .Y(_476_)
        );
        
        NOR2X1 _1253_ (
            .A(Ain12b_11_bF$buf1),
            .B(_454_),
            .Y(_477_)
        );
        
        OAI21X1 _1254_ (
            .A(_477_),
            .B(_455_),
            .C(_474_),
            .Y(_478_)
        );
        
        NAND2X1 _1255_ (
            .A(_478_),
            .B(_476_),
            .Y(_479_)
        );
        
        AOI21X1 _1256_ (
            .A(_466_),
            .B(_457_),
            .C(_479_),
            .Y(_480_)
        );
        
        NAND3X1 _1257_ (
            .A(_457_),
            .B(_479_),
            .C(_466_),
            .Y(_481_)
        );
        
        NAND2X1 _1258_ (
            .A(_186_),
            .B(_481_),
            .Y(_482_)
        );
        
        OAI22X1 _1259_ (
            .A(_154_),
            .B(LoadCtl_6_bF$buf0),
            .C(_480_),
            .D(_482_),
            .Y(_13_)
        );
        
        INVX1 _1260_ (
            .A(Ain0[0]),
            .Y(_483_)
        );
        
        INVX1 _1261_ (
            .A(_190_),
            .Y(_484_)
        );
        
        NAND2X1 _1262_ (
            .A(Stg_0_bF$buf5),
            .B(Stg_1_bF$buf3),
            .Y(_485_)
        );
        
        OAI21X1 _1263_ (
            .A(_183__bF$buf3),
            .B(_484_),
            .C(_485_),
            .Y(_486_)
        );
        
        NOR2X1 _1264_ (
            .A(_483_),
            .B(_486_),
            .Y(_487_)
        );
        
        AND2X2 _1265_ (
            .A(_486_),
            .B(_483_),
            .Y(_488_)
        );
        
        OR2X2 _1266_ (
            .A(_488_),
            .B(_487_),
            .Y(_489_)
        );
        
        NAND2X1 _1267_ (
            .A(Acalc[0]),
            .B(_188__bF$buf0),
            .Y(_490_)
        );
        
        OAI21X1 _1268_ (
            .A(_188__bF$buf4),
            .B(_489_),
            .C(_490_),
            .Y(_14_)
        );
        
        NAND2X1 _1269_ (
            .A(Acalc[1]),
            .B(_188__bF$buf3),
            .Y(_491_)
        );
        
        INVX2 _1270_ (
            .A(Stg_0_bF$buf4),
            .Y(_492_)
        );
        
        OAI21X1 _1271_ (
            .A(Stg_1_bF$buf2),
            .B(_492_),
            .C(Stg_2_bF$buf4),
            .Y(_493_)
        );
        
        OAI21X1 _1272_ (
            .A(Stg_2_bF$buf3),
            .B(_492_),
            .C(_493_),
            .Y(_494_)
        );
        
        OAI21X1 _1273_ (
            .A(Ain12b_11_bF$buf0),
            .B(_486_),
            .C(_494_),
            .Y(_495_)
        );
        
        OAI21X1 _1274_ (
            .A(Ain12b_11_bF$buf4),
            .B(_494_),
            .C(_495_),
            .Y(_496_)
        );
        
        OR2X2 _1275_ (
            .A(_496_),
            .B(Ain0[1]),
            .Y(_497_)
        );
        
        NAND2X1 _1276_ (
            .A(Ain0[1]),
            .B(_496_),
            .Y(_498_)
        );
        
        NAND2X1 _1277_ (
            .A(_498_),
            .B(_497_),
            .Y(_499_)
        );
        
        NOR2X1 _1278_ (
            .A(_487_),
            .B(_499_),
            .Y(_500_)
        );
        
        NAND2X1 _1279_ (
            .A(_487_),
            .B(_499_),
            .Y(_501_)
        );
        
        NAND2X1 _1280_ (
            .A(LoadCtl_6_bF$buf4),
            .B(_501_),
            .Y(_502_)
        );
        
        OAI21X1 _1281_ (
            .A(_500_),
            .B(_502_),
            .C(_491_),
            .Y(_15_)
        );
        
        NAND2X1 _1282_ (
            .A(Acalc[2]),
            .B(_188__bF$buf2),
            .Y(_503_)
        );
        
        INVX1 _1283_ (
            .A(Ain0[1]),
            .Y(_504_)
        );
        
        OAI21X1 _1284_ (
            .A(_504_),
            .B(_496_),
            .C(_501_),
            .Y(_505_)
        );
        
        OAI21X1 _1285_ (
            .A(_492_),
            .B(_164__bF$buf4),
            .C(Ain12b_11_bF$buf3),
            .Y(_506_)
        );
        
        NAND3X1 _1286_ (
            .A(Stg_2_bF$buf2),
            .B(_484_),
            .C(_506_),
            .Y(_507_)
        );
        
        OAI21X1 _1287_ (
            .A(Stg_2_bF$buf1),
            .B(_506_),
            .C(_507_),
            .Y(_508_)
        );
        
        NAND2X1 _1288_ (
            .A(Ain1[0]),
            .B(_508_),
            .Y(_509_)
        );
        
        OR2X2 _1289_ (
            .A(_508_),
            .B(Ain1[0]),
            .Y(_510_)
        );
        
        NAND2X1 _1290_ (
            .A(_509_),
            .B(_510_),
            .Y(_511_)
        );
        
        INVX1 _1291_ (
            .A(_511_),
            .Y(_512_)
        );
        
        NOR2X1 _1292_ (
            .A(_512_),
            .B(_505_),
            .Y(_513_)
        );
        
        NAND2X1 _1293_ (
            .A(_512_),
            .B(_505_),
            .Y(_514_)
        );
        
        NAND2X1 _1294_ (
            .A(LoadCtl_6_bF$buf3),
            .B(_514_),
            .Y(_515_)
        );
        
        OAI21X1 _1295_ (
            .A(_513_),
            .B(_515_),
            .C(_503_),
            .Y(_16_)
        );
        
        NAND2X1 _1296_ (
            .A(_509_),
            .B(_514_),
            .Y(_516_)
        );
        
        INVX1 _1297_ (
            .A(_516_),
            .Y(_517_)
        );
        
        INVX1 _1298_ (
            .A(Ain1[1]),
            .Y(_518_)
        );
        
        OAI21X1 _1299_ (
            .A(Stg_0_bF$buf3),
            .B(_164__bF$buf3),
            .C(Stg_2_bF$buf0),
            .Y(_519_)
        );
        
        NAND2X1 _1300_ (
            .A(_201__bF$buf3),
            .B(_519_),
            .Y(_520_)
        );
        
        OAI21X1 _1301_ (
            .A(Stg_2_bF$buf4),
            .B(Stg_1_bF$buf1),
            .C(Ain12b_11_bF$buf2),
            .Y(_521_)
        );
        
        OAI21X1 _1302_ (
            .A(_492_),
            .B(_521_),
            .C(_520_),
            .Y(_522_)
        );
        
        NOR2X1 _1303_ (
            .A(_518_),
            .B(_522_),
            .Y(_523_)
        );
        
        NAND2X1 _1304_ (
            .A(_518_),
            .B(_522_),
            .Y(_524_)
        );
        
        INVX1 _1305_ (
            .A(_524_),
            .Y(_525_)
        );
        
        OAI21X1 _1306_ (
            .A(_523_),
            .B(_525_),
            .C(_517_),
            .Y(_526_)
        );
        
        INVX1 _1307_ (
            .A(_523_),
            .Y(_527_)
        );
        
        NAND3X1 _1308_ (
            .A(_527_),
            .B(_524_),
            .C(_516_),
            .Y(_528_)
        );
        
        NAND2X1 _1309_ (
            .A(_528_),
            .B(_526_),
            .Y(_529_)
        );
        
        NAND2X1 _1310_ (
            .A(Acalc[3]),
            .B(_188__bF$buf1),
            .Y(_530_)
        );
        
        OAI21X1 _1311_ (
            .A(_188__bF$buf0),
            .B(_529_),
            .C(_530_),
            .Y(_17_)
        );
        
        NAND2X1 _1312_ (
            .A(Acalc[4]),
            .B(_188__bF$buf4),
            .Y(_531_)
        );
        
        NOR2X1 _1313_ (
            .A(Ain12b_11_bF$buf1),
            .B(_494_),
            .Y(_532_)
        );
        
        NAND3X1 _1314_ (
            .A(Stg_0_bF$buf2),
            .B(_183__bF$buf2),
            .C(_164__bF$buf2),
            .Y(_533_)
        );
        
        AOI21X1 _1315_ (
            .A(_493_),
            .B(_533_),
            .C(_201__bF$buf2),
            .Y(_534_)
        );
        
        NOR2X1 _1316_ (
            .A(_534_),
            .B(_532_),
            .Y(_535_)
        );
        
        NAND2X1 _1317_ (
            .A(Ain12b[4]),
            .B(_535_),
            .Y(_536_)
        );
        
        INVX1 _1318_ (
            .A(Ain12b[4]),
            .Y(_537_)
        );
        
        OAI21X1 _1319_ (
            .A(_534_),
            .B(_532_),
            .C(_537_),
            .Y(_538_)
        );
        
        OAI21X1 _1320_ (
            .A(_525_),
            .B(_517_),
            .C(_527_),
            .Y(_539_)
        );
        
        AOI21X1 _1321_ (
            .A(_536_),
            .B(_538_),
            .C(_539_),
            .Y(_540_)
        );
        
        NAND2X1 _1322_ (
            .A(_538_),
            .B(_536_),
            .Y(_541_)
        );
        
        INVX1 _1323_ (
            .A(_539_),
            .Y(_542_)
        );
        
        OAI21X1 _1324_ (
            .A(_541_),
            .B(_542_),
            .C(LoadCtl_6_bF$buf2),
            .Y(_543_)
        );
        
        OAI21X1 _1325_ (
            .A(_540_),
            .B(_543_),
            .C(_531_),
            .Y(_18_)
        );
        
        NAND2X1 _1326_ (
            .A(Acalc[5]),
            .B(_188__bF$buf3),
            .Y(_544_)
        );
        
        OAI21X1 _1327_ (
            .A(_541_),
            .B(_542_),
            .C(_536_),
            .Y(_545_)
        );
        
        OAI21X1 _1328_ (
            .A(_190_),
            .B(_292_),
            .C(_201__bF$buf1),
            .Y(_546_)
        );
        
        INVX1 _1329_ (
            .A(_546_),
            .Y(_547_)
        );
        
        OAI21X1 _1330_ (
            .A(Stg_0_bF$buf1),
            .B(Stg_1_bF$buf0),
            .C(_184_),
            .Y(_548_)
        );
        
        NOR2X1 _1331_ (
            .A(_201__bF$buf0),
            .B(_548_),
            .Y(_549_)
        );
        
        NOR2X1 _1332_ (
            .A(_549_),
            .B(_547_),
            .Y(_550_)
        );
        
        AND2X2 _1333_ (
            .A(_550_),
            .B(Ain12b[5]),
            .Y(_551_)
        );
        
        INVX1 _1334_ (
            .A(_551_),
            .Y(_552_)
        );
        
        INVX1 _1335_ (
            .A(Ain12b[5]),
            .Y(_553_)
        );
        
        OAI21X1 _1336_ (
            .A(_549_),
            .B(_547_),
            .C(_553_),
            .Y(_554_)
        );
        
        NAND2X1 _1337_ (
            .A(_554_),
            .B(_552_),
            .Y(_555_)
        );
        
        INVX1 _1338_ (
            .A(_555_),
            .Y(_556_)
        );
        
        NOR2X1 _1339_ (
            .A(_556_),
            .B(_545_),
            .Y(_557_)
        );
        
        NAND2X1 _1340_ (
            .A(_556_),
            .B(_545_),
            .Y(_558_)
        );
        
        NAND2X1 _1341_ (
            .A(LoadCtl_6_bF$buf1),
            .B(_558_),
            .Y(_559_)
        );
        
        OAI21X1 _1342_ (
            .A(_557_),
            .B(_559_),
            .C(_544_),
            .Y(_19_)
        );
        
        NOR2X1 _1343_ (
            .A(_541_),
            .B(_555_),
            .Y(_560_)
        );
        
        OAI21X1 _1344_ (
            .A(_536_),
            .B(_555_),
            .C(_552_),
            .Y(_561_)
        );
        
        AOI21X1 _1345_ (
            .A(_539_),
            .B(_560_),
            .C(_561_),
            .Y(_562_)
        );
        
        OAI21X1 _1346_ (
            .A(Stg_2_bF$buf3),
            .B(_485_),
            .C(_191_),
            .Y(_563_)
        );
        
        NOR2X1 _1347_ (
            .A(_201__bF$buf6),
            .B(_563_),
            .Y(_564_)
        );
        
        AND2X2 _1348_ (
            .A(_563_),
            .B(_201__bF$buf5),
            .Y(_565_)
        );
        
        NOR2X1 _1349_ (
            .A(_564_),
            .B(_565_),
            .Y(_566_)
        );
        
        NAND2X1 _1350_ (
            .A(Ain12b[6]),
            .B(_566_),
            .Y(_567_)
        );
        
        INVX1 _1351_ (
            .A(Ain12b[6]),
            .Y(_568_)
        );
        
        OAI21X1 _1352_ (
            .A(_564_),
            .B(_565_),
            .C(_568_),
            .Y(_569_)
        );
        
        NAND2X1 _1353_ (
            .A(_569_),
            .B(_567_),
            .Y(_570_)
        );
        
        AND2X2 _1354_ (
            .A(_562_),
            .B(_570_),
            .Y(_571_)
        );
        
        OAI21X1 _1355_ (
            .A(_570_),
            .B(_562_),
            .C(LoadCtl_6_bF$buf0),
            .Y(_572_)
        );
        
        OAI22X1 _1356_ (
            .A(_110_),
            .B(LoadCtl_6_bF$buf4),
            .C(_572_),
            .D(_571_),
            .Y(_20_)
        );
        
        OAI21X1 _1357_ (
            .A(_570_),
            .B(_562_),
            .C(_567_),
            .Y(_573_)
        );
        
        NAND3X1 _1358_ (
            .A(_183__bF$buf1),
            .B(_492_),
            .C(_201__bF$buf4),
            .Y(_574_)
        );
        
        OAI21X1 _1359_ (
            .A(Stg_2_bF$buf2),
            .B(Stg_0_bF$buf0),
            .C(Ain12b_11_bF$buf0),
            .Y(_575_)
        );
        
        NAND2X1 _1360_ (
            .A(_575_),
            .B(_574_),
            .Y(_576_)
        );
        
        INVX1 _1361_ (
            .A(_576_),
            .Y(_577_)
        );
        
        NAND2X1 _1362_ (
            .A(Ain12b[7]),
            .B(_577_),
            .Y(_578_)
        );
        
        INVX1 _1363_ (
            .A(_578_),
            .Y(_579_)
        );
        
        NOR2X1 _1364_ (
            .A(Ain12b[7]),
            .B(_577_),
            .Y(_580_)
        );
        
        NOR2X1 _1365_ (
            .A(_580_),
            .B(_579_),
            .Y(_581_)
        );
        
        INVX1 _1366_ (
            .A(_581_),
            .Y(_582_)
        );
        
        OR2X2 _1367_ (
            .A(_573_),
            .B(_582_),
            .Y(_583_)
        );
        
        AOI21X1 _1368_ (
            .A(_573_),
            .B(_582_),
            .C(_188__bF$buf2),
            .Y(_584_)
        );
        
        AOI22X1 _1369_ (
            .A(_124_),
            .B(_188__bF$buf1),
            .C(_583_),
            .D(_584_),
            .Y(_21_)
        );
        
        NAND2X1 _1370_ (
            .A(Acalc[8]),
            .B(_188__bF$buf0),
            .Y(_585_)
        );
        
        NAND2X1 _1371_ (
            .A(_201__bF$buf3),
            .B(_292_),
            .Y(_586_)
        );
        
        NAND2X1 _1372_ (
            .A(_521_),
            .B(_586_),
            .Y(_587_)
        );
        
        INVX1 _1373_ (
            .A(_587_),
            .Y(_588_)
        );
        
        NAND2X1 _1374_ (
            .A(Ain12b[8]),
            .B(_588_),
            .Y(_589_)
        );
        
        INVX1 _1375_ (
            .A(Ain12b[8]),
            .Y(_590_)
        );
        
        NAND2X1 _1376_ (
            .A(_590_),
            .B(_587_),
            .Y(_591_)
        );
        
        NAND2X1 _1377_ (
            .A(_591_),
            .B(_589_),
            .Y(_592_)
        );
        
        INVX1 _1378_ (
            .A(_592_),
            .Y(_593_)
        );
        
        OAI21X1 _1379_ (
            .A(_580_),
            .B(_567_),
            .C(_578_),
            .Y(_594_)
        );
        
        OR2X2 _1380_ (
            .A(_570_),
            .B(_582_),
            .Y(_595_)
        );
        
        INVX1 _1381_ (
            .A(_595_),
            .Y(_596_)
        );
        
        AOI21X1 _1382_ (
            .A(_561_),
            .B(_596_),
            .C(_594_),
            .Y(_597_)
        );
        
        NAND2X1 _1383_ (
            .A(_596_),
            .B(_560_),
            .Y(_598_)
        );
        
        OAI21X1 _1384_ (
            .A(_598_),
            .B(_542_),
            .C(_597_),
            .Y(_599_)
        );
        
        NOR2X1 _1385_ (
            .A(_593_),
            .B(_599_),
            .Y(_600_)
        );
        
        INVX1 _1386_ (
            .A(_599_),
            .Y(_601_)
        );
        
        OAI21X1 _1387_ (
            .A(_592_),
            .B(_601_),
            .C(LoadCtl_6_bF$buf3),
            .Y(_602_)
        );
        
        OAI21X1 _1388_ (
            .A(_600_),
            .B(_602_),
            .C(_585_),
            .Y(_22_)
        );
        
        NAND2X1 _1389_ (
            .A(Acalc[9]),
            .B(_188__bF$buf4),
            .Y(_603_)
        );
        
        INVX1 _1390_ (
            .A(_589_),
            .Y(_604_)
        );
        
        AOI21X1 _1391_ (
            .A(_599_),
            .B(_593_),
            .C(_604_),
            .Y(_605_)
        );
        
        INVX1 _1392_ (
            .A(Ain12b[9]),
            .Y(_606_)
        );
        
        NAND2X1 _1393_ (
            .A(Ain12b_11_bF$buf4),
            .B(_606_),
            .Y(_607_)
        );
        
        NAND2X1 _1394_ (
            .A(Ain12b[9]),
            .B(_201__bF$buf2),
            .Y(_608_)
        );
        
        NAND2X1 _1395_ (
            .A(_607_),
            .B(_608_),
            .Y(_609_)
        );
        
        AND2X2 _1396_ (
            .A(_605_),
            .B(_609_),
            .Y(_610_)
        );
        
        OAI21X1 _1397_ (
            .A(_609_),
            .B(_605_),
            .C(LoadCtl_6_bF$buf2),
            .Y(_611_)
        );
        
        OAI21X1 _1398_ (
            .A(_611_),
            .B(_610_),
            .C(_603_),
            .Y(_23_)
        );
        
        OAI21X1 _1399_ (
            .A(_609_),
            .B(_589_),
            .C(_608_),
            .Y(_612_)
        );
        
        OR2X2 _1400_ (
            .A(_592_),
            .B(_609_),
            .Y(_613_)
        );
        
        INVX1 _1401_ (
            .A(_613_),
            .Y(_614_)
        );
        
        AOI21X1 _1402_ (
            .A(_599_),
            .B(_614_),
            .C(_612_),
            .Y(_615_)
        );
        
        INVX1 _1403_ (
            .A(Ain12b[10]),
            .Y(_616_)
        );
        
        NAND2X1 _1404_ (
            .A(Ain12b_11_bF$buf3),
            .B(_616_),
            .Y(_617_)
        );
        
        NAND2X1 _1405_ (
            .A(Ain12b[10]),
            .B(_201__bF$buf1),
            .Y(_618_)
        );
        
        NAND2X1 _1406_ (
            .A(_617_),
            .B(_618_),
            .Y(_619_)
        );
        
        AND2X2 _1407_ (
            .A(_615_),
            .B(_619_),
            .Y(_620_)
        );
        
        OAI21X1 _1408_ (
            .A(_619_),
            .B(_615_),
            .C(LoadCtl_6_bF$buf1),
            .Y(_621_)
        );
        
        OAI22X1 _1409_ (
            .A(_106_),
            .B(LoadCtl_6_bF$buf0),
            .C(_621_),
            .D(_620_),
            .Y(_24_)
        );
        
        NAND2X1 _1410_ (
            .A(Acalc[11]),
            .B(_188__bF$buf3),
            .Y(_622_)
        );
        
        OAI21X1 _1411_ (
            .A(_619_),
            .B(_615_),
            .C(_618_),
            .Y(_623_)
        );
        
        OAI21X1 _1412_ (
            .A(_188__bF$buf2),
            .B(_623_),
            .C(_622_),
            .Y(_25_)
        );
        
        NAND3X1 _1413_ (
            .A(LoadCtl[5]),
            .B(_137_),
            .C(_109_),
            .Y(_624_)
        );
        
        NOR2X1 _1414_ (
            .A(_117_),
            .B(_624_),
            .Y(_625_)
        );
        
        NAND2X1 _1415_ (
            .A(Xin[0]),
            .B(_625_),
            .Y(_626_)
        );
        
        OAI21X1 _1416_ (
            .A(_458_),
            .B(_625_),
            .C(_626_),
            .Y(_26_)
        );
        
        NAND2X1 _1417_ (
            .A(Xin[1]),
            .B(_625_),
            .Y(_627_)
        );
        
        OAI21X1 _1418_ (
            .A(_471_),
            .B(_625_),
            .C(_627_),
            .Y(_27_)
        );
        
        NOR2X1 _1419_ (
            .A(_137_),
            .B(_117_),
            .Y(_628_)
        );
        
        AND2X2 _1420_ (
            .A(_628_),
            .B(_109_),
            .Y(_629_)
        );
        
        NAND2X1 _1421_ (
            .A(Xin[0]),
            .B(_629_),
            .Y(_630_)
        );
        
        OAI21X1 _1422_ (
            .A(_422_),
            .B(_629_),
            .C(_630_),
            .Y(_28_)
        );
        
        NAND2X1 _1423_ (
            .A(Xin[1]),
            .B(_629_),
            .Y(_631_)
        );
        
        OAI21X1 _1424_ (
            .A(_441_),
            .B(_629_),
            .C(_631_),
            .Y(_29_)
        );
        
        NOR2X1 _1425_ (
            .A(_113_),
            .B(_117_),
            .Y(_632_)
        );
        
        NAND2X1 _1426_ (
            .A(Xin[0]),
            .B(_632_),
            .Y(_633_)
        );
        
        OAI21X1 _1427_ (
            .A(_172_),
            .B(_632_),
            .C(_633_),
            .Y(_30_)
        );
        
        NAND2X1 _1428_ (
            .A(Xin[1]),
            .B(_632_),
            .Y(_634_)
        );
        
        OAI21X1 _1429_ (
            .A(_209_),
            .B(_632_),
            .C(_634_),
            .Y(_31_)
        );
        
        NOR2X1 _1430_ (
            .A(_112_),
            .B(_117_),
            .Y(_635_)
        );
        
        NAND2X1 _1431_ (
            .A(Xin[0]),
            .B(_635_),
            .Y(_636_)
        );
        
        OAI21X1 _1432_ (
            .A(_175_),
            .B(_635_),
            .C(_636_),
            .Y(_32_)
        );
        
        NAND2X1 _1433_ (
            .A(Xin[1]),
            .B(_635_),
            .Y(_637_)
        );
        
        OAI21X1 _1434_ (
            .A(_212_),
            .B(_635_),
            .C(_637_),
            .Y(_33_)
        );
        
        NAND2X1 _1435_ (
            .A(Xin[0]),
            .B(_119_),
            .Y(_638_)
        );
        
        OAI21X1 _1436_ (
            .A(_165_),
            .B(_119_),
            .C(_638_),
            .Y(_34_)
        );
        
        NAND2X1 _1437_ (
            .A(Xin[1]),
            .B(_119_),
            .Y(_639_)
        );
        
        OAI21X1 _1438_ (
            .A(_202_),
            .B(_119_),
            .C(_639_),
            .Y(_35_)
        );
        
        NAND2X1 _1439_ (
            .A(LoadCtl_0_bF$buf3),
            .B(Xin[0]),
            .Y(_640_)
        );
        
        OAI21X1 _1440_ (
            .A(LoadCtl_0_bF$buf2),
            .B(_168_),
            .C(_640_),
            .Y(_36_)
        );
        
        NAND2X1 _1441_ (
            .A(LoadCtl_0_bF$buf1),
            .B(Xin[1]),
            .Y(_641_)
        );
        
        OAI21X1 _1442_ (
            .A(LoadCtl_0_bF$buf0),
            .B(_205_),
            .C(_641_),
            .Y(_37_)
        );
        
        NAND2X1 _1443_ (
            .A(Yin[0]),
            .B(_625_),
            .Y(_642_)
        );
        
        OAI21X1 _1444_ (
            .A(_311_),
            .B(_625_),
            .C(_642_),
            .Y(_38_)
        );
        
        NAND2X1 _1445_ (
            .A(Yin[1]),
            .B(_625_),
            .Y(_643_)
        );
        
        OAI21X1 _1446_ (
            .A(_356_),
            .B(_625_),
            .C(_643_),
            .Y(_39_)
        );
        
        INVX1 _1447_ (
            .A(Yin12b[8]),
            .Y(_644_)
        );
        
        NAND2X1 _1448_ (
            .A(Yin[0]),
            .B(_629_),
            .Y(_645_)
        );
        
        OAI21X1 _1449_ (
            .A(_644_),
            .B(_629_),
            .C(_645_),
            .Y(_40_)
        );
        
        NAND2X1 _1450_ (
            .A(Yin[1]),
            .B(_629_),
            .Y(_646_)
        );
        
        OAI21X1 _1451_ (
            .A(_284_),
            .B(_629_),
            .C(_646_),
            .Y(_41_)
        );
        
        NAND2X1 _1452_ (
            .A(Yin[0]),
            .B(_632_),
            .Y(_647_)
        );
        
        OAI21X1 _1453_ (
            .A(_241_),
            .B(_632_),
            .C(_647_),
            .Y(_42_)
        );
        
        NAND2X1 _1454_ (
            .A(Yin[1]),
            .B(_632_),
            .Y(_648_)
        );
        
        OAI21X1 _1455_ (
            .A(_262_),
            .B(_632_),
            .C(_648_),
            .Y(_43_)
        );
        
        NAND2X1 _1456_ (
            .A(Yin[0]),
            .B(_635_),
            .Y(_649_)
        );
        
        OAI21X1 _1457_ (
            .A(_244_),
            .B(_635_),
            .C(_649_),
            .Y(_44_)
        );
        
        NAND2X1 _1458_ (
            .A(Yin[1]),
            .B(_635_),
            .Y(_650_)
        );
        
        OAI21X1 _1459_ (
            .A(_265_),
            .B(_635_),
            .C(_650_),
            .Y(_45_)
        );
        
        NAND2X1 _1460_ (
            .A(Yin[0]),
            .B(_119_),
            .Y(_651_)
        );
        
        OAI21X1 _1461_ (
            .A(_234_),
            .B(_119_),
            .C(_651_),
            .Y(_46_)
        );
        
        NAND2X1 _1462_ (
            .A(Yin[1]),
            .B(_119_),
            .Y(_652_)
        );
        
        OAI21X1 _1463_ (
            .A(_256_),
            .B(_119_),
            .C(_652_),
            .Y(_47_)
        );
        
        NAND2X1 _1464_ (
            .A(LoadCtl_0_bF$buf3),
            .B(Yin[0]),
            .Y(_653_)
        );
        
        OAI21X1 _1465_ (
            .A(LoadCtl_0_bF$buf2),
            .B(_163_),
            .C(_653_),
            .Y(_48_)
        );
        
        NAND2X1 _1466_ (
            .A(LoadCtl_0_bF$buf1),
            .B(Yin[1]),
            .Y(_654_)
        );
        
        OAI21X1 _1467_ (
            .A(LoadCtl_0_bF$buf0),
            .B(_200_),
            .C(_654_),
            .Y(_49_)
        );
        
        NAND2X1 _1468_ (
            .A(Ain[0]),
            .B(_625_),
            .Y(_655_)
        );
        
        OAI21X1 _1469_ (
            .A(_616_),
            .B(_625_),
            .C(_655_),
            .Y(_50_)
        );
        
        NAND2X1 _1470_ (
            .A(Ain[1]),
            .B(_625_),
            .Y(_656_)
        );
        
        OAI21X1 _1471_ (
            .A(_201__bF$buf0),
            .B(_625_),
            .C(_656_),
            .Y(_51_)
        );
        
        NAND2X1 _1472_ (
            .A(Ain[0]),
            .B(_629_),
            .Y(_657_)
        );
        
        OAI21X1 _1473_ (
            .A(_590_),
            .B(_629_),
            .C(_657_),
            .Y(_52_)
        );
        
        NAND2X1 _1474_ (
            .A(Ain[1]),
            .B(_629_),
            .Y(_658_)
        );
        
        OAI21X1 _1475_ (
            .A(_606_),
            .B(_629_),
            .C(_658_),
            .Y(_53_)
        );
        
        NAND2X1 _1476_ (
            .A(Ain[0]),
            .B(_632_),
            .Y(_659_)
        );
        
        OAI21X1 _1477_ (
            .A(_568_),
            .B(_632_),
            .C(_659_),
            .Y(_54_)
        );
        
        INVX1 _1478_ (
            .A(Ain[1]),
            .Y(_660_)
        );
        
        NOR2X1 _1479_ (
            .A(Ain12b[7]),
            .B(_632_),
            .Y(_661_)
        );
        
        AOI21X1 _1480_ (
            .A(_660_),
            .B(_632_),
            .C(_661_),
            .Y(_55_)
        );
        
        NAND2X1 _1481_ (
            .A(Ain[0]),
            .B(_635_),
            .Y(_662_)
        );
        
        OAI21X1 _1482_ (
            .A(_537_),
            .B(_635_),
            .C(_662_),
            .Y(_56_)
        );
        
        NAND2X1 _1483_ (
            .A(Ain[1]),
            .B(_635_),
            .Y(_663_)
        );
        
        OAI21X1 _1484_ (
            .A(_553_),
            .B(_635_),
            .C(_663_),
            .Y(_57_)
        );
        
        INVX1 _1485_ (
            .A(Ain[0]),
            .Y(_664_)
        );
        
        INVX1 _1486_ (
            .A(_119_),
            .Y(_665_)
        );
        
        OAI21X1 _1487_ (
            .A(LoadCtl_0_bF$buf3),
            .B(_118_),
            .C(Ain1[0]),
            .Y(_666_)
        );
        
        OAI21X1 _1488_ (
            .A(_664_),
            .B(_665_),
            .C(_666_),
            .Y(_58_)
        );
        
        OAI21X1 _1489_ (
            .A(LoadCtl_0_bF$buf2),
            .B(_118_),
            .C(Ain1[1]),
            .Y(_667_)
        );
        
        OAI21X1 _1490_ (
            .A(_660_),
            .B(_665_),
            .C(_667_),
            .Y(_59_)
        );
        
        NAND2X1 _1491_ (
            .A(LoadCtl_0_bF$buf1),
            .B(Ain[0]),
            .Y(_668_)
        );
        
        OAI21X1 _1492_ (
            .A(LoadCtl_0_bF$buf0),
            .B(_483_),
            .C(_668_),
            .Y(_60_)
        );
        
        NAND2X1 _1493_ (
            .A(LoadCtl_0_bF$buf3),
            .B(Ain[1]),
            .Y(_669_)
        );
        
        OAI21X1 _1494_ (
            .A(LoadCtl_0_bF$buf2),
            .B(_504_),
            .C(_669_),
            .Y(_61_)
        );
        
        INVX1 _1495_ (
            .A(_860_),
            .Y(_670_)
        );
        
        NAND2X1 _1496_ (
            .A(LoadCtl_6_bF$buf4),
            .B(ISin),
            .Y(_671_)
        );
        
        OAI21X1 _1497_ (
            .A(LoadCtl_6_bF$buf3),
            .B(_670_),
            .C(_671_),
            .Y(_62_)
        );
        
        NAND2X1 _1498_ (
            .A(Ycalc[2]),
            .B(_188__bF$buf1),
            .Y(_672_)
        );
        
        AOI21X1 _1499_ (
            .A(_181_),
            .B(_228_),
            .C(_226_),
            .Y(_673_)
        );
        
        NAND2X1 _1500_ (
            .A(_199_),
            .B(_224_),
            .Y(_674_)
        );
        
        MUX2X1 _1501_ (
            .A(Xin12b[9]),
            .B(Xin12b[8]),
            .S(Stg_0_bF$buf6),
            .Y(_675_)
        );
        
        MUX2X1 _1502_ (
            .A(_675_),
            .B(_196_),
            .S(Stg_1_bF$buf3),
            .Y(_676_)
        );
        
        OAI22X1 _1503_ (
            .A(_184_),
            .B(_193_),
            .C(_197_),
            .D(_289_),
            .Y(_677_)
        );
        
        AOI21X1 _1504_ (
            .A(Stg_2_bF$buf1),
            .B(_676_),
            .C(_677_),
            .Y(_678_)
        );
        
        NAND3X1 _1505_ (
            .A(_201__bF$buf6),
            .B(_678_),
            .C(_674_),
            .Y(_679_)
        );
        
        NAND2X1 _1506_ (
            .A(_492_),
            .B(_165_),
            .Y(_680_)
        );
        
        NAND2X1 _1507_ (
            .A(Stg_0_bF$buf5),
            .B(_202_),
            .Y(_681_)
        );
        
        NAND3X1 _1508_ (
            .A(Stg_1_bF$buf2),
            .B(_681_),
            .C(_680_),
            .Y(_682_)
        );
        
        NAND2X1 _1509_ (
            .A(_164__bF$buf1),
            .B(_170_),
            .Y(_683_)
        );
        
        NAND3X1 _1510_ (
            .A(_183__bF$buf0),
            .B(_682_),
            .C(_683_),
            .Y(_684_)
        );
        
        NAND2X1 _1511_ (
            .A(_492_),
            .B(_175_),
            .Y(_685_)
        );
        
        NAND2X1 _1512_ (
            .A(Stg_0_bF$buf4),
            .B(_212_),
            .Y(_686_)
        );
        
        NAND3X1 _1513_ (
            .A(_164__bF$buf0),
            .B(_686_),
            .C(_685_),
            .Y(_687_)
        );
        
        NAND2X1 _1514_ (
            .A(Stg_1_bF$buf1),
            .B(_174_),
            .Y(_688_)
        );
        
        NAND3X1 _1515_ (
            .A(Stg_2_bF$buf0),
            .B(_687_),
            .C(_688_),
            .Y(_689_)
        );
        
        NAND2X1 _1516_ (
            .A(Stg_1_bF$buf0),
            .B(_204_),
            .Y(_690_)
        );
        
        NAND2X1 _1517_ (
            .A(_164__bF$buf4),
            .B(_207_),
            .Y(_691_)
        );
        
        NAND3X1 _1518_ (
            .A(_183__bF$buf3),
            .B(_690_),
            .C(_691_),
            .Y(_692_)
        );
        
        NAND2X1 _1519_ (
            .A(_164__bF$buf3),
            .B(_214_),
            .Y(_693_)
        );
        
        NAND2X1 _1520_ (
            .A(Stg_1_bF$buf3),
            .B(_211_),
            .Y(_694_)
        );
        
        NAND3X1 _1521_ (
            .A(Stg_2_bF$buf4),
            .B(_693_),
            .C(_694_),
            .Y(_695_)
        );
        
        AOI22X1 _1522_ (
            .A(_684_),
            .B(_689_),
            .C(_692_),
            .D(_695_),
            .Y(_696_)
        );
        
        INVX1 _1523_ (
            .A(_678_),
            .Y(_697_)
        );
        
        OAI21X1 _1524_ (
            .A(Ain12b_11_bF$buf2),
            .B(_696_),
            .C(_697_),
            .Y(_698_)
        );
        
        AOI21X1 _1525_ (
            .A(_698_),
            .B(_679_),
            .C(Yin1[0]),
            .Y(_699_)
        );
        
        NAND3X1 _1526_ (
            .A(Yin1[0]),
            .B(_679_),
            .C(_698_),
            .Y(_700_)
        );
        
        INVX1 _1527_ (
            .A(_700_),
            .Y(_701_)
        );
        
        OR2X2 _1528_ (
            .A(_701_),
            .B(_699_),
            .Y(_702_)
        );
        
        NOR2X1 _1529_ (
            .A(_673_),
            .B(_702_),
            .Y(_703_)
        );
        
        INVX1 _1530_ (
            .A(_703_),
            .Y(_704_)
        );
        
        OAI21X1 _1531_ (
            .A(_699_),
            .B(_701_),
            .C(_673_),
            .Y(_705_)
        );
        
        AOI21X1 _1532_ (
            .A(_704_),
            .B(_705_),
            .C(_192_),
            .Y(_706_)
        );
        
        OAI21X1 _1533_ (
            .A(Stg_1_bF$buf2),
            .B(_574_),
            .C(LoadCtl_6_bF$buf2),
            .Y(_707_)
        );
        
        OAI21X1 _1534_ (
            .A(_707_),
            .B(_706_),
            .C(_672_),
            .Y(_63_)
        );
        
        INVX1 _1535_ (
            .A(Ycalc[3]),
            .Y(_708_)
        );
        
        INVX2 _1536_ (
            .A(_707_),
            .Y(_709_)
        );
        
        OAI21X1 _1537_ (
            .A(_699_),
            .B(_673_),
            .C(_700_),
            .Y(_710_)
        );
        
        INVX1 _1538_ (
            .A(_710_),
            .Y(_711_)
        );
        
        NAND3X1 _1539_ (
            .A(_678_),
            .B(_199_),
            .C(_224_),
            .Y(_712_)
        );
        
        NAND2X1 _1540_ (
            .A(Stg_0_bF$buf3),
            .B(Xin12b[10]),
            .Y(_713_)
        );
        
        OAI21X1 _1541_ (
            .A(Stg_0_bF$buf2),
            .B(_441_),
            .C(_713_),
            .Y(_714_)
        );
        
        NAND2X1 _1542_ (
            .A(_164__bF$buf2),
            .B(_221_),
            .Y(_715_)
        );
        
        OAI21X1 _1543_ (
            .A(_164__bF$buf1),
            .B(_714_),
            .C(_715_),
            .Y(_716_)
        );
        
        OAI22X1 _1544_ (
            .A(_184_),
            .B(_218_),
            .C(_222_),
            .D(_289_),
            .Y(_717_)
        );
        
        INVX1 _1545_ (
            .A(_717_),
            .Y(_718_)
        );
        
        OAI21X1 _1546_ (
            .A(_183__bF$buf2),
            .B(_716_),
            .C(_718_),
            .Y(_719_)
        );
        
        NAND3X1 _1547_ (
            .A(_201__bF$buf5),
            .B(_719_),
            .C(_712_),
            .Y(_720_)
        );
        
        INVX1 _1548_ (
            .A(_712_),
            .Y(_721_)
        );
        
        NAND2X1 _1549_ (
            .A(Stg_0_bF$buf1),
            .B(_458_),
            .Y(_722_)
        );
        
        OAI21X1 _1550_ (
            .A(Stg_0_bF$buf0),
            .B(Xin12b[9]),
            .C(_722_),
            .Y(_723_)
        );
        
        NAND2X1 _1551_ (
            .A(_164__bF$buf0),
            .B(_211_),
            .Y(_724_)
        );
        
        OAI21X1 _1552_ (
            .A(_164__bF$buf4),
            .B(_723_),
            .C(_724_),
            .Y(_725_)
        );
        
        AOI21X1 _1553_ (
            .A(_725_),
            .B(Stg_2_bF$buf3),
            .C(_717_),
            .Y(_726_)
        );
        
        OAI21X1 _1554_ (
            .A(Ain12b_11_bF$buf1),
            .B(_721_),
            .C(_726_),
            .Y(_727_)
        );
        
        NAND2X1 _1555_ (
            .A(_720_),
            .B(_727_),
            .Y(_728_)
        );
        
        NAND2X1 _1556_ (
            .A(Yin1[1]),
            .B(_728_),
            .Y(_729_)
        );
        
        NOR2X1 _1557_ (
            .A(Yin1[1]),
            .B(_728_),
            .Y(_730_)
        );
        
        INVX1 _1558_ (
            .A(_730_),
            .Y(_731_)
        );
        
        NAND2X1 _1559_ (
            .A(_729_),
            .B(_731_),
            .Y(_732_)
        );
        
        AOI21X1 _1560_ (
            .A(_732_),
            .B(_711_),
            .C(_192_),
            .Y(_733_)
        );
        
        OAI21X1 _1561_ (
            .A(_711_),
            .B(_732_),
            .C(_733_),
            .Y(_734_)
        );
        
        AOI22X1 _1562_ (
            .A(_708_),
            .B(_188__bF$buf0),
            .C(_734_),
            .D(_709_),
            .Y(_64_)
        );
        
        NAND3X1 _1563_ (
            .A(_678_),
            .B(_726_),
            .C(_696_),
            .Y(_735_)
        );
        
        NAND2X1 _1564_ (
            .A(Stg_0_bF$buf6),
            .B(Xin12b[11]),
            .Y(_736_)
        );
        
        OAI21X1 _1565_ (
            .A(Stg_0_bF$buf5),
            .B(_458_),
            .C(_736_),
            .Y(_737_)
        );
        
        NAND2X1 _1566_ (
            .A(Stg_1_bF$buf1),
            .B(_737_),
            .Y(_738_)
        );
        
        OAI21X1 _1567_ (
            .A(Stg_1_bF$buf0),
            .B(_675_),
            .C(_738_),
            .Y(_739_)
        );
        
        NAND2X1 _1568_ (
            .A(Stg_2_bF$buf2),
            .B(_739_),
            .Y(_740_)
        );
        
        OAI21X1 _1569_ (
            .A(Stg_2_bF$buf1),
            .B(_178_),
            .C(_740_),
            .Y(_741_)
        );
        
        NAND3X1 _1570_ (
            .A(_201__bF$buf4),
            .B(_741_),
            .C(_735_),
            .Y(_742_)
        );
        
        NOR2X1 _1571_ (
            .A(_719_),
            .B(_712_),
            .Y(_743_)
        );
        
        INVX1 _1572_ (
            .A(_741_),
            .Y(_744_)
        );
        
        OAI21X1 _1573_ (
            .A(Ain12b_11_bF$buf0),
            .B(_743_),
            .C(_744_),
            .Y(_745_)
        );
        
        NAND3X1 _1574_ (
            .A(_244_),
            .B(_742_),
            .C(_745_),
            .Y(_746_)
        );
        
        INVX1 _1575_ (
            .A(_742_),
            .Y(_747_)
        );
        
        AOI21X1 _1576_ (
            .A(_735_),
            .B(_201__bF$buf3),
            .C(_741_),
            .Y(_748_)
        );
        
        OAI21X1 _1577_ (
            .A(_748_),
            .B(_747_),
            .C(Yin12b[4]),
            .Y(_749_)
        );
        
        NAND2X1 _1578_ (
            .A(_746_),
            .B(_749_),
            .Y(_750_)
        );
        
        OAI21X1 _1579_ (
            .A(Yin1[1]),
            .B(_728_),
            .C(_710_),
            .Y(_751_)
        );
        
        AND2X2 _1580_ (
            .A(_751_),
            .B(_729_),
            .Y(_752_)
        );
        
        AOI21X1 _1581_ (
            .A(_752_),
            .B(_750_),
            .C(_192_),
            .Y(_753_)
        );
        
        OAI21X1 _1582_ (
            .A(_750_),
            .B(_752_),
            .C(_753_),
            .Y(_754_)
        );
        
        AOI22X1 _1583_ (
            .A(_133_),
            .B(_188__bF$buf4),
            .C(_754_),
            .D(_709_),
            .Y(_65_)
        );
        
        AOI21X1 _1584_ (
            .A(_751_),
            .B(_729_),
            .C(_750_),
            .Y(_755_)
        );
        
        INVX1 _1585_ (
            .A(_755_),
            .Y(_756_)
        );
        
        NOR2X1 _1586_ (
            .A(_164__bF$buf3),
            .B(_471_),
            .Y(_757_)
        );
        
        AOI21X1 _1587_ (
            .A(_164__bF$buf2),
            .B(_714_),
            .C(_757_),
            .Y(_758_)
        );
        
        NAND2X1 _1588_ (
            .A(_183__bF$buf1),
            .B(_223_),
            .Y(_759_)
        );
        
        OAI21X1 _1589_ (
            .A(_183__bF$buf0),
            .B(_758_),
            .C(_759_),
            .Y(_760_)
        );
        
        INVX1 _1590_ (
            .A(_760_),
            .Y(_761_)
        );
        
        OAI21X1 _1591_ (
            .A(_741_),
            .B(_735_),
            .C(_201__bF$buf2),
            .Y(_762_)
        );
        
        NOR2X1 _1592_ (
            .A(_761_),
            .B(_762_),
            .Y(_763_)
        );
        
        INVX1 _1593_ (
            .A(_763_),
            .Y(_764_)
        );
        
        NAND2X1 _1594_ (
            .A(_761_),
            .B(_762_),
            .Y(_765_)
        );
        
        NAND3X1 _1595_ (
            .A(_265_),
            .B(_765_),
            .C(_764_),
            .Y(_766_)
        );
        
        INVX1 _1596_ (
            .A(_765_),
            .Y(_767_)
        );
        
        OAI21X1 _1597_ (
            .A(_763_),
            .B(_767_),
            .C(Yin12b[5]),
            .Y(_768_)
        );
        
        AND2X2 _1598_ (
            .A(_766_),
            .B(_768_),
            .Y(_769_)
        );
        
        AOI21X1 _1599_ (
            .A(_756_),
            .B(_749_),
            .C(_769_),
            .Y(_770_)
        );
        
        NAND3X1 _1600_ (
            .A(_749_),
            .B(_769_),
            .C(_756_),
            .Y(_771_)
        );
        
        OAI21X1 _1601_ (
            .A(Stg_2_bF$buf0),
            .B(_484_),
            .C(_771_),
            .Y(_772_)
        );
        
        OAI21X1 _1602_ (
            .A(_770_),
            .B(_772_),
            .C(_709_),
            .Y(_773_)
        );
        
        OAI21X1 _1603_ (
            .A(_142_),
            .B(LoadCtl_6_bF$buf1),
            .C(_773_),
            .Y(_66_)
        );
        
        NAND3X1 _1604_ (
            .A(_744_),
            .B(_761_),
            .C(_743_),
            .Y(_774_)
        );
        
        AOI21X1 _1605_ (
            .A(_164__bF$buf1),
            .B(_737_),
            .C(_757_),
            .Y(_775_)
        );
        
        NAND2X1 _1606_ (
            .A(_183__bF$buf3),
            .B(_676_),
            .Y(_776_)
        );
        
        OAI21X1 _1607_ (
            .A(_183__bF$buf2),
            .B(_775_),
            .C(_776_),
            .Y(_777_)
        );
        
        NAND3X1 _1608_ (
            .A(_201__bF$buf1),
            .B(_777_),
            .C(_774_),
            .Y(_778_)
        );
        
        NOR3X1 _1609_ (
            .A(_741_),
            .B(_760_),
            .C(_735_),
            .Y(_779_)
        );
        
        INVX1 _1610_ (
            .A(_777_),
            .Y(_780_)
        );
        
        OAI21X1 _1611_ (
            .A(Ain12b_11_bF$buf4),
            .B(_779_),
            .C(_780_),
            .Y(_781_)
        );
        
        NAND3X1 _1612_ (
            .A(_241_),
            .B(_778_),
            .C(_781_),
            .Y(_782_)
        );
        
        NAND3X1 _1613_ (
            .A(_201__bF$buf0),
            .B(_780_),
            .C(_774_),
            .Y(_783_)
        );
        
        OAI21X1 _1614_ (
            .A(Ain12b_11_bF$buf3),
            .B(_779_),
            .C(_777_),
            .Y(_784_)
        );
        
        NAND3X1 _1615_ (
            .A(Yin12b[6]),
            .B(_783_),
            .C(_784_),
            .Y(_785_)
        );
        
        NAND2X1 _1616_ (
            .A(_782_),
            .B(_785_),
            .Y(_786_)
        );
        
        NAND2X1 _1617_ (
            .A(_749_),
            .B(_768_),
            .Y(_787_)
        );
        
        OAI21X1 _1618_ (
            .A(_787_),
            .B(_755_),
            .C(_766_),
            .Y(_788_)
        );
        
        AOI21X1 _1619_ (
            .A(_788_),
            .B(_786_),
            .C(_192_),
            .Y(_789_)
        );
        
        OAI21X1 _1620_ (
            .A(_786_),
            .B(_788_),
            .C(_789_),
            .Y(_790_)
        );
        
        AOI22X1 _1621_ (
            .A(_132_),
            .B(_188__bF$buf3),
            .C(_790_),
            .D(_709_),
            .Y(_67_)
        );
        
        INVX1 _1622_ (
            .A(_785_),
            .Y(_791_)
        );
        
        AND2X2 _1623_ (
            .A(_749_),
            .B(_746_),
            .Y(_792_)
        );
        
        NAND3X1 _1624_ (
            .A(_768_),
            .B(_766_),
            .C(_792_),
            .Y(_793_)
        );
        
        INVX1 _1625_ (
            .A(_749_),
            .Y(_794_)
        );
        
        AOI21X1 _1626_ (
            .A(_764_),
            .B(_765_),
            .C(_265_),
            .Y(_795_)
        );
        
        AOI21X1 _1627_ (
            .A(_794_),
            .B(_766_),
            .C(_795_),
            .Y(_796_)
        );
        
        OAI21X1 _1628_ (
            .A(_793_),
            .B(_752_),
            .C(_796_),
            .Y(_797_)
        );
        
        AOI21X1 _1629_ (
            .A(_797_),
            .B(_782_),
            .C(_791_),
            .Y(_798_)
        );
        
        NAND2X1 _1630_ (
            .A(_780_),
            .B(_779_),
            .Y(_799_)
        );
        
        NOR2X1 _1631_ (
            .A(_183__bF$buf1),
            .B(_471_),
            .Y(_800_)
        );
        
        AOI21X1 _1632_ (
            .A(_725_),
            .B(_183__bF$buf0),
            .C(_800_),
            .Y(_801_)
        );
        
        NAND3X1 _1633_ (
            .A(_201__bF$buf6),
            .B(_801_),
            .C(_799_),
            .Y(_802_)
        );
        
        INVX1 _1634_ (
            .A(_801_),
            .Y(_803_)
        );
        
        OAI21X1 _1635_ (
            .A(_777_),
            .B(_774_),
            .C(_201__bF$buf5),
            .Y(_804_)
        );
        
        NAND2X1 _1636_ (
            .A(_803_),
            .B(_804_),
            .Y(_805_)
        );
        
        AOI21X1 _1637_ (
            .A(_805_),
            .B(_802_),
            .C(Yin12b[7]),
            .Y(_806_)
        );
        
        NAND3X1 _1638_ (
            .A(_201__bF$buf4),
            .B(_803_),
            .C(_799_),
            .Y(_807_)
        );
        
        NAND2X1 _1639_ (
            .A(_801_),
            .B(_804_),
            .Y(_808_)
        );
        
        AOI21X1 _1640_ (
            .A(_808_),
            .B(_807_),
            .C(_262_),
            .Y(_809_)
        );
        
        NOR2X1 _1641_ (
            .A(_806_),
            .B(_809_),
            .Y(_810_)
        );
        
        NOR2X1 _1642_ (
            .A(_810_),
            .B(_798_),
            .Y(_811_)
        );
        
        NAND2X1 _1643_ (
            .A(_810_),
            .B(_798_),
            .Y(_812_)
        );
        
        OAI21X1 _1644_ (
            .A(Stg_2_bF$buf4),
            .B(_484_),
            .C(_812_),
            .Y(_813_)
        );
        
        OAI21X1 _1645_ (
            .A(_201__bF$buf3),
            .B(_191_),
            .C(LoadCtl_6_bF$buf0),
            .Y(_814_)
        );
        
        INVX1 _1646_ (
            .A(_814_),
            .Y(_815_)
        );
        
        OAI21X1 _1647_ (
            .A(_811_),
            .B(_813_),
            .C(_815_),
            .Y(_816_)
        );
        
        OAI21X1 _1648_ (
            .A(_141_),
            .B(LoadCtl_6_bF$buf4),
            .C(_816_),
            .Y(_68_)
        );
        
        INVX1 _1649_ (
            .A(Ycalc[8]),
            .Y(_817_)
        );
        
        NAND3X1 _1650_ (
            .A(_262_),
            .B(_807_),
            .C(_808_),
            .Y(_818_)
        );
        
        AOI21X1 _1651_ (
            .A(_791_),
            .B(_818_),
            .C(_809_),
            .Y(_819_)
        );
        
        AND2X2 _1652_ (
            .A(_782_),
            .B(_785_),
            .Y(_820_)
        );
        
        NAND3X1 _1653_ (
            .A(Yin12b[7]),
            .B(_802_),
            .C(_805_),
            .Y(_821_)
        );
        
        NAND3X1 _1654_ (
            .A(_818_),
            .B(_821_),
            .C(_820_),
            .Y(_822_)
        );
        
        OAI21X1 _1655_ (
            .A(_822_),
            .B(_788_),
            .C(_819_),
            .Y(_823_)
        );
        
        NAND3X1 _1656_ (
            .A(_780_),
            .B(_801_),
            .C(_779_),
            .Y(_824_)
        );
        
        INVX1 _1657_ (
            .A(_739_),
            .Y(_825_)
        );
        
        INVX1 _1658_ (
            .A(_800_),
            .Y(_826_)
        );
        
        OAI21X1 _1659_ (
            .A(Stg_2_bF$buf3),
            .B(_825_),
            .C(_826_),
            .Y(_827_)
        );
        
        INVX1 _1660_ (
            .A(_827_),
            .Y(_828_)
        );
        
        NAND3X1 _1661_ (
            .A(_201__bF$buf2),
            .B(_828_),
            .C(_824_),
            .Y(_829_)
        );
        
        INVX1 _1662_ (
            .A(_829_),
            .Y(_830_)
        );
        
        AOI21X1 _1663_ (
            .A(_824_),
            .B(_201__bF$buf1),
            .C(_828_),
            .Y(_831_)
        );
        
        OAI21X1 _1664_ (
            .A(_831_),
            .B(_830_),
            .C(_644_),
            .Y(_832_)
        );
        
        OAI21X1 _1665_ (
            .A(_803_),
            .B(_799_),
            .C(_201__bF$buf0),
            .Y(_833_)
        );
        
        NAND2X1 _1666_ (
            .A(_827_),
            .B(_833_),
            .Y(_834_)
        );
        
        NAND3X1 _1667_ (
            .A(Yin12b[8]),
            .B(_829_),
            .C(_834_),
            .Y(_835_)
        );
        
        AND2X2 _1668_ (
            .A(_832_),
            .B(_835_),
            .Y(_836_)
        );
        
        AND2X2 _1669_ (
            .A(_823_),
            .B(_836_),
            .Y(_837_)
        );
        
        OAI21X1 _1670_ (
            .A(_836_),
            .B(_823_),
            .C(_191_),
            .Y(_838_)
        );
        
        OR2X2 _1671_ (
            .A(_837_),
            .B(_838_),
            .Y(_839_)
        );
        
        AOI22X1 _1672_ (
            .A(_817_),
            .B(_188__bF$buf2),
            .C(_839_),
            .D(_815_),
            .Y(_69_)
        );
        
        INVX1 _1673_ (
            .A(_835_),
            .Y(_840_)
        );
        
        NOR2X1 _1674_ (
            .A(_840_),
            .B(_837_),
            .Y(_841_)
        );
        
        NOR2X1 _1675_ (
            .A(_827_),
            .B(_824_),
            .Y(_842_)
        );
        
        OAI21X1 _1676_ (
            .A(Stg_2_bF$buf2),
            .B(_758_),
            .C(_826_),
            .Y(_843_)
        );
        
        INVX1 _1677_ (
            .A(_843_),
            .Y(_844_)
        );
        
        OAI21X1 _1678_ (
            .A(Ain12b_11_bF$buf2),
            .B(_842_),
            .C(_844_),
            .Y(_845_)
        );
        
        NOR2X1 _1679_ (
            .A(_777_),
            .B(_774_),
            .Y(_846_)
        );
        
        NAND3X1 _1680_ (
            .A(_801_),
            .B(_828_),
            .C(_846_),
            .Y(_847_)
        );
        
        NAND3X1 _1681_ (
            .A(_201__bF$buf6),
            .B(_843_),
            .C(_847_),
            .Y(_848_)
        );
        
        NAND3X1 _1682_ (
            .A(_284_),
            .B(_848_),
            .C(_845_),
            .Y(_849_)
        );
        
        AOI21X1 _1683_ (
            .A(_847_),
            .B(_201__bF$buf5),
            .C(_843_),
            .Y(_850_)
        );
        
        OAI21X1 _1684_ (
            .A(_827_),
            .B(_824_),
            .C(_201__bF$buf4),
            .Y(_851_)
        );
        
        NOR2X1 _1685_ (
            .A(_844_),
            .B(_851_),
            .Y(_852_)
        );
        
        OAI21X1 _1686_ (
            .A(_850_),
            .B(_852_),
            .C(Yin12b[9]),
            .Y(_853_)
        );
        
        AND2X2 _1687_ (
            .A(_853_),
            .B(_849_),
            .Y(_854_)
        );
        
        AND2X2 _1688_ (
            .A(_841_),
            .B(_854_),
            .Y(_855_)
        );
        
        OAI21X1 _1689_ (
            .A(_854_),
            .B(_841_),
            .C(_191_),
            .Y(_856_)
        );
        
        OAI21X1 _1690_ (
            .A(_856_),
            .B(_855_),
            .C(_709_),
            .Y(_857_)
        );
        
        OAI21X1 _1691_ (
            .A(_138_),
            .B(LoadCtl_6_bF$buf3),
            .C(_857_),
            .Y(_70_)
        );
        
        OAI21X1 _1692_ (
            .A(Stg_2_bF$buf1),
            .B(_775_),
            .C(_826_),
            .Y(_858_)
        );
        
        INVX1 _1693_ (
            .A(_858_),
            .Y(_73_)
        );
        
        OAI21X1 _1694_ (
            .A(_843_),
            .B(_847_),
            .C(_201__bF$buf3),
            .Y(_74_)
        );
        
        OR2X2 _1695_ (
            .A(_74_),
            .B(_73_),
            .Y(_75_)
        );
        
        NAND2X1 _1696_ (
            .A(_844_),
            .B(_842_),
            .Y(_76_)
        );
        
        AOI21X1 _1697_ (
            .A(_76_),
            .B(_201__bF$buf2),
            .C(_858_),
            .Y(_77_)
        );
        
        INVX1 _1698_ (
            .A(_77_),
            .Y(_78_)
        );
        
        NAND3X1 _1699_ (
            .A(_311_),
            .B(_75_),
            .C(_78_),
            .Y(_79_)
        );
        
        NOR2X1 _1700_ (
            .A(_73_),
            .B(_74_),
            .Y(_80_)
        );
        
        OAI21X1 _1701_ (
            .A(_77_),
            .B(_80_),
            .C(Yin12b[10]),
            .Y(_81_)
        );
        
        NAND2X1 _1702_ (
            .A(_81_),
            .B(_79_),
            .Y(_82_)
        );
        
        AOI21X1 _1703_ (
            .A(_845_),
            .B(_848_),
            .C(_284_),
            .Y(_83_)
        );
        
        AOI21X1 _1704_ (
            .A(_840_),
            .B(_849_),
            .C(_83_),
            .Y(_84_)
        );
        
        NAND3X1 _1705_ (
            .A(_836_),
            .B(_854_),
            .C(_823_),
            .Y(_85_)
        );
        
        AOI21X1 _1706_ (
            .A(_85_),
            .B(_84_),
            .C(_82_),
            .Y(_86_)
        );
        
        AND2X2 _1707_ (
            .A(_79_),
            .B(_81_),
            .Y(_87_)
        );
        
        OAI21X1 _1708_ (
            .A(_785_),
            .B(_806_),
            .C(_821_),
            .Y(_88_)
        );
        
        NOR3X1 _1709_ (
            .A(_786_),
            .B(_806_),
            .C(_809_),
            .Y(_89_)
        );
        
        AOI21X1 _1710_ (
            .A(_89_),
            .B(_797_),
            .C(_88_),
            .Y(_90_)
        );
        
        NAND3X1 _1711_ (
            .A(_849_),
            .B(_853_),
            .C(_836_),
            .Y(_91_)
        );
        
        OAI21X1 _1712_ (
            .A(_91_),
            .B(_90_),
            .C(_84_),
            .Y(_92_)
        );
        
        OAI21X1 _1713_ (
            .A(_87_),
            .B(_92_),
            .C(_191_),
            .Y(_93_)
        );
        
        OR2X2 _1714_ (
            .A(_93_),
            .B(_86_),
            .Y(_94_)
        );
        
        AOI22X1 _1715_ (
            .A(_129_),
            .B(_188__bF$buf1),
            .C(_94_),
            .D(_709_),
            .Y(_71_)
        );
        
        NAND2X1 _1716_ (
            .A(Ycalc[11]),
            .B(_188__bF$buf0),
            .Y(_95_)
        );
        
        INVX1 _1717_ (
            .A(_81_),
            .Y(_96_)
        );
        
        OAI21X1 _1718_ (
            .A(_858_),
            .B(_76_),
            .C(_201__bF$buf1),
            .Y(_97_)
        );
        
        NAND2X1 _1719_ (
            .A(_475_),
            .B(_97_),
            .Y(_98_)
        );
        
        OR2X2 _1720_ (
            .A(_97_),
            .B(_475_),
            .Y(_99_)
        );
        
        NAND2X1 _1721_ (
            .A(_98_),
            .B(_99_),
            .Y(_100_)
        );
        
        INVX1 _1722_ (
            .A(_100_),
            .Y(_101_)
        );
        
        NOR3X1 _1723_ (
            .A(_96_),
            .B(_101_),
            .C(_86_),
            .Y(_102_)
        );
        
        AOI21X1 _1724_ (
            .A(_92_),
            .B(_87_),
            .C(_96_),
            .Y(_103_)
        );
        
        OAI21X1 _1725_ (
            .A(_100_),
            .B(_103_),
            .C(_191_),
            .Y(_104_)
        );
        
        OAI21X1 _1726_ (
            .A(_102_),
            .B(_104_),
            .C(_709_),
            .Y(_105_)
        );
        
        NAND2X1 _1727_ (
            .A(_95_),
            .B(_105_),
            .Y(_72_)
        );
        
        DFFPOSX1 _1728_ (
            .CLK(clk_bF$buf7),
            .D(_0_),
            .Q(Ycalc[0])
        );
        
        DFFPOSX1 _1729_ (
            .CLK(clk_bF$buf6),
            .D(_1_),
            .Q(Ycalc[1])
        );
        
        DFFPOSX1 _1730_ (
            .CLK(clk_bF$buf5),
            .D(_2_),
            .Q(Xcalc[0])
        );
        
        DFFPOSX1 _1731_ (
            .CLK(clk_bF$buf4),
            .D(_3_),
            .Q(Xcalc[1])
        );
        
        DFFPOSX1 _1732_ (
            .CLK(clk_bF$buf3),
            .D(_4_),
            .Q(Xcalc[2])
        );
        
        DFFPOSX1 _1733_ (
            .CLK(clk_bF$buf2),
            .D(_5_),
            .Q(Xcalc[3])
        );
        
        DFFPOSX1 _1734_ (
            .CLK(clk_bF$buf1),
            .D(_6_),
            .Q(Xcalc[4])
        );
        
        DFFPOSX1 _1735_ (
            .CLK(clk_bF$buf0),
            .D(_7_),
            .Q(Xcalc[5])
        );
        
        DFFPOSX1 _1736_ (
            .CLK(clk_bF$buf7),
            .D(_8_),
            .Q(Xcalc[6])
        );
        
        DFFPOSX1 _1737_ (
            .CLK(clk_bF$buf6),
            .D(_9_),
            .Q(Xcalc[7])
        );
        
        DFFPOSX1 _1738_ (
            .CLK(clk_bF$buf5),
            .D(_10_),
            .Q(Xcalc[8])
        );
        
        DFFPOSX1 _1739_ (
            .CLK(clk_bF$buf4),
            .D(_11_),
            .Q(Xcalc[9])
        );
        
        DFFPOSX1 _1740_ (
            .CLK(clk_bF$buf3),
            .D(_12_),
            .Q(Xcalc[10])
        );
        
        DFFPOSX1 _1741_ (
            .CLK(clk_bF$buf2),
            .D(_13_),
            .Q(Xcalc[11])
        );
        
        DFFPOSX1 _1742_ (
            .CLK(clk_bF$buf1),
            .D(_14_),
            .Q(Acalc[0])
        );
        
        DFFPOSX1 _1743_ (
            .CLK(clk_bF$buf0),
            .D(_15_),
            .Q(Acalc[1])
        );
        
        DFFPOSX1 _1744_ (
            .CLK(clk_bF$buf7),
            .D(_16_),
            .Q(Acalc[2])
        );
        
        DFFPOSX1 _1745_ (
            .CLK(clk_bF$buf6),
            .D(_17_),
            .Q(Acalc[3])
        );
        
        DFFPOSX1 _1746_ (
            .CLK(clk_bF$buf5),
            .D(_18_),
            .Q(Acalc[4])
        );
        
        DFFPOSX1 _1747_ (
            .CLK(clk_bF$buf4),
            .D(_19_),
            .Q(Acalc[5])
        );
        
        DFFPOSX1 _1748_ (
            .CLK(clk_bF$buf3),
            .D(_20_),
            .Q(Acalc[6])
        );
        
        DFFPOSX1 _1749_ (
            .CLK(clk_bF$buf2),
            .D(_21_),
            .Q(Acalc[7])
        );
        
        DFFPOSX1 _1750_ (
            .CLK(clk_bF$buf1),
            .D(_22_),
            .Q(Acalc[8])
        );
        
        DFFPOSX1 _1751_ (
            .CLK(clk_bF$buf0),
            .D(_23_),
            .Q(Acalc[9])
        );
        
        DFFPOSX1 _1752_ (
            .CLK(clk_bF$buf7),
            .D(_24_),
            .Q(Acalc[10])
        );
        
        DFFPOSX1 _1753_ (
            .CLK(clk_bF$buf6),
            .D(_25_),
            .Q(Acalc[11])
        );
        
        DFFPOSX1 _1754_ (
            .CLK(clk_bF$buf5),
            .D(_26_),
            .Q(Xin12b[10])
        );
        
        DFFPOSX1 _1755_ (
            .CLK(clk_bF$buf4),
            .D(_27_),
            .Q(Xin12b[11])
        );
        
        DFFPOSX1 _1756_ (
            .CLK(clk_bF$buf3),
            .D(_28_),
            .Q(Xin12b[8])
        );
        
        DFFPOSX1 _1757_ (
            .CLK(clk_bF$buf2),
            .D(_29_),
            .Q(Xin12b[9])
        );
        
        DFFPOSX1 _1758_ (
            .CLK(clk_bF$buf1),
            .D(_30_),
            .Q(Xin12b[6])
        );
        
        DFFPOSX1 _1759_ (
            .CLK(clk_bF$buf0),
            .D(_31_),
            .Q(Xin12b[7])
        );
        
        DFFPOSX1 _1760_ (
            .CLK(clk_bF$buf7),
            .D(_32_),
            .Q(Xin12b[4])
        );
        
        DFFPOSX1 _1761_ (
            .CLK(clk_bF$buf6),
            .D(_33_),
            .Q(Xin12b[5])
        );
        
        DFFPOSX1 _1762_ (
            .CLK(clk_bF$buf5),
            .D(_34_),
            .Q(Xin1[0])
        );
        
        DFFPOSX1 _1763_ (
            .CLK(clk_bF$buf4),
            .D(_35_),
            .Q(Xin1[1])
        );
        
        DFFPOSX1 _1764_ (
            .CLK(clk_bF$buf3),
            .D(_36_),
            .Q(Xin0[0])
        );
        
        DFFPOSX1 _1765_ (
            .CLK(clk_bF$buf2),
            .D(_37_),
            .Q(Xin0[1])
        );
        
        DFFPOSX1 _1766_ (
            .CLK(clk_bF$buf1),
            .D(_38_),
            .Q(Yin12b[10])
        );
        
        DFFPOSX1 _1767_ (
            .CLK(clk_bF$buf0),
            .D(_39_),
            .Q(Yin12b[11])
        );
        
        DFFPOSX1 _1768_ (
            .CLK(clk_bF$buf7),
            .D(_40_),
            .Q(Yin12b[8])
        );
        
        DFFPOSX1 _1769_ (
            .CLK(clk_bF$buf6),
            .D(_41_),
            .Q(Yin12b[9])
        );
        
        DFFPOSX1 _1770_ (
            .CLK(clk_bF$buf5),
            .D(_42_),
            .Q(Yin12b[6])
        );
        
        DFFPOSX1 _1771_ (
            .CLK(clk_bF$buf4),
            .D(_43_),
            .Q(Yin12b[7])
        );
        
        DFFPOSX1 _1772_ (
            .CLK(clk_bF$buf3),
            .D(_44_),
            .Q(Yin12b[4])
        );
        
        DFFPOSX1 _1773_ (
            .CLK(clk_bF$buf2),
            .D(_45_),
            .Q(Yin12b[5])
        );
        
        DFFPOSX1 _1774_ (
            .CLK(clk_bF$buf1),
            .D(_46_),
            .Q(Yin1[0])
        );
        
        DFFPOSX1 _1775_ (
            .CLK(clk_bF$buf0),
            .D(_47_),
            .Q(Yin1[1])
        );
        
        DFFPOSX1 _1776_ (
            .CLK(clk_bF$buf7),
            .D(_48_),
            .Q(Yin0[0])
        );
        
        DFFPOSX1 _1777_ (
            .CLK(clk_bF$buf6),
            .D(_49_),
            .Q(Yin0[1])
        );
        
        DFFPOSX1 _1778_ (
            .CLK(clk_bF$buf5),
            .D(_50_),
            .Q(Ain12b[10])
        );
        
        DFFPOSX1 _1779_ (
            .CLK(clk_bF$buf4),
            .D(_51_),
            .Q(Ain12b[11])
        );
        
        DFFPOSX1 _1780_ (
            .CLK(clk_bF$buf3),
            .D(_52_),
            .Q(Ain12b[8])
        );
        
        DFFPOSX1 _1781_ (
            .CLK(clk_bF$buf2),
            .D(_53_),
            .Q(Ain12b[9])
        );
        
        DFFPOSX1 _1782_ (
            .CLK(clk_bF$buf1),
            .D(_54_),
            .Q(Ain12b[6])
        );
        
        DFFPOSX1 _1783_ (
            .CLK(clk_bF$buf0),
            .D(_55_),
            .Q(Ain12b[7])
        );
        
        DFFPOSX1 _1784_ (
            .CLK(clk_bF$buf7),
            .D(_56_),
            .Q(Ain12b[4])
        );
        
        DFFPOSX1 _1785_ (
            .CLK(clk_bF$buf6),
            .D(_57_),
            .Q(Ain12b[5])
        );
        
        DFFPOSX1 _1786_ (
            .CLK(clk_bF$buf5),
            .D(_58_),
            .Q(Ain1[0])
        );
        
        DFFPOSX1 _1787_ (
            .CLK(clk_bF$buf4),
            .D(_59_),
            .Q(Ain1[1])
        );
        
        DFFPOSX1 _1788_ (
            .CLK(clk_bF$buf3),
            .D(_60_),
            .Q(Ain0[0])
        );
        
        DFFPOSX1 _1789_ (
            .CLK(clk_bF$buf2),
            .D(_61_),
            .Q(Ain0[1])
        );
        
        DFFPOSX1 _1790_ (
            .CLK(clk_bF$buf1),
            .D(Rdy),
            .Q(LoadCtl[0])
        );
        
        DFFPOSX1 _1791_ (
            .CLK(clk_bF$buf0),
            .D(LoadCtl_0_bF$buf1),
            .Q(LoadCtl[1])
        );
        
        DFFPOSX1 _1792_ (
            .CLK(clk_bF$buf7),
            .D(LoadCtl[1]),
            .Q(LoadCtl[2])
        );
        
        DFFPOSX1 _1793_ (
            .CLK(clk_bF$buf6),
            .D(LoadCtl[2]),
            .Q(LoadCtl[3])
        );
        
        DFFPOSX1 _1794_ (
            .CLK(clk_bF$buf5),
            .D(LoadCtl[3]),
            .Q(LoadCtl[4])
        );
        
        DFFPOSX1 _1795_ (
            .CLK(clk_bF$buf4),
            .D(LoadCtl[4]),
            .Q(LoadCtl[5])
        );
        
        DFFPOSX1 _1796_ (
            .CLK(clk_bF$buf3),
            .D(LoadCtl[5]),
            .Q(LoadCtl[6])
        );
        
        DFFPOSX1 _1797_ (
            .CLK(clk_bF$buf2),
            .D(_62_),
            .Q(_860_)
        );
        
        DFFPOSX1 _1798_ (
            .CLK(clk_bF$buf1),
            .D(_63_),
            .Q(Ycalc[2])
        );
        
        DFFPOSX1 _1799_ (
            .CLK(clk_bF$buf0),
            .D(_64_),
            .Q(Ycalc[3])
        );
        
        DFFPOSX1 _1800_ (
            .CLK(clk_bF$buf7),
            .D(_65_),
            .Q(Ycalc[4])
        );
        
        DFFPOSX1 _1801_ (
            .CLK(clk_bF$buf6),
            .D(_66_),
            .Q(Ycalc[5])
        );
        
        DFFPOSX1 _1802_ (
            .CLK(clk_bF$buf5),
            .D(_67_),
            .Q(Ycalc[6])
        );
        
        DFFPOSX1 _1803_ (
            .CLK(clk_bF$buf4),
            .D(_68_),
            .Q(Ycalc[7])
        );
        
        DFFPOSX1 _1804_ (
            .CLK(clk_bF$buf3),
            .D(_69_),
            .Q(Ycalc[8])
        );
        
        DFFPOSX1 _1805_ (
            .CLK(clk_bF$buf2),
            .D(_70_),
            .Q(Ycalc[9])
        );
        
        DFFPOSX1 _1806_ (
            .CLK(clk_bF$buf1),
            .D(_71_),
            .Q(Ycalc[10])
        );
        
        DFFPOSX1 _1807_ (
            .CLK(clk_bF$buf0),
            .D(_72_),
            .Q(Ycalc[11])
        );
        
        BUFX2 _1808_ (
            .A(_859_[0]),
            .Y(Aout[0])
        );
        
        BUFX2 _1809_ (
            .A(_859_[1]),
            .Y(Aout[1])
        );
        
        BUFX2 _1810_ (
            .A(_860_),
            .Y(ISout)
        );
        
        BUFX2 _1811_ (
            .A(LoadCtl_6_bF$buf2),
            .Y(Vld)
        );
        
        BUFX2 _1812_ (
            .A(_861_[0]),
            .Y(Xout[0])
        );
        
        BUFX2 _1813_ (
            .A(_861_[1]),
            .Y(Xout[1])
        );
        
        BUFX2 _1814_ (
            .A(_862_[0]),
            .Y(Yout[0])
        );
        
        BUFX2 _1815_ (
            .A(_862_[1]),
            .Y(Yout[1])
        );
        
        INVX1 _863_ (
            .A(Acalc[10]),
            .Y(_106_)
        );
        
        NAND2X1 _864_ (
            .A(LoadCtl[4]),
            .B(Acalc[8]),
            .Y(_107_)
        );
        
        OAI21X1 _865_ (
            .A(LoadCtl[4]),
            .B(_106_),
            .C(_107_),
            .Y(_108_)
        );
        
        NOR2X1 _866_ (
            .A(LoadCtl[3]),
            .B(LoadCtl[2]),
            .Y(_109_)
        );
        
        INVX1 _867_ (
            .A(Acalc[6]),
            .Y(_110_)
        );
        
        NAND2X1 _868_ (
            .A(LoadCtl[2]),
            .B(Acalc[4]),
            .Y(_111_)
        );
        
        INVX2 _869_ (
            .A(LoadCtl[2]),
            .Y(_112_)
        );
        
        NAND2X1 _870_ (
            .A(LoadCtl[3]),
            .B(_112_),
            .Y(_113_)
        );
        
        OAI21X1 _871_ (
            .A(_110_),
            .B(_113_),
            .C(_111_),
            .Y(_114_)
        );
        
        AOI21X1 _872_ (
            .A(_108_),
            .B(_109_),
            .C(_114_),
            .Y(_115_)
        );
        
        NOR2X1 _873_ (
            .A(LoadCtl_0_bF$buf0),
            .B(LoadCtl[1]),
            .Y(_116_)
        );
        
        INVX2 _874_ (
            .A(_116_),
            .Y(_117_)
        );
        
        INVX1 _875_ (
            .A(LoadCtl[1]),
            .Y(_118_)
        );
        
        NOR2X1 _876_ (
            .A(LoadCtl_0_bF$buf3),
            .B(_118_),
            .Y(_119_)
        );
        
        AOI22X1 _877_ (
            .A(LoadCtl_0_bF$buf2),
            .B(Acalc[0]),
            .C(_119_),
            .D(Acalc[2]),
            .Y(_120_)
        );
        
        OAI21X1 _878_ (
            .A(_117_),
            .B(_115_),
            .C(_120_),
            .Y(_859_[0])
        );
        
        INVX1 _879_ (
            .A(Acalc[11]),
            .Y(_121_)
        );
        
        NAND2X1 _880_ (
            .A(LoadCtl[4]),
            .B(Acalc[9]),
            .Y(_122_)
        );
        
        OAI21X1 _881_ (
            .A(LoadCtl[4]),
            .B(_121_),
            .C(_122_),
            .Y(_123_)
        );
        
        INVX1 _882_ (
            .A(Acalc[7]),
            .Y(_124_)
        );
        
        NAND2X1 _883_ (
            .A(LoadCtl[2]),
            .B(Acalc[5]),
            .Y(_125_)
        );
        
        OAI21X1 _884_ (
            .A(_124_),
            .B(_113_),
            .C(_125_),
            .Y(_126_)
        );
        
        AOI21X1 _885_ (
            .A(_109_),
            .B(_123_),
            .C(_126_),
            .Y(_127_)
        );
        
        AOI22X1 _886_ (
            .A(LoadCtl_0_bF$buf1),
            .B(Acalc[1]),
            .C(_119_),
            .D(Acalc[3]),
            .Y(_128_)
        );
        
        OAI21X1 _887_ (
            .A(_117_),
            .B(_127_),
            .C(_128_),
            .Y(_859_[1])
        );
        
        INVX1 _888_ (
            .A(Ycalc[10]),
            .Y(_129_)
        );
        
        NAND2X1 _889_ (
            .A(LoadCtl[4]),
            .B(Ycalc[8]),
            .Y(_130_)
        );
        
        OAI21X1 _890_ (
            .A(LoadCtl[4]),
            .B(_129_),
            .C(_130_),
            .Y(_131_)
        );
        
        INVX1 _891_ (
            .A(Ycalc[6]),
            .Y(_132_)
        );
        
        INVX1 _892_ (
            .A(Ycalc[4]),
            .Y(_133_)
        );
        
        OAI22X1 _893_ (
            .A(_112_),
            .B(_133_),
            .C(_132_),
            .D(_113_),
            .Y(_134_)
        );
        
        AOI21X1 _894_ (
            .A(_109_),
            .B(_131_),
            .C(_134_),
            .Y(_135_)
        );
        
        AOI22X1 _895_ (
            .A(LoadCtl_0_bF$buf0),
            .B(Ycalc[0]),
            .C(_119_),
            .D(Ycalc[2]),
            .Y(_136_)
        );
        
        OAI21X1 _896_ (
            .A(_117_),
            .B(_135_),
            .C(_136_),
            .Y(_862_[0])
        );
        
        INVX1 _897_ (
            .A(LoadCtl[4]),
            .Y(_137_)
        );
        
        INVX1 _898_ (
            .A(Ycalc[9]),
            .Y(_138_)
        );
        
        NAND2X1 _899_ (
            .A(Ycalc[11]),
            .B(_137_),
            .Y(_139_)
        );
        
        OAI21X1 _900_ (
            .A(_137_),
            .B(_138_),
            .C(_139_),
            .Y(_140_)
        );
        
        INVX1 _901_ (
            .A(Ycalc[7]),
            .Y(_141_)
        );
        
        INVX1 _902_ (
            .A(Ycalc[5]),
            .Y(_142_)
        );
        
        OAI22X1 _903_ (
            .A(_112_),
            .B(_142_),
            .C(_141_),
            .D(_113_),
            .Y(_143_)
        );
        
        AOI21X1 _904_ (
            .A(_109_),
            .B(_140_),
            .C(_143_),
            .Y(_144_)
        );
        
        AOI22X1 _905_ (
            .A(LoadCtl_0_bF$buf3),
            .B(Ycalc[1]),
            .C(_119_),
            .D(Ycalc[3]),
            .Y(_145_)
        );
        
        OAI21X1 _906_ (
            .A(_117_),
            .B(_144_),
            .C(_145_),
            .Y(_862_[1])
        );
        
        INVX1 _907_ (
            .A(Xcalc[10]),
            .Y(_146_)
        );
        
        NAND2X1 _908_ (
            .A(LoadCtl[4]),
            .B(Xcalc[8]),
            .Y(_147_)
        );
        
        OAI21X1 _909_ (
            .A(LoadCtl[4]),
            .B(_146_),
            .C(_147_),
            .Y(_148_)
        );
        
        INVX1 _910_ (
            .A(Xcalc[6]),
            .Y(_149_)
        );
        
        INVX1 _911_ (
            .A(Xcalc[4]),
            .Y(_150_)
        );
        
        OAI22X1 _912_ (
            .A(_112_),
            .B(_150_),
            .C(_149_),
            .D(_113_),
            .Y(_151_)
        );
        
        AOI21X1 _913_ (
            .A(_109_),
            .B(_148_),
            .C(_151_),
            .Y(_152_)
        );
        
        AOI22X1 _914_ (
            .A(LoadCtl_0_bF$buf2),
            .B(Xcalc[0]),
            .C(_119_),
            .D(Xcalc[2]),
            .Y(_153_)
        );
        
        OAI21X1 _915_ (
            .A(_117_),
            .B(_152_),
            .C(_153_),
            .Y(_861_[0])
        );
        
        INVX1 _916_ (
            .A(Xcalc[11]),
            .Y(_154_)
        );
        
        NAND2X1 _917_ (
            .A(LoadCtl[4]),
            .B(Xcalc[9]),
            .Y(_155_)
        );
        
        OAI21X1 _918_ (
            .A(LoadCtl[4]),
            .B(_154_),
            .C(_155_),
            .Y(_156_)
        );
        
        INVX1 _919_ (
            .A(Xcalc[7]),
            .Y(_157_)
        );
        
        INVX1 _920_ (
            .A(Xcalc[5]),
            .Y(_158_)
        );
        
        OAI22X1 _921_ (
            .A(_112_),
            .B(_158_),
            .C(_157_),
            .D(_113_),
            .Y(_159_)
        );
        
        AOI21X1 _922_ (
            .A(_109_),
            .B(_156_),
            .C(_159_),
            .Y(_160_)
        );
        
        AOI22X1 _923_ (
            .A(LoadCtl_0_bF$buf1),
            .B(Xcalc[1]),
            .C(_119_),
            .D(Xcalc[3]),
            .Y(_161_)
        );
        
        OAI21X1 _924_ (
            .A(_117_),
            .B(_160_),
            .C(_161_),
            .Y(_861_[1])
        );
        
        INVX1 _925_ (
            .A(Ycalc[0]),
            .Y(_162_)
        );
        
        INVX1 _926_ (
            .A(Yin0[0]),
            .Y(_163_)
        );
        
        INVX8 _927_ (
            .A(Stg_1_bF$buf3),
            .Y(_164_)
        );
        
        INVX1 _928_ (
            .A(Xin1[0]),
            .Y(_165_)
        );
        
        NAND2X1 _929_ (
            .A(Stg_0_bF$buf4),
            .B(Xin1[1]),
            .Y(_166_)
        );
        
        OAI21X1 _930_ (
            .A(Stg_0_bF$buf3),
            .B(_165_),
            .C(_166_),
            .Y(_167_)
        );
        
        INVX1 _931_ (
            .A(Xin0[0]),
            .Y(_168_)
        );
        
        NAND2X1 _932_ (
            .A(Xin0[1]),
            .B(Stg_0_bF$buf2),
            .Y(_169_)
        );
        
        OAI21X1 _933_ (
            .A(Stg_0_bF$buf1),
            .B(_168_),
            .C(_169_),
            .Y(_170_)
        );
        
        MUX2X1 _934_ (
            .A(_170_),
            .B(_167_),
            .S(_164__bF$buf0),
            .Y(_171_)
        );
        
        INVX1 _935_ (
            .A(Xin12b[6]),
            .Y(_172_)
        );
        
        NAND2X1 _936_ (
            .A(Stg_0_bF$buf0),
            .B(Xin12b[7]),
            .Y(_173_)
        );
        
        OAI21X1 _937_ (
            .A(Stg_0_bF$buf6),
            .B(_172_),
            .C(_173_),
            .Y(_174_)
        );
        
        INVX1 _938_ (
            .A(Xin12b[4]),
            .Y(_175_)
        );
        
        NAND2X1 _939_ (
            .A(Stg_0_bF$buf5),
            .B(Xin12b[5]),
            .Y(_176_)
        );
        
        OAI21X1 _940_ (
            .A(Stg_0_bF$buf4),
            .B(_175_),
            .C(_176_),
            .Y(_177_)
        );
        
        MUX2X1 _941_ (
            .A(_177_),
            .B(_174_),
            .S(_164__bF$buf4),
            .Y(_178_)
        );
        
        MUX2X1 _942_ (
            .A(_178_),
            .B(_171_),
            .S(Stg_2_bF$buf0),
            .Y(_179_)
        );
        
        NOR2X1 _943_ (
            .A(_163_),
            .B(_179_),
            .Y(_180_)
        );
        
        NAND2X1 _944_ (
            .A(_163_),
            .B(_179_),
            .Y(_181_)
        );
        
        INVX1 _945_ (
            .A(_181_),
            .Y(_182_)
        );
        
        INVX4 _946_ (
            .A(Stg_2_bF$buf4),
            .Y(_183_)
        );
        
        NAND2X1 _947_ (
            .A(_183__bF$buf3),
            .B(_164__bF$buf3),
            .Y(_184_)
        );
        
        OAI21X1 _948_ (
            .A(Stg_0_bF$buf3),
            .B(_184_),
            .C(LoadCtl_6_bF$buf1),
            .Y(_185_)
        );
        
        INVX2 _949_ (
            .A(_185_),
            .Y(_186_)
        );
        
        OAI21X1 _950_ (
            .A(_180_),
            .B(_182_),
            .C(_186_),
            .Y(_187_)
        );
        
        OAI21X1 _951_ (
            .A(_162_),
            .B(LoadCtl_6_bF$buf0),
            .C(_187_),
            .Y(_0_)
        );
        
        INVX8 _952_ (
            .A(LoadCtl_6_bF$buf4),
            .Y(_188_)
        );
        
        NAND2X1 _953_ (
            .A(Ycalc[1]),
            .B(_188__bF$buf4),
            .Y(_189_)
        );
        
        NOR2X1 _954_ (
            .A(Stg_0_bF$buf2),
            .B(Stg_1_bF$buf2),
            .Y(_190_)
        );
        
        NAND2X1 _955_ (
            .A(_183__bF$buf2),
            .B(_190_),
            .Y(_191_)
        );
        
        INVX2 _956_ (
            .A(_191_),
            .Y(_192_)
        );
        
        MUX2X1 _957_ (
            .A(Xin1[1]),
            .B(Xin1[0]),
            .S(Stg_0_bF$buf1),
            .Y(_193_)
        );
        
        MUX2X1 _958_ (
            .A(Xin0[1]),
            .B(Xin0[0]),
            .S(Stg_0_bF$buf0),
            .Y(_194_)
        );
        
        MUX2X1 _959_ (
            .A(_194_),
            .B(_193_),
            .S(_164__bF$buf2),
            .Y(_195_)
        );
        
        MUX2X1 _960_ (
            .A(Xin12b[7]),
            .B(Xin12b[6]),
            .S(Stg_0_bF$buf6),
            .Y(_196_)
        );
        
        MUX2X1 _961_ (
            .A(Xin12b[5]),
            .B(Xin12b[4]),
            .S(Stg_0_bF$buf5),
            .Y(_197_)
        );
        
        MUX2X1 _962_ (
            .A(_197_),
            .B(_196_),
            .S(_164__bF$buf1),
            .Y(_198_)
        );
        
        MUX2X1 _963_ (
            .A(_198_),
            .B(_195_),
            .S(Stg_2_bF$buf3),
            .Y(_199_)
        );
        
        INVX1 _964_ (
            .A(Yin0[1]),
            .Y(_200_)
        );
        
        INVX8 _965_ (
            .A(Ain12b_11_bF$buf1),
            .Y(_201_)
        );
        
        INVX1 _966_ (
            .A(Xin1[1]),
            .Y(_202_)
        );
        
        NAND2X1 _967_ (
            .A(Stg_0_bF$buf4),
            .B(Xin12b[4]),
            .Y(_203_)
        );
        
        OAI21X1 _968_ (
            .A(Stg_0_bF$buf3),
            .B(_202_),
            .C(_203_),
            .Y(_204_)
        );
        
        INVX1 _969_ (
            .A(Xin0[1]),
            .Y(_205_)
        );
        
        NAND2X1 _970_ (
            .A(Stg_0_bF$buf2),
            .B(Xin1[0]),
            .Y(_206_)
        );
        
        OAI21X1 _971_ (
            .A(Stg_0_bF$buf1),
            .B(_205_),
            .C(_206_),
            .Y(_207_)
        );
        
        MUX2X1 _972_ (
            .A(_207_),
            .B(_204_),
            .S(_164__bF$buf0),
            .Y(_208_)
        );
        
        INVX1 _973_ (
            .A(Xin12b[7]),
            .Y(_209_)
        );
        
        NAND2X1 _974_ (
            .A(Stg_0_bF$buf0),
            .B(Xin12b[8]),
            .Y(_210_)
        );
        
        OAI21X1 _975_ (
            .A(Stg_0_bF$buf6),
            .B(_209_),
            .C(_210_),
            .Y(_211_)
        );
        
        INVX1 _976_ (
            .A(Xin12b[5]),
            .Y(_212_)
        );
        
        NAND2X1 _977_ (
            .A(Stg_0_bF$buf5),
            .B(Xin12b[6]),
            .Y(_213_)
        );
        
        OAI21X1 _978_ (
            .A(Stg_0_bF$buf4),
            .B(_212_),
            .C(_213_),
            .Y(_214_)
        );
        
        MUX2X1 _979_ (
            .A(_214_),
            .B(_211_),
            .S(_164__bF$buf4),
            .Y(_215_)
        );
        
        MUX2X1 _980_ (
            .A(_215_),
            .B(_208_),
            .S(Stg_2_bF$buf2),
            .Y(_216_)
        );
        
        NAND3X1 _981_ (
            .A(_201__bF$buf0),
            .B(_179_),
            .C(_216_),
            .Y(_217_)
        );
        
        MUX2X1 _982_ (
            .A(Xin12b[4]),
            .B(Xin1[1]),
            .S(Stg_0_bF$buf3),
            .Y(_218_)
        );
        
        MUX2X1 _983_ (
            .A(Xin1[0]),
            .B(Xin0[1]),
            .S(Stg_0_bF$buf2),
            .Y(_219_)
        );
        
        MUX2X1 _984_ (
            .A(_219_),
            .B(_218_),
            .S(_164__bF$buf3),
            .Y(_220_)
        );
        
        MUX2X1 _985_ (
            .A(Xin12b[8]),
            .B(Xin12b[7]),
            .S(Stg_0_bF$buf1),
            .Y(_221_)
        );
        
        MUX2X1 _986_ (
            .A(Xin12b[6]),
            .B(Xin12b[5]),
            .S(Stg_0_bF$buf0),
            .Y(_222_)
        );
        
        MUX2X1 _987_ (
            .A(_222_),
            .B(_221_),
            .S(_164__bF$buf2),
            .Y(_223_)
        );
        
        MUX2X1 _988_ (
            .A(_223_),
            .B(_220_),
            .S(Stg_2_bF$buf1),
            .Y(_224_)
        );
        
        OAI21X1 _989_ (
            .A(Ain12b_11_bF$buf0),
            .B(_199_),
            .C(_224_),
            .Y(_225_)
        );
        
        AOI21X1 _990_ (
            .A(_225_),
            .B(_217_),
            .C(_200_),
            .Y(_226_)
        );
        
        INVX1 _991_ (
            .A(_226_),
            .Y(_227_)
        );
        
        NAND3X1 _992_ (
            .A(_200_),
            .B(_217_),
            .C(_225_),
            .Y(_228_)
        );
        
        AND2X2 _993_ (
            .A(_227_),
            .B(_228_),
            .Y(_229_)
        );
        
        OAI21X1 _994_ (
            .A(Yin0[0]),
            .B(_199_),
            .C(_229_),
            .Y(_230_)
        );
        
        OR2X2 _995_ (
            .A(_229_),
            .B(_181_),
            .Y(_231_)
        );
        
        AOI21X1 _996_ (
            .A(_231_),
            .B(_230_),
            .C(_192_),
            .Y(_232_)
        );
        
        OAI21X1 _997_ (
            .A(_188__bF$buf3),
            .B(_232_),
            .C(_189_),
            .Y(_1_)
        );
        
        NAND2X1 _998_ (
            .A(Xcalc[0]),
            .B(_188__bF$buf2),
            .Y(_233_)
        );
        
        INVX1 _999_ (
            .A(Yin1[0]),
            .Y(_234_)
        );
        
        endmodule
        
