magic
tech scmos
magscale 1 2
timestamp 1740695740
<< metal1 >>
rect -62 4818 -2 5058
rect 5050 5042 5142 5058
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 3577 4737 3593 4743
rect 3577 4663 3583 4737
rect 3577 4657 3593 4663
rect 5082 4578 5142 5042
rect 5050 4562 5142 4578
rect 1607 4497 1633 4503
rect 2087 4477 2233 4483
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 3407 4177 3553 4183
rect 5082 4098 5142 4562
rect 5050 4082 5142 4098
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 5082 3618 5142 4082
rect 5050 3602 5142 3618
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 5082 3138 5142 3602
rect 5050 3122 5142 3138
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 1087 2717 1253 2723
rect 5082 2658 5142 3122
rect 5050 2642 5142 2658
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 4087 2317 4193 2323
rect 5082 2178 5142 2642
rect 5050 2162 5142 2178
rect 2867 2037 2933 2043
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 1427 1837 1573 1843
rect 5082 1698 5142 2162
rect 5050 1682 5142 1698
rect 2547 1597 2753 1603
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 5082 1218 5142 1682
rect 5050 1202 5142 1218
rect -62 962 30 978
rect -62 498 -2 962
rect 5082 738 5142 1202
rect 5050 722 5142 738
rect 1467 657 1533 663
rect -62 482 30 498
rect -62 18 -2 482
rect 5082 258 5142 722
rect 5050 242 5142 258
rect -62 2 30 18
rect 5082 2 5142 242
<< m2contact >>
rect 3593 4733 3607 4747
rect 3593 4653 3607 4667
rect 1593 4493 1607 4507
rect 1633 4493 1647 4507
rect 2073 4473 2087 4487
rect 2233 4473 2247 4487
rect 3393 4173 3407 4187
rect 3553 4173 3567 4187
rect 1073 2713 1087 2727
rect 1253 2713 1267 2727
rect 4073 2313 4087 2327
rect 4193 2313 4207 2327
rect 2853 2033 2867 2047
rect 2933 2033 2947 2047
rect 1413 1833 1427 1847
rect 1573 1833 1587 1847
rect 2533 1593 2547 1607
rect 2753 1593 2767 1607
rect 1453 653 1467 667
rect 1533 653 1547 667
<< metal2 >>
rect 3476 5096 3503 5103
rect 556 4956 583 4963
rect 536 4907 543 4943
rect 576 4927 583 4956
rect 696 4963 703 4973
rect 676 4956 703 4963
rect 576 4903 583 4913
rect 576 4896 603 4903
rect 236 4676 243 4893
rect 516 4696 523 4713
rect 276 4676 303 4683
rect 236 4447 243 4463
rect 296 4247 303 4676
rect 536 4623 543 4683
rect 556 4647 563 4703
rect 576 4667 583 4683
rect 596 4667 603 4896
rect 536 4616 563 4623
rect 316 4467 323 4493
rect 256 4216 263 4233
rect 276 4047 283 4213
rect 276 3996 283 4033
rect 316 4007 323 4453
rect 436 4207 443 4473
rect 456 4456 483 4463
rect 456 4447 463 4456
rect 496 4436 503 4473
rect 516 4456 523 4473
rect 556 4443 563 4616
rect 576 4447 583 4473
rect 536 4436 563 4443
rect 536 4216 543 4233
rect 576 4207 583 4433
rect 516 4016 523 4033
rect 276 3716 283 3733
rect 256 3607 263 3703
rect 96 3516 103 3593
rect 156 3523 163 3533
rect 136 3516 163 3523
rect 96 3207 103 3223
rect 136 3167 143 3223
rect 156 3167 163 3516
rect 316 3467 323 3993
rect 536 3763 543 4033
rect 676 4003 683 4956
rect 776 4707 783 4963
rect 1076 4956 1103 4963
rect 1096 4947 1103 4956
rect 1216 4956 1223 4973
rect 1316 4963 1323 4973
rect 1296 4956 1323 4963
rect 816 4687 823 4703
rect 856 4696 863 4933
rect 736 4247 743 4493
rect 776 4427 783 4673
rect 796 4667 803 4683
rect 836 4643 843 4683
rect 1056 4667 1063 4943
rect 816 4636 843 4643
rect 816 4456 823 4636
rect 736 4203 743 4233
rect 736 4196 763 4203
rect 776 4047 783 4223
rect 816 4216 823 4413
rect 616 3996 643 4003
rect 656 3996 683 4003
rect 516 3756 543 3763
rect 516 3743 523 3756
rect 496 3736 523 3743
rect 216 3216 223 3453
rect 436 3447 443 3733
rect 496 3527 503 3736
rect 636 3687 643 3996
rect 676 3547 683 3996
rect 736 3787 743 4003
rect 836 3987 843 4443
rect 1036 4423 1043 4473
rect 1056 4456 1063 4493
rect 1096 4456 1103 4473
rect 1076 4436 1083 4453
rect 1136 4443 1143 4633
rect 1156 4607 1163 4663
rect 1416 4547 1423 4643
rect 1376 4507 1383 4513
rect 1476 4507 1483 4693
rect 1376 4476 1383 4493
rect 1476 4487 1483 4493
rect 1116 4436 1143 4443
rect 1036 4416 1063 4423
rect 996 3956 1003 3993
rect 1016 3987 1023 4213
rect 1056 3963 1063 4416
rect 1136 4223 1143 4233
rect 1116 4216 1143 4223
rect 1136 4007 1143 4216
rect 1396 4216 1403 4233
rect 1276 4027 1283 4213
rect 1247 3996 1263 4003
rect 1036 3956 1063 3963
rect 816 3727 823 3753
rect 1076 3736 1083 3773
rect 1116 3736 1123 3753
rect 616 3516 643 3523
rect 656 3516 663 3533
rect 456 3467 463 3483
rect 496 3447 503 3483
rect 76 2263 83 3053
rect 256 3023 263 3313
rect 456 3247 463 3433
rect 516 3243 523 3493
rect 496 3236 523 3243
rect 247 3016 263 3023
rect 356 3023 363 3153
rect 356 3016 383 3023
rect 96 2667 103 2743
rect 136 2723 143 2743
rect 216 2736 243 2743
rect 156 2723 163 2733
rect 136 2716 163 2723
rect 76 2256 103 2263
rect 136 2083 143 2263
rect 156 2083 163 2716
rect 236 2687 243 2736
rect 256 2707 263 3016
rect 336 2667 343 2743
rect 376 2727 383 2733
rect 256 2556 263 2653
rect 296 2556 303 2573
rect 236 2536 243 2553
rect 216 2256 243 2263
rect 236 2247 243 2256
rect 96 2076 123 2083
rect 136 2076 163 2083
rect 116 1767 123 2076
rect 156 1327 163 2076
rect 216 2007 223 2083
rect 276 2067 283 2533
rect 316 2267 323 2553
rect 216 1843 223 1993
rect 196 1836 223 1843
rect 196 1803 203 1836
rect 196 1796 223 1803
rect 236 1576 243 1783
rect 256 1596 263 1753
rect 236 1116 243 1273
rect 216 1083 223 1103
rect 216 1076 243 1083
rect 236 867 243 1076
rect 36 816 43 853
rect 76 343 83 853
rect 136 823 143 833
rect 116 816 143 823
rect 116 343 123 816
rect 236 636 243 853
rect 316 827 323 1773
rect 336 1287 343 1793
rect 356 1587 363 2053
rect 376 1327 383 2693
rect 416 1347 423 3233
rect 476 3207 483 3223
rect 636 3207 643 3516
rect 736 3307 743 3523
rect 756 3267 763 3713
rect 736 3236 743 3253
rect 656 3056 683 3063
rect 456 2736 463 2753
rect 616 2727 623 2743
rect 456 2283 463 2673
rect 536 2556 543 2653
rect 636 2587 643 3013
rect 676 3007 683 3056
rect 696 2736 703 2773
rect 716 2547 723 3213
rect 756 3207 763 3223
rect 796 3027 803 3693
rect 836 3687 843 3703
rect 1236 3687 1243 3993
rect 1276 3963 1283 4013
rect 1276 3956 1303 3963
rect 1056 3516 1063 3553
rect 896 3016 903 3493
rect 1036 3403 1043 3503
rect 1016 3396 1043 3403
rect 876 2987 883 3003
rect 836 2576 843 2953
rect 916 2947 923 2993
rect 936 2763 943 3013
rect 1016 2987 1023 3396
rect 1076 3256 1083 3293
rect 936 2756 963 2763
rect 856 2707 863 2753
rect 1036 2723 1043 2753
rect 1096 2727 1103 3253
rect 1116 3003 1123 3273
rect 1176 3263 1183 3533
rect 1196 3516 1203 3533
rect 1176 3256 1203 3263
rect 1196 3223 1203 3256
rect 1176 3207 1183 3223
rect 1196 3216 1223 3223
rect 1296 3216 1303 3693
rect 1356 3667 1363 3703
rect 1356 3527 1363 3653
rect 1456 3056 1463 3073
rect 1116 2996 1143 3003
rect 1116 2787 1123 2996
rect 1176 2807 1183 3003
rect 1176 2747 1183 2793
rect 1276 2756 1283 2773
rect 1316 2756 1323 2793
rect 1016 2716 1043 2723
rect 556 2536 583 2543
rect 456 2276 483 2283
rect 436 2107 443 2273
rect 536 2247 543 2253
rect 576 2247 583 2536
rect 856 2287 863 2693
rect 1016 2287 1023 2716
rect 1076 2543 1083 2713
rect 1116 2576 1143 2583
rect 1096 2556 1103 2573
rect 1056 2536 1083 2543
rect 1136 2527 1143 2576
rect 1176 2547 1183 2733
rect 1256 2727 1263 2743
rect 1036 2296 1063 2303
rect 1036 2263 1043 2296
rect 476 2083 483 2233
rect 756 2147 763 2253
rect 796 2247 803 2263
rect 1036 2256 1063 2263
rect 456 2076 483 2083
rect 476 1787 483 2076
rect 516 1807 523 2093
rect 796 2076 823 2083
rect 556 1787 563 1803
rect 456 1147 463 1593
rect 536 1576 543 1783
rect 676 1747 683 1783
rect 556 1596 563 1733
rect 456 1116 463 1133
rect 516 1096 523 1153
rect 576 1107 583 1333
rect 476 963 483 1093
rect 476 956 503 963
rect 276 636 283 813
rect 456 367 463 653
rect 496 607 503 956
rect 616 836 623 1313
rect 656 1167 663 1323
rect 676 1116 683 1293
rect 696 1083 703 1593
rect 716 1307 723 1783
rect 816 1647 823 2076
rect 856 1576 863 1813
rect 896 1607 903 2073
rect 896 1563 903 1593
rect 876 1556 903 1563
rect 836 1347 843 1553
rect 796 1303 803 1313
rect 776 1296 803 1303
rect 836 1127 843 1333
rect 696 1076 723 1083
rect 576 603 583 813
rect 716 747 723 1076
rect 756 823 763 833
rect 856 827 863 1333
rect 916 1303 923 2093
rect 1056 2056 1063 2256
rect 1036 1987 1043 2043
rect 1036 1667 1043 1763
rect 1036 1347 1043 1653
rect 1076 1627 1083 2043
rect 1116 1616 1143 1623
rect 1076 1583 1083 1613
rect 1076 1576 1103 1583
rect 1136 1567 1143 1616
rect 1196 1347 1203 2713
rect 1316 2503 1323 2573
rect 1396 2556 1403 2773
rect 1436 2747 1443 3023
rect 1336 2536 1363 2543
rect 1336 2527 1343 2536
rect 1316 2496 1343 2503
rect 1336 2276 1343 2496
rect 1356 2267 1363 2536
rect 1316 2107 1323 2243
rect 1316 2047 1323 2063
rect 1356 1807 1363 1973
rect 1336 1563 1343 1753
rect 1336 1556 1363 1563
rect 1396 1556 1403 1653
rect 1416 1607 1423 1833
rect 1476 1647 1483 4473
rect 1556 4003 1563 4533
rect 1576 4267 1583 4933
rect 1856 4927 1863 4943
rect 1656 4676 1683 4683
rect 1676 4647 1683 4676
rect 1596 4467 1603 4493
rect 1616 4483 1623 4533
rect 1636 4507 1643 4643
rect 1736 4627 1743 4893
rect 1896 4887 1903 4973
rect 3136 4956 3163 4963
rect 1896 4683 1903 4873
rect 1956 4687 1963 4953
rect 2356 4923 2363 4933
rect 2096 4687 2103 4923
rect 2136 4887 2143 4923
rect 2356 4916 2383 4923
rect 2616 4707 2623 4953
rect 2976 4707 2983 4923
rect 1896 4676 1923 4683
rect 1616 4476 1643 4483
rect 1696 4456 1703 4513
rect 1536 3996 1563 4003
rect 1596 4003 1603 4453
rect 1616 4147 1623 4203
rect 1596 3996 1623 4003
rect 1536 3787 1543 3996
rect 1556 3536 1563 3693
rect 1536 3467 1543 3503
rect 1536 3267 1543 3453
rect 1616 3307 1623 3996
rect 1676 3927 1683 4183
rect 1656 3716 1683 3723
rect 1676 3687 1683 3716
rect 1736 3707 1743 4613
rect 1896 4527 1903 4676
rect 2456 4676 2483 4683
rect 2516 4676 2523 4693
rect 2456 4667 2463 4676
rect 1976 4627 1983 4663
rect 2156 4643 2163 4653
rect 2196 4647 2203 4663
rect 2156 4636 2183 4643
rect 1896 4187 1903 4513
rect 1936 4476 1943 4493
rect 1956 4476 1983 4483
rect 1956 4467 1963 4476
rect 1916 4216 1923 4233
rect 1956 4227 1963 4453
rect 2076 4247 2083 4473
rect 2236 4463 2243 4473
rect 2236 4456 2263 4463
rect 2516 4456 2523 4473
rect 2556 4456 2563 4513
rect 1936 4187 1943 4203
rect 1836 3976 1843 4013
rect 1876 3976 1883 3993
rect 1856 3967 1863 3973
rect 1976 3967 1983 4233
rect 2196 4223 2203 4433
rect 2196 4216 2223 4223
rect 2116 4147 2123 4213
rect 1636 3667 1643 3683
rect 1676 3567 1683 3673
rect 1816 3496 1823 3913
rect 1876 3727 1883 3933
rect 1796 3267 1803 3483
rect 1836 3463 1843 3483
rect 1816 3456 1843 3463
rect 1576 3227 1583 3243
rect 1556 3207 1563 3223
rect 1696 3016 1703 3213
rect 1736 3003 1743 3233
rect 1676 2967 1683 3003
rect 1716 2996 1743 3003
rect 1716 2987 1723 2996
rect 1536 2687 1543 2743
rect 1576 2707 1583 2743
rect 1636 2576 1643 2673
rect 1416 1576 1423 1593
rect 896 1296 923 1303
rect 916 1087 923 1296
rect 1036 1096 1043 1313
rect 1016 867 1023 1083
rect 1116 867 1123 1333
rect 1196 1316 1203 1333
rect 1436 1307 1443 1323
rect 1216 1147 1223 1303
rect 1216 1107 1223 1133
rect 1456 1127 1463 1343
rect 1496 1336 1503 2293
rect 1116 836 1123 853
rect 736 807 743 823
rect 756 816 783 823
rect 776 636 783 733
rect 816 636 823 793
rect 956 636 963 673
rect 996 667 1003 833
rect 1096 747 1103 823
rect 1136 687 1143 823
rect 996 636 1003 653
rect 1136 627 1143 643
rect 796 607 803 623
rect 556 596 583 603
rect 476 376 483 593
rect 496 347 503 353
rect 76 336 103 343
rect 116 336 143 343
rect 216 336 243 343
rect 136 167 143 336
rect 236 187 243 336
rect 516 307 523 383
rect 1036 376 1063 383
rect 336 156 343 173
rect 516 167 523 293
rect 536 167 543 363
rect 716 176 723 193
rect 756 187 763 343
rect 796 307 803 343
rect 1016 176 1023 333
rect 1036 327 1043 376
rect 736 156 763 163
rect 1116 156 1123 293
rect 1176 167 1183 653
rect 1196 367 1203 853
rect 1216 636 1223 653
rect 1236 627 1243 873
rect 1396 856 1403 1093
rect 1256 636 1263 673
rect 1156 156 1173 163
rect 536 147 543 153
rect 756 147 763 156
rect 1276 163 1283 673
rect 1456 667 1463 1113
rect 1356 376 1383 383
rect 1376 347 1383 376
rect 1416 167 1423 373
rect 1236 147 1243 163
rect 1276 156 1303 163
rect 1476 107 1483 1133
rect 1516 1107 1523 2093
rect 1576 2056 1583 2293
rect 1596 2247 1603 2283
rect 1676 2263 1683 2553
rect 1656 2256 1683 2263
rect 1636 2047 1643 2073
rect 1676 2047 1683 2256
rect 1696 2087 1703 2273
rect 1596 1887 1603 2043
rect 1576 1816 1583 1833
rect 1616 1816 1643 1823
rect 1636 1703 1643 1816
rect 1616 1696 1643 1703
rect 1536 1307 1543 1593
rect 1616 1327 1623 1696
rect 1696 1576 1703 1613
rect 1716 1303 1723 2973
rect 1756 2727 1763 3253
rect 1796 3187 1803 3223
rect 1816 3187 1823 3456
rect 1876 3223 1883 3713
rect 1936 3487 1943 3703
rect 1956 3687 1963 3723
rect 1856 3216 1883 3223
rect 2016 3207 2023 3223
rect 2036 3067 2043 3693
rect 1776 1847 1783 2953
rect 1816 2767 1823 2993
rect 1856 2743 1863 3013
rect 1856 2736 1883 2743
rect 1876 2547 1883 2736
rect 1896 2587 1903 2723
rect 1916 2536 1923 2573
rect 1936 2556 1943 2593
rect 1956 2583 1963 3053
rect 2036 3036 2043 3053
rect 1956 2576 1983 2583
rect 1976 2567 1983 2576
rect 1796 2103 1803 2233
rect 1796 2096 1823 2103
rect 1796 1887 1803 2096
rect 1856 2063 1863 2313
rect 1916 2296 1923 2313
rect 2056 2287 2063 3953
rect 2096 3216 2103 4013
rect 2116 3963 2123 4133
rect 2216 4027 2223 4216
rect 2316 4207 2323 4413
rect 2576 4247 2583 4443
rect 2416 4187 2423 4213
rect 2436 4183 2443 4233
rect 2496 4216 2503 4233
rect 2436 4176 2463 4183
rect 2456 3987 2463 4176
rect 2616 4003 2623 4693
rect 2856 4676 2863 4693
rect 2776 4663 2783 4673
rect 2776 4656 2803 4663
rect 2896 4663 2903 4673
rect 2876 4656 2903 4663
rect 3016 4627 3023 4663
rect 3096 4656 3123 4663
rect 3116 4647 3123 4656
rect 3156 4627 3163 4956
rect 3456 4956 3483 4963
rect 3496 4956 3503 5096
rect 4416 5047 4423 5103
rect 3756 4963 3763 4973
rect 3596 4956 3623 4963
rect 3656 4956 3683 4963
rect 3736 4956 3763 4963
rect 3216 4927 3223 4953
rect 3476 4707 3483 4956
rect 3596 4747 3603 4956
rect 2676 4207 2683 4473
rect 2856 4456 2863 4473
rect 2896 4456 2903 4493
rect 3016 4487 3023 4593
rect 3236 4507 3243 4693
rect 3576 4683 3583 4713
rect 3576 4676 3603 4683
rect 3636 4676 3643 4693
rect 3607 4656 3623 4663
rect 3656 4647 3663 4663
rect 3676 4627 3683 4956
rect 3896 4643 3903 4683
rect 3896 4636 3923 4643
rect 3136 4476 3143 4493
rect 2816 4427 2823 4453
rect 2696 4227 2703 4413
rect 2716 4216 2743 4223
rect 2716 4207 2723 4216
rect 2756 4187 2763 4203
rect 2616 3996 2643 4003
rect 2116 3956 2143 3963
rect 2176 3927 2183 3963
rect 2196 3763 2203 3973
rect 2176 3756 2203 3763
rect 2176 3723 2183 3756
rect 2176 3716 2203 3723
rect 2116 3687 2123 3713
rect 2116 3516 2123 3673
rect 2176 3547 2183 3716
rect 2216 3687 2223 3703
rect 2356 3496 2363 3513
rect 2356 3187 2363 3243
rect 2396 3236 2403 3253
rect 2456 3227 2463 3973
rect 2496 3667 2503 3703
rect 2496 3467 2503 3653
rect 2616 3607 2623 3996
rect 2656 3967 2663 3983
rect 2956 3747 2963 3963
rect 2756 3716 2783 3723
rect 2816 3716 2823 3733
rect 2756 3687 2763 3716
rect 2796 3667 2803 3683
rect 2736 3516 2763 3523
rect 2956 3516 2983 3523
rect 2996 3516 3003 3593
rect 2756 3507 2763 3516
rect 2656 3496 2683 3503
rect 2656 3487 2663 3496
rect 2476 3207 2483 3233
rect 2096 3067 2103 3173
rect 2076 2787 2083 3033
rect 2096 3027 2103 3053
rect 2476 3043 2483 3193
rect 2556 3087 2563 3293
rect 2636 3236 2643 3313
rect 2716 3167 2723 3493
rect 2556 3043 2563 3073
rect 2316 3036 2343 3043
rect 2156 2776 2163 2813
rect 2096 2747 2103 2763
rect 2096 2263 2103 2633
rect 2216 2556 2223 2573
rect 2276 2563 2283 2973
rect 2256 2556 2283 2563
rect 2176 2536 2203 2543
rect 2036 2227 2043 2263
rect 2076 2256 2103 2263
rect 2156 2256 2163 2273
rect 1856 2056 1883 2063
rect 1736 1347 1743 1553
rect 1776 1336 1783 1573
rect 1716 1296 1743 1303
rect 1536 1096 1543 1293
rect 1596 1116 1623 1123
rect 1516 787 1523 1093
rect 1616 1087 1623 1116
rect 1616 827 1623 1073
rect 1516 647 1523 773
rect 1536 636 1543 653
rect 1576 636 1583 813
rect 1716 787 1723 823
rect 1596 376 1603 673
rect 1636 376 1663 383
rect 1616 327 1623 363
rect 1656 347 1663 376
rect 1736 207 1743 1296
rect 1836 1127 1843 1873
rect 1856 1307 1863 1803
rect 1876 1767 1883 1823
rect 1916 1816 1943 1823
rect 1936 1767 1943 1816
rect 1916 1596 1923 1633
rect 1796 1096 1803 1113
rect 1836 1096 1843 1113
rect 1836 847 1843 1053
rect 1816 636 1823 753
rect 1856 603 1863 653
rect 1876 643 1883 1333
rect 1936 1007 1943 1573
rect 2036 1303 2043 2093
rect 2096 1827 2103 2133
rect 2156 2076 2163 2213
rect 2176 2127 2183 2536
rect 2236 2287 2243 2533
rect 2276 2247 2283 2556
rect 2296 2547 2303 3013
rect 2336 2987 2343 3036
rect 2396 3036 2423 3043
rect 2456 3036 2483 3043
rect 2536 3036 2563 3043
rect 2396 3007 2403 3036
rect 2356 2776 2383 2783
rect 2416 2776 2443 2783
rect 2356 2707 2363 2776
rect 2436 2607 2443 2776
rect 2476 2647 2483 3036
rect 2776 3016 2783 3173
rect 2856 3007 2863 3253
rect 2976 3227 2983 3516
rect 3016 3047 3023 4473
rect 3236 4467 3243 4493
rect 3616 4487 3623 4613
rect 3436 4476 3463 4483
rect 3376 4456 3383 4473
rect 3456 4467 3463 4476
rect 3676 4483 3683 4493
rect 3656 4476 3683 4483
rect 3236 4003 3243 4313
rect 3276 4216 3283 4233
rect 3316 4216 3343 4223
rect 3336 4167 3343 4216
rect 3416 4207 3423 4453
rect 3396 4187 3403 4193
rect 3216 3996 3243 4003
rect 3216 3967 3223 3996
rect 3136 3716 3143 3733
rect 3056 3703 3063 3713
rect 3056 3696 3083 3703
rect 3176 3703 3183 3713
rect 3156 3696 3183 3703
rect 3156 3516 3163 3533
rect 3196 3267 3203 3733
rect 3296 3547 3303 3703
rect 3296 3487 3303 3533
rect 3336 3447 3343 4153
rect 3496 3976 3503 4213
rect 3556 4187 3563 4223
rect 3596 4216 3603 4233
rect 3576 4187 3583 4203
rect 3536 4003 3543 4013
rect 3616 4007 3623 4473
rect 3856 4216 3863 4233
rect 3876 4107 3883 4203
rect 3536 3996 3563 4003
rect 3536 3963 3543 3996
rect 3647 3996 3663 4003
rect 3676 3996 3683 4093
rect 3476 3747 3483 3963
rect 3516 3956 3543 3963
rect 3376 3696 3403 3703
rect 3396 3687 3403 3696
rect 3656 3487 3663 3996
rect 3916 3767 3923 4636
rect 3956 4627 3963 4663
rect 3996 4647 4003 4943
rect 4156 4667 4163 4953
rect 4256 4687 4263 4943
rect 3996 4507 4003 4633
rect 4176 4456 4183 4683
rect 4236 4647 4243 4663
rect 4236 4627 4243 4633
rect 4236 4447 4243 4613
rect 4156 4327 4163 4443
rect 4196 4227 4203 4433
rect 4096 4216 4123 4223
rect 3856 3736 3883 3743
rect 3916 3736 3943 3743
rect 3756 3487 3763 3503
rect 3756 3327 3763 3453
rect 3636 3256 3663 3263
rect 3056 3223 3063 3253
rect 3036 3216 3063 3223
rect 3076 3043 3083 3153
rect 3076 3036 3103 3043
rect 2756 2947 2763 3003
rect 2676 2767 2683 2783
rect 2716 2776 2743 2783
rect 2656 2747 2663 2763
rect 2696 2743 2703 2763
rect 2676 2736 2703 2743
rect 2476 2576 2483 2593
rect 2496 2556 2503 2693
rect 2676 2547 2683 2736
rect 2736 2727 2743 2776
rect 2696 2556 2703 2633
rect 2796 2563 2803 2613
rect 2776 2556 2803 2563
rect 2456 2287 2463 2303
rect 2196 2076 2203 2133
rect 2116 2056 2143 2063
rect 2116 1807 2123 2056
rect 2196 1816 2203 1833
rect 2236 1607 2243 2113
rect 2396 2096 2403 2273
rect 2436 2127 2443 2283
rect 2476 2247 2483 2283
rect 2676 2076 2683 2293
rect 2716 2287 2723 2303
rect 2696 2267 2703 2283
rect 2696 2047 2703 2063
rect 2396 1807 2403 1993
rect 2396 1783 2403 1793
rect 2396 1776 2423 1783
rect 2176 1596 2203 1603
rect 2016 1296 2043 1303
rect 1936 867 1943 993
rect 2016 887 2023 1296
rect 2056 1167 2063 1293
rect 2096 1116 2103 1133
rect 2156 1107 2163 1593
rect 2176 1587 2183 1596
rect 2296 1347 2303 1593
rect 2436 1567 2443 1763
rect 2336 1336 2343 1553
rect 2316 1147 2323 1323
rect 2456 1307 2463 1633
rect 2476 1627 2483 2033
rect 2736 1867 2743 2253
rect 2856 2047 2863 2993
rect 2976 2743 2983 3033
rect 3096 3007 3103 3036
rect 3296 3036 3323 3043
rect 3016 2743 3023 2753
rect 3096 2747 3103 2993
rect 3236 2763 3243 2833
rect 3296 2807 3303 3036
rect 3336 2847 3343 3243
rect 3356 3047 3363 3213
rect 3236 2756 3263 2763
rect 3296 2756 3303 2773
rect 2956 2736 2983 2743
rect 2996 2736 3023 2743
rect 2916 2263 2923 2633
rect 2896 2256 2923 2263
rect 2936 2096 2943 2233
rect 2956 2107 2963 2736
rect 2996 2547 3003 2736
rect 3336 2743 3343 2793
rect 3316 2736 3343 2743
rect 3456 2647 3463 2743
rect 3356 2576 3363 2613
rect 3096 2556 3123 2563
rect 3116 2547 3123 2556
rect 3016 2536 3043 2543
rect 3016 2527 3023 2536
rect 3076 2287 3083 2533
rect 2476 1596 2483 1613
rect 2496 1347 2503 1583
rect 2536 1576 2543 1593
rect 2496 1287 2503 1333
rect 2596 1267 2603 1303
rect 2316 1127 2323 1133
rect 2016 856 2043 863
rect 1956 807 1963 843
rect 1996 767 2003 843
rect 2036 827 2043 856
rect 1876 636 1903 643
rect 1896 607 1903 636
rect 2116 616 2123 1103
rect 2256 887 2263 1093
rect 2456 1027 2463 1083
rect 2256 856 2263 873
rect 1836 596 1863 603
rect 2156 603 2163 653
rect 2136 596 2163 603
rect 1876 167 1883 343
rect 1916 327 1923 343
rect 1896 127 1903 323
rect 2056 156 2063 353
rect 2096 327 2103 593
rect 2196 323 2203 853
rect 2276 647 2283 833
rect 2396 616 2403 833
rect 2376 367 2383 603
rect 2476 343 2483 353
rect 2456 336 2483 343
rect 2176 316 2203 323
rect 2176 167 2183 316
rect 2196 156 2203 293
rect 2036 127 2043 143
rect 2496 127 2503 373
rect 2516 267 2523 1013
rect 2536 856 2543 873
rect 2576 856 2603 863
rect 2556 627 2563 843
rect 2596 827 2603 856
rect 2556 607 2563 613
rect 2616 407 2623 1833
rect 2676 1763 2683 1793
rect 2676 1756 2703 1763
rect 2736 1167 2743 1853
rect 2756 1607 2763 1793
rect 2816 1596 2823 1813
rect 2856 1596 2863 1613
rect 2756 1567 2763 1593
rect 2776 1576 2803 1583
rect 2776 1547 2783 1576
rect 2836 1567 2843 1583
rect 2896 1303 2903 1333
rect 2876 1296 2903 1303
rect 2676 1096 2683 1153
rect 2696 1076 2703 1093
rect 2736 1076 2763 1083
rect 2636 616 2663 623
rect 2636 567 2643 616
rect 2676 596 2683 633
rect 2736 603 2743 1053
rect 2756 1047 2763 1076
rect 2796 843 2803 1253
rect 2916 1007 2923 1093
rect 2796 836 2823 843
rect 2856 827 2863 843
rect 2716 596 2743 603
rect 2676 356 2683 553
rect 2796 336 2823 343
rect 2696 267 2703 323
rect 1776 107 1783 123
rect 2516 123 2523 193
rect 2816 156 2823 336
rect 2836 307 2843 343
rect 2856 156 2863 413
rect 2916 367 2923 653
rect 2936 387 2943 2033
rect 3016 1816 3043 1823
rect 3036 1787 3043 1816
rect 3056 1616 3083 1623
rect 2976 1147 2983 1613
rect 3056 1547 3063 1616
rect 3116 1563 3123 2513
rect 3236 2283 3243 2293
rect 3236 2276 3263 2283
rect 3196 2076 3203 2133
rect 3236 2076 3243 2253
rect 3316 2247 3323 2263
rect 3436 2263 3443 2633
rect 3436 2256 3463 2263
rect 3476 2243 3483 2773
rect 3536 2736 3543 3253
rect 3656 3207 3663 3256
rect 3736 3147 3743 3223
rect 3636 3047 3643 3053
rect 3576 2987 3583 3003
rect 3456 2236 3483 2243
rect 3196 1763 3203 1813
rect 3276 1796 3283 1813
rect 3436 1807 3443 1833
rect 3456 1807 3463 2236
rect 3476 2043 3483 2133
rect 3556 2043 3563 2933
rect 3636 2607 3643 3033
rect 3756 2667 3763 3313
rect 3856 3307 3863 3736
rect 3896 3467 3903 3503
rect 3776 2647 3783 3223
rect 3856 3216 3883 3223
rect 3876 3187 3883 3216
rect 3936 3207 3943 3736
rect 4096 3287 4103 4216
rect 4236 3996 4243 4153
rect 4276 3996 4283 4973
rect 4476 4663 4483 5103
rect 4716 5047 4723 5103
rect 4516 4956 4523 5033
rect 4556 4956 4563 4973
rect 4456 4476 4463 4663
rect 4476 4656 4503 4663
rect 4756 4663 4763 5103
rect 4816 4956 4823 5033
rect 5036 4727 5043 5103
rect 5036 4696 5063 4703
rect 4756 4656 4783 4663
rect 4496 4487 4503 4633
rect 4296 3976 4323 3983
rect 4316 3727 4323 3976
rect 4196 3716 4223 3723
rect 4136 3487 4143 3703
rect 4176 3496 4183 3673
rect 3896 3036 3903 3133
rect 3836 2767 3843 3033
rect 4056 2767 4063 3233
rect 4076 3207 4083 3223
rect 3796 2727 3803 2763
rect 3876 2743 3883 2753
rect 3596 2556 3623 2563
rect 3636 2556 3643 2593
rect 3736 2556 3743 2573
rect 3616 2307 3623 2556
rect 3796 2287 3803 2653
rect 3816 2587 3823 2743
rect 3856 2736 3883 2743
rect 4076 2587 4083 2723
rect 4156 2627 4163 3483
rect 4176 3036 4183 3053
rect 3876 2563 3883 2573
rect 3856 2556 3883 2563
rect 4096 2556 4103 2593
rect 4136 2556 4163 2563
rect 3936 2276 3943 2553
rect 3776 2063 3783 2233
rect 3816 2096 3823 2253
rect 4076 2103 4083 2313
rect 4076 2096 4103 2103
rect 3776 2056 3803 2063
rect 3476 2036 3503 2043
rect 3196 1756 3223 1763
rect 3136 1567 3143 1583
rect 3096 1556 3123 1563
rect 2976 1116 2983 1133
rect 3016 1116 3023 1353
rect 3056 1307 3063 1533
rect 3096 1243 3103 1556
rect 3456 1563 3463 1593
rect 3436 1556 3463 1563
rect 3416 1336 3423 1353
rect 3116 1267 3123 1323
rect 3196 1307 3203 1333
rect 3096 1236 3123 1243
rect 2996 623 3003 1073
rect 3116 856 3123 1236
rect 3196 843 3203 1153
rect 3176 836 3203 843
rect 3256 787 3263 1313
rect 3276 1096 3283 1253
rect 3316 1096 3323 1113
rect 3356 1083 3363 1333
rect 3336 1076 3363 1083
rect 3376 823 3383 1073
rect 3416 836 3423 1113
rect 3476 843 3483 1253
rect 3496 1087 3503 2036
rect 3536 2036 3563 2043
rect 3536 1843 3543 2036
rect 3516 1836 3543 1843
rect 3456 836 3483 843
rect 3376 816 3403 823
rect 2976 616 3003 623
rect 2976 427 2983 616
rect 2916 336 2923 353
rect 3076 343 3083 673
rect 3176 656 3203 663
rect 3176 587 3183 656
rect 3236 623 3243 733
rect 3256 643 3263 773
rect 3256 636 3283 643
rect 3356 636 3363 673
rect 3376 667 3383 816
rect 3436 807 3443 823
rect 3396 636 3423 643
rect 3216 616 3243 623
rect 3416 607 3423 636
rect 3056 336 3083 343
rect 3056 307 3063 336
rect 3096 307 3103 343
rect 2836 127 2843 143
rect 2516 116 2533 123
rect 2576 107 2583 123
rect 3036 -24 3043 73
rect 3076 -24 3083 93
rect 3136 87 3143 123
rect 3176 87 3183 573
rect 3436 363 3443 513
rect 3416 356 3443 363
rect 3396 156 3403 293
rect 3436 156 3443 356
rect 3416 127 3423 143
rect 3516 47 3523 1836
rect 3576 1816 3583 1833
rect 3816 1767 3823 1803
rect 3856 1796 3863 1853
rect 4056 1787 4063 2063
rect 3836 1767 3843 1783
rect 3976 1767 3983 1783
rect 4016 1767 4023 1783
rect 4096 1776 4103 2096
rect 3676 1547 3683 1583
rect 3656 1327 3663 1513
rect 3696 1327 3703 1343
rect 3796 1327 3803 1613
rect 3916 1596 3923 1613
rect 3676 1267 3683 1323
rect 3696 1307 3703 1313
rect 3596 1096 3603 1113
rect 3556 -24 3563 393
rect 3576 107 3583 1083
rect 3616 647 3623 1073
rect 3676 787 3683 803
rect 3716 787 3723 1323
rect 3796 1296 3803 1313
rect 3836 1107 3843 1533
rect 3916 1287 3923 1303
rect 3876 1116 3883 1273
rect 3916 1116 3943 1123
rect 3856 1096 3863 1113
rect 3936 1087 3943 1116
rect 3736 847 3743 1053
rect 3916 856 3943 863
rect 3976 856 4003 863
rect 3736 667 3743 833
rect 3916 827 3923 856
rect 3776 607 3783 633
rect 3916 527 3923 813
rect 3996 807 4003 856
rect 4076 603 4083 1073
rect 4116 627 4123 2273
rect 4156 1827 4163 2556
rect 4196 2327 4203 3273
rect 4216 3247 4223 3716
rect 4376 3687 4383 4473
rect 4436 4456 4443 4473
rect 4676 4467 4683 4493
rect 4707 4476 4723 4483
rect 4436 4196 4443 4253
rect 4456 4167 4463 4183
rect 4696 4183 4703 4473
rect 4776 4456 4803 4463
rect 4696 4176 4723 4183
rect 4416 3743 4423 4153
rect 4556 3996 4563 4153
rect 4616 4003 4623 4173
rect 4596 3996 4623 4003
rect 4396 3736 4423 3743
rect 4396 3487 4403 3736
rect 4436 3496 4443 3673
rect 4416 3287 4423 3483
rect 4476 3267 4483 3533
rect 4256 2556 4263 2593
rect 4276 2307 4283 3253
rect 4476 3207 4483 3253
rect 4476 3056 4483 3173
rect 4336 2763 4343 2813
rect 4336 2756 4363 2763
rect 4396 2756 4403 3033
rect 4456 3007 4463 3013
rect 4376 2607 4383 2743
rect 4396 2563 4403 2573
rect 4376 2556 4403 2563
rect 4176 2087 4183 2293
rect 4176 1807 4183 2073
rect 4216 2067 4223 2283
rect 4276 2256 4283 2293
rect 4336 2263 4343 2553
rect 4416 2527 4423 2743
rect 4336 2256 4363 2263
rect 4316 2076 4323 2253
rect 4356 2107 4363 2256
rect 4336 2027 4343 2063
rect 4176 1627 4183 1793
rect 4176 1567 4183 1613
rect 4136 1116 4143 1133
rect 4176 1116 4183 1353
rect 4256 1336 4263 1353
rect 4196 1096 4223 1103
rect 4216 1067 4223 1096
rect 4256 836 4263 853
rect 4296 827 4303 2013
rect 4396 1963 4403 2073
rect 4396 1956 4423 1963
rect 4416 1787 4423 1956
rect 4436 1787 4443 2093
rect 4496 2076 4503 2093
rect 4336 1547 4343 1783
rect 4436 1767 4443 1773
rect 4436 1607 4443 1753
rect 4476 1567 4483 1593
rect 4376 1287 4383 1303
rect 4516 1303 4523 3733
rect 4576 3707 4583 3993
rect 4616 3707 4623 3996
rect 4496 1296 4523 1303
rect 4416 687 4423 1293
rect 4456 1096 4463 1273
rect 4496 1083 4503 1093
rect 4516 1087 4523 1296
rect 4436 1047 4443 1083
rect 4476 1076 4503 1083
rect 4476 856 4503 863
rect 4476 847 4483 856
rect 4596 847 4603 3433
rect 4636 2743 4643 3693
rect 4716 3547 4723 3703
rect 4676 3516 4683 3533
rect 4736 3523 4743 3693
rect 4796 3687 4803 4456
rect 4856 3996 4883 4003
rect 4876 3967 4883 3996
rect 4716 3516 4743 3523
rect 4716 3223 4723 3293
rect 4656 3216 4683 3223
rect 4696 3216 4723 3223
rect 4616 2736 4643 2743
rect 4636 2583 4643 2736
rect 4656 2607 4663 2743
rect 4676 2727 4683 3216
rect 4696 3003 4703 3193
rect 4696 2996 4723 3003
rect 4756 2627 4763 3003
rect 4636 2576 4663 2583
rect 4636 2527 4643 2543
rect 4656 1843 4663 2576
rect 4696 2087 4703 2613
rect 4716 2296 4723 2313
rect 4756 2307 4763 2593
rect 4776 2287 4783 3493
rect 4896 3227 4903 3513
rect 4936 3483 4943 4693
rect 4956 4167 4963 4183
rect 4976 3516 5003 3523
rect 4976 3487 4983 3516
rect 4936 3476 4963 3483
rect 4916 2743 4923 3253
rect 4936 3047 4943 3223
rect 4956 3067 4963 3476
rect 5016 3107 5023 4683
rect 5036 4476 5043 4653
rect 5056 3087 5063 4696
rect 4896 2736 4923 2743
rect 4636 1836 4663 1843
rect 4516 827 4523 843
rect 4416 623 4423 673
rect 4416 616 4443 623
rect 4016 587 4023 603
rect 4056 596 4083 603
rect 3716 376 3723 393
rect 3656 123 3663 373
rect 3996 356 4003 373
rect 4096 347 4103 593
rect 3976 327 3983 343
rect 4116 327 4123 343
rect 4236 336 4243 393
rect 4436 347 4443 616
rect 4456 376 4483 383
rect 4456 343 4463 376
rect 4456 336 4483 343
rect 4016 156 4043 163
rect 4036 147 4043 156
rect 4156 156 4163 333
rect 4456 167 4463 336
rect 4476 176 4483 336
rect 4496 183 4503 363
rect 4496 176 4523 183
rect 3996 127 4003 143
rect 4516 127 4523 176
rect 3656 116 3673 123
rect 3716 87 3723 123
rect 3596 -24 3603 33
rect 4636 -24 4643 1836
rect 4696 1816 4703 2073
rect 4836 2056 4843 2533
rect 4876 2267 4883 2673
rect 4916 2556 4923 2713
rect 4936 2687 4943 2743
rect 4956 2607 4963 3053
rect 4956 2556 4963 2593
rect 4936 2527 4943 2543
rect 4716 1603 4723 1813
rect 4796 1707 4803 1783
rect 4696 1596 4723 1603
rect 4756 1596 4763 1693
rect 4816 1607 4823 2043
rect 4916 1787 4923 2313
rect 4976 2307 4983 3073
rect 5056 3036 5063 3053
rect 5036 3007 5043 3023
rect 4936 2247 4943 2273
rect 4956 2263 4963 2293
rect 4956 2256 4983 2263
rect 4956 2047 4963 2256
rect 4696 1567 4703 1596
rect 4696 1303 4703 1553
rect 4736 1527 4743 1583
rect 4696 1296 4723 1303
rect 4716 1127 4723 1296
rect 4776 1247 4783 1323
rect 4836 1287 4843 1773
rect 4976 1563 4983 1773
rect 4976 1556 5003 1563
rect 5056 1307 5063 2293
rect 5076 2287 5083 3093
rect 4936 1287 4943 1303
rect 4756 1087 4763 1113
rect 5016 1096 5023 1233
rect 4736 1076 4753 1083
rect 5056 1083 5063 1293
rect 5036 1076 5063 1083
rect 4776 856 4803 863
rect 4776 823 4783 856
rect 4776 816 4803 823
rect 4696 607 4703 623
rect 4736 407 4743 653
rect 4736 376 4743 393
rect 4796 367 4803 816
rect 4976 616 4983 853
rect 4996 323 5003 603
rect 5036 356 5043 373
rect 4996 316 5023 323
rect 4776 136 4783 253
rect 5016 247 5023 316
rect 4816 123 4823 133
rect 4796 116 4823 123
rect 4956 27 4963 233
rect 4996 27 5003 123
rect 4956 -24 4963 13
<< m3contact >>
rect 693 4973 707 4987
rect 1213 4973 1227 4987
rect 1313 4973 1327 4987
rect 1533 4973 1547 4987
rect 1793 4973 1807 4987
rect 1893 4973 1907 4987
rect 513 4953 527 4967
rect 213 4933 227 4947
rect 493 4933 507 4947
rect 193 4913 207 4927
rect 233 4913 247 4927
rect 653 4953 667 4967
rect 573 4913 587 4927
rect 233 4893 247 4907
rect 533 4893 547 4907
rect 513 4713 527 4727
rect 253 4493 267 4507
rect 233 4433 247 4447
rect 573 4653 587 4667
rect 593 4653 607 4667
rect 553 4633 567 4647
rect 313 4493 327 4507
rect 433 4473 447 4487
rect 493 4473 507 4487
rect 513 4473 527 4487
rect 313 4453 327 4467
rect 253 4233 267 4247
rect 293 4233 307 4247
rect 213 4213 227 4227
rect 273 4213 287 4227
rect 233 4193 247 4207
rect 273 4033 287 4047
rect 253 4013 267 4027
rect 233 3993 247 4007
rect 453 4433 467 4447
rect 573 4473 587 4487
rect 573 4433 587 4447
rect 533 4233 547 4247
rect 493 4213 507 4227
rect 433 4193 447 4207
rect 513 4193 527 4207
rect 573 4193 587 4207
rect 513 4033 527 4047
rect 533 4033 547 4047
rect 313 3993 327 4007
rect 273 3733 287 3747
rect 233 3713 247 3727
rect 293 3693 307 3707
rect 93 3593 107 3607
rect 253 3593 267 3607
rect 153 3533 167 3547
rect 93 3193 107 3207
rect 213 3513 227 3527
rect 493 3973 507 3987
rect 1033 4953 1047 4967
rect 1173 4953 1187 4967
rect 1813 4953 1827 4967
rect 853 4933 867 4947
rect 1013 4933 1027 4947
rect 773 4693 787 4707
rect 773 4673 787 4687
rect 733 4493 747 4507
rect 813 4673 827 4687
rect 793 4653 807 4667
rect 1093 4933 1107 4947
rect 1553 4933 1567 4947
rect 1573 4933 1587 4947
rect 1473 4693 1487 4707
rect 1393 4673 1407 4687
rect 1053 4653 1067 4667
rect 1113 4653 1127 4667
rect 1133 4633 1147 4647
rect 1053 4493 1067 4507
rect 1033 4473 1047 4487
rect 793 4433 807 4447
rect 773 4413 787 4427
rect 813 4413 827 4427
rect 733 4233 747 4247
rect 793 4193 807 4207
rect 773 4033 787 4047
rect 433 3733 447 3747
rect 213 3453 227 3467
rect 313 3453 327 3467
rect 553 3733 567 3747
rect 533 3713 547 3727
rect 633 3673 647 3687
rect 1093 4473 1107 4487
rect 1073 4453 1087 4467
rect 1153 4593 1167 4607
rect 1413 4533 1427 4547
rect 1373 4513 1387 4527
rect 1553 4533 1567 4547
rect 1373 4493 1387 4507
rect 1473 4493 1487 4507
rect 1413 4473 1427 4487
rect 1473 4473 1487 4487
rect 1013 4213 1027 4227
rect 993 3993 1007 4007
rect 833 3973 847 3987
rect 973 3973 987 3987
rect 1013 3973 1027 3987
rect 1133 4233 1147 4247
rect 1393 4233 1407 4247
rect 1073 4213 1087 4227
rect 1093 4193 1107 4207
rect 1273 4213 1287 4227
rect 1353 4213 1367 4227
rect 1373 4193 1387 4207
rect 1273 4013 1287 4027
rect 1133 3993 1147 4007
rect 1233 3993 1247 4007
rect 733 3773 747 3787
rect 1073 3773 1087 3787
rect 813 3753 827 3767
rect 1113 3753 1127 3767
rect 753 3713 767 3727
rect 813 3713 827 3727
rect 853 3713 867 3727
rect 1093 3713 1107 3727
rect 653 3533 667 3547
rect 673 3533 687 3547
rect 493 3513 507 3527
rect 473 3493 487 3507
rect 513 3493 527 3507
rect 453 3453 467 3467
rect 433 3433 447 3447
rect 453 3433 467 3447
rect 493 3433 507 3447
rect 253 3313 267 3327
rect 133 3153 147 3167
rect 153 3153 167 3167
rect 73 3053 87 3067
rect 233 3013 247 3027
rect 413 3233 427 3247
rect 453 3233 467 3247
rect 353 3153 367 3167
rect 153 2733 167 2747
rect 93 2653 107 2667
rect 253 2693 267 2707
rect 233 2673 247 2687
rect 373 2733 387 2747
rect 373 2713 387 2727
rect 373 2693 387 2707
rect 253 2653 267 2667
rect 333 2653 347 2667
rect 233 2553 247 2567
rect 293 2573 307 2587
rect 313 2553 327 2567
rect 273 2533 287 2547
rect 233 2233 247 2247
rect 113 1753 127 1767
rect 313 2253 327 2267
rect 273 2053 287 2067
rect 353 2053 367 2067
rect 213 1993 227 2007
rect 253 1793 267 1807
rect 333 1793 347 1807
rect 273 1773 287 1787
rect 313 1773 327 1787
rect 253 1753 267 1767
rect 293 1593 307 1607
rect 273 1573 287 1587
rect 153 1313 167 1327
rect 233 1313 247 1327
rect 233 1273 247 1287
rect 33 853 47 867
rect 73 853 87 867
rect 233 853 247 867
rect 133 833 147 847
rect 153 813 167 827
rect 353 1573 367 1587
rect 433 3213 447 3227
rect 733 3293 747 3307
rect 793 3693 807 3707
rect 733 3253 747 3267
rect 753 3253 767 3267
rect 773 3233 787 3247
rect 713 3213 727 3227
rect 473 3193 487 3207
rect 633 3193 647 3207
rect 633 3013 647 3027
rect 453 2753 467 2767
rect 573 2733 587 2747
rect 613 2713 627 2727
rect 453 2673 467 2687
rect 433 2273 447 2287
rect 533 2653 547 2667
rect 493 2553 507 2567
rect 673 2993 687 3007
rect 693 2773 707 2787
rect 633 2573 647 2587
rect 753 3193 767 3207
rect 1313 3993 1327 4007
rect 1293 3693 1307 3707
rect 833 3673 847 3687
rect 1233 3673 1247 3687
rect 1053 3553 1067 3567
rect 1013 3513 1027 3527
rect 1173 3533 1187 3547
rect 1193 3533 1207 3547
rect 1153 3513 1167 3527
rect 893 3493 907 3507
rect 993 3493 1007 3507
rect 793 3013 807 3027
rect 933 3013 947 3027
rect 913 2993 927 3007
rect 873 2973 887 2987
rect 833 2953 847 2967
rect 913 2933 927 2947
rect 853 2753 867 2767
rect 1073 3293 1087 3307
rect 1033 3253 1047 3267
rect 1113 3273 1127 3287
rect 1093 3253 1107 3267
rect 1053 3233 1067 3247
rect 1013 2973 1027 2987
rect 993 2753 1007 2767
rect 1033 2753 1047 2767
rect 973 2733 987 2747
rect 1013 2733 1027 2747
rect 1273 3513 1287 3527
rect 1393 3693 1407 3707
rect 1373 3673 1387 3687
rect 1353 3653 1367 3667
rect 1353 3513 1367 3527
rect 1173 3193 1187 3207
rect 1453 3073 1467 3087
rect 1153 3013 1167 3027
rect 1173 2793 1187 2807
rect 1313 2793 1327 2807
rect 1113 2773 1127 2787
rect 1273 2773 1287 2787
rect 1393 2773 1407 2787
rect 1173 2733 1187 2747
rect 853 2693 867 2707
rect 513 2533 527 2547
rect 513 2273 527 2287
rect 493 2253 507 2267
rect 533 2253 547 2267
rect 713 2533 727 2547
rect 813 2533 827 2547
rect 1093 2713 1107 2727
rect 1093 2573 1107 2587
rect 1293 2733 1307 2747
rect 1333 2733 1347 2747
rect 1193 2713 1207 2727
rect 1173 2533 1187 2547
rect 1133 2513 1147 2527
rect 773 2273 787 2287
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 1013 2273 1027 2287
rect 753 2253 767 2267
rect 1093 2293 1107 2307
rect 1073 2273 1087 2287
rect 473 2233 487 2247
rect 533 2233 547 2247
rect 573 2233 587 2247
rect 433 2093 447 2107
rect 793 2233 807 2247
rect 753 2133 767 2147
rect 513 2093 527 2107
rect 913 2093 927 2107
rect 493 2053 507 2067
rect 753 2073 767 2087
rect 513 1793 527 1807
rect 473 1773 487 1787
rect 493 1773 507 1787
rect 453 1593 467 1607
rect 413 1333 427 1347
rect 373 1313 387 1327
rect 333 1273 347 1287
rect 553 1773 567 1787
rect 553 1733 567 1747
rect 673 1733 687 1747
rect 593 1593 607 1607
rect 693 1593 707 1607
rect 573 1573 587 1587
rect 573 1333 587 1347
rect 633 1333 647 1347
rect 673 1333 687 1347
rect 513 1153 527 1167
rect 453 1133 467 1147
rect 493 1113 507 1127
rect 473 1093 487 1107
rect 613 1313 627 1327
rect 573 1093 587 1107
rect 473 833 487 847
rect 273 813 287 827
rect 313 813 327 827
rect 253 653 267 667
rect 453 653 467 667
rect 673 1293 687 1307
rect 653 1153 667 1167
rect 633 1113 647 1127
rect 793 1773 807 1787
rect 893 2073 907 2087
rect 853 1813 867 1827
rect 813 1633 827 1647
rect 893 1593 907 1607
rect 833 1553 847 1567
rect 833 1333 847 1347
rect 853 1333 867 1347
rect 793 1313 807 1327
rect 713 1293 727 1307
rect 813 1293 827 1307
rect 753 1113 767 1127
rect 833 1113 847 1127
rect 573 813 587 827
rect 533 613 547 627
rect 473 593 487 607
rect 493 593 507 607
rect 513 593 527 607
rect 753 833 767 847
rect 1033 1973 1047 1987
rect 1053 1793 1067 1807
rect 1033 1653 1047 1667
rect 1073 1613 1087 1627
rect 1133 1553 1147 1567
rect 1313 2573 1327 2587
rect 1353 2573 1367 2587
rect 1433 2733 1447 2747
rect 1333 2513 1347 2527
rect 1373 2533 1387 2547
rect 1353 2253 1367 2267
rect 1293 2093 1307 2107
rect 1313 2093 1327 2107
rect 1313 2033 1327 2047
rect 1353 1973 1367 1987
rect 1293 1813 1307 1827
rect 1333 1813 1347 1827
rect 1273 1793 1287 1807
rect 1313 1793 1327 1807
rect 1353 1793 1367 1807
rect 1333 1753 1347 1767
rect 1393 1653 1407 1667
rect 1373 1573 1387 1587
rect 1853 4913 1867 4927
rect 1733 4893 1747 4907
rect 1613 4533 1627 4547
rect 1673 4633 1687 4647
rect 1953 4953 1967 4967
rect 2613 4953 2627 4967
rect 2653 4953 2667 4967
rect 2693 4953 2707 4967
rect 3093 4953 3107 4967
rect 1893 4873 1907 4887
rect 2113 4933 2127 4947
rect 2353 4933 2367 4947
rect 2393 4933 2407 4947
rect 2413 4913 2427 4927
rect 2133 4873 2147 4887
rect 2673 4933 2687 4947
rect 2713 4933 2727 4947
rect 2953 4933 2967 4947
rect 2933 4913 2947 4927
rect 2513 4693 2527 4707
rect 2613 4693 2627 4707
rect 2853 4693 2867 4707
rect 2973 4693 2987 4707
rect 1733 4613 1747 4627
rect 1693 4513 1707 4527
rect 1673 4473 1687 4487
rect 1593 4453 1607 4467
rect 1653 4453 1667 4467
rect 1573 4253 1587 4267
rect 1573 4013 1587 4027
rect 1653 4193 1667 4207
rect 1633 4173 1647 4187
rect 1613 4133 1627 4147
rect 1533 3773 1547 3787
rect 1553 3693 1567 3707
rect 1533 3453 1547 3467
rect 1673 3913 1687 3927
rect 1953 4673 1967 4687
rect 2093 4673 2107 4687
rect 2233 4673 2247 4687
rect 1933 4653 1947 4667
rect 2153 4653 2167 4667
rect 2453 4653 2467 4667
rect 2533 4653 2547 4667
rect 2193 4633 2207 4647
rect 2493 4633 2507 4647
rect 1973 4613 1987 4627
rect 1893 4513 1907 4527
rect 2553 4513 2567 4527
rect 1933 4493 1947 4507
rect 2513 4473 2527 4487
rect 1953 4453 1967 4467
rect 1913 4233 1927 4247
rect 2213 4453 2227 4467
rect 2193 4433 2207 4447
rect 2233 4433 2247 4447
rect 2273 4433 2287 4447
rect 2533 4433 2547 4447
rect 1973 4233 1987 4247
rect 2073 4233 2087 4247
rect 1953 4213 1967 4227
rect 1893 4173 1907 4187
rect 1933 4173 1947 4187
rect 1833 4013 1847 4027
rect 1873 3993 1887 4007
rect 1853 3973 1867 3987
rect 2113 4213 2127 4227
rect 2153 4213 2167 4227
rect 2313 4413 2327 4427
rect 2173 4193 2187 4207
rect 2113 4133 2127 4147
rect 2093 4013 2107 4027
rect 1853 3953 1867 3967
rect 1893 3953 1907 3967
rect 1973 3953 1987 3967
rect 2053 3953 2067 3967
rect 1873 3933 1887 3947
rect 1813 3913 1827 3927
rect 1733 3693 1747 3707
rect 1673 3673 1687 3687
rect 1633 3653 1647 3667
rect 1673 3553 1687 3567
rect 1873 3713 1887 3727
rect 1913 3713 1927 3727
rect 1613 3293 1627 3307
rect 1533 3253 1547 3267
rect 1753 3253 1767 3267
rect 1793 3253 1807 3267
rect 1533 3233 1547 3247
rect 1733 3233 1747 3247
rect 1513 3213 1527 3227
rect 1573 3213 1587 3227
rect 1693 3213 1707 3227
rect 1553 3193 1567 3207
rect 1713 2973 1727 2987
rect 1673 2953 1687 2967
rect 1553 2713 1567 2727
rect 1573 2693 1587 2707
rect 1533 2673 1547 2687
rect 1633 2673 1647 2687
rect 1673 2553 1687 2567
rect 1653 2533 1667 2547
rect 1493 2293 1507 2307
rect 1573 2293 1587 2307
rect 1473 1633 1487 1647
rect 1413 1593 1427 1607
rect 1033 1333 1047 1347
rect 1113 1333 1127 1347
rect 1193 1333 1207 1347
rect 1033 1313 1047 1327
rect 913 1073 927 1087
rect 1053 1073 1067 1087
rect 1153 1313 1167 1327
rect 1173 1293 1187 1307
rect 1433 1293 1447 1307
rect 1213 1133 1227 1147
rect 1293 1133 1307 1147
rect 1513 2093 1527 2107
rect 1473 1313 1487 1327
rect 1473 1133 1487 1147
rect 1453 1113 1467 1127
rect 1213 1093 1227 1107
rect 1273 1093 1287 1107
rect 1393 1093 1407 1107
rect 1233 873 1247 887
rect 1013 853 1027 867
rect 1113 853 1127 867
rect 1193 853 1207 867
rect 993 833 1007 847
rect 1153 833 1167 847
rect 853 813 867 827
rect 733 793 747 807
rect 813 793 827 807
rect 713 733 727 747
rect 773 733 787 747
rect 953 673 967 687
rect 1093 733 1107 747
rect 1133 673 1147 687
rect 993 653 1007 667
rect 1173 653 1187 667
rect 1073 633 1087 647
rect 833 613 847 627
rect 1133 613 1147 627
rect 793 593 807 607
rect 453 353 467 367
rect 493 353 507 367
rect 493 333 507 347
rect 513 293 527 307
rect 233 173 247 187
rect 333 173 347 187
rect 133 153 147 167
rect 713 193 727 207
rect 773 313 787 327
rect 1013 333 1027 347
rect 793 293 807 307
rect 753 173 767 187
rect 1073 333 1087 347
rect 1033 313 1047 327
rect 1113 293 1127 307
rect 373 153 387 167
rect 453 153 467 167
rect 513 153 527 167
rect 533 153 547 167
rect 693 153 707 167
rect 1213 653 1227 667
rect 1433 853 1447 867
rect 1413 833 1427 847
rect 1253 673 1267 687
rect 1273 673 1287 687
rect 1233 613 1247 627
rect 1193 353 1207 367
rect 1173 153 1187 167
rect 1313 373 1327 387
rect 1333 353 1347 367
rect 1413 373 1427 387
rect 1373 333 1387 347
rect 1373 153 1387 167
rect 1413 153 1427 167
rect 213 133 227 147
rect 533 133 547 147
rect 753 133 767 147
rect 993 133 1007 147
rect 1233 133 1247 147
rect 1633 2273 1647 2287
rect 1613 2253 1627 2267
rect 1693 2273 1707 2287
rect 1593 2233 1607 2247
rect 1633 2073 1647 2087
rect 1693 2073 1707 2087
rect 1553 2033 1567 2047
rect 1633 2033 1647 2047
rect 1673 2033 1687 2047
rect 1593 1873 1607 1887
rect 1593 1793 1607 1807
rect 1533 1593 1547 1607
rect 1693 1613 1707 1627
rect 1653 1573 1667 1587
rect 1633 1553 1647 1567
rect 1673 1553 1687 1567
rect 1613 1313 1627 1327
rect 1533 1293 1547 1307
rect 1833 3253 1847 3267
rect 1893 3693 1907 3707
rect 2033 3693 2047 3707
rect 1953 3673 1967 3687
rect 1933 3473 1947 3487
rect 1973 3213 1987 3227
rect 2013 3193 2027 3207
rect 1793 3173 1807 3187
rect 1813 3173 1827 3187
rect 1953 3053 1967 3067
rect 2033 3053 2047 3067
rect 1853 3013 1867 3027
rect 1813 2993 1827 3007
rect 1773 2953 1787 2967
rect 1753 2713 1767 2727
rect 1813 2753 1827 2767
rect 1833 2753 1847 2767
rect 1933 2593 1947 2607
rect 1893 2573 1907 2587
rect 1913 2573 1927 2587
rect 1873 2533 1887 2547
rect 1993 3033 2007 3047
rect 1973 3013 1987 3027
rect 2013 3013 2027 3027
rect 1973 2553 1987 2567
rect 1953 2533 1967 2547
rect 1853 2313 1867 2327
rect 1913 2313 1927 2327
rect 1793 2233 1807 2247
rect 1833 2073 1847 2087
rect 1873 2293 1887 2307
rect 2073 3493 2087 3507
rect 2433 4233 2447 4247
rect 2493 4233 2507 4247
rect 2573 4233 2587 4247
rect 2413 4213 2427 4227
rect 2313 4193 2327 4207
rect 2413 4173 2427 4187
rect 2453 4213 2467 4227
rect 2473 4193 2487 4207
rect 2213 4013 2227 4027
rect 2433 4013 2447 4027
rect 2773 4673 2787 4687
rect 2813 4673 2827 4687
rect 2893 4673 2907 4687
rect 2833 4653 2847 4667
rect 2973 4653 2987 4667
rect 3113 4633 3127 4647
rect 3213 4953 3227 4967
rect 4413 5033 4427 5047
rect 3753 4973 3767 4987
rect 3973 4973 3987 4987
rect 4233 4973 4247 4987
rect 4273 4973 4287 4987
rect 3213 4913 3227 4927
rect 3573 4713 3587 4727
rect 3233 4693 3247 4707
rect 3473 4693 3487 4707
rect 3013 4613 3027 4627
rect 3153 4613 3167 4627
rect 3013 4593 3027 4607
rect 2893 4493 2907 4507
rect 2673 4473 2687 4487
rect 2853 4473 2867 4487
rect 2813 4453 2827 4467
rect 3353 4673 3367 4687
rect 3633 4693 3647 4707
rect 3333 4633 3347 4647
rect 3653 4633 3667 4647
rect 4153 4953 4167 4967
rect 3933 4673 3947 4687
rect 3913 4653 3927 4667
rect 3613 4613 3627 4627
rect 3673 4613 3687 4627
rect 3133 4493 3147 4507
rect 3233 4493 3247 4507
rect 3013 4473 3027 4487
rect 3093 4473 3107 4487
rect 2833 4433 2847 4447
rect 2873 4433 2887 4447
rect 2693 4413 2707 4427
rect 2813 4413 2827 4427
rect 2693 4213 2707 4227
rect 2773 4213 2787 4227
rect 2673 4193 2687 4207
rect 2713 4193 2727 4207
rect 2793 4193 2807 4207
rect 2753 4173 2767 4187
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 2413 3973 2427 3987
rect 2453 3973 2467 3987
rect 2173 3913 2187 3927
rect 2113 3713 2127 3727
rect 2113 3673 2127 3687
rect 2233 3713 2247 3727
rect 2253 3693 2267 3707
rect 2213 3673 2227 3687
rect 2133 3533 2147 3547
rect 2173 3533 2187 3547
rect 2353 3513 2367 3527
rect 2393 3493 2407 3507
rect 2373 3473 2387 3487
rect 2413 3473 2427 3487
rect 2393 3253 2407 3267
rect 2533 3713 2547 3727
rect 2473 3673 2487 3687
rect 2493 3653 2507 3667
rect 2673 3993 2687 4007
rect 2693 3973 2707 3987
rect 2973 3973 2987 3987
rect 2653 3953 2667 3967
rect 2993 3953 3007 3967
rect 2813 3733 2827 3747
rect 2953 3733 2967 3747
rect 2833 3693 2847 3707
rect 2753 3673 2767 3687
rect 2793 3653 2807 3667
rect 2613 3593 2627 3607
rect 2993 3593 3007 3607
rect 2693 3513 2707 3527
rect 2713 3493 2727 3507
rect 2753 3493 2767 3507
rect 2653 3473 2667 3487
rect 2493 3453 2507 3467
rect 2633 3313 2647 3327
rect 2553 3293 2567 3307
rect 2473 3233 2487 3247
rect 2373 3213 2387 3227
rect 2413 3213 2427 3227
rect 2453 3213 2467 3227
rect 2473 3193 2487 3207
rect 2093 3173 2107 3187
rect 2353 3173 2367 3187
rect 2093 3053 2107 3067
rect 2293 3053 2307 3067
rect 2073 3033 2087 3047
rect 2273 3033 2287 3047
rect 2853 3253 2867 3267
rect 2773 3233 2787 3247
rect 2773 3173 2787 3187
rect 2713 3153 2727 3167
rect 2553 3073 2567 3087
rect 2093 3013 2107 3027
rect 2293 3013 2307 3027
rect 2273 2973 2287 2987
rect 2153 2813 2167 2827
rect 2073 2773 2087 2787
rect 2113 2773 2127 2787
rect 2133 2753 2147 2767
rect 2093 2733 2107 2747
rect 2093 2633 2107 2647
rect 1893 2273 1907 2287
rect 2053 2273 2067 2287
rect 2213 2573 2227 2587
rect 2153 2273 2167 2287
rect 2033 2213 2047 2227
rect 2153 2213 2167 2227
rect 2093 2133 2107 2147
rect 2033 2093 2047 2107
rect 1793 1873 1807 1887
rect 1833 1873 1847 1887
rect 1773 1833 1787 1847
rect 1773 1573 1787 1587
rect 1733 1553 1747 1567
rect 1733 1333 1747 1347
rect 1753 1313 1767 1327
rect 1513 1093 1527 1107
rect 1553 1113 1567 1127
rect 1573 1093 1587 1107
rect 1613 1073 1627 1087
rect 1573 813 1587 827
rect 1613 813 1627 827
rect 1673 813 1687 827
rect 1513 773 1527 787
rect 1553 653 1567 667
rect 1513 633 1527 647
rect 1693 793 1707 807
rect 1713 773 1727 787
rect 1593 673 1607 687
rect 1653 333 1667 347
rect 1613 313 1627 327
rect 1893 1793 1907 1807
rect 1873 1753 1887 1767
rect 1933 1753 1947 1767
rect 1913 1633 1927 1647
rect 1953 1593 1967 1607
rect 1933 1573 1947 1587
rect 1873 1333 1887 1347
rect 1853 1293 1867 1307
rect 1793 1113 1807 1127
rect 1833 1113 1847 1127
rect 1813 1073 1827 1087
rect 1853 1073 1867 1087
rect 1833 1053 1847 1067
rect 1833 833 1847 847
rect 1813 753 1827 767
rect 1853 653 1867 667
rect 2233 2533 2247 2547
rect 2233 2273 2247 2287
rect 2393 2993 2407 3007
rect 2333 2973 2347 2987
rect 2393 2753 2407 2767
rect 2353 2693 2367 2707
rect 2973 3213 2987 3227
rect 3673 4493 3687 4507
rect 3873 4493 3887 4507
rect 3373 4473 3387 4487
rect 3393 4473 3407 4487
rect 3233 4453 3247 4467
rect 3533 4473 3547 4487
rect 3573 4473 3587 4487
rect 3613 4473 3627 4487
rect 3413 4453 3427 4467
rect 3453 4453 3467 4467
rect 3233 4313 3247 4327
rect 3033 4193 3047 4207
rect 3053 4153 3067 4167
rect 3093 3993 3107 4007
rect 3133 3993 3147 4007
rect 3273 4233 3287 4247
rect 3293 4193 3307 4207
rect 3593 4233 3607 4247
rect 3493 4213 3507 4227
rect 3393 4193 3407 4207
rect 3413 4193 3427 4207
rect 3333 4153 3347 4167
rect 3213 3953 3227 3967
rect 3133 3733 3147 3747
rect 3193 3733 3207 3747
rect 3053 3713 3067 3727
rect 3093 3713 3107 3727
rect 3173 3713 3187 3727
rect 3113 3693 3127 3707
rect 3153 3533 3167 3547
rect 3113 3513 3127 3527
rect 3253 3693 3267 3707
rect 3293 3533 3307 3547
rect 3233 3513 3247 3527
rect 3293 3473 3307 3487
rect 3533 4193 3547 4207
rect 3573 4173 3587 4187
rect 3533 4013 3547 4027
rect 3893 4453 3907 4467
rect 3853 4233 3867 4247
rect 3893 4213 3907 4227
rect 3673 4093 3687 4107
rect 3873 4093 3887 4107
rect 3613 3993 3627 4007
rect 3633 3993 3647 4007
rect 3473 3733 3487 3747
rect 3613 3713 3627 3727
rect 3393 3673 3407 3687
rect 3593 3673 3607 3687
rect 3473 3533 3487 3547
rect 3493 3493 3507 3507
rect 4153 4653 4167 4667
rect 3993 4633 4007 4647
rect 3953 4613 3967 4627
rect 3993 4493 4007 4507
rect 4213 4673 4227 4687
rect 4253 4673 4267 4687
rect 4193 4653 4207 4667
rect 4233 4633 4247 4647
rect 4233 4613 4247 4627
rect 4193 4433 4207 4447
rect 4233 4433 4247 4447
rect 4153 4313 4167 4327
rect 3973 4013 3987 4027
rect 3993 3973 4007 3987
rect 3913 3753 3927 3767
rect 3653 3473 3667 3487
rect 3753 3473 3767 3487
rect 3753 3453 3767 3467
rect 3333 3433 3347 3447
rect 3753 3313 3767 3327
rect 3053 3253 3067 3267
rect 3193 3253 3207 3267
rect 3313 3253 3327 3267
rect 3353 3253 3367 3267
rect 3533 3253 3547 3267
rect 3593 3253 3607 3267
rect 3073 3213 3087 3227
rect 3073 3153 3087 3167
rect 2973 3033 2987 3047
rect 3013 3033 3027 3047
rect 3033 3033 3047 3047
rect 2793 2993 2807 3007
rect 2853 2993 2867 3007
rect 2753 2933 2767 2947
rect 2673 2753 2687 2767
rect 2653 2733 2667 2747
rect 2493 2693 2507 2707
rect 2473 2633 2487 2647
rect 2433 2593 2447 2607
rect 2473 2593 2487 2607
rect 2653 2553 2667 2567
rect 2733 2713 2747 2727
rect 2693 2633 2707 2647
rect 2793 2613 2807 2627
rect 2293 2533 2307 2547
rect 2533 2533 2547 2547
rect 2673 2533 2687 2547
rect 2413 2293 2427 2307
rect 2673 2293 2687 2307
rect 2393 2273 2407 2287
rect 2273 2233 2287 2247
rect 2193 2133 2207 2147
rect 2173 2113 2187 2127
rect 2233 2113 2247 2127
rect 2093 1813 2107 1827
rect 2173 2053 2187 2067
rect 2193 1833 2207 1847
rect 2153 1813 2167 1827
rect 2113 1793 2127 1807
rect 2173 1793 2187 1807
rect 2453 2273 2467 2287
rect 2473 2233 2487 2247
rect 2433 2113 2447 2127
rect 2753 2293 2767 2307
rect 2713 2273 2727 2287
rect 2733 2273 2747 2287
rect 2693 2253 2707 2267
rect 2733 2253 2747 2267
rect 2813 2253 2827 2267
rect 2713 2073 2727 2087
rect 2413 2053 2427 2067
rect 2653 2053 2667 2067
rect 2473 2033 2487 2047
rect 2693 2033 2707 2047
rect 2393 1993 2407 2007
rect 2393 1793 2407 1807
rect 2453 1773 2467 1787
rect 2153 1593 2167 1607
rect 1933 993 1947 1007
rect 2053 1293 2067 1307
rect 2053 1153 2067 1167
rect 2093 1133 2107 1147
rect 2133 1113 2147 1127
rect 2233 1593 2247 1607
rect 2253 1593 2267 1607
rect 2293 1593 2307 1607
rect 2173 1573 2187 1587
rect 2213 1553 2227 1567
rect 2453 1633 2467 1647
rect 2333 1553 2347 1567
rect 2433 1553 2447 1567
rect 2293 1333 2307 1347
rect 3093 2993 3107 3007
rect 3013 2753 3027 2767
rect 3233 2833 3247 2847
rect 3353 3213 3367 3227
rect 3353 3033 3367 3047
rect 3333 2833 3347 2847
rect 3293 2793 3307 2807
rect 3333 2793 3347 2807
rect 3293 2773 3307 2787
rect 2913 2633 2927 2647
rect 2933 2253 2947 2267
rect 2933 2233 2947 2247
rect 3093 2733 3107 2747
rect 3273 2733 3287 2747
rect 3473 2773 3487 2787
rect 3413 2733 3427 2747
rect 3433 2633 3447 2647
rect 3453 2633 3467 2647
rect 3353 2613 3367 2627
rect 3053 2553 3067 2567
rect 2993 2533 3007 2547
rect 3073 2533 3087 2547
rect 3113 2533 3127 2547
rect 3333 2533 3347 2547
rect 3013 2513 3027 2527
rect 3113 2513 3127 2527
rect 3073 2273 3087 2287
rect 2953 2093 2967 2107
rect 2953 2053 2967 2067
rect 2733 1853 2747 1867
rect 2613 1833 2627 1847
rect 2473 1613 2487 1627
rect 2513 1593 2527 1607
rect 2493 1333 2507 1347
rect 2453 1293 2467 1307
rect 2553 1293 2567 1307
rect 2493 1273 2507 1287
rect 2593 1253 2607 1267
rect 2313 1133 2327 1147
rect 2313 1113 2327 1127
rect 2013 873 2027 887
rect 1933 853 1947 867
rect 1973 853 1987 867
rect 1953 793 1967 807
rect 2033 813 2047 827
rect 1993 753 2007 767
rect 2153 1093 2167 1107
rect 2253 1093 2267 1107
rect 2433 1093 2447 1107
rect 2413 1073 2427 1087
rect 2453 1013 2467 1027
rect 2513 1013 2527 1027
rect 2253 873 2267 887
rect 2193 853 2207 867
rect 2293 853 2307 867
rect 2153 653 2167 667
rect 1893 593 1907 607
rect 2093 593 2107 607
rect 2053 353 2067 367
rect 1733 193 1747 207
rect 1873 153 1887 167
rect 1753 133 1767 147
rect 1913 313 1927 327
rect 2013 153 2027 167
rect 2153 353 2167 367
rect 2093 313 2107 327
rect 2273 833 2287 847
rect 2393 833 2407 847
rect 2273 633 2287 647
rect 2413 593 2427 607
rect 2493 373 2507 387
rect 2373 353 2387 367
rect 2473 353 2487 367
rect 2413 333 2427 347
rect 2433 313 2447 327
rect 2193 293 2207 307
rect 2153 153 2167 167
rect 2173 153 2187 167
rect 2273 153 2287 167
rect 1993 133 2007 147
rect 2533 873 2547 887
rect 2593 813 2607 827
rect 2553 613 2567 627
rect 2553 593 2567 607
rect 2673 1793 2687 1807
rect 2713 1793 2727 1807
rect 2813 1813 2827 1827
rect 2753 1793 2767 1807
rect 2753 1593 2767 1607
rect 2853 1613 2867 1627
rect 2753 1553 2767 1567
rect 2833 1553 2847 1567
rect 2773 1533 2787 1547
rect 2893 1333 2907 1347
rect 2833 1293 2847 1307
rect 2853 1273 2867 1287
rect 2793 1253 2807 1267
rect 2673 1153 2687 1167
rect 2733 1153 2747 1167
rect 2693 1093 2707 1107
rect 2713 1093 2727 1107
rect 2733 1053 2747 1067
rect 2673 633 2687 647
rect 2693 613 2707 627
rect 2753 1033 2767 1047
rect 2913 1093 2927 1107
rect 2913 993 2927 1007
rect 2833 853 2847 867
rect 2873 853 2887 867
rect 2853 813 2867 827
rect 2913 653 2927 667
rect 2633 553 2647 567
rect 2673 553 2687 567
rect 2613 393 2627 407
rect 2853 413 2867 427
rect 2513 253 2527 267
rect 2693 253 2707 267
rect 2513 193 2527 207
rect 1733 113 1747 127
rect 1893 113 1907 127
rect 2033 113 2047 127
rect 2493 113 2507 127
rect 2833 293 2847 307
rect 2973 1813 2987 1827
rect 2993 1793 3007 1807
rect 3033 1773 3047 1787
rect 2973 1613 2987 1627
rect 3093 1593 3107 1607
rect 3233 2293 3247 2307
rect 3293 2273 3307 2287
rect 3233 2253 3247 2267
rect 3273 2253 3287 2267
rect 3193 2133 3207 2147
rect 3413 2253 3427 2267
rect 3313 2233 3327 2247
rect 3613 3233 3627 3247
rect 3653 3193 3667 3207
rect 3733 3133 3747 3147
rect 3633 3053 3647 3067
rect 3633 3033 3647 3047
rect 3593 3013 3607 3027
rect 3613 2993 3627 3007
rect 3573 2973 3587 2987
rect 3553 2933 3567 2947
rect 3533 2253 3547 2267
rect 3213 2053 3227 2067
rect 3253 2053 3267 2067
rect 3433 1833 3447 1847
rect 3193 1813 3207 1827
rect 3273 1813 3287 1827
rect 3473 2133 3487 2147
rect 3513 2053 3527 2067
rect 3893 3713 3907 3727
rect 3893 3453 3907 3467
rect 3853 3293 3867 3307
rect 3753 2653 3767 2667
rect 4153 4213 4167 4227
rect 4193 4213 4207 4227
rect 4133 4193 4147 4207
rect 4233 4153 4247 4167
rect 4513 5033 4527 5047
rect 4713 5033 4727 5047
rect 4553 4973 4567 4987
rect 4373 4473 4387 4487
rect 4433 4473 4447 4487
rect 4733 4653 4747 4667
rect 4813 5033 4827 5047
rect 4773 4953 4787 4967
rect 5033 4713 5047 4727
rect 4933 4693 4947 4707
rect 4993 4693 5007 4707
rect 4493 4633 4507 4647
rect 4673 4493 4687 4507
rect 4493 4473 4507 4487
rect 4253 3973 4267 3987
rect 4153 3713 4167 3727
rect 4173 3693 4187 3707
rect 4173 3673 4187 3687
rect 4133 3473 4147 3487
rect 4093 3273 4107 3287
rect 4053 3233 4067 3247
rect 4093 3233 4107 3247
rect 4133 3233 4147 3247
rect 3933 3193 3947 3207
rect 3873 3173 3887 3187
rect 3893 3133 3907 3147
rect 3833 3033 3847 3047
rect 3933 3033 3947 3047
rect 3873 3013 3887 3027
rect 3913 3013 3927 3027
rect 4113 3213 4127 3227
rect 4073 3193 4087 3207
rect 3833 2753 3847 2767
rect 3873 2753 3887 2767
rect 4053 2753 4067 2767
rect 4093 2753 4107 2767
rect 3793 2713 3807 2727
rect 3793 2653 3807 2667
rect 3773 2633 3787 2647
rect 3633 2593 3647 2607
rect 3733 2573 3747 2587
rect 3773 2553 3787 2567
rect 3613 2293 3627 2307
rect 4193 3473 4207 3487
rect 4193 3273 4207 3287
rect 4173 3053 4187 3067
rect 4153 2613 4167 2627
rect 4093 2593 4107 2607
rect 3813 2573 3827 2587
rect 3873 2573 3887 2587
rect 4073 2573 4087 2587
rect 3933 2553 3947 2567
rect 3793 2273 3807 2287
rect 3813 2253 3827 2267
rect 3773 2233 3787 2247
rect 4113 2273 4127 2287
rect 3433 1793 3447 1807
rect 3453 1793 3467 1807
rect 3233 1773 3247 1787
rect 3453 1593 3467 1607
rect 3413 1573 3427 1587
rect 3053 1533 3067 1547
rect 3013 1353 3027 1367
rect 2973 1133 2987 1147
rect 3053 1293 3067 1307
rect 3133 1553 3147 1567
rect 3393 1553 3407 1567
rect 3413 1353 3427 1367
rect 3193 1333 3207 1347
rect 3353 1333 3367 1347
rect 3453 1333 3467 1347
rect 3153 1313 3167 1327
rect 3253 1313 3267 1327
rect 3133 1293 3147 1307
rect 3173 1293 3187 1307
rect 3193 1293 3207 1307
rect 3113 1253 3127 1267
rect 2993 1093 3007 1107
rect 3033 1093 3047 1107
rect 2993 1073 3007 1087
rect 2953 653 2967 667
rect 3193 1153 3207 1167
rect 3153 853 3167 867
rect 3133 833 3147 847
rect 3273 1253 3287 1267
rect 3313 1113 3327 1127
rect 3293 1073 3307 1087
rect 3433 1313 3447 1327
rect 3473 1253 3487 1267
rect 3413 1113 3427 1127
rect 3373 1073 3387 1087
rect 3853 1853 3867 1867
rect 3493 1073 3507 1087
rect 3253 773 3267 787
rect 3233 733 3247 747
rect 3073 673 3087 687
rect 2973 413 2987 427
rect 2933 373 2947 387
rect 2913 353 2927 367
rect 2973 333 2987 347
rect 3353 673 3367 687
rect 3433 793 3447 807
rect 3373 653 3387 667
rect 3413 593 3427 607
rect 3173 573 3187 587
rect 3053 293 3067 307
rect 3093 293 3107 307
rect 2553 133 2567 147
rect 2793 133 2807 147
rect 3113 133 3127 147
rect 2533 113 2547 127
rect 2833 113 2847 127
rect 3093 113 3107 127
rect 1473 93 1487 107
rect 1773 93 1787 107
rect 2573 93 2587 107
rect 3073 93 3087 107
rect 3033 73 3047 87
rect 3433 513 3447 527
rect 3393 313 3407 327
rect 3393 293 3407 307
rect 3373 133 3387 147
rect 3413 113 3427 127
rect 3133 73 3147 87
rect 3173 73 3187 87
rect 3573 1833 3587 1847
rect 3533 1813 3547 1827
rect 3553 1793 3567 1807
rect 3873 1773 3887 1787
rect 4053 1773 4067 1787
rect 3813 1753 3827 1767
rect 3833 1753 3847 1767
rect 3973 1753 3987 1767
rect 4013 1753 4027 1767
rect 3653 1613 3667 1627
rect 3793 1613 3807 1627
rect 3913 1613 3927 1627
rect 3673 1533 3687 1547
rect 3653 1513 3667 1527
rect 3733 1333 3747 1347
rect 3953 1593 3967 1607
rect 3933 1573 3947 1587
rect 3973 1573 3987 1587
rect 3833 1533 3847 1547
rect 3653 1313 3667 1327
rect 3693 1313 3707 1327
rect 3693 1293 3707 1307
rect 3673 1253 3687 1267
rect 3593 1113 3607 1127
rect 3553 393 3567 407
rect 3513 33 3527 47
rect 3613 1073 3627 1087
rect 3693 833 3707 847
rect 3793 1313 3807 1327
rect 3873 1293 3887 1307
rect 3873 1273 3887 1287
rect 3913 1273 3927 1287
rect 3853 1113 3867 1127
rect 3833 1093 3847 1107
rect 3893 1093 3907 1107
rect 3933 1073 3947 1087
rect 4073 1073 4087 1087
rect 3733 1053 3747 1067
rect 3733 833 3747 847
rect 3673 773 3687 787
rect 3713 773 3727 787
rect 3953 833 3967 847
rect 3913 813 3927 827
rect 3733 653 3747 667
rect 3613 633 3627 647
rect 3693 633 3707 647
rect 3733 633 3747 647
rect 3773 633 3787 647
rect 3713 613 3727 627
rect 3753 613 3767 627
rect 3773 593 3787 607
rect 3993 793 4007 807
rect 4033 613 4047 627
rect 4313 3713 4327 3727
rect 4693 4473 4707 4487
rect 4753 4473 4767 4487
rect 4473 4453 4487 4467
rect 4673 4453 4687 4467
rect 4433 4253 4447 4267
rect 4393 4193 4407 4207
rect 4413 4173 4427 4187
rect 4613 4173 4627 4187
rect 4673 4173 4687 4187
rect 4733 4453 4747 4467
rect 4413 4153 4427 4167
rect 4453 4153 4467 4167
rect 4553 4153 4567 4167
rect 4573 3993 4587 4007
rect 4373 3673 4387 3687
rect 4453 3733 4467 3747
rect 4513 3733 4527 3747
rect 4433 3713 4447 3727
rect 4433 3673 4447 3687
rect 4473 3533 4487 3547
rect 4393 3473 4407 3487
rect 4453 3473 4467 3487
rect 4413 3273 4427 3287
rect 4273 3253 4287 3267
rect 4393 3253 4407 3267
rect 4433 3253 4447 3267
rect 4473 3253 4487 3267
rect 4213 3233 4227 3247
rect 4213 3033 4227 3047
rect 4253 2593 4267 2607
rect 4413 3233 4427 3247
rect 4473 3193 4487 3207
rect 4473 3173 4487 3187
rect 4393 3033 4407 3047
rect 4333 2813 4347 2827
rect 4453 3013 4467 3027
rect 4453 2993 4467 3007
rect 4373 2593 4387 2607
rect 4393 2573 4407 2587
rect 4293 2553 4307 2567
rect 4333 2553 4347 2567
rect 4173 2293 4187 2307
rect 4193 2293 4207 2307
rect 4233 2293 4247 2307
rect 4273 2293 4287 2307
rect 4173 2073 4187 2087
rect 4153 1813 4167 1827
rect 4313 2253 4327 2267
rect 4413 2513 4427 2527
rect 4393 2253 4407 2267
rect 4353 2093 4367 2107
rect 4433 2093 4447 2107
rect 4493 2093 4507 2107
rect 4353 2073 4367 2087
rect 4393 2073 4407 2087
rect 4213 2053 4227 2067
rect 4293 2053 4307 2067
rect 4293 2013 4307 2027
rect 4333 2013 4347 2027
rect 4173 1793 4187 1807
rect 4173 1613 4187 1627
rect 4233 1573 4247 1587
rect 4173 1553 4187 1567
rect 4213 1553 4227 1567
rect 4253 1553 4267 1567
rect 4173 1353 4187 1367
rect 4253 1353 4267 1367
rect 4133 1133 4147 1147
rect 4213 1333 4227 1347
rect 4233 1313 4247 1327
rect 4153 1093 4167 1107
rect 4213 1053 4227 1067
rect 4253 853 4267 867
rect 4353 1793 4367 1807
rect 4393 1793 4407 1807
rect 4453 2073 4467 2087
rect 4373 1773 4387 1787
rect 4413 1773 4427 1787
rect 4433 1773 4447 1787
rect 4433 1753 4447 1767
rect 4353 1593 4367 1607
rect 4393 1593 4407 1607
rect 4433 1593 4447 1607
rect 4473 1593 4487 1607
rect 4473 1553 4487 1567
rect 4333 1533 4347 1547
rect 4413 1293 4427 1307
rect 4573 3693 4587 3707
rect 4613 3693 4627 3707
rect 4633 3693 4647 3707
rect 4673 3693 4687 3707
rect 4593 3433 4607 3447
rect 4573 2073 4587 2087
rect 4373 1273 4387 1287
rect 4213 813 4227 827
rect 4293 813 4307 827
rect 4193 793 4207 807
rect 4453 1273 4467 1287
rect 4493 1093 4507 1107
rect 4513 1073 4527 1087
rect 4433 1033 4447 1047
rect 4533 853 4547 867
rect 4733 3693 4747 3707
rect 4673 3533 4687 3547
rect 4713 3533 4727 3547
rect 4813 3993 4827 4007
rect 4873 3953 4887 3967
rect 4793 3673 4807 3687
rect 4893 3513 4907 3527
rect 4693 3493 4707 3507
rect 4733 3493 4747 3507
rect 4773 3493 4787 3507
rect 4713 3293 4727 3307
rect 4613 2573 4627 2587
rect 4693 3193 4707 3207
rect 4733 3013 4747 3027
rect 4673 2713 4687 2727
rect 4693 2613 4707 2627
rect 4753 2613 4767 2627
rect 4653 2593 4667 2607
rect 4633 2513 4647 2527
rect 4753 2593 4767 2607
rect 4713 2313 4727 2327
rect 4753 2293 4767 2307
rect 4993 4473 5007 4487
rect 4993 4173 5007 4187
rect 4953 4153 4967 4167
rect 4953 3693 4967 3707
rect 4993 3693 5007 3707
rect 4953 3513 4967 3527
rect 4913 3253 4927 3267
rect 4893 3213 4907 3227
rect 4973 3473 4987 3487
rect 4973 3213 4987 3227
rect 5033 4653 5047 4667
rect 5013 3093 5027 3107
rect 5073 3093 5087 3107
rect 4973 3073 4987 3087
rect 5053 3073 5067 3087
rect 4953 3053 4967 3067
rect 4933 3033 4947 3047
rect 4913 2713 4927 2727
rect 4873 2673 4887 2687
rect 4833 2533 4847 2547
rect 4733 2273 4747 2287
rect 4773 2273 4787 2287
rect 4693 2073 4707 2087
rect 4473 833 4487 847
rect 4593 833 4607 847
rect 4513 813 4527 827
rect 4413 673 4427 687
rect 4113 613 4127 627
rect 4293 613 4307 627
rect 4093 593 4107 607
rect 4013 573 4027 587
rect 3913 513 3927 527
rect 3713 393 3727 407
rect 3653 373 3667 387
rect 3673 373 3687 387
rect 3993 373 4007 387
rect 3693 353 3707 367
rect 3953 353 3967 367
rect 4233 393 4247 407
rect 4013 333 4027 347
rect 4093 333 4107 347
rect 4153 333 4167 347
rect 4433 333 4447 347
rect 4513 373 4527 387
rect 3973 313 3987 327
rect 4113 313 4127 327
rect 3973 153 3987 167
rect 4113 153 4127 167
rect 4233 153 4247 167
rect 4453 153 4467 167
rect 3693 133 3707 147
rect 3953 133 3967 147
rect 4033 133 4047 147
rect 4493 133 4507 147
rect 3673 113 3687 127
rect 3573 93 3587 107
rect 3993 113 4007 127
rect 4513 113 4527 127
rect 3713 73 3727 87
rect 3593 33 3607 47
rect 4653 1813 4667 1827
rect 4933 2673 4947 2687
rect 4953 2593 4967 2607
rect 4893 2533 4907 2547
rect 4933 2513 4947 2527
rect 4913 2313 4927 2327
rect 4873 2253 4887 2267
rect 4713 1813 4727 1827
rect 4673 1793 4687 1807
rect 4753 1693 4767 1707
rect 4793 1693 4807 1707
rect 4853 2033 4867 2047
rect 5053 3053 5067 3067
rect 5013 3033 5027 3047
rect 4993 3013 5007 3027
rect 5033 2993 5047 3007
rect 4953 2293 4967 2307
rect 4973 2293 4987 2307
rect 5053 2293 5067 2307
rect 4933 2273 4947 2287
rect 4993 2273 5007 2287
rect 5033 2273 5047 2287
rect 4933 2233 4947 2247
rect 5013 2253 5027 2267
rect 4953 2033 4967 2047
rect 4833 1773 4847 1787
rect 4913 1773 4927 1787
rect 4973 1773 4987 1787
rect 4813 1593 4827 1607
rect 4693 1553 4707 1567
rect 4773 1573 4787 1587
rect 4733 1513 4747 1527
rect 4733 1313 4747 1327
rect 4753 1293 4767 1307
rect 5013 1573 5027 1587
rect 5033 1553 5047 1567
rect 5073 2273 5087 2287
rect 4893 1293 4907 1307
rect 5013 1293 5027 1307
rect 5053 1293 5067 1307
rect 4833 1273 4847 1287
rect 4933 1273 4947 1287
rect 4773 1233 4787 1247
rect 5013 1233 5027 1247
rect 4713 1113 4727 1127
rect 4753 1113 4767 1127
rect 4713 1093 4727 1107
rect 4693 1073 4707 1087
rect 4753 1073 4767 1087
rect 4993 1073 5007 1087
rect 4833 853 4847 867
rect 4973 853 4987 867
rect 4813 833 4827 847
rect 4673 653 4687 667
rect 4733 653 4747 667
rect 4693 593 4707 607
rect 4733 393 4747 407
rect 4773 373 4787 387
rect 4953 593 4967 607
rect 4753 353 4767 367
rect 4793 353 4807 367
rect 5033 373 5047 387
rect 4773 253 4787 267
rect 4953 233 4967 247
rect 5013 233 5027 247
rect 4813 133 4827 147
rect 4753 113 4767 127
rect 5013 133 5027 147
rect 5033 113 5047 127
rect 4953 13 4967 27
rect 4993 13 5007 27
<< metal3 >>
rect 4427 5036 4513 5044
rect 4727 5036 4813 5044
rect 707 4976 1213 4984
rect 1327 4976 1533 4984
rect 1807 4976 1893 4984
rect 3767 4976 3973 4984
rect 3996 4976 4233 4984
rect 527 4956 653 4964
rect 1047 4956 1173 4964
rect 1827 4956 1953 4964
rect 2627 4956 2653 4964
rect 2707 4956 3093 4964
rect 3996 4964 4004 4976
rect 4287 4976 4553 4984
rect 3227 4956 4004 4964
rect 4167 4956 4773 4964
rect 227 4936 493 4944
rect 867 4936 1013 4944
rect 1107 4936 1553 4944
rect 1567 4936 1573 4944
rect 2127 4936 2353 4944
rect 2407 4936 2673 4944
rect 2727 4936 2953 4944
rect -24 4916 193 4924
rect 247 4916 573 4924
rect 1867 4916 2413 4924
rect 2947 4916 3213 4924
rect 247 4896 533 4904
rect 547 4896 1733 4904
rect 1907 4876 2133 4884
rect 527 4716 3573 4724
rect 787 4696 1473 4704
rect 2527 4696 2613 4704
rect 2627 4696 2853 4704
rect 2867 4696 2973 4704
rect 3247 4696 3473 4704
rect 3487 4696 3633 4704
rect 4947 4696 4993 4704
rect 787 4676 813 4684
rect 1407 4676 1953 4684
rect 1967 4676 2093 4684
rect 2247 4676 2773 4684
rect 2907 4676 3353 4684
rect 3367 4676 3933 4684
rect 4227 4676 4253 4684
rect 587 4656 593 4664
rect 607 4656 793 4664
rect 807 4656 1053 4664
rect 1067 4656 1113 4664
rect 1947 4656 2153 4664
rect 2167 4656 2453 4664
rect 2816 4664 2824 4673
rect 5036 4667 5044 4713
rect 2547 4656 2824 4664
rect 2847 4656 2973 4664
rect 3927 4656 4153 4664
rect 4207 4656 4733 4664
rect 567 4636 1133 4644
rect 1687 4636 2193 4644
rect 2207 4636 2493 4644
rect 3127 4636 3333 4644
rect 3667 4636 3993 4644
rect 4247 4636 4493 4644
rect 1747 4616 1973 4624
rect 3027 4616 3153 4624
rect 3167 4616 3613 4624
rect 3627 4616 3673 4624
rect 3967 4616 4233 4624
rect 1167 4596 3013 4604
rect 1427 4536 1553 4544
rect 1567 4536 1613 4544
rect 1387 4516 1693 4524
rect 1907 4516 2553 4524
rect 267 4496 313 4504
rect 747 4496 1053 4504
rect 1067 4496 1373 4504
rect 1487 4496 1933 4504
rect 2907 4496 3133 4504
rect 3147 4496 3233 4504
rect 3687 4496 3873 4504
rect 4007 4496 4673 4504
rect 447 4476 493 4484
rect 527 4476 573 4484
rect 1047 4476 1093 4484
rect 1427 4476 1473 4484
rect 1687 4476 2513 4484
rect 2687 4476 2853 4484
rect 3027 4476 3093 4484
rect 3216 4476 3373 4484
rect 327 4456 1073 4464
rect 1607 4456 1653 4464
rect 1967 4456 2213 4464
rect 2516 4456 2813 4464
rect 247 4436 453 4444
rect 587 4436 793 4444
rect 2207 4436 2233 4444
rect 2516 4444 2524 4456
rect 3216 4464 3224 4476
rect 3407 4476 3533 4484
rect 3587 4476 3613 4484
rect 4387 4476 4433 4484
rect 4507 4476 4693 4484
rect 4767 4476 4993 4484
rect 2856 4456 3224 4464
rect 2287 4436 2524 4444
rect 2856 4444 2864 4456
rect 3247 4456 3413 4464
rect 3467 4456 3893 4464
rect 3907 4456 4473 4464
rect 4687 4456 4733 4464
rect 2847 4436 2864 4444
rect 4207 4436 4233 4444
rect 787 4416 813 4424
rect 2536 4424 2544 4433
rect 2327 4416 2693 4424
rect 2876 4424 2884 4433
rect 2827 4416 2884 4424
rect 3247 4316 4153 4324
rect 1587 4256 4433 4264
rect 267 4236 293 4244
rect 307 4236 533 4244
rect 547 4236 733 4244
rect 1147 4236 1393 4244
rect 1927 4236 1973 4244
rect 1987 4236 2073 4244
rect 2447 4236 2493 4244
rect 2587 4236 3273 4244
rect 3607 4236 3853 4244
rect 227 4216 273 4224
rect 507 4216 644 4224
rect 247 4196 433 4204
rect 527 4196 573 4204
rect 636 4204 644 4216
rect 1027 4216 1073 4224
rect 1287 4216 1353 4224
rect 1967 4216 2113 4224
rect 2127 4216 2153 4224
rect 2427 4216 2453 4224
rect 2707 4216 2773 4224
rect 3507 4216 3893 4224
rect 4167 4216 4193 4224
rect 636 4196 793 4204
rect 807 4196 1093 4204
rect 1387 4196 1653 4204
rect 2187 4196 2313 4204
rect 2487 4196 2673 4204
rect 2727 4196 2784 4204
rect 1647 4176 1893 4184
rect 1947 4176 2413 4184
rect 2427 4176 2753 4184
rect 2776 4184 2784 4196
rect 2807 4196 3033 4204
rect 3307 4196 3393 4204
rect 3427 4196 3533 4204
rect 4147 4196 4393 4204
rect 2776 4176 3573 4184
rect 4427 4176 4604 4184
rect 3067 4156 3333 4164
rect 4247 4156 4413 4164
rect 4427 4156 4453 4164
rect 4467 4156 4553 4164
rect 4596 4164 4604 4176
rect 4627 4176 4673 4184
rect 5116 4184 5124 4204
rect 5007 4176 5124 4184
rect 4596 4156 4953 4164
rect 1627 4136 2113 4144
rect 3687 4096 3873 4104
rect 287 4036 513 4044
rect 527 4036 533 4044
rect 547 4036 773 4044
rect 267 4016 1273 4024
rect 1587 4016 1833 4024
rect 2107 4016 2213 4024
rect 2227 4016 2433 4024
rect 3547 4016 3973 4024
rect 247 3996 313 4004
rect 1007 3996 1133 4004
rect 1147 3996 1233 4004
rect 1327 3996 1873 4004
rect 2687 3996 3093 4004
rect 3147 3996 3613 4004
rect 3627 3996 3633 4004
rect 4587 3996 4813 4004
rect 507 3976 833 3984
rect 847 3976 973 3984
rect 1027 3976 1853 3984
rect 2167 3976 2193 3984
rect 2427 3976 2453 3984
rect 2707 3976 2973 3984
rect 4007 3976 4253 3984
rect 1907 3956 1973 3964
rect 2067 3956 2653 3964
rect 3007 3956 3213 3964
rect 4887 3956 5124 3964
rect 1856 3944 1864 3953
rect 1856 3936 1873 3944
rect 1687 3916 1813 3924
rect 1827 3916 2173 3924
rect 747 3776 1073 3784
rect 1087 3776 1533 3784
rect 827 3756 1113 3764
rect 287 3736 433 3744
rect 447 3736 553 3744
rect 2827 3736 2953 3744
rect 2967 3736 3133 3744
rect 3147 3736 3193 3744
rect 3207 3736 3473 3744
rect 247 3716 533 3724
rect 767 3716 813 3724
rect 867 3716 1093 3724
rect 1887 3716 1913 3724
rect 2127 3716 2233 3724
rect 2547 3716 3053 3724
rect 3187 3716 3613 3724
rect 3627 3716 3884 3724
rect 307 3696 793 3704
rect 1307 3696 1393 3704
rect 1407 3696 1553 3704
rect 1747 3696 1893 3704
rect 1907 3696 2033 3704
rect 2047 3696 2253 3704
rect 3096 3704 3104 3713
rect 2847 3696 3104 3704
rect 3127 3696 3253 3704
rect 3876 3704 3884 3716
rect 3916 3724 3924 3753
rect 4467 3736 4513 3744
rect 3907 3716 3924 3724
rect 4327 3716 4433 3724
rect 4156 3704 4164 3713
rect 3876 3696 4164 3704
rect 4187 3696 4573 3704
rect 4627 3696 4633 3704
rect 4647 3696 4673 3704
rect 4747 3696 4953 3704
rect 5116 3704 5124 3724
rect 5007 3696 5124 3704
rect 647 3676 833 3684
rect 1247 3676 1373 3684
rect 1687 3676 1953 3684
rect 1967 3676 2113 3684
rect 2227 3676 2473 3684
rect 2487 3676 2753 3684
rect 3407 3676 3593 3684
rect 4187 3676 4373 3684
rect 4447 3676 4793 3684
rect 1367 3656 1633 3664
rect 2507 3656 2793 3664
rect 107 3596 253 3604
rect 2627 3596 2993 3604
rect 1067 3556 1673 3564
rect 167 3536 653 3544
rect 667 3536 673 3544
rect 687 3536 1173 3544
rect 1187 3536 1193 3544
rect 2147 3536 2173 3544
rect 3167 3536 3293 3544
rect 3316 3536 3473 3544
rect 227 3516 493 3524
rect 1027 3516 1153 3524
rect 1287 3516 1353 3524
rect 2367 3516 2424 3524
rect 487 3496 513 3504
rect 907 3496 993 3504
rect 2087 3496 2393 3504
rect 2416 3504 2424 3516
rect 2707 3516 3113 3524
rect 3316 3524 3324 3536
rect 4487 3536 4673 3544
rect 4687 3536 4713 3544
rect 3247 3516 3324 3524
rect 4907 3516 4953 3524
rect 2416 3496 2713 3504
rect 2767 3496 3493 3504
rect 3507 3496 4693 3504
rect 4747 3496 4773 3504
rect 1947 3476 2373 3484
rect 2427 3476 2653 3484
rect 3307 3476 3653 3484
rect 3667 3476 3753 3484
rect 4147 3476 4193 3484
rect 4207 3476 4393 3484
rect 4407 3476 4453 3484
rect 4987 3476 5124 3484
rect 227 3456 313 3464
rect 327 3456 453 3464
rect 1547 3456 2493 3464
rect 3767 3456 3893 3464
rect 447 3436 453 3444
rect 467 3436 493 3444
rect 3347 3436 4593 3444
rect 267 3316 2633 3324
rect 2647 3316 3753 3324
rect 747 3296 1073 3304
rect 1087 3296 1613 3304
rect 2567 3296 3853 3304
rect 4727 3296 5124 3304
rect 1127 3276 4093 3284
rect 4207 3276 4413 3284
rect 747 3256 753 3264
rect 767 3256 1033 3264
rect 1047 3256 1093 3264
rect 1516 3256 1533 3264
rect 427 3236 453 3244
rect 787 3236 1053 3244
rect 1516 3227 1524 3256
rect 1767 3256 1793 3264
rect 1807 3256 1833 3264
rect 2407 3256 2853 3264
rect 3067 3256 3193 3264
rect 3207 3256 3313 3264
rect 3367 3256 3533 3264
rect 3547 3256 3593 3264
rect 4036 3256 4144 3264
rect 1547 3236 1733 3244
rect 2487 3236 2773 3244
rect 4036 3244 4044 3256
rect 4136 3247 4144 3256
rect 4287 3256 4393 3264
rect 4447 3256 4473 3264
rect 4927 3256 5124 3264
rect 3627 3236 4044 3244
rect 4067 3236 4093 3244
rect 4227 3236 4413 3244
rect 447 3216 713 3224
rect 1587 3216 1693 3224
rect 1987 3216 2373 3224
rect 2427 3216 2453 3224
rect 2987 3216 3073 3224
rect 3087 3216 3353 3224
rect 4127 3216 4893 3224
rect 4987 3216 5124 3224
rect 107 3196 473 3204
rect 647 3196 753 3204
rect 1187 3196 1553 3204
rect 2027 3196 2473 3204
rect 3667 3196 3933 3204
rect 3947 3196 4073 3204
rect 4087 3196 4473 3204
rect 4487 3196 4693 3204
rect 1807 3176 1813 3184
rect 1827 3176 2093 3184
rect 2367 3176 2773 3184
rect 3887 3176 4473 3184
rect 147 3156 153 3164
rect 167 3156 353 3164
rect 2727 3156 3073 3164
rect 3747 3136 3893 3144
rect 5027 3096 5073 3104
rect 1467 3076 2553 3084
rect 4987 3076 5053 3084
rect -24 3056 73 3064
rect 1967 3056 2033 3064
rect 2107 3056 2293 3064
rect 3647 3056 4173 3064
rect 4967 3056 5053 3064
rect 2007 3036 2073 3044
rect 2987 3036 3013 3044
rect 3027 3036 3033 3044
rect 3367 3036 3633 3044
rect 3847 3036 3933 3044
rect 3947 3036 4213 3044
rect 4227 3036 4393 3044
rect 4947 3036 5013 3044
rect -24 3016 233 3024
rect 647 3016 793 3024
rect 947 3016 1153 3024
rect 1867 3016 1973 3024
rect 2027 3016 2093 3024
rect 2276 3024 2284 3033
rect 2276 3016 2293 3024
rect 3607 3016 3873 3024
rect 3927 3016 4453 3024
rect 4747 3016 4993 3024
rect 687 2996 913 3004
rect 1827 2996 2393 3004
rect 2807 2996 2853 3004
rect 3107 2996 3613 3004
rect 4467 2996 5033 3004
rect 887 2976 1013 2984
rect 1027 2976 1713 2984
rect 2287 2976 2333 2984
rect 2347 2976 3573 2984
rect 847 2956 1673 2964
rect 1687 2956 1773 2964
rect 927 2936 2753 2944
rect 2767 2936 3553 2944
rect 3247 2836 3333 2844
rect 2167 2816 4333 2824
rect 1187 2796 1313 2804
rect 1327 2796 3293 2804
rect 3307 2796 3333 2804
rect 707 2776 1113 2784
rect 1287 2776 1393 2784
rect 2087 2776 2113 2784
rect 3307 2776 3473 2784
rect 467 2756 853 2764
rect 1007 2756 1033 2764
rect 1316 2756 1813 2764
rect 167 2736 373 2744
rect 587 2736 973 2744
rect 1027 2736 1173 2744
rect 1316 2744 1324 2756
rect 1847 2756 2133 2764
rect 2407 2756 2673 2764
rect 3027 2756 3833 2764
rect 3887 2756 4053 2764
rect 4067 2756 4093 2764
rect 1307 2736 1324 2744
rect 1347 2736 1433 2744
rect 2107 2736 2653 2744
rect 2667 2736 3093 2744
rect 3287 2736 3413 2744
rect 387 2716 613 2724
rect 1107 2716 1193 2724
rect 1567 2716 1753 2724
rect 2747 2716 3793 2724
rect 4687 2716 4913 2724
rect 267 2696 373 2704
rect 867 2696 1573 2704
rect 1587 2696 2353 2704
rect 2367 2696 2493 2704
rect 247 2676 453 2684
rect 467 2676 1533 2684
rect 1547 2676 1633 2684
rect 4887 2676 4933 2684
rect 107 2656 253 2664
rect 347 2656 533 2664
rect 3767 2656 3793 2664
rect 2107 2636 2473 2644
rect 2487 2636 2693 2644
rect 2707 2636 2913 2644
rect 2927 2636 3433 2644
rect 3447 2636 3453 2644
rect 3467 2636 3773 2644
rect 2807 2616 3353 2624
rect 3367 2616 4153 2624
rect 4707 2616 4753 2624
rect 1947 2596 2433 2604
rect 2447 2596 2473 2604
rect 3647 2596 4093 2604
rect 4267 2596 4373 2604
rect 4667 2596 4753 2604
rect 4767 2596 4953 2604
rect 307 2576 633 2584
rect 1107 2576 1313 2584
rect 1327 2576 1353 2584
rect 1907 2576 1913 2584
rect 1927 2576 2213 2584
rect 3747 2576 3813 2584
rect 3887 2576 4073 2584
rect 4407 2576 4613 2584
rect 247 2556 313 2564
rect 507 2556 544 2564
rect 287 2536 513 2544
rect 536 2544 544 2556
rect 1687 2556 1973 2564
rect 2667 2556 3053 2564
rect 3787 2556 3933 2564
rect 3947 2556 4293 2564
rect 4307 2556 4333 2564
rect 536 2536 713 2544
rect 727 2536 813 2544
rect 1187 2536 1373 2544
rect 1667 2536 1873 2544
rect 1887 2536 1953 2544
rect 2247 2536 2293 2544
rect 2547 2536 2673 2544
rect 3007 2536 3073 2544
rect 3127 2536 3333 2544
rect 4847 2536 4893 2544
rect 1147 2516 1333 2524
rect 3027 2516 3113 2524
rect 4427 2516 4633 2524
rect 4647 2516 4933 2524
rect 1867 2316 1913 2324
rect 4727 2316 4913 2324
rect 1107 2296 1493 2304
rect 1587 2296 1873 2304
rect 2427 2296 2664 2304
rect 447 2276 513 2284
rect 527 2276 773 2284
rect 827 2276 853 2284
rect 1027 2276 1073 2284
rect 1647 2276 1693 2284
rect 1907 2276 2053 2284
rect 2167 2276 2233 2284
rect 2247 2276 2393 2284
rect 2407 2276 2453 2284
rect 2656 2284 2664 2296
rect 2687 2296 2744 2304
rect 2736 2287 2744 2296
rect 2767 2296 3233 2304
rect 3627 2296 4173 2304
rect 4187 2296 4193 2304
rect 4247 2296 4273 2304
rect 4767 2296 4953 2304
rect 4987 2296 5053 2304
rect 2656 2276 2713 2284
rect 3087 2276 3293 2284
rect 3807 2276 4113 2284
rect 4747 2276 4773 2284
rect 4947 2276 4993 2284
rect 5047 2276 5073 2284
rect 327 2256 493 2264
rect 547 2256 753 2264
rect 1367 2256 1613 2264
rect 2707 2256 2733 2264
rect 2947 2256 3233 2264
rect 3287 2256 3413 2264
rect 3547 2256 3813 2264
rect 4327 2256 4393 2264
rect 4887 2256 5013 2264
rect 247 2236 473 2244
rect 487 2236 533 2244
rect 587 2236 793 2244
rect 1607 2236 1793 2244
rect 2287 2236 2473 2244
rect 2816 2244 2824 2253
rect 2487 2236 2933 2244
rect 3327 2236 3773 2244
rect 3787 2236 4933 2244
rect 2047 2216 2153 2224
rect 767 2136 2093 2144
rect 2107 2136 2193 2144
rect 2207 2136 3193 2144
rect 3207 2136 3473 2144
rect 2187 2116 2233 2124
rect 2247 2116 2433 2124
rect 447 2096 513 2104
rect 927 2096 1293 2104
rect 1327 2096 1513 2104
rect 2047 2096 2953 2104
rect 4367 2096 4433 2104
rect 4447 2096 4493 2104
rect 767 2076 893 2084
rect 1647 2076 1693 2084
rect 1707 2076 1833 2084
rect 4187 2076 4353 2084
rect 4407 2076 4453 2084
rect 4587 2076 4693 2084
rect 287 2056 353 2064
rect 367 2056 493 2064
rect 2187 2056 2413 2064
rect 2427 2056 2653 2064
rect 2716 2064 2724 2073
rect 2716 2056 2953 2064
rect 2967 2056 3213 2064
rect 3267 2056 3513 2064
rect 4227 2056 4293 2064
rect 1327 2036 1553 2044
rect 1567 2036 1633 2044
rect 1687 2036 2473 2044
rect 2487 2036 2693 2044
rect 4867 2036 4953 2044
rect 4307 2016 4333 2024
rect 227 1996 2393 2004
rect 1047 1976 1353 1984
rect 1607 1876 1793 1884
rect 1807 1876 1833 1884
rect 2747 1856 3853 1864
rect 1787 1836 2193 1844
rect 2207 1836 2613 1844
rect 3447 1836 3573 1844
rect 867 1816 1293 1824
rect 1347 1816 1904 1824
rect 1896 1807 1904 1816
rect 2107 1816 2153 1824
rect 2827 1816 2973 1824
rect 2987 1816 3193 1824
rect 3287 1816 3533 1824
rect 4167 1816 4653 1824
rect 4667 1816 4713 1824
rect 267 1796 333 1804
rect 347 1796 513 1804
rect 1067 1796 1273 1804
rect 1327 1796 1353 1804
rect 1367 1796 1593 1804
rect 2127 1796 2173 1804
rect 2407 1796 2673 1804
rect 2727 1796 2753 1804
rect 3007 1796 3433 1804
rect 3467 1796 3553 1804
rect 4187 1796 4353 1804
rect 4407 1796 4673 1804
rect 287 1776 313 1784
rect 327 1776 473 1784
rect 487 1776 493 1784
rect 567 1776 793 1784
rect 807 1776 2453 1784
rect 2467 1776 3033 1784
rect 3047 1776 3233 1784
rect 3887 1776 4053 1784
rect 4387 1776 4413 1784
rect 4447 1776 4833 1784
rect 4927 1776 4973 1784
rect 127 1756 253 1764
rect 1347 1756 1873 1764
rect 1947 1756 3813 1764
rect 3847 1756 3973 1764
rect 4027 1756 4433 1764
rect 567 1736 673 1744
rect 4767 1696 4793 1704
rect 1047 1656 1393 1664
rect 827 1636 1473 1644
rect 1487 1636 1913 1644
rect 1927 1636 2453 1644
rect 1087 1616 1693 1624
rect 2487 1616 2853 1624
rect 2867 1616 2973 1624
rect 3667 1616 3793 1624
rect 3927 1616 4173 1624
rect 307 1596 453 1604
rect 607 1596 693 1604
rect 907 1596 1413 1604
rect 1427 1596 1533 1604
rect 1967 1596 2153 1604
rect 2167 1596 2233 1604
rect 2267 1596 2293 1604
rect 2527 1596 2744 1604
rect 287 1576 353 1584
rect 367 1576 573 1584
rect 1667 1576 1773 1584
rect 1787 1576 1933 1584
rect 1947 1576 2173 1584
rect 2736 1584 2744 1596
rect 2767 1596 3093 1604
rect 3396 1596 3453 1604
rect 3396 1584 3404 1596
rect 3967 1596 4353 1604
rect 4407 1596 4433 1604
rect 4487 1596 4813 1604
rect 2736 1576 3404 1584
rect 3427 1576 3933 1584
rect 3987 1576 4233 1584
rect 4787 1576 5013 1584
rect 847 1556 1133 1564
rect 1376 1564 1384 1573
rect 1376 1556 1633 1564
rect 1687 1556 1733 1564
rect 2227 1556 2333 1564
rect 2347 1556 2433 1564
rect 2767 1556 2833 1564
rect 3147 1556 3393 1564
rect 4187 1556 4213 1564
rect 4267 1556 4473 1564
rect 4707 1556 5033 1564
rect 2787 1536 3053 1544
rect 3687 1536 3833 1544
rect 3847 1536 4333 1544
rect 3667 1516 4733 1524
rect 3027 1356 3413 1364
rect 4187 1356 4253 1364
rect 427 1336 573 1344
rect 587 1336 633 1344
rect 687 1336 833 1344
rect 867 1336 1033 1344
rect 1127 1336 1193 1344
rect 1747 1336 1873 1344
rect 2307 1336 2493 1344
rect 2907 1336 3193 1344
rect 3367 1336 3453 1344
rect 3747 1336 4213 1344
rect 167 1316 233 1324
rect 247 1316 364 1324
rect 356 1304 364 1316
rect 387 1316 613 1324
rect 807 1316 844 1324
rect 356 1296 673 1304
rect 687 1296 713 1304
rect 727 1296 813 1304
rect 836 1304 844 1316
rect 1047 1316 1153 1324
rect 1487 1316 1613 1324
rect 1627 1316 1753 1324
rect 2836 1316 3153 1324
rect 2836 1307 2844 1316
rect 3167 1316 3253 1324
rect 3447 1316 3653 1324
rect 3707 1316 3793 1324
rect 4247 1316 4733 1324
rect 836 1296 1173 1304
rect 1447 1296 1533 1304
rect 1867 1296 2053 1304
rect 2467 1296 2553 1304
rect 3067 1296 3133 1304
rect 3187 1296 3193 1304
rect 3207 1296 3693 1304
rect 3887 1296 4413 1304
rect 4767 1296 4893 1304
rect 5027 1296 5053 1304
rect 247 1276 333 1284
rect 2507 1276 2853 1284
rect 3887 1276 3913 1284
rect 4387 1276 4453 1284
rect 4847 1276 4933 1284
rect 2607 1256 2793 1264
rect 2807 1256 3113 1264
rect 3127 1256 3273 1264
rect 3287 1256 3473 1264
rect 3487 1256 3673 1264
rect 4787 1236 5013 1244
rect 527 1156 653 1164
rect 2067 1156 2673 1164
rect 2687 1156 2733 1164
rect 2747 1156 3193 1164
rect 467 1136 1213 1144
rect 1307 1136 1473 1144
rect 2107 1136 2313 1144
rect 2987 1136 4133 1144
rect 507 1116 633 1124
rect 767 1116 833 1124
rect 847 1116 1453 1124
rect 1567 1116 1793 1124
rect 1847 1116 2133 1124
rect 2327 1116 3313 1124
rect 3327 1116 3413 1124
rect 3607 1116 3853 1124
rect 4727 1116 4753 1124
rect 487 1096 573 1104
rect 1227 1096 1273 1104
rect 1407 1096 1513 1104
rect 1527 1096 1573 1104
rect 2167 1096 2253 1104
rect 2447 1096 2693 1104
rect 2927 1096 2993 1104
rect 3847 1096 3893 1104
rect 3907 1096 4153 1104
rect 4507 1096 4713 1104
rect 927 1076 1053 1084
rect 1067 1076 1613 1084
rect 1867 1076 2413 1084
rect 1816 1064 1824 1073
rect 1816 1056 1833 1064
rect 2716 1064 2724 1093
rect 3036 1084 3044 1093
rect 3007 1076 3044 1084
rect 3307 1076 3373 1084
rect 3507 1076 3613 1084
rect 3627 1076 3933 1084
rect 3947 1076 4073 1084
rect 4527 1076 4693 1084
rect 4767 1076 4993 1084
rect 2716 1056 2733 1064
rect 3747 1056 4213 1064
rect 2767 1036 4433 1044
rect 2467 1016 2513 1024
rect 1947 996 2913 1004
rect 1247 876 2013 884
rect 2267 876 2533 884
rect 47 856 73 864
rect 87 856 233 864
rect 1027 856 1113 864
rect 1127 856 1193 864
rect 1207 856 1433 864
rect 1947 856 1973 864
rect 2207 856 2293 864
rect 2307 856 2833 864
rect 2887 856 3153 864
rect 4267 856 4533 864
rect 4847 856 4973 864
rect 147 836 473 844
rect 487 836 753 844
rect 767 836 993 844
rect 1167 836 1413 844
rect 1847 836 2273 844
rect 2407 836 3133 844
rect 3707 836 3733 844
rect 3967 836 4473 844
rect 4607 836 4813 844
rect 167 816 273 824
rect 287 816 313 824
rect 587 816 853 824
rect 867 816 1573 824
rect 1627 816 1673 824
rect 2047 816 2593 824
rect 2607 816 2853 824
rect 3927 816 4213 824
rect 4307 816 4513 824
rect 747 796 813 804
rect 1707 796 1953 804
rect 3447 796 3993 804
rect 4007 796 4193 804
rect 1527 776 1713 784
rect 3267 776 3673 784
rect 3687 776 3713 784
rect 1827 756 1993 764
rect 727 736 773 744
rect 787 736 1093 744
rect 1107 736 3233 744
rect 967 676 1133 684
rect 1267 676 1273 684
rect 1287 676 1593 684
rect 3087 676 3353 684
rect 3367 676 4413 684
rect 267 656 453 664
rect 1007 656 1173 664
rect 1187 656 1213 664
rect 1567 656 1853 664
rect 1867 656 2153 664
rect 2927 656 2953 664
rect 2967 656 3373 664
rect 3716 656 3733 664
rect 1087 636 1513 644
rect 2287 636 2673 644
rect 3627 636 3693 644
rect 3716 627 3724 656
rect 4687 656 4733 664
rect 3747 636 3773 644
rect 547 616 833 624
rect 1147 616 1233 624
rect 2567 616 2693 624
rect 3767 616 4033 624
rect 4127 616 4293 624
rect 487 596 493 604
rect 507 596 513 604
rect 527 596 793 604
rect 1907 596 2093 604
rect 2427 596 2553 604
rect 3427 596 3773 604
rect 4107 596 4693 604
rect 4707 596 4953 604
rect 3187 576 4013 584
rect 2647 556 2673 564
rect 3447 516 3913 524
rect 2867 416 2973 424
rect 2627 396 3553 404
rect 3567 396 3713 404
rect 4247 396 4733 404
rect 1327 376 1413 384
rect 2507 376 2933 384
rect 2947 376 3653 384
rect 3667 376 3673 384
rect 3687 376 3993 384
rect 4527 376 4773 384
rect 4787 376 5033 384
rect 467 356 493 364
rect 1207 356 1333 364
rect 2067 356 2153 364
rect 2167 356 2373 364
rect 2487 356 2913 364
rect 3707 356 3953 364
rect 4767 356 4793 364
rect 507 336 1013 344
rect 1087 336 1373 344
rect 1387 336 1653 344
rect 2427 336 2973 344
rect 4027 336 4093 344
rect 4167 336 4433 344
rect 787 316 1033 324
rect 1627 316 1913 324
rect 2107 316 2433 324
rect 2976 324 2984 333
rect 2976 316 3393 324
rect 3987 316 4113 324
rect 527 296 793 304
rect 807 296 1113 304
rect 2207 296 2833 304
rect 2847 296 3053 304
rect 3107 296 3393 304
rect 2527 256 2693 264
rect 2707 256 4773 264
rect 4967 236 5013 244
rect 727 196 1733 204
rect 1747 196 2513 204
rect 247 176 333 184
rect 347 176 753 184
rect 147 156 373 164
rect 467 156 513 164
rect 547 156 693 164
rect 1187 156 1373 164
rect 1396 156 1413 164
rect 227 136 533 144
rect 767 136 993 144
rect 1396 144 1404 156
rect 1427 156 1873 164
rect 2027 156 2153 164
rect 2187 156 2273 164
rect 3987 156 4113 164
rect 4247 156 4453 164
rect 1247 136 1404 144
rect 1767 136 1993 144
rect 2567 136 2793 144
rect 3127 136 3373 144
rect 3707 136 3953 144
rect 4047 136 4493 144
rect 4507 136 4804 144
rect 1747 116 1893 124
rect 1907 116 2033 124
rect 2047 116 2493 124
rect 2547 116 2833 124
rect 2847 116 3093 124
rect 3107 116 3413 124
rect 3687 116 3993 124
rect 4527 116 4753 124
rect 4796 124 4804 136
rect 4827 136 5013 144
rect 4796 116 5033 124
rect 1487 96 1773 104
rect 1787 96 2573 104
rect 2587 96 3073 104
rect 3087 96 3573 104
rect 3047 76 3133 84
rect 3147 76 3173 84
rect 3187 76 3713 84
rect 3527 36 3593 44
rect 4967 16 4993 24
use INVX1  _273_
timestamp 0
transform -1 0 4490 0 -1 3130
box -6 -8 66 248
use NAND2X1  _274_
timestamp 0
transform -1 0 4770 0 -1 3130
box -6 -8 86 248
use OAI21X1  _275_
timestamp 0
transform -1 0 5070 0 -1 3130
box -6 -8 106 248
use INVX1  _276_
timestamp 0
transform -1 0 3830 0 -1 2170
box -6 -8 66 248
use NAND2X1  _277_
timestamp 0
transform 1 0 4990 0 1 4570
box -6 -8 86 248
use OAI21X1  _278_
timestamp 0
transform 1 0 4970 0 1 2170
box -6 -8 106 248
use INVX1  _279_
timestamp 0
transform 1 0 4610 0 -1 2650
box -6 -8 66 248
use NAND2X1  _280_
timestamp 0
transform -1 0 4870 0 -1 2170
box -6 -8 86 248
use OAI21X1  _281_
timestamp 0
transform -1 0 4970 0 -1 2650
box -6 -8 106 248
use INVX1  _282_
timestamp 0
transform 1 0 4070 0 1 2650
box -6 -8 66 248
use NAND2X1  _283_
timestamp 0
transform -1 0 3650 0 1 3130
box -6 -8 86 248
use OAI21X1  _284_
timestamp 0
transform 1 0 4070 0 1 3130
box -6 -8 106 248
use INVX1  _285_
timestamp 0
transform 1 0 3470 0 -1 3610
box -6 -8 66 248
use NAND2X1  _286_
timestamp 0
transform -1 0 4770 0 1 2170
box -6 -8 86 248
use OAI21X1  _287_
timestamp 0
transform 1 0 4670 0 -1 3610
box -6 -8 106 248
use INVX1  _288_
timestamp 0
transform 1 0 3590 0 1 3610
box -6 -8 66 248
use NAND2X1  _289_
timestamp 0
transform -1 0 4450 0 1 3130
box -6 -8 86 248
use OAI21X1  _290_
timestamp 0
transform 1 0 4130 0 1 3610
box -6 -8 106 248
use INVX1  _291_
timestamp 0
transform 1 0 1530 0 -1 5050
box -6 -8 66 248
use NAND2X1  _292_
timestamp 0
transform -1 0 4170 0 1 4090
box -6 -8 86 248
use OAI21X1  _293_
timestamp 0
transform -1 0 4470 0 1 4090
box -6 -8 106 248
use INVX1  _294_
timestamp 0
transform 1 0 3970 0 -1 5050
box -6 -8 66 248
use NAND2X1  _295_
timestamp 0
transform -1 0 4470 0 -1 3610
box -6 -8 86 248
use OAI21X1  _296_
timestamp 0
transform 1 0 4710 0 -1 4570
box -6 -8 106 248
use INVX1  _297_
timestamp 0
transform 1 0 4230 0 -1 5050
box -6 -8 66 248
use NAND2X1  _298_
timestamp 0
transform -1 0 4210 0 -1 4570
box -6 -8 86 248
use OAI21X1  _299_
timestamp 0
transform -1 0 4250 0 1 4570
box -6 -8 106 248
use INVX1  _300_
timestamp 0
transform 1 0 3330 0 1 4570
box -6 -8 66 248
use NAND2X1  _301_
timestamp 0
transform -1 0 3930 0 1 3610
box -6 -8 86 248
use OAI21X1  _302_
timestamp 0
transform -1 0 3970 0 1 4570
box -6 -8 106 248
use INVX1  _303_
timestamp 0
transform 1 0 3870 0 -1 4570
box -6 -8 66 248
use NAND2X1  _304_
timestamp 0
transform -1 0 4210 0 -1 3610
box -6 -8 86 248
use OAI21X1  _305_
timestamp 0
transform -1 0 4510 0 -1 4570
box -6 -8 106 248
use INVX1  _306_
timestamp 0
transform 1 0 3970 0 -1 4090
box -6 -8 66 248
use NAND2X1  _307_
timestamp 0
transform 1 0 4410 0 1 3610
box -6 -8 86 248
use OAI21X1  _308_
timestamp 0
transform 1 0 4230 0 -1 4090
box -6 -8 106 248
use INVX1  _309_
timestamp 0
transform -1 0 850 0 -1 2650
box -6 -8 66 248
use INVX1  _310_
timestamp 0
transform -1 0 250 0 -1 250
box -6 -8 66 248
use NOR2X1  _311_
timestamp 0
transform -1 0 290 0 -1 730
box -6 -8 86 248
use NAND3X1  _312_
timestamp 0
transform -1 0 550 0 1 250
box -6 -8 106 248
use NAND2X1  _313_
timestamp 0
transform 1 0 450 0 -1 3610
box -6 -8 86 248
use OAI21X1  _314_
timestamp 0
transform 1 0 430 0 1 3130
box -6 -8 106 248
use INVX1  _315_
timestamp 0
transform 1 0 1630 0 1 3610
box -6 -8 66 248
use INVX1  _316_
timestamp 0
transform -1 0 1030 0 -1 250
box -6 -8 66 248
use NOR2X1  _317_
timestamp 0
transform 1 0 690 0 -1 250
box -6 -8 86 248
use NAND2X1  _318_
timestamp 0
transform -1 0 930 0 -1 3130
box -6 -8 86 248
use OAI21X1  _319_
timestamp 0
transform -1 0 1070 0 -1 3610
box -6 -8 106 248
use INVX1  _320_
timestamp 0
transform -1 0 1570 0 -1 3610
box -6 -8 66 248
use NAND2X1  _321_
timestamp 0
transform 1 0 1670 0 -1 3130
box -6 -8 86 248
use OAI21X1  _322_
timestamp 0
transform 1 0 1510 0 1 3130
box -6 -8 106 248
use INVX1  _323_
timestamp 0
transform -1 0 670 0 -1 3130
box -6 -8 66 248
use INVX2  _324_
timestamp 0
transform 1 0 210 0 -1 1210
box -6 -8 66 248
use OR2X2  _325_
timestamp 0
transform 1 0 430 0 -1 2170
box -6 -8 106 248
use OAI21X1  _326_
timestamp 0
transform -1 0 550 0 1 2170
box -6 -8 106 248
use OAI21X1  _327_
timestamp 0
transform -1 0 310 0 -1 2650
box -6 -8 106 248
use OAI21X1  _328_
timestamp 0
transform 1 0 750 0 1 2170
box -6 -8 106 248
use OAI21X1  _329_
timestamp 0
transform 1 0 490 0 -1 2650
box -6 -8 106 248
use INVX1  _330_
timestamp 0
transform 1 0 2930 0 -1 2170
box -6 -8 66 248
use NAND2X1  _331_
timestamp 0
transform 1 0 3490 0 -1 2170
box -6 -8 86 248
use OAI21X1  _332_
timestamp 0
transform 1 0 3190 0 -1 2170
box -6 -8 106 248
use INVX1  _333_
timestamp 0
transform 1 0 2390 0 -1 2170
box -6 -8 66 248
use NAND2X1  _334_
timestamp 0
transform 1 0 2150 0 1 1690
box -6 -8 86 248
use OAI21X1  _335_
timestamp 0
transform -1 0 2210 0 -1 2170
box -6 -8 106 248
use INVX4  _336_
timestamp 0
transform -1 0 290 0 1 4570
box -6 -8 86 248
use NAND2X1  _337_
timestamp 0
transform 1 0 190 0 -1 5050
box -6 -8 86 248
use OAI21X1  _338_
timestamp 0
transform -1 0 570 0 -1 5050
box -6 -8 106 248
use INVX1  _339_
timestamp 0
transform 1 0 3650 0 -1 1690
box -6 -8 66 248
use INVX8  _340_
timestamp 0
transform -1 0 4250 0 -1 3130
box -6 -8 126 248
use NAND2X1  _341_
timestamp 0
transform -1 0 4710 0 1 1690
box -6 -8 86 248
use OAI21X1  _342_
timestamp 0
transform 1 0 4330 0 1 1690
box -6 -8 106 248
use NAND3X1  _343_
timestamp 0
transform 1 0 3670 0 1 1210
box -6 -8 106 248
use INVX1  _344_
timestamp 0
transform 1 0 3670 0 1 730
box -6 -8 66 248
use OAI21X1  _345_
timestamp 0
transform 1 0 4130 0 -1 1210
box -6 -8 106 248
use NAND2X1  _346_
timestamp 0
transform 1 0 4210 0 1 1210
box -6 -8 86 248
use NAND2X1  _347_
timestamp 0
transform -1 0 5050 0 -1 1210
box -6 -8 86 248
use OAI21X1  _348_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 106 248
use INVX1  _349_
timestamp 0
transform 1 0 2690 0 1 1690
box -6 -8 66 248
use OAI21X1  _350_
timestamp 0
transform -1 0 3190 0 1 1210
box -6 -8 106 248
use OR2X2  _351_
timestamp 0
transform 1 0 3070 0 -1 1690
box -6 -8 106 248
use NOR2X1  _352_
timestamp 0
transform -1 0 2890 0 1 1210
box -6 -8 86 248
use OAI21X1  _353_
timestamp 0
transform 1 0 2470 0 -1 1690
box -6 -8 106 248
use NAND2X1  _354_
timestamp 0
transform -1 0 3450 0 -1 1690
box -6 -8 86 248
use NAND2X1  _355_
timestamp 0
transform -1 0 4270 0 -1 1690
box -6 -8 86 248
use OAI21X1  _356_
timestamp 0
transform 1 0 3910 0 -1 1690
box -6 -8 106 248
use OAI21X1  _357_
timestamp 0
transform -1 0 2870 0 -1 1690
box -6 -8 106 248
use NAND2X1  _358_
timestamp 0
transform -1 0 3030 0 1 1690
box -6 -8 86 248
use OR2X2  _359_
timestamp 0
transform 1 0 3210 0 1 1690
box -6 -8 106 248
use NAND2X1  _360_
timestamp 0
transform -1 0 3590 0 1 1690
box -6 -8 86 248
use NAND2X1  _361_
timestamp 0
transform -1 0 3370 0 1 3130
box -6 -8 86 248
use OAI21X1  _362_
timestamp 0
transform -1 0 3330 0 1 2650
box -6 -8 106 248
use NOR2X1  _363_
timestamp 0
transform 1 0 2410 0 1 1690
box -6 -8 86 248
use NAND2X1  _364_
timestamp 0
transform 1 0 2290 0 1 1210
box -6 -8 86 248
use NAND3X1  _365_
timestamp 0
transform 1 0 3270 0 -1 1210
box -6 -8 106 248
use INVX1  _366_
timestamp 0
transform 1 0 2950 0 -1 730
box -6 -8 66 248
use AND2X2  _367_
timestamp 0
transform -1 0 2270 0 -1 1690
box -6 -8 106 248
use OAI21X1  _368_
timestamp 0
transform 1 0 2970 0 -1 1210
box -6 -8 106 248
use NAND2X1  _369_
timestamp 0
transform -1 0 3470 0 1 1210
box -6 -8 86 248
use NAND2X1  _370_
timestamp 0
transform 1 0 4990 0 -1 1690
box -6 -8 86 248
use OAI21X1  _371_
timestamp 0
transform 1 0 4710 0 -1 1690
box -6 -8 106 248
use INVX1  _372_
timestamp 0
transform 1 0 3390 0 1 250
box -6 -8 66 248
use OAI21X1  _373_
timestamp 0
transform 1 0 3390 0 1 730
box -6 -8 106 248
use OR2X2  _374_
timestamp 0
transform 1 0 4190 0 1 730
box -6 -8 106 248
use NAND2X1  _375_
timestamp 0
transform 1 0 3930 0 1 730
box -6 -8 86 248
use NAND2X1  _376_
timestamp 0
transform 1 0 4490 0 1 730
box -6 -8 86 248
use NAND2X1  _377_
timestamp 0
transform -1 0 4250 0 1 2170
box -6 -8 86 248
use OAI21X1  _378_
timestamp 0
transform -1 0 4370 0 -1 2170
box -6 -8 106 248
use NOR2X1  _379_
timestamp 0
transform -1 0 2470 0 1 250
box -6 -8 86 248
use NAND2X1  _380_
timestamp 0
transform 1 0 1730 0 1 1210
box -6 -8 86 248
use NAND3X1  _381_
timestamp 0
transform 1 0 1430 0 1 1210
box -6 -8 106 248
use INVX1  _382_
timestamp 0
transform -1 0 1130 0 -1 1690
box -6 -8 66 248
use NAND2X1  _383_
timestamp 0
transform 1 0 1570 0 1 1690
box -6 -8 86 248
use NAND2X1  _384_
timestamp 0
transform -1 0 1090 0 -1 2170
box -6 -8 86 248
use NAND2X1  _385_
timestamp 0
transform -1 0 1110 0 1 2170
box -6 -8 86 248
use NAND2X1  _386_
timestamp 0
transform 1 0 1130 0 -1 3130
box -6 -8 86 248
use OAI21X1  _387_
timestamp 0
transform -1 0 1030 0 1 2650
box -6 -8 106 248
use INVX1  _388_
timestamp 0
transform -1 0 4090 0 -1 2170
box -6 -8 66 248
use NAND3X1  _389_
timestamp 0
transform -1 0 1710 0 -1 1690
box -6 -8 106 248
use NAND3X1  _390_
timestamp 0
transform -1 0 1430 0 -1 1690
box -6 -8 106 248
use INVX1  _391_
timestamp 0
transform 1 0 1030 0 1 1690
box -6 -8 66 248
use NAND2X1  _392_
timestamp 0
transform -1 0 890 0 -1 1690
box -6 -8 86 248
use NAND3X1  _393_
timestamp 0
transform 1 0 1270 0 1 1690
box -6 -8 106 248
use NAND3X1  _394_
timestamp 0
transform 1 0 1850 0 1 1690
box -6 -8 106 248
use OAI21X1  _395_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 106 248
use INVX1  _396_
timestamp 0
transform 1 0 1290 0 -1 2170
box -6 -8 66 248
use NOR2X1  _397_
timestamp 0
transform 1 0 1530 0 -1 730
box -6 -8 86 248
use NAND2X1  _398_
timestamp 0
transform 1 0 2090 0 -1 730
box -6 -8 86 248
use OAI21X1  _399_
timestamp 0
transform 1 0 2090 0 -1 1210
box -6 -8 106 248
use OR2X2  _400_
timestamp 0
transform 1 0 1810 0 -1 2170
box -6 -8 106 248
use NAND2X1  _401_
timestamp 0
transform 1 0 1550 0 -1 2170
box -6 -8 86 248
use NAND2X1  _402_
timestamp 0
transform 1 0 1870 0 1 2170
box -6 -8 86 248
use NAND2X1  _403_
timestamp 0
transform -1 0 3010 0 -1 4090
box -6 -8 86 248
use OAI21X1  _404_
timestamp 0
transform 1 0 2630 0 -1 4090
box -6 -8 106 248
use INVX1  _405_
timestamp 0
transform -1 0 1470 0 -1 3130
box -6 -8 66 248
use INVX1  _406_
timestamp 0
transform 1 0 1310 0 1 2170
box -6 -8 66 248
use OAI21X1  _407_
timestamp 0
transform -1 0 1670 0 1 2170
box -6 -8 106 248
use OR2X2  _408_
timestamp 0
transform -1 0 1130 0 -1 2650
box -6 -8 106 248
use AOI21X1  _409_
timestamp 0
transform 1 0 1330 0 -1 2650
box -6 -8 106 248
use AOI22X1  _410_
timestamp 0
transform -1 0 1350 0 1 2650
box -6 -8 126 248
use INVX1  _411_
timestamp 0
transform -1 0 3370 0 -1 2650
box -6 -8 66 248
use AND2X2  _412_
timestamp 0
transform -1 0 1890 0 -1 730
box -6 -8 106 248
use NOR2X1  _413_
timestamp 0
transform 1 0 1670 0 1 730
box -6 -8 86 248
use NAND3X1  _414_
timestamp 0
transform 1 0 1950 0 1 730
box -6 -8 106 248
use NAND3X1  _415_
timestamp 0
transform 1 0 2810 0 1 730
box -6 -8 106 248
use INVX1  _416_
timestamp 0
transform -1 0 2190 0 1 250
box -6 -8 66 248
use NAND2X1  _417_
timestamp 0
transform 1 0 2530 0 1 730
box -6 -8 86 248
use NAND2X1  _418_
timestamp 0
transform 1 0 2370 0 -1 730
box -6 -8 86 248
use NAND3X1  _419_
timestamp 0
transform -1 0 3190 0 1 730
box -6 -8 106 248
use OAI21X1  _420_
timestamp 0
transform -1 0 3110 0 -1 2650
box -6 -8 106 248
use NAND2X1  _421_
timestamp 0
transform 1 0 4690 0 -1 1210
box -6 -8 86 248
use INVX1  _422_
timestamp 0
transform 1 0 4470 0 -1 250
box -6 -8 66 248
use NAND2X1  _423_
timestamp 0
transform 1 0 4990 0 -1 250
box -6 -8 86 248
use INVX1  _424_
timestamp 0
transform 1 0 5010 0 1 250
box -6 -8 66 248
use NAND2X1  _425_
timestamp 0
transform 1 0 4470 0 1 250
box -6 -8 86 248
use NAND2X1  _426_
timestamp 0
transform -1 0 4810 0 -1 250
box -6 -8 86 248
use INVX1  _427_
timestamp 0
transform -1 0 2710 0 1 250
box -6 -8 66 248
use NAND2X1  _428_
timestamp 0
transform 1 0 2250 0 1 730
box -6 -8 86 248
use NAND3X1  _429_
timestamp 0
transform 1 0 2650 0 -1 730
box -6 -8 106 248
use OAI21X1  _430_
timestamp 0
transform -1 0 1610 0 -1 1210
box -6 -8 106 248
use NAND3X1  _431_
timestamp 0
transform 1 0 1790 0 -1 1210
box -6 -8 106 248
use NAND2X1  _432_
timestamp 0
transform -1 0 2470 0 -1 1210
box -6 -8 86 248
use NAND3X1  _433_
timestamp 0
transform 1 0 2670 0 -1 1210
box -6 -8 106 248
use NAND2X1  _434_
timestamp 0
transform -1 0 4490 0 -1 1210
box -6 -8 86 248
use NAND2X1  _435_
timestamp 0
transform 1 0 3570 0 -1 3130
box -6 -8 86 248
use OAI21X1  _436_
timestamp 0
transform -1 0 3950 0 -1 3130
box -6 -8 106 248
use NAND3X1  _437_
timestamp 0
transform -1 0 2490 0 1 2170
box -6 -8 106 248
use OAI21X1  _438_
timestamp 0
transform -1 0 2730 0 -1 2170
box -6 -8 106 248
use NAND3X1  _439_
timestamp 0
transform 1 0 2690 0 1 2170
box -6 -8 106 248
use OAI21X1  _440_
timestamp 0
transform -1 0 3330 0 1 2170
box -6 -8 106 248
use INVX1  _441_
timestamp 0
transform 1 0 1630 0 -1 2650
box -6 -8 66 248
use OAI21X1  _442_
timestamp 0
transform -1 0 2270 0 -1 2650
box -6 -8 106 248
use OR2X2  _443_
timestamp 0
transform -1 0 1910 0 1 2650
box -6 -8 106 248
use NOR2X1  _444_
timestamp 0
transform -1 0 2330 0 -1 3130
box -6 -8 86 248
use OAI21X1  _445_
timestamp 0
transform -1 0 2050 0 -1 3130
box -6 -8 106 248
use NAND3X1  _446_
timestamp 0
transform 1 0 2090 0 1 2650
box -6 -8 106 248
use OAI21X1  _447_
timestamp 0
transform -1 0 4430 0 1 2650
box -6 -8 106 248
use OAI21X1  _448_
timestamp 0
transform -1 0 1990 0 -1 2650
box -6 -8 106 248
use NAND2X1  _449_
timestamp 0
transform 1 0 2370 0 1 2650
box -6 -8 86 248
use OR2X2  _450_
timestamp 0
transform 1 0 2470 0 -1 2650
box -6 -8 106 248
use NAND3X1  _451_
timestamp 0
transform 1 0 2650 0 1 2650
box -6 -8 106 248
use OAI21X1  _452_
timestamp 0
transform -1 0 3870 0 1 2650
box -6 -8 106 248
use NOR2X1  _453_
timestamp 0
transform 1 0 1530 0 1 2650
box -6 -8 86 248
use NAND2X1  _454_
timestamp 0
transform -1 0 1850 0 -1 3610
box -6 -8 86 248
use NAND2X1  _455_
timestamp 0
transform 1 0 2130 0 -1 4090
box -6 -8 86 248
use OR2X2  _456_
timestamp 0
transform -1 0 2150 0 -1 3610
box -6 -8 106 248
use AND2X2  _457_
timestamp 0
transform 1 0 1790 0 1 3130
box -6 -8 106 248
use OAI21X1  _458_
timestamp 0
transform 1 0 1890 0 1 3610
box -6 -8 106 248
use NAND3X1  _459_
timestamp 0
transform 1 0 2350 0 -1 3610
box -6 -8 106 248
use OAI21X1  _460_
timestamp 0
transform -1 0 2750 0 -1 3610
box -6 -8 106 248
use OAI21X1  _461_
timestamp 0
transform -1 0 2270 0 1 3610
box -6 -8 106 248
use OR2X2  _462_
timestamp 0
transform 1 0 2470 0 1 3610
box -6 -8 106 248
use AOI21X1  _463_
timestamp 0
transform 1 0 2770 0 1 3610
box -6 -8 106 248
use AOI22X1  _464_
timestamp 0
transform -1 0 3170 0 1 3610
box -6 -8 126 248
use NOR2X1  _465_
timestamp 0
transform 1 0 1350 0 1 3610
box -6 -8 86 248
use NAND2X1  _466_
timestamp 0
transform -1 0 1130 0 1 4090
box -6 -8 86 248
use NAND3X1  _467_
timestamp 0
transform 1 0 750 0 1 4090
box -6 -8 106 248
use INVX1  _468_
timestamp 0
transform -1 0 530 0 -1 4090
box -6 -8 66 248
use NAND2X1  _469_
timestamp 0
transform -1 0 550 0 1 4090
box -6 -8 86 248
use NAND2X1  _470_
timestamp 0
transform -1 0 850 0 -1 4570
box -6 -8 86 248
use NAND3X1  _471_
timestamp 0
transform 1 0 790 0 1 4570
box -6 -8 106 248
use OAI21X1  _472_
timestamp 0
transform -1 0 1090 0 -1 5050
box -6 -8 106 248
use NAND3X1  _473_
timestamp 0
transform 1 0 970 0 -1 4090
box -6 -8 106 248
use NAND3X1  _474_
timestamp 0
transform 1 0 1050 0 -1 4570
box -6 -8 106 248
use INVX1  _475_
timestamp 0
transform -1 0 270 0 -1 4570
box -6 -8 66 248
use NAND2X1  _476_
timestamp 0
transform -1 0 270 0 1 4090
box -6 -8 86 248
use NAND3X1  _477_
timestamp 0
transform 1 0 470 0 -1 4570
box -6 -8 106 248
use NAND3X1  _478_
timestamp 0
transform -1 0 590 0 1 4570
box -6 -8 106 248
use OAI21X1  _479_
timestamp 0
transform -1 0 3670 0 1 4570
box -6 -8 106 248
use INVX1  _480_
timestamp 0
transform -1 0 1430 0 1 4570
box -6 -8 66 248
use NOR2X1  _481_
timestamp 0
transform -1 0 290 0 -1 4090
box -6 -8 86 248
use NAND2X1  _482_
timestamp 0
transform -1 0 1410 0 1 4090
box -6 -8 86 248
use OAI21X1  _483_
timestamp 0
transform -1 0 1690 0 1 4090
box -6 -8 106 248
use OR2X2  _484_
timestamp 0
transform 1 0 1790 0 -1 5050
box -6 -8 106 248
use NAND2X1  _485_
timestamp 0
transform 1 0 2090 0 -1 5050
box -6 -8 86 248
use NAND2X1  _486_
timestamp 0
transform 1 0 2370 0 -1 5050
box -6 -8 86 248
use NAND2X1  _487_
timestamp 0
transform 1 0 2930 0 -1 5050
box -6 -8 86 248
use OAI21X1  _488_
timestamp 0
transform 1 0 2650 0 -1 5050
box -6 -8 106 248
use INVX1  _489_
timestamp 0
transform 1 0 1630 0 1 4570
box -6 -8 66 248
use OAI21X1  _490_
timestamp 0
transform -1 0 1990 0 1 4570
box -6 -8 106 248
use OR2X2  _491_
timestamp 0
transform 1 0 2170 0 1 4570
box -6 -8 106 248
use AOI21X1  _492_
timestamp 0
transform 1 0 2470 0 1 4570
box -6 -8 106 248
use AOI22X1  _493_
timestamp 0
transform -1 0 2890 0 1 4570
box -6 -8 126 248
use AND2X2  _494_
timestamp 0
transform 1 0 1250 0 -1 4090
box -6 -8 106 248
use NOR2X1  _495_
timestamp 0
transform 1 0 1550 0 -1 4090
box -6 -8 86 248
use NAND3X1  _496_
timestamp 0
transform 1 0 1830 0 -1 4090
box -6 -8 106 248
use NAND3X1  _497_
timestamp 0
transform 1 0 2210 0 -1 4570
box -6 -8 106 248
use INVX1  _498_
timestamp 0
transform -1 0 2450 0 -1 4090
box -6 -8 66 248
use NAND2X1  _499_
timestamp 0
transform -1 0 1970 0 1 4090
box -6 -8 86 248
use NAND2X1  _500_
timestamp 0
transform -1 0 2510 0 1 4090
box -6 -8 86 248
use NAND3X1  _501_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 106 248
use OAI21X1  _502_
timestamp 0
transform -1 0 3450 0 -1 4570
box -6 -8 106 248
use NAND2X1  _503_
timestamp 0
transform -1 0 3530 0 -1 4090
box -6 -8 86 248
use INVX1  _504_
timestamp 0
transform 1 0 4670 0 -1 730
box -6 -8 66 248
use NAND2X1  _505_
timestamp 0
transform -1 0 5010 0 -1 730
box -6 -8 86 248
use NAND2X1  _506_
timestamp 0
transform 1 0 4730 0 1 250
box -6 -8 86 248
use NAND2X1  _507_
timestamp 0
transform -1 0 4850 0 1 730
box -6 -8 86 248
use INVX1  _508_
timestamp 0
transform -1 0 3070 0 1 4090
box -6 -8 66 248
use NAND2X1  _509_
timestamp 0
transform 1 0 2150 0 1 4090
box -6 -8 86 248
use NAND3X1  _510_
timestamp 0
transform -1 0 2810 0 1 4090
box -6 -8 106 248
use OAI21X1  _511_
timestamp 0
transform 1 0 1630 0 -1 4570
box -6 -8 106 248
use NAND3X1  _512_
timestamp 0
transform 1 0 2510 0 -1 4570
box -6 -8 106 248
use NAND2X1  _513_
timestamp 0
transform -1 0 3330 0 1 4090
box -6 -8 86 248
use NAND3X1  _514_
timestamp 0
transform 1 0 3530 0 1 4090
box -6 -8 106 248
use NAND2X1  _515_
timestamp 0
transform -1 0 3910 0 1 4090
box -6 -8 86 248
use NOR2X1  _516_
timestamp 0
transform 1 0 750 0 1 250
box -6 -8 86 248
use AND2X2  _517_
timestamp 0
transform 1 0 1010 0 1 250
box -6 -8 106 248
use NAND2X1  _518_
timestamp 0
transform 1 0 1590 0 1 250
box -6 -8 86 248
use NOR2X1  _519_
timestamp 0
transform 1 0 1870 0 1 250
box -6 -8 86 248
use NAND2X1  _520_
timestamp 0
transform -1 0 1790 0 -1 250
box -6 -8 86 248
use OAI21X1  _521_
timestamp 0
transform -1 0 2070 0 -1 250
box -6 -8 106 248
use NAND2X1  _522_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 86 248
use OAI21X1  _523_
timestamp 0
transform -1 0 4030 0 -1 250
box -6 -8 106 248
use INVX1  _524_
timestamp 0
transform -1 0 1310 0 -1 1210
box -6 -8 66 248
use NAND2X1  _525_
timestamp 0
transform 1 0 1310 0 1 250
box -6 -8 86 248
use NAND2X1  _526_
timestamp 0
transform -1 0 1070 0 -1 1210
box -6 -8 86 248
use OAI21X1  _527_
timestamp 0
transform -1 0 1230 0 1 1210
box -6 -8 106 248
use INVX1  _528_
timestamp 0
transform 1 0 3190 0 -1 730
box -6 -8 66 248
use NAND2X1  _529_
timestamp 0
transform 1 0 1390 0 1 730
box -6 -8 86 248
use OAI21X1  _530_
timestamp 0
transform 1 0 1090 0 1 730
box -6 -8 106 248
use NAND2X1  _531_
timestamp 0
transform -1 0 690 0 1 1210
box -6 -8 86 248
use OAI21X1  _532_
timestamp 0
transform 1 0 450 0 -1 1210
box -6 -8 106 248
use NAND2X1  _533_
timestamp 0
transform -1 0 570 0 -1 730
box -6 -8 86 248
use OAI21X1  _534_
timestamp 0
transform 1 0 770 0 -1 730
box -6 -8 106 248
use NAND2X1  _535_
timestamp 0
transform -1 0 2590 0 -1 250
box -6 -8 86 248
use OAI21X1  _536_
timestamp 0
transform -1 0 2870 0 -1 250
box -6 -8 106 248
use NAND2X1  _537_
timestamp 0
transform -1 0 3150 0 -1 250
box -6 -8 86 248
use OAI21X1  _538_
timestamp 0
transform -1 0 3450 0 -1 250
box -6 -8 106 248
use OAI21X1  _539_
timestamp 0
transform -1 0 290 0 1 1690
box -6 -8 106 248
use OAI21X1  _540_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _541_
timestamp 0
transform 1 0 490 0 1 1690
box -6 -8 106 248
use OAI21X1  _542_
timestamp 0
transform -1 0 610 0 -1 1690
box -6 -8 106 248
use NAND2X1  _543_
timestamp 0
transform -1 0 3630 0 -1 1210
box -6 -8 86 248
use OAI21X1  _544_
timestamp 0
transform -1 0 3930 0 -1 1210
box -6 -8 106 248
use NAND2X1  _545_
timestamp 0
transform -1 0 4070 0 -1 730
box -6 -8 86 248
use OAI21X1  _546_
timestamp 0
transform 1 0 3690 0 -1 730
box -6 -8 106 248
use NAND2X1  _547_
timestamp 0
transform 1 0 2750 0 -1 3130
box -6 -8 86 248
use OAI21X1  _548_
timestamp 0
transform -1 0 2430 0 1 3130
box -6 -8 106 248
use NAND2X1  _549_
timestamp 0
transform -1 0 3730 0 1 250
box -6 -8 86 248
use OAI21X1  _550_
timestamp 0
transform -1 0 4030 0 1 250
box -6 -8 106 248
use NAND2X1  _551_
timestamp 0
transform 1 0 1070 0 1 3610
box -6 -8 86 248
use OAI21X1  _552_
timestamp 0
transform 1 0 790 0 1 3610
box -6 -8 106 248
use NAND2X1  _553_
timestamp 0
transform -1 0 1090 0 1 3130
box -6 -8 86 248
use OAI21X1  _554_
timestamp 0
transform 1 0 710 0 1 3130
box -6 -8 106 248
use NAND2X1  _555_
timestamp 0
transform 1 0 510 0 1 3610
box -6 -8 86 248
use OAI21X1  _556_
timestamp 0
transform -1 0 310 0 1 3610
box -6 -8 106 248
use DFFPOSX1  _557_
timestamp 0
transform 1 0 570 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _558_
timestamp 0
transform 1 0 4370 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _559_
timestamp 0
transform 1 0 4810 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _560_
timestamp 0
transform 1 0 4270 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _561_
timestamp 0
transform 1 0 3330 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _562_
timestamp 0
transform 1 0 4710 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _563_
timestamp 0
transform -1 0 4490 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _564_
timestamp 0
transform 1 0 490 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _565_
timestamp 0
transform 1 0 3890 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _566_
timestamp 0
transform 1 0 3010 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _567_
timestamp 0
transform 1 0 2330 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _568_
timestamp 0
transform 1 0 2570 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _569_
timestamp 0
transform 1 0 4290 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _570_
timestamp 0
transform 1 0 3650 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _571_
timestamp 0
transform 1 0 3330 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _572_
timestamp 0
transform 1 0 4170 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _573_
timestamp 0
transform 1 0 3650 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _574_
timestamp 0
transform 1 0 3030 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _575_
timestamp 0
transform 1 0 3170 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _576_
timestamp 0
transform 1 0 1090 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _577_
timestamp 0
transform 1 0 3530 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _578_
timestamp 0
transform 1 0 3010 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _579_
timestamp 0
transform 1 0 2890 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _580_
timestamp 0
transform 1 0 3450 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _581_
timestamp 0
transform -1 0 3770 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _582_
timestamp 0
transform 1 0 2070 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _583_
timestamp 0
transform 1 0 4030 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _584_
timestamp 0
transform 1 0 690 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _585_
timestamp 0
transform 1 0 870 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _586_
timestamp 0
transform 1 0 550 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _587_
timestamp 0
transform 1 0 650 0 1 730
box -6 -8 246 248
use DFFPOSX1  _588_
timestamp 0
transform 1 0 2710 0 1 250
box -6 -8 246 248
use DFFPOSX1  _589_
timestamp 0
transform -1 0 3190 0 1 250
box -6 -8 246 248
use DFFPOSX1  _590_
timestamp 0
transform 1 0 10 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _591_
timestamp 0
transform 1 0 590 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _592_
timestamp 0
transform -1 0 4010 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _593_
timestamp 0
transform -1 0 3490 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _594_
timestamp 0
transform 1 0 1890 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _595_
timestamp 0
transform 1 0 4030 0 1 250
box -6 -8 246 248
use DFFPOSX1  _596_
timestamp 0
transform 1 0 530 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _597_
timestamp 0
transform 1 0 530 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _598_
timestamp 0
transform 1 0 10 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _599_
timestamp 0
transform 1 0 10 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _600_
timestamp 0
transform 1 0 1070 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _601_
timestamp 0
transform 1 0 1090 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _602_
timestamp 0
transform 1 0 10 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _603_
timestamp 0
transform 1 0 250 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _604_
timestamp 0
transform -1 0 3030 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _605_
timestamp 0
transform 1 0 1950 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _606_
timestamp 0
transform 1 0 10 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _607_
timestamp 0
transform -1 0 250 0 1 730
box -6 -8 246 248
use DFFPOSX1  _608_
timestamp 0
transform 1 0 10 0 1 250
box -6 -8 246 248
use DFFPOSX1  _609_
timestamp 0
transform 1 0 250 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _610_
timestamp 0
transform 1 0 1030 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _611_
timestamp 0
transform -1 0 1510 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _612_
timestamp 0
transform -1 0 1350 0 -1 730
box -6 -8 246 248
use BUFX2  _613_
timestamp 0
transform 1 0 4930 0 1 3130
box -6 -8 86 248
use BUFX2  _614_
timestamp 0
transform -1 0 4950 0 1 2650
box -6 -8 86 248
use BUFX2  _615_
timestamp 0
transform 1 0 4450 0 1 4570
box -6 -8 86 248
use BUFX2  _616_
timestamp 0
transform -1 0 4570 0 -1 5050
box -6 -8 86 248
use BUFX2  _617_
timestamp 0
transform 1 0 4650 0 1 3130
box -6 -8 86 248
use BUFX2  _618_
timestamp 0
transform 1 0 4950 0 -1 3610
box -6 -8 86 248
use BUFX2  _619_
timestamp 0
transform 1 0 4950 0 1 3610
box -6 -8 86 248
use BUFX2  _620_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 86 248
use BUFX2  _621_
timestamp 0
transform 1 0 4950 0 1 4090
box -6 -8 86 248
use BUFX2  _622_
timestamp 0
transform 1 0 4990 0 -1 4570
box -6 -8 86 248
use BUFX2  _623_
timestamp 0
transform 1 0 4730 0 1 4570
box -6 -8 86 248
use BUFX2  _624_
timestamp 0
transform 1 0 4770 0 -1 5050
box -6 -8 86 248
use BUFX2  _625_
timestamp 0
transform 1 0 3450 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 4610 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 4610 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 4670 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform 1 0 4670 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform -1 0 1430 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 1930 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 1910 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 2550 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert15
timestamp 0
transform -1 0 810 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 2950 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 2010 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform 1 0 3090 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 1170 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 3030 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 4090 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 3370 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 3650 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform -1 0 3090 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 2950 0 -1 3610
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert0
timestamp 0
transform -1 0 3930 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert1
timestamp 0
transform -1 0 410 0 1 1210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert2
timestamp 0
transform 1 0 210 0 -1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert3
timestamp 0
transform 1 0 2610 0 1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert4
timestamp 0
transform 1 0 4270 0 -1 730
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert5
timestamp 0
transform -1 0 650 0 1 730
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert6
timestamp 0
transform 1 0 3770 0 1 2170
box -6 -8 206 248
use FILL  FILL72750x10950
timestamp 0
transform 1 0 4850 0 1 730
box -6 -8 26 248
use FILL  FILL72750x72150
timestamp 0
transform -1 0 4870 0 -1 5050
box -6 -8 26 248
use FILL  FILL73050x10950
timestamp 0
transform 1 0 4870 0 1 730
box -6 -8 26 248
use FILL  FILL73050x28950
timestamp 0
transform -1 0 4890 0 -1 2170
box -6 -8 26 248
use FILL  FILL73050x72150
timestamp 0
transform -1 0 4890 0 -1 5050
box -6 -8 26 248
use FILL  FILL73350x10950
timestamp 0
transform 1 0 4890 0 1 730
box -6 -8 26 248
use FILL  FILL73350x28950
timestamp 0
transform -1 0 4910 0 -1 2170
box -6 -8 26 248
use FILL  FILL73350x57750
timestamp 0
transform -1 0 4910 0 -1 4090
box -6 -8 26 248
use FILL  FILL73350x72150
timestamp 0
transform -1 0 4910 0 -1 5050
box -6 -8 26 248
use FILL  FILL73650x10950
timestamp 0
transform 1 0 4910 0 1 730
box -6 -8 26 248
use FILL  FILL73650x28950
timestamp 0
transform -1 0 4930 0 -1 2170
box -6 -8 26 248
use FILL  FILL73650x57750
timestamp 0
transform -1 0 4930 0 -1 4090
box -6 -8 26 248
use FILL  FILL73650x72150
timestamp 0
transform -1 0 4930 0 -1 5050
box -6 -8 26 248
use FILL  FILL73950x10950
timestamp 0
transform 1 0 4930 0 1 730
box -6 -8 26 248
use FILL  FILL73950x28950
timestamp 0
transform -1 0 4950 0 -1 2170
box -6 -8 26 248
use FILL  FILL73950x57750
timestamp 0
transform -1 0 4950 0 -1 4090
box -6 -8 26 248
use FILL  FILL73950x72150
timestamp 0
transform -1 0 4950 0 -1 5050
box -6 -8 26 248
use FILL  FILL74250x10950
timestamp 0
transform 1 0 4950 0 1 730
box -6 -8 26 248
use FILL  FILL74250x25350
timestamp 0
transform 1 0 4950 0 1 1690
box -6 -8 26 248
use FILL  FILL74250x28950
timestamp 0
transform -1 0 4970 0 -1 2170
box -6 -8 26 248
use FILL  FILL74250x39750
timestamp 0
transform 1 0 4950 0 1 2650
box -6 -8 26 248
use FILL  FILL74250x57750
timestamp 0
transform -1 0 4970 0 -1 4090
box -6 -8 26 248
use FILL  FILL74250x72150
timestamp 0
transform -1 0 4970 0 -1 5050
box -6 -8 26 248
use FILL  FILL74550x10950
timestamp 0
transform 1 0 4970 0 1 730
box -6 -8 26 248
use FILL  FILL74550x25350
timestamp 0
transform 1 0 4970 0 1 1690
box -6 -8 26 248
use FILL  FILL74550x28950
timestamp 0
transform -1 0 4990 0 -1 2170
box -6 -8 26 248
use FILL  FILL74550x36150
timestamp 0
transform -1 0 4990 0 -1 2650
box -6 -8 26 248
use FILL  FILL74550x39750
timestamp 0
transform 1 0 4970 0 1 2650
box -6 -8 26 248
use FILL  FILL74550x57750
timestamp 0
transform -1 0 4990 0 -1 4090
box -6 -8 26 248
use FILL  FILL74550x72150
timestamp 0
transform -1 0 4990 0 -1 5050
box -6 -8 26 248
use FILL  FILL74850x10950
timestamp 0
transform 1 0 4990 0 1 730
box -6 -8 26 248
use FILL  FILL74850x25350
timestamp 0
transform 1 0 4990 0 1 1690
box -6 -8 26 248
use FILL  FILL74850x28950
timestamp 0
transform -1 0 5010 0 -1 2170
box -6 -8 26 248
use FILL  FILL74850x36150
timestamp 0
transform -1 0 5010 0 -1 2650
box -6 -8 26 248
use FILL  FILL74850x39750
timestamp 0
transform 1 0 4990 0 1 2650
box -6 -8 26 248
use FILL  FILL74850x57750
timestamp 0
transform -1 0 5010 0 -1 4090
box -6 -8 26 248
use FILL  FILL74850x72150
timestamp 0
transform -1 0 5010 0 -1 5050
box -6 -8 26 248
use FILL  FILL75150x7350
timestamp 0
transform -1 0 5030 0 -1 730
box -6 -8 26 248
use FILL  FILL75150x10950
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 26 248
use FILL  FILL75150x25350
timestamp 0
transform 1 0 5010 0 1 1690
box -6 -8 26 248
use FILL  FILL75150x28950
timestamp 0
transform -1 0 5030 0 -1 2170
box -6 -8 26 248
use FILL  FILL75150x36150
timestamp 0
transform -1 0 5030 0 -1 2650
box -6 -8 26 248
use FILL  FILL75150x39750
timestamp 0
transform 1 0 5010 0 1 2650
box -6 -8 26 248
use FILL  FILL75150x46950
timestamp 0
transform 1 0 5010 0 1 3130
box -6 -8 26 248
use FILL  FILL75150x57750
timestamp 0
transform -1 0 5030 0 -1 4090
box -6 -8 26 248
use FILL  FILL75150x72150
timestamp 0
transform -1 0 5030 0 -1 5050
box -6 -8 26 248
use FILL  FILL75450x7350
timestamp 0
transform -1 0 5050 0 -1 730
box -6 -8 26 248
use FILL  FILL75450x10950
timestamp 0
transform 1 0 5030 0 1 730
box -6 -8 26 248
use FILL  FILL75450x25350
timestamp 0
transform 1 0 5030 0 1 1690
box -6 -8 26 248
use FILL  FILL75450x28950
timestamp 0
transform -1 0 5050 0 -1 2170
box -6 -8 26 248
use FILL  FILL75450x36150
timestamp 0
transform -1 0 5050 0 -1 2650
box -6 -8 26 248
use FILL  FILL75450x39750
timestamp 0
transform 1 0 5030 0 1 2650
box -6 -8 26 248
use FILL  FILL75450x46950
timestamp 0
transform 1 0 5030 0 1 3130
box -6 -8 26 248
use FILL  FILL75450x50550
timestamp 0
transform -1 0 5050 0 -1 3610
box -6 -8 26 248
use FILL  FILL75450x54150
timestamp 0
transform 1 0 5030 0 1 3610
box -6 -8 26 248
use FILL  FILL75450x57750
timestamp 0
transform -1 0 5050 0 -1 4090
box -6 -8 26 248
use FILL  FILL75450x61350
timestamp 0
transform 1 0 5030 0 1 4090
box -6 -8 26 248
use FILL  FILL75450x72150
timestamp 0
transform -1 0 5050 0 -1 5050
box -6 -8 26 248
use FILL  FILL75750x7350
timestamp 0
transform -1 0 5070 0 -1 730
box -6 -8 26 248
use FILL  FILL75750x10950
timestamp 0
transform 1 0 5050 0 1 730
box -6 -8 26 248
use FILL  FILL75750x14550
timestamp 0
transform -1 0 5070 0 -1 1210
box -6 -8 26 248
use FILL  FILL75750x18150
timestamp 0
transform 1 0 5050 0 1 1210
box -6 -8 26 248
use FILL  FILL75750x25350
timestamp 0
transform 1 0 5050 0 1 1690
box -6 -8 26 248
use FILL  FILL75750x28950
timestamp 0
transform -1 0 5070 0 -1 2170
box -6 -8 26 248
use FILL  FILL75750x36150
timestamp 0
transform -1 0 5070 0 -1 2650
box -6 -8 26 248
use FILL  FILL75750x39750
timestamp 0
transform 1 0 5050 0 1 2650
box -6 -8 26 248
use FILL  FILL75750x46950
timestamp 0
transform 1 0 5050 0 1 3130
box -6 -8 26 248
use FILL  FILL75750x50550
timestamp 0
transform -1 0 5070 0 -1 3610
box -6 -8 26 248
use FILL  FILL75750x54150
timestamp 0
transform 1 0 5050 0 1 3610
box -6 -8 26 248
use FILL  FILL75750x57750
timestamp 0
transform -1 0 5070 0 -1 4090
box -6 -8 26 248
use FILL  FILL75750x61350
timestamp 0
transform 1 0 5050 0 1 4090
box -6 -8 26 248
use FILL  FILL75750x72150
timestamp 0
transform -1 0 5070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__273_
timestamp 0
transform -1 0 4270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__274_
timestamp 0
transform -1 0 4510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__275_
timestamp 0
transform -1 0 4790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__276_
timestamp 0
transform -1 0 3590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__277_
timestamp 0
transform 1 0 4810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__278_
timestamp 0
transform 1 0 4770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__279_
timestamp 0
transform 1 0 4410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__280_
timestamp 0
transform -1 0 4630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__281_
timestamp 0
transform -1 0 4690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__282_
timestamp 0
transform 1 0 3870 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__283_
timestamp 0
transform -1 0 3390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__284_
timestamp 0
transform 1 0 3890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__285_
timestamp 0
transform 1 0 3270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__286_
timestamp 0
transform -1 0 4510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__287_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__288_
timestamp 0
transform 1 0 3410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__289_
timestamp 0
transform -1 0 4190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__290_
timestamp 0
transform 1 0 3930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__291_
timestamp 0
transform 1 0 1330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__292_
timestamp 0
transform -1 0 3930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__293_
timestamp 0
transform -1 0 4190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__294_
timestamp 0
transform 1 0 3770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__295_
timestamp 0
transform -1 0 4230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__296_
timestamp 0
transform 1 0 4510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__297_
timestamp 0
transform 1 0 4030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__298_
timestamp 0
transform -1 0 3950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__299_
timestamp 0
transform -1 0 3990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__300_
timestamp 0
transform 1 0 3130 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__301_
timestamp 0
transform -1 0 3670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__302_
timestamp 0
transform -1 0 3690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__303_
timestamp 0
transform 1 0 3690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__304_
timestamp 0
transform -1 0 3950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__305_
timestamp 0
transform -1 0 4230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__306_
timestamp 0
transform 1 0 3770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__307_
timestamp 0
transform 1 0 4230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__308_
timestamp 0
transform 1 0 4030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__309_
timestamp 0
transform -1 0 610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__310_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__311_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__312_
timestamp 0
transform -1 0 270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__313_
timestamp 0
transform 1 0 250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__314_
timestamp 0
transform 1 0 250 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__315_
timestamp 0
transform 1 0 1430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__316_
timestamp 0
transform -1 0 790 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__317_
timestamp 0
transform 1 0 490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__318_
timestamp 0
transform -1 0 690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__319_
timestamp 0
transform -1 0 790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__320_
timestamp 0
transform -1 0 1330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__321_
timestamp 0
transform 1 0 1470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__322_
timestamp 0
transform 1 0 1330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__323_
timestamp 0
transform -1 0 430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__324_
timestamp 0
transform 1 0 10 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__325_
timestamp 0
transform 1 0 250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__326_
timestamp 0
transform -1 0 270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__327_
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__328_
timestamp 0
transform 1 0 550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__329_
timestamp 0
transform 1 0 310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__330_
timestamp 0
transform 1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__331_
timestamp 0
transform 1 0 3290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__332_
timestamp 0
transform 1 0 2990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__333_
timestamp 0
transform 1 0 2210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__334_
timestamp 0
transform 1 0 1950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__335_
timestamp 0
transform -1 0 1930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__336_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__337_
timestamp 0
transform 1 0 10 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__338_
timestamp 0
transform -1 0 290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__339_
timestamp 0
transform 1 0 3450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__340_
timestamp 0
transform -1 0 3970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__341_
timestamp 0
transform -1 0 4450 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__342_
timestamp 0
transform 1 0 4130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__343_
timestamp 0
transform 1 0 3470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__344_
timestamp 0
transform 1 0 3490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__345_
timestamp 0
transform 1 0 3930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__346_
timestamp 0
transform 1 0 4010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__347_
timestamp 0
transform -1 0 4790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__348_
timestamp 0
transform 1 0 4530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__349_
timestamp 0
transform 1 0 2490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__350_
timestamp 0
transform -1 0 2910 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__351_
timestamp 0
transform 1 0 2870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__352_
timestamp 0
transform -1 0 2650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__353_
timestamp 0
transform 1 0 2270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__354_
timestamp 0
transform -1 0 3190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__355_
timestamp 0
transform -1 0 4030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__356_
timestamp 0
transform 1 0 3710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__357_
timestamp 0
transform -1 0 2590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__358_
timestamp 0
transform -1 0 2770 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__359_
timestamp 0
transform 1 0 3030 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__360_
timestamp 0
transform -1 0 3330 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__361_
timestamp 0
transform -1 0 3110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__362_
timestamp 0
transform -1 0 3050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__363_
timestamp 0
transform 1 0 2230 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__364_
timestamp 0
transform 1 0 2090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__365_
timestamp 0
transform 1 0 3070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__366_
timestamp 0
transform 1 0 2750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__367_
timestamp 0
transform -1 0 2010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__368_
timestamp 0
transform 1 0 2770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__369_
timestamp 0
transform -1 0 3210 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__370_
timestamp 0
transform 1 0 4810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__371_
timestamp 0
transform 1 0 4510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__372_
timestamp 0
transform 1 0 3190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__373_
timestamp 0
transform 1 0 3190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__374_
timestamp 0
transform 1 0 4010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__375_
timestamp 0
transform 1 0 3730 0 1 730
box -6 -8 26 248
use FILL  FILL_0__376_
timestamp 0
transform 1 0 4290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__377_
timestamp 0
transform -1 0 3990 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__378_
timestamp 0
transform -1 0 4110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__379_
timestamp 0
transform -1 0 2210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__380_
timestamp 0
transform 1 0 1530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__381_
timestamp 0
transform 1 0 1230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__382_
timestamp 0
transform -1 0 910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__383_
timestamp 0
transform 1 0 1370 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__384_
timestamp 0
transform -1 0 830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__385_
timestamp 0
transform -1 0 870 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__386_
timestamp 0
transform 1 0 930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__387_
timestamp 0
transform -1 0 750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__388_
timestamp 0
transform -1 0 3850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__389_
timestamp 0
transform -1 0 1450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__390_
timestamp 0
transform -1 0 1150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__391_
timestamp 0
transform 1 0 830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__392_
timestamp 0
transform -1 0 630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__393_
timestamp 0
transform 1 0 1090 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__394_
timestamp 0
transform 1 0 1650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__395_
timestamp 0
transform -1 0 3610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__396_
timestamp 0
transform 1 0 1090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__397_
timestamp 0
transform 1 0 1350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__398_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__399_
timestamp 0
transform 1 0 1890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__400_
timestamp 0
transform 1 0 1630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__401_
timestamp 0
transform 1 0 1350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__402_
timestamp 0
transform 1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__403_
timestamp 0
transform -1 0 2750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__404_
timestamp 0
transform 1 0 2450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__405_
timestamp 0
transform -1 0 1230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__406_
timestamp 0
transform 1 0 1110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__407_
timestamp 0
transform -1 0 1390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__408_
timestamp 0
transform -1 0 870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__409_
timestamp 0
transform 1 0 1130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__410_
timestamp 0
transform -1 0 1050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__411_
timestamp 0
transform -1 0 3130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__412_
timestamp 0
transform -1 0 1630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__413_
timestamp 0
transform 1 0 1470 0 1 730
box -6 -8 26 248
use FILL  FILL_0__414_
timestamp 0
transform 1 0 1750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__415_
timestamp 0
transform 1 0 2610 0 1 730
box -6 -8 26 248
use FILL  FILL_0__416_
timestamp 0
transform -1 0 1970 0 1 250
box -6 -8 26 248
use FILL  FILL_0__417_
timestamp 0
transform 1 0 2330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__418_
timestamp 0
transform 1 0 2170 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__419_
timestamp 0
transform -1 0 2930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__420_
timestamp 0
transform -1 0 2830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__421_
timestamp 0
transform 1 0 4490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__422_
timestamp 0
transform 1 0 4270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__423_
timestamp 0
transform 1 0 4810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__424_
timestamp 0
transform 1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__425_
timestamp 0
transform 1 0 4270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__426_
timestamp 0
transform -1 0 4550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__427_
timestamp 0
transform -1 0 2490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__428_
timestamp 0
transform 1 0 2050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__429_
timestamp 0
transform 1 0 2450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__430_
timestamp 0
transform -1 0 1330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__431_
timestamp 0
transform 1 0 1610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__432_
timestamp 0
transform -1 0 2210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__433_
timestamp 0
transform 1 0 2470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__434_
timestamp 0
transform -1 0 4250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__435_
timestamp 0
transform 1 0 3370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__436_
timestamp 0
transform -1 0 3670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__437_
timestamp 0
transform -1 0 2210 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__438_
timestamp 0
transform -1 0 2470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__439_
timestamp 0
transform 1 0 2490 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__440_
timestamp 0
transform -1 0 3050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__441_
timestamp 0
transform 1 0 1430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__442_
timestamp 0
transform -1 0 2010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__443_
timestamp 0
transform -1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__444_
timestamp 0
transform -1 0 2070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__445_
timestamp 0
transform -1 0 1770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__446_
timestamp 0
transform 1 0 1910 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__447_
timestamp 0
transform -1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__448_
timestamp 0
transform -1 0 1710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__449_
timestamp 0
transform 1 0 2190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__450_
timestamp 0
transform 1 0 2270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__451_
timestamp 0
transform 1 0 2450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__452_
timestamp 0
transform -1 0 3590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__453_
timestamp 0
transform 1 0 1350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__454_
timestamp 0
transform -1 0 1590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__455_
timestamp 0
transform 1 0 1930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__456_
timestamp 0
transform -1 0 1870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__457_
timestamp 0
transform 1 0 1610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__458_
timestamp 0
transform 1 0 1690 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__459_
timestamp 0
transform 1 0 2150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__460_
timestamp 0
transform -1 0 2470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__461_
timestamp 0
transform -1 0 2010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__462_
timestamp 0
transform 1 0 2270 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__463_
timestamp 0
transform 1 0 2570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__464_
timestamp 0
transform -1 0 2890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__465_
timestamp 0
transform 1 0 1150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__466_
timestamp 0
transform -1 0 870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__467_
timestamp 0
transform 1 0 550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__468_
timestamp 0
transform -1 0 310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__469_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__470_
timestamp 0
transform -1 0 590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__471_
timestamp 0
transform 1 0 590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__472_
timestamp 0
transform -1 0 830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__473_
timestamp 0
transform 1 0 770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__474_
timestamp 0
transform 1 0 850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__475_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__476_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__477_
timestamp 0
transform 1 0 270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__478_
timestamp 0
transform -1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__479_
timestamp 0
transform -1 0 3410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__480_
timestamp 0
transform -1 0 1190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__481_
timestamp 0
transform -1 0 30 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__482_
timestamp 0
transform -1 0 1150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__483_
timestamp 0
transform -1 0 1430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__484_
timestamp 0
transform 1 0 1590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__485_
timestamp 0
transform 1 0 1890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__486_
timestamp 0
transform 1 0 2170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__487_
timestamp 0
transform 1 0 2750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__488_
timestamp 0
transform 1 0 2450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__489_
timestamp 0
transform 1 0 1430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__490_
timestamp 0
transform -1 0 1710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__491_
timestamp 0
transform 1 0 1990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__492_
timestamp 0
transform 1 0 2270 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__493_
timestamp 0
transform -1 0 2590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__494_
timestamp 0
transform 1 0 1070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__495_
timestamp 0
transform 1 0 1350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__496_
timestamp 0
transform 1 0 1630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__497_
timestamp 0
transform 1 0 2010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__498_
timestamp 0
transform -1 0 2230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__499_
timestamp 0
transform -1 0 1710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__500_
timestamp 0
transform -1 0 2250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__501_
timestamp 0
transform -1 0 2630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__502_
timestamp 0
transform -1 0 3190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__503_
timestamp 0
transform -1 0 3270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__504_
timestamp 0
transform 1 0 4470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__505_
timestamp 0
transform -1 0 4750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__506_
timestamp 0
transform 1 0 4550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__507_
timestamp 0
transform -1 0 4590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__508_
timestamp 0
transform -1 0 2830 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__509_
timestamp 0
transform 1 0 1970 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__510_
timestamp 0
transform -1 0 2530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__511_
timestamp 0
transform 1 0 1430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__512_
timestamp 0
transform 1 0 2310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__513_
timestamp 0
transform -1 0 3090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__514_
timestamp 0
transform 1 0 3330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__515_
timestamp 0
transform -1 0 3650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__516_
timestamp 0
transform 1 0 550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__517_
timestamp 0
transform 1 0 830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__518_
timestamp 0
transform 1 0 1390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__519_
timestamp 0
transform 1 0 1670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__520_
timestamp 0
transform -1 0 1530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__521_
timestamp 0
transform -1 0 1810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__522_
timestamp 0
transform -1 0 3470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__523_
timestamp 0
transform -1 0 3750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__524_
timestamp 0
transform -1 0 1090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__525_
timestamp 0
transform 1 0 1110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__526_
timestamp 0
transform -1 0 810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__527_
timestamp 0
transform -1 0 950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__528_
timestamp 0
transform 1 0 3010 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__529_
timestamp 0
transform 1 0 1190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__530_
timestamp 0
transform 1 0 890 0 1 730
box -6 -8 26 248
use FILL  FILL_0__531_
timestamp 0
transform -1 0 430 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__532_
timestamp 0
transform 1 0 270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__533_
timestamp 0
transform -1 0 310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__534_
timestamp 0
transform 1 0 570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__535_
timestamp 0
transform -1 0 2330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__536_
timestamp 0
transform -1 0 2610 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__537_
timestamp 0
transform -1 0 2890 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__538_
timestamp 0
transform -1 0 3170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__539_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__540_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__541_
timestamp 0
transform 1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__542_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__543_
timestamp 0
transform -1 0 3390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__544_
timestamp 0
transform -1 0 3650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__545_
timestamp 0
transform -1 0 3810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__546_
timestamp 0
transform 1 0 3490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__547_
timestamp 0
transform 1 0 2570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__548_
timestamp 0
transform -1 0 2150 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__549_
timestamp 0
transform -1 0 3470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__550_
timestamp 0
transform -1 0 3750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__551_
timestamp 0
transform 1 0 890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__552_
timestamp 0
transform 1 0 590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__553_
timestamp 0
transform -1 0 830 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__554_
timestamp 0
transform 1 0 530 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__555_
timestamp 0
transform 1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__556_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__613_
timestamp 0
transform 1 0 4730 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__614_
timestamp 0
transform -1 0 4710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__615_
timestamp 0
transform 1 0 4250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__616_
timestamp 0
transform -1 0 4310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__617_
timestamp 0
transform 1 0 4450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__618_
timestamp 0
transform 1 0 4770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__619_
timestamp 0
transform 1 0 4750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__620_
timestamp 0
transform 1 0 4610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__621_
timestamp 0
transform 1 0 4750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__622_
timestamp 0
transform 1 0 4810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__623_
timestamp 0
transform 1 0 4530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__624_
timestamp 0
transform 1 0 4570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__625_
timestamp 0
transform 1 0 3250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 4430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 4350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 4470 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform 1 0 4490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform -1 0 1170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 1730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 1710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 2370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 1810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform 1 0 2910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 2830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 3890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 3130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 3390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform -1 0 2830 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 2750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert0
timestamp 0
transform -1 0 3550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert1
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert2
timestamp 0
transform 1 0 10 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert3
timestamp 0
transform 1 0 2430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert4
timestamp 0
transform 1 0 4070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert5
timestamp 0
transform -1 0 270 0 1 730
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert6
timestamp 0
transform 1 0 3570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__273_
timestamp 0
transform -1 0 4290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__274_
timestamp 0
transform -1 0 4530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__275_
timestamp 0
transform -1 0 4810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__276_
timestamp 0
transform -1 0 3610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__277_
timestamp 0
transform 1 0 4830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__278_
timestamp 0
transform 1 0 4790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__279_
timestamp 0
transform 1 0 4430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__280_
timestamp 0
transform -1 0 4650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__281_
timestamp 0
transform -1 0 4710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__282_
timestamp 0
transform 1 0 3890 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__283_
timestamp 0
transform -1 0 3410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__284_
timestamp 0
transform 1 0 3910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__285_
timestamp 0
transform 1 0 3290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__286_
timestamp 0
transform -1 0 4530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__287_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__288_
timestamp 0
transform 1 0 3430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__289_
timestamp 0
transform -1 0 4210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__290_
timestamp 0
transform 1 0 3950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__291_
timestamp 0
transform 1 0 1350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__292_
timestamp 0
transform -1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__293_
timestamp 0
transform -1 0 4210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__294_
timestamp 0
transform 1 0 3790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__295_
timestamp 0
transform -1 0 4250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__296_
timestamp 0
transform 1 0 4530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__297_
timestamp 0
transform 1 0 4050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__298_
timestamp 0
transform -1 0 3970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__299_
timestamp 0
transform -1 0 4010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__300_
timestamp 0
transform 1 0 3150 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__301_
timestamp 0
transform -1 0 3690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__302_
timestamp 0
transform -1 0 3710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__303_
timestamp 0
transform 1 0 3710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__304_
timestamp 0
transform -1 0 3970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__305_
timestamp 0
transform -1 0 4250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__306_
timestamp 0
transform 1 0 3790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__307_
timestamp 0
transform 1 0 4250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__308_
timestamp 0
transform 1 0 4050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__309_
timestamp 0
transform -1 0 630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__310_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__311_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__312_
timestamp 0
transform -1 0 290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__313_
timestamp 0
transform 1 0 270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__314_
timestamp 0
transform 1 0 270 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__315_
timestamp 0
transform 1 0 1450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__316_
timestamp 0
transform -1 0 810 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__317_
timestamp 0
transform 1 0 510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__318_
timestamp 0
transform -1 0 710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__319_
timestamp 0
transform -1 0 810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__320_
timestamp 0
transform -1 0 1350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__321_
timestamp 0
transform 1 0 1490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__322_
timestamp 0
transform 1 0 1350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__323_
timestamp 0
transform -1 0 450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__324_
timestamp 0
transform 1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__325_
timestamp 0
transform 1 0 270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__326_
timestamp 0
transform -1 0 290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__327_
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__328_
timestamp 0
transform 1 0 570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__329_
timestamp 0
transform 1 0 330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__330_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__331_
timestamp 0
transform 1 0 3310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__332_
timestamp 0
transform 1 0 3010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__333_
timestamp 0
transform 1 0 2230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__334_
timestamp 0
transform 1 0 1970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__335_
timestamp 0
transform -1 0 1950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__336_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__337_
timestamp 0
transform 1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__338_
timestamp 0
transform -1 0 310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__339_
timestamp 0
transform 1 0 3470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__340_
timestamp 0
transform -1 0 3990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__341_
timestamp 0
transform -1 0 4470 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__342_
timestamp 0
transform 1 0 4150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__343_
timestamp 0
transform 1 0 3490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__344_
timestamp 0
transform 1 0 3510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__345_
timestamp 0
transform 1 0 3950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__346_
timestamp 0
transform 1 0 4030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__347_
timestamp 0
transform -1 0 4810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__348_
timestamp 0
transform 1 0 4550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__349_
timestamp 0
transform 1 0 2510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__350_
timestamp 0
transform -1 0 2930 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__351_
timestamp 0
transform 1 0 2890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__352_
timestamp 0
transform -1 0 2670 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__353_
timestamp 0
transform 1 0 2290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__354_
timestamp 0
transform -1 0 3210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__355_
timestamp 0
transform -1 0 4050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__356_
timestamp 0
transform 1 0 3730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__357_
timestamp 0
transform -1 0 2610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__358_
timestamp 0
transform -1 0 2790 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__359_
timestamp 0
transform 1 0 3050 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__360_
timestamp 0
transform -1 0 3350 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__361_
timestamp 0
transform -1 0 3130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__362_
timestamp 0
transform -1 0 3070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__363_
timestamp 0
transform 1 0 2250 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__364_
timestamp 0
transform 1 0 2110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__365_
timestamp 0
transform 1 0 3090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__366_
timestamp 0
transform 1 0 2770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__367_
timestamp 0
transform -1 0 2030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__368_
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__369_
timestamp 0
transform -1 0 3230 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__370_
timestamp 0
transform 1 0 4830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__371_
timestamp 0
transform 1 0 4530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__372_
timestamp 0
transform 1 0 3210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__373_
timestamp 0
transform 1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__374_
timestamp 0
transform 1 0 4030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__375_
timestamp 0
transform 1 0 3750 0 1 730
box -6 -8 26 248
use FILL  FILL_1__376_
timestamp 0
transform 1 0 4310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__377_
timestamp 0
transform -1 0 4010 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__378_
timestamp 0
transform -1 0 4130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__379_
timestamp 0
transform -1 0 2230 0 1 250
box -6 -8 26 248
use FILL  FILL_1__380_
timestamp 0
transform 1 0 1550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__381_
timestamp 0
transform 1 0 1250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__382_
timestamp 0
transform -1 0 930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__383_
timestamp 0
transform 1 0 1390 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__384_
timestamp 0
transform -1 0 850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__385_
timestamp 0
transform -1 0 890 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__386_
timestamp 0
transform 1 0 950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__387_
timestamp 0
transform -1 0 770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__388_
timestamp 0
transform -1 0 3870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__389_
timestamp 0
transform -1 0 1470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__390_
timestamp 0
transform -1 0 1170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__391_
timestamp 0
transform 1 0 850 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__392_
timestamp 0
transform -1 0 650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__393_
timestamp 0
transform 1 0 1110 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__394_
timestamp 0
transform 1 0 1670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__395_
timestamp 0
transform -1 0 3630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__396_
timestamp 0
transform 1 0 1110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__397_
timestamp 0
transform 1 0 1370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__398_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__399_
timestamp 0
transform 1 0 1910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__400_
timestamp 0
transform 1 0 1650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__401_
timestamp 0
transform 1 0 1370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__402_
timestamp 0
transform 1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__403_
timestamp 0
transform -1 0 2770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__404_
timestamp 0
transform 1 0 2470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__405_
timestamp 0
transform -1 0 1250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__406_
timestamp 0
transform 1 0 1130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__407_
timestamp 0
transform -1 0 1410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__408_
timestamp 0
transform -1 0 890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__409_
timestamp 0
transform 1 0 1150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__410_
timestamp 0
transform -1 0 1070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__411_
timestamp 0
transform -1 0 3150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__412_
timestamp 0
transform -1 0 1650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__413_
timestamp 0
transform 1 0 1490 0 1 730
box -6 -8 26 248
use FILL  FILL_1__414_
timestamp 0
transform 1 0 1770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__415_
timestamp 0
transform 1 0 2630 0 1 730
box -6 -8 26 248
use FILL  FILL_1__416_
timestamp 0
transform -1 0 1990 0 1 250
box -6 -8 26 248
use FILL  FILL_1__417_
timestamp 0
transform 1 0 2350 0 1 730
box -6 -8 26 248
use FILL  FILL_1__418_
timestamp 0
transform 1 0 2190 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__419_
timestamp 0
transform -1 0 2950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__420_
timestamp 0
transform -1 0 2850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__421_
timestamp 0
transform 1 0 4510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__422_
timestamp 0
transform 1 0 4290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__423_
timestamp 0
transform 1 0 4830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__424_
timestamp 0
transform 1 0 4830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__425_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__426_
timestamp 0
transform -1 0 4570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__427_
timestamp 0
transform -1 0 2510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__428_
timestamp 0
transform 1 0 2070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__429_
timestamp 0
transform 1 0 2470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__430_
timestamp 0
transform -1 0 1350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__431_
timestamp 0
transform 1 0 1630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__432_
timestamp 0
transform -1 0 2230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__433_
timestamp 0
transform 1 0 2490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__434_
timestamp 0
transform -1 0 4270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__435_
timestamp 0
transform 1 0 3390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__436_
timestamp 0
transform -1 0 3690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__437_
timestamp 0
transform -1 0 2230 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__438_
timestamp 0
transform -1 0 2490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__439_
timestamp 0
transform 1 0 2510 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__440_
timestamp 0
transform -1 0 3070 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__441_
timestamp 0
transform 1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__442_
timestamp 0
transform -1 0 2030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__443_
timestamp 0
transform -1 0 1650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__444_
timestamp 0
transform -1 0 2090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__445_
timestamp 0
transform -1 0 1790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__446_
timestamp 0
transform 1 0 1930 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__447_
timestamp 0
transform -1 0 4170 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__448_
timestamp 0
transform -1 0 1730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__449_
timestamp 0
transform 1 0 2210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__450_
timestamp 0
transform 1 0 2290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__451_
timestamp 0
transform 1 0 2470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__452_
timestamp 0
transform -1 0 3610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__453_
timestamp 0
transform 1 0 1370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__454_
timestamp 0
transform -1 0 1610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__455_
timestamp 0
transform 1 0 1950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__456_
timestamp 0
transform -1 0 1890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__457_
timestamp 0
transform 1 0 1630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__458_
timestamp 0
transform 1 0 1710 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__459_
timestamp 0
transform 1 0 2170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__460_
timestamp 0
transform -1 0 2490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__461_
timestamp 0
transform -1 0 2030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__462_
timestamp 0
transform 1 0 2290 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__463_
timestamp 0
transform 1 0 2590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__464_
timestamp 0
transform -1 0 2910 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__465_
timestamp 0
transform 1 0 1170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__466_
timestamp 0
transform -1 0 890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__467_
timestamp 0
transform 1 0 570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__468_
timestamp 0
transform -1 0 330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__469_
timestamp 0
transform -1 0 310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__470_
timestamp 0
transform -1 0 610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__471_
timestamp 0
transform 1 0 610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__472_
timestamp 0
transform -1 0 850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__473_
timestamp 0
transform 1 0 790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__474_
timestamp 0
transform 1 0 870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__475_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__476_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__477_
timestamp 0
transform 1 0 290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__478_
timestamp 0
transform -1 0 330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__479_
timestamp 0
transform -1 0 3430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__480_
timestamp 0
transform -1 0 1210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__481_
timestamp 0
transform -1 0 50 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__482_
timestamp 0
transform -1 0 1170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__483_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__484_
timestamp 0
transform 1 0 1610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__485_
timestamp 0
transform 1 0 1910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__486_
timestamp 0
transform 1 0 2190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__487_
timestamp 0
transform 1 0 2770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__488_
timestamp 0
transform 1 0 2470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__489_
timestamp 0
transform 1 0 1450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__490_
timestamp 0
transform -1 0 1730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__491_
timestamp 0
transform 1 0 2010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__492_
timestamp 0
transform 1 0 2290 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__493_
timestamp 0
transform -1 0 2610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__494_
timestamp 0
transform 1 0 1090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__495_
timestamp 0
transform 1 0 1370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__496_
timestamp 0
transform 1 0 1650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__497_
timestamp 0
transform 1 0 2030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__498_
timestamp 0
transform -1 0 2250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__499_
timestamp 0
transform -1 0 1730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__500_
timestamp 0
transform -1 0 2270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__501_
timestamp 0
transform -1 0 2650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__502_
timestamp 0
transform -1 0 3210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__503_
timestamp 0
transform -1 0 3290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__504_
timestamp 0
transform 1 0 4490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__505_
timestamp 0
transform -1 0 4770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__506_
timestamp 0
transform 1 0 4570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__507_
timestamp 0
transform -1 0 4610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__508_
timestamp 0
transform -1 0 2850 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__509_
timestamp 0
transform 1 0 1990 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__510_
timestamp 0
transform -1 0 2550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__511_
timestamp 0
transform 1 0 1450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__512_
timestamp 0
transform 1 0 2330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__513_
timestamp 0
transform -1 0 3110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__514_
timestamp 0
transform 1 0 3350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__515_
timestamp 0
transform -1 0 3670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__516_
timestamp 0
transform 1 0 570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__517_
timestamp 0
transform 1 0 850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__518_
timestamp 0
transform 1 0 1410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__519_
timestamp 0
transform 1 0 1690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__520_
timestamp 0
transform -1 0 1550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__521_
timestamp 0
transform -1 0 1830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__522_
timestamp 0
transform -1 0 3490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__523_
timestamp 0
transform -1 0 3770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__524_
timestamp 0
transform -1 0 1110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__525_
timestamp 0
transform 1 0 1130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__526_
timestamp 0
transform -1 0 830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__527_
timestamp 0
transform -1 0 970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__528_
timestamp 0
transform 1 0 3030 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__529_
timestamp 0
transform 1 0 1210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__530_
timestamp 0
transform 1 0 910 0 1 730
box -6 -8 26 248
use FILL  FILL_1__531_
timestamp 0
transform -1 0 450 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__532_
timestamp 0
transform 1 0 290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__533_
timestamp 0
transform -1 0 330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__534_
timestamp 0
transform 1 0 590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__535_
timestamp 0
transform -1 0 2350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__536_
timestamp 0
transform -1 0 2630 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__537_
timestamp 0
transform -1 0 2910 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__538_
timestamp 0
transform -1 0 3190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__539_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__540_
timestamp 0
transform -1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__541_
timestamp 0
transform 1 0 310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__542_
timestamp 0
transform -1 0 350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__543_
timestamp 0
transform -1 0 3410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__544_
timestamp 0
transform -1 0 3670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__545_
timestamp 0
transform -1 0 3830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__546_
timestamp 0
transform 1 0 3510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__547_
timestamp 0
transform 1 0 2590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__548_
timestamp 0
transform -1 0 2170 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__549_
timestamp 0
transform -1 0 3490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__550_
timestamp 0
transform -1 0 3770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__551_
timestamp 0
transform 1 0 910 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__552_
timestamp 0
transform 1 0 610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__553_
timestamp 0
transform -1 0 850 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__554_
timestamp 0
transform 1 0 550 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__555_
timestamp 0
transform 1 0 330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__556_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__613_
timestamp 0
transform 1 0 4750 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__614_
timestamp 0
transform -1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__615_
timestamp 0
transform 1 0 4270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__616_
timestamp 0
transform -1 0 4330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__617_
timestamp 0
transform 1 0 4470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__618_
timestamp 0
transform 1 0 4790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__619_
timestamp 0
transform 1 0 4770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__620_
timestamp 0
transform 1 0 4630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__621_
timestamp 0
transform 1 0 4770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__622_
timestamp 0
transform 1 0 4830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__623_
timestamp 0
transform 1 0 4550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__624_
timestamp 0
transform 1 0 4590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__625_
timestamp 0
transform 1 0 3270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 4450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 4370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 4490 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform 1 0 4510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform -1 0 1190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 1750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 1730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 2390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform -1 0 570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 2770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 1830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform 1 0 2930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform -1 0 930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 2850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 3910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 3150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform -1 0 3410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform -1 0 2850 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 2770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert0
timestamp 0
transform -1 0 3570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert1
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert2
timestamp 0
transform 1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert3
timestamp 0
transform 1 0 2450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert4
timestamp 0
transform 1 0 4090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert5
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert6
timestamp 0
transform 1 0 3590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__273_
timestamp 0
transform -1 0 4310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__274_
timestamp 0
transform -1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__275_
timestamp 0
transform -1 0 4830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__276_
timestamp 0
transform -1 0 3630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__277_
timestamp 0
transform 1 0 4850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__278_
timestamp 0
transform 1 0 4810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__279_
timestamp 0
transform 1 0 4450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__280_
timestamp 0
transform -1 0 4670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__281_
timestamp 0
transform -1 0 4730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__282_
timestamp 0
transform 1 0 3910 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__283_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__284_
timestamp 0
transform 1 0 3930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__285_
timestamp 0
transform 1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__286_
timestamp 0
transform -1 0 4550 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__287_
timestamp 0
transform 1 0 4510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__288_
timestamp 0
transform 1 0 3450 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__289_
timestamp 0
transform -1 0 4230 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__290_
timestamp 0
transform 1 0 3970 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__291_
timestamp 0
transform 1 0 1370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__292_
timestamp 0
transform -1 0 3970 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__293_
timestamp 0
transform -1 0 4230 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__294_
timestamp 0
transform 1 0 3810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__295_
timestamp 0
transform -1 0 4270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__296_
timestamp 0
transform 1 0 4550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__297_
timestamp 0
transform 1 0 4070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__298_
timestamp 0
transform -1 0 3990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__299_
timestamp 0
transform -1 0 4030 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__300_
timestamp 0
transform 1 0 3170 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__301_
timestamp 0
transform -1 0 3710 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__302_
timestamp 0
transform -1 0 3730 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__303_
timestamp 0
transform 1 0 3730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__304_
timestamp 0
transform -1 0 3990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__305_
timestamp 0
transform -1 0 4270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__306_
timestamp 0
transform 1 0 3810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__307_
timestamp 0
transform 1 0 4270 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__308_
timestamp 0
transform 1 0 4070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__309_
timestamp 0
transform -1 0 650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__310_
timestamp 0
transform -1 0 70 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__311_
timestamp 0
transform -1 0 70 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__312_
timestamp 0
transform -1 0 310 0 1 250
box -6 -8 26 248
use FILL  FILL_2__313_
timestamp 0
transform 1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__314_
timestamp 0
transform 1 0 290 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__315_
timestamp 0
transform 1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__316_
timestamp 0
transform -1 0 830 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__317_
timestamp 0
transform 1 0 530 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__318_
timestamp 0
transform -1 0 730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__319_
timestamp 0
transform -1 0 830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__320_
timestamp 0
transform -1 0 1370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__321_
timestamp 0
transform 1 0 1510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__322_
timestamp 0
transform 1 0 1370 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__323_
timestamp 0
transform -1 0 470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__324_
timestamp 0
transform 1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__325_
timestamp 0
transform 1 0 290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__326_
timestamp 0
transform -1 0 310 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__327_
timestamp 0
transform -1 0 70 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__328_
timestamp 0
transform 1 0 590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__329_
timestamp 0
transform 1 0 350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__330_
timestamp 0
transform 1 0 2770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__331_
timestamp 0
transform 1 0 3330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__332_
timestamp 0
transform 1 0 3030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__333_
timestamp 0
transform 1 0 2250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__334_
timestamp 0
transform 1 0 1990 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__335_
timestamp 0
transform -1 0 1970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__336_
timestamp 0
transform -1 0 70 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__337_
timestamp 0
transform 1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__338_
timestamp 0
transform -1 0 330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__339_
timestamp 0
transform 1 0 3490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__340_
timestamp 0
transform -1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__341_
timestamp 0
transform -1 0 4490 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__342_
timestamp 0
transform 1 0 4170 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__343_
timestamp 0
transform 1 0 3510 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__344_
timestamp 0
transform 1 0 3530 0 1 730
box -6 -8 26 248
use FILL  FILL_2__345_
timestamp 0
transform 1 0 3970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__346_
timestamp 0
transform 1 0 4050 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__347_
timestamp 0
transform -1 0 4830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__348_
timestamp 0
transform 1 0 4570 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__349_
timestamp 0
transform 1 0 2530 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__350_
timestamp 0
transform -1 0 2950 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__351_
timestamp 0
transform 1 0 2910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__352_
timestamp 0
transform -1 0 2690 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__353_
timestamp 0
transform 1 0 2310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__354_
timestamp 0
transform -1 0 3230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__355_
timestamp 0
transform -1 0 4070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__356_
timestamp 0
transform 1 0 3750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__357_
timestamp 0
transform -1 0 2630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__358_
timestamp 0
transform -1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__359_
timestamp 0
transform 1 0 3070 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__360_
timestamp 0
transform -1 0 3370 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__361_
timestamp 0
transform -1 0 3150 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__362_
timestamp 0
transform -1 0 3090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__363_
timestamp 0
transform 1 0 2270 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__364_
timestamp 0
transform 1 0 2130 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__365_
timestamp 0
transform 1 0 3110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__366_
timestamp 0
transform 1 0 2790 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__367_
timestamp 0
transform -1 0 2050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__368_
timestamp 0
transform 1 0 2810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__369_
timestamp 0
transform -1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__370_
timestamp 0
transform 1 0 4850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__371_
timestamp 0
transform 1 0 4550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__372_
timestamp 0
transform 1 0 3230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__373_
timestamp 0
transform 1 0 3230 0 1 730
box -6 -8 26 248
use FILL  FILL_2__374_
timestamp 0
transform 1 0 4050 0 1 730
box -6 -8 26 248
use FILL  FILL_2__375_
timestamp 0
transform 1 0 3770 0 1 730
box -6 -8 26 248
use FILL  FILL_2__376_
timestamp 0
transform 1 0 4330 0 1 730
box -6 -8 26 248
use FILL  FILL_2__377_
timestamp 0
transform -1 0 4030 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__378_
timestamp 0
transform -1 0 4150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__379_
timestamp 0
transform -1 0 2250 0 1 250
box -6 -8 26 248
use FILL  FILL_2__380_
timestamp 0
transform 1 0 1570 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__381_
timestamp 0
transform 1 0 1270 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__382_
timestamp 0
transform -1 0 950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__383_
timestamp 0
transform 1 0 1410 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__384_
timestamp 0
transform -1 0 870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__385_
timestamp 0
transform -1 0 910 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__386_
timestamp 0
transform 1 0 970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__387_
timestamp 0
transform -1 0 790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__388_
timestamp 0
transform -1 0 3890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__389_
timestamp 0
transform -1 0 1490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__390_
timestamp 0
transform -1 0 1190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__391_
timestamp 0
transform 1 0 870 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__392_
timestamp 0
transform -1 0 670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__393_
timestamp 0
transform 1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__394_
timestamp 0
transform 1 0 1690 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__395_
timestamp 0
transform -1 0 3650 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__396_
timestamp 0
transform 1 0 1130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__397_
timestamp 0
transform 1 0 1390 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__398_
timestamp 0
transform 1 0 1930 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__399_
timestamp 0
transform 1 0 1930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__400_
timestamp 0
transform 1 0 1670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__401_
timestamp 0
transform 1 0 1390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__402_
timestamp 0
transform 1 0 1710 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__403_
timestamp 0
transform -1 0 2790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__404_
timestamp 0
transform 1 0 2490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__405_
timestamp 0
transform -1 0 1270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__406_
timestamp 0
transform 1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__407_
timestamp 0
transform -1 0 1430 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__408_
timestamp 0
transform -1 0 910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__409_
timestamp 0
transform 1 0 1170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__410_
timestamp 0
transform -1 0 1090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__411_
timestamp 0
transform -1 0 3170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__412_
timestamp 0
transform -1 0 1670 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__413_
timestamp 0
transform 1 0 1510 0 1 730
box -6 -8 26 248
use FILL  FILL_2__414_
timestamp 0
transform 1 0 1790 0 1 730
box -6 -8 26 248
use FILL  FILL_2__415_
timestamp 0
transform 1 0 2650 0 1 730
box -6 -8 26 248
use FILL  FILL_2__416_
timestamp 0
transform -1 0 2010 0 1 250
box -6 -8 26 248
use FILL  FILL_2__417_
timestamp 0
transform 1 0 2370 0 1 730
box -6 -8 26 248
use FILL  FILL_2__418_
timestamp 0
transform 1 0 2210 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__419_
timestamp 0
transform -1 0 2970 0 1 730
box -6 -8 26 248
use FILL  FILL_2__420_
timestamp 0
transform -1 0 2870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__421_
timestamp 0
transform 1 0 4530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__422_
timestamp 0
transform 1 0 4310 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__423_
timestamp 0
transform 1 0 4850 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__424_
timestamp 0
transform 1 0 4850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__425_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 26 248
use FILL  FILL_2__426_
timestamp 0
transform -1 0 4590 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__427_
timestamp 0
transform -1 0 2530 0 1 250
box -6 -8 26 248
use FILL  FILL_2__428_
timestamp 0
transform 1 0 2090 0 1 730
box -6 -8 26 248
use FILL  FILL_2__429_
timestamp 0
transform 1 0 2490 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__430_
timestamp 0
transform -1 0 1370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__431_
timestamp 0
transform 1 0 1650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__432_
timestamp 0
transform -1 0 2250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__433_
timestamp 0
transform 1 0 2510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__434_
timestamp 0
transform -1 0 4290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__435_
timestamp 0
transform 1 0 3410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__436_
timestamp 0
transform -1 0 3710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__437_
timestamp 0
transform -1 0 2250 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__438_
timestamp 0
transform -1 0 2510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__439_
timestamp 0
transform 1 0 2530 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__440_
timestamp 0
transform -1 0 3090 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__441_
timestamp 0
transform 1 0 1470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__442_
timestamp 0
transform -1 0 2050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__443_
timestamp 0
transform -1 0 1670 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__444_
timestamp 0
transform -1 0 2110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__445_
timestamp 0
transform -1 0 1810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__446_
timestamp 0
transform 1 0 1950 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__447_
timestamp 0
transform -1 0 4190 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__448_
timestamp 0
transform -1 0 1750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__449_
timestamp 0
transform 1 0 2230 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__450_
timestamp 0
transform 1 0 2310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__451_
timestamp 0
transform 1 0 2490 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__452_
timestamp 0
transform -1 0 3630 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__453_
timestamp 0
transform 1 0 1390 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__454_
timestamp 0
transform -1 0 1630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__455_
timestamp 0
transform 1 0 1970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__456_
timestamp 0
transform -1 0 1910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__457_
timestamp 0
transform 1 0 1650 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__458_
timestamp 0
transform 1 0 1730 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__459_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__460_
timestamp 0
transform -1 0 2510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__461_
timestamp 0
transform -1 0 2050 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__462_
timestamp 0
transform 1 0 2310 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__463_
timestamp 0
transform 1 0 2610 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__464_
timestamp 0
transform -1 0 2930 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__465_
timestamp 0
transform 1 0 1190 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__466_
timestamp 0
transform -1 0 910 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__467_
timestamp 0
transform 1 0 590 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__468_
timestamp 0
transform -1 0 350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__469_
timestamp 0
transform -1 0 330 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__470_
timestamp 0
transform -1 0 630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__471_
timestamp 0
transform 1 0 630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__472_
timestamp 0
transform -1 0 870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__473_
timestamp 0
transform 1 0 810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__474_
timestamp 0
transform 1 0 890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__475_
timestamp 0
transform -1 0 70 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__476_
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__477_
timestamp 0
transform 1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__478_
timestamp 0
transform -1 0 350 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__479_
timestamp 0
transform -1 0 3450 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__480_
timestamp 0
transform -1 0 1230 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__481_
timestamp 0
transform -1 0 70 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__482_
timestamp 0
transform -1 0 1190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__483_
timestamp 0
transform -1 0 1470 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__484_
timestamp 0
transform 1 0 1630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__485_
timestamp 0
transform 1 0 1930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__486_
timestamp 0
transform 1 0 2210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__487_
timestamp 0
transform 1 0 2790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__488_
timestamp 0
transform 1 0 2490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__489_
timestamp 0
transform 1 0 1470 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__490_
timestamp 0
transform -1 0 1750 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__491_
timestamp 0
transform 1 0 2030 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__492_
timestamp 0
transform 1 0 2310 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__493_
timestamp 0
transform -1 0 2630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__494_
timestamp 0
transform 1 0 1110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__495_
timestamp 0
transform 1 0 1390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__496_
timestamp 0
transform 1 0 1670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__497_
timestamp 0
transform 1 0 2050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__498_
timestamp 0
transform -1 0 2270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__499_
timestamp 0
transform -1 0 1750 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__500_
timestamp 0
transform -1 0 2290 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__501_
timestamp 0
transform -1 0 2670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__502_
timestamp 0
transform -1 0 3230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__503_
timestamp 0
transform -1 0 3310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__504_
timestamp 0
transform 1 0 4510 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__505_
timestamp 0
transform -1 0 4790 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__506_
timestamp 0
transform 1 0 4590 0 1 250
box -6 -8 26 248
use FILL  FILL_2__507_
timestamp 0
transform -1 0 4630 0 1 730
box -6 -8 26 248
use FILL  FILL_2__508_
timestamp 0
transform -1 0 2870 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__509_
timestamp 0
transform 1 0 2010 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__510_
timestamp 0
transform -1 0 2570 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__511_
timestamp 0
transform 1 0 1470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__512_
timestamp 0
transform 1 0 2350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__513_
timestamp 0
transform -1 0 3130 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__514_
timestamp 0
transform 1 0 3370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__515_
timestamp 0
transform -1 0 3690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__516_
timestamp 0
transform 1 0 590 0 1 250
box -6 -8 26 248
use FILL  FILL_2__517_
timestamp 0
transform 1 0 870 0 1 250
box -6 -8 26 248
use FILL  FILL_2__518_
timestamp 0
transform 1 0 1430 0 1 250
box -6 -8 26 248
use FILL  FILL_2__519_
timestamp 0
transform 1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_2__520_
timestamp 0
transform -1 0 1570 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__521_
timestamp 0
transform -1 0 1850 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__522_
timestamp 0
transform -1 0 3510 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__523_
timestamp 0
transform -1 0 3790 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__524_
timestamp 0
transform -1 0 1130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__525_
timestamp 0
transform 1 0 1150 0 1 250
box -6 -8 26 248
use FILL  FILL_2__526_
timestamp 0
transform -1 0 850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__527_
timestamp 0
transform -1 0 990 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__528_
timestamp 0
transform 1 0 3050 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__529_
timestamp 0
transform 1 0 1230 0 1 730
box -6 -8 26 248
use FILL  FILL_2__530_
timestamp 0
transform 1 0 930 0 1 730
box -6 -8 26 248
use FILL  FILL_2__531_
timestamp 0
transform -1 0 470 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__532_
timestamp 0
transform 1 0 310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__533_
timestamp 0
transform -1 0 350 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__534_
timestamp 0
transform 1 0 610 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__535_
timestamp 0
transform -1 0 2370 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__536_
timestamp 0
transform -1 0 2650 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__537_
timestamp 0
transform -1 0 2930 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__538_
timestamp 0
transform -1 0 3210 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__539_
timestamp 0
transform -1 0 70 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__540_
timestamp 0
transform -1 0 70 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__541_
timestamp 0
transform 1 0 330 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__542_
timestamp 0
transform -1 0 370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__543_
timestamp 0
transform -1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__544_
timestamp 0
transform -1 0 3690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__545_
timestamp 0
transform -1 0 3850 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__546_
timestamp 0
transform 1 0 3530 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__547_
timestamp 0
transform 1 0 2610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__548_
timestamp 0
transform -1 0 2190 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__549_
timestamp 0
transform -1 0 3510 0 1 250
box -6 -8 26 248
use FILL  FILL_2__550_
timestamp 0
transform -1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__551_
timestamp 0
transform 1 0 930 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__552_
timestamp 0
transform 1 0 630 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__553_
timestamp 0
transform -1 0 870 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__554_
timestamp 0
transform 1 0 570 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__555_
timestamp 0
transform 1 0 350 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__556_
timestamp 0
transform -1 0 70 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__613_
timestamp 0
transform 1 0 4770 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__614_
timestamp 0
transform -1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__615_
timestamp 0
transform 1 0 4290 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__616_
timestamp 0
transform -1 0 4350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__617_
timestamp 0
transform 1 0 4490 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__618_
timestamp 0
transform 1 0 4810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__619_
timestamp 0
transform 1 0 4790 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__620_
timestamp 0
transform 1 0 4650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__621_
timestamp 0
transform 1 0 4790 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__622_
timestamp 0
transform 1 0 4850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__623_
timestamp 0
transform 1 0 4570 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__624_
timestamp 0
transform 1 0 4610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__625_
timestamp 0
transform 1 0 3290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform 1 0 4470 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 4390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert9
timestamp 0
transform 1 0 4510 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform 1 0 4530 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform -1 0 1210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 1770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 1750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 2410 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform -1 0 590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 2790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform 1 0 2950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform -1 0 950 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 2870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform 1 0 3930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 3170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform -1 0 3430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform -1 0 2870 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform 1 0 2790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert0
timestamp 0
transform -1 0 3590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert1
timestamp 0
transform -1 0 70 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert2
timestamp 0
transform 1 0 50 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert3
timestamp 0
transform 1 0 2470 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert4
timestamp 0
transform 1 0 4110 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert5
timestamp 0
transform -1 0 310 0 1 730
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert6
timestamp 0
transform 1 0 3610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__273_
timestamp 0
transform -1 0 4330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__274_
timestamp 0
transform -1 0 4570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__275_
timestamp 0
transform -1 0 4850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__276_
timestamp 0
transform -1 0 3650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__277_
timestamp 0
transform 1 0 4870 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__278_
timestamp 0
transform 1 0 4830 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__279_
timestamp 0
transform 1 0 4470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__280_
timestamp 0
transform -1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__281_
timestamp 0
transform -1 0 4750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__282_
timestamp 0
transform 1 0 3930 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__283_
timestamp 0
transform -1 0 3450 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__284_
timestamp 0
transform 1 0 3950 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__285_
timestamp 0
transform 1 0 3330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__286_
timestamp 0
transform -1 0 4570 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__287_
timestamp 0
transform 1 0 4530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__288_
timestamp 0
transform 1 0 3470 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__289_
timestamp 0
transform -1 0 4250 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__290_
timestamp 0
transform 1 0 3990 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__291_
timestamp 0
transform 1 0 1390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__292_
timestamp 0
transform -1 0 3990 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__293_
timestamp 0
transform -1 0 4250 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__294_
timestamp 0
transform 1 0 3830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__295_
timestamp 0
transform -1 0 4290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__296_
timestamp 0
transform 1 0 4570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__297_
timestamp 0
transform 1 0 4090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__298_
timestamp 0
transform -1 0 4010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__299_
timestamp 0
transform -1 0 4050 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__300_
timestamp 0
transform 1 0 3190 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__301_
timestamp 0
transform -1 0 3730 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__302_
timestamp 0
transform -1 0 3750 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__303_
timestamp 0
transform 1 0 3750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__304_
timestamp 0
transform -1 0 4010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__305_
timestamp 0
transform -1 0 4290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__306_
timestamp 0
transform 1 0 3830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__307_
timestamp 0
transform 1 0 4290 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__308_
timestamp 0
transform 1 0 4090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__309_
timestamp 0
transform -1 0 670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__310_
timestamp 0
transform -1 0 90 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__311_
timestamp 0
transform -1 0 90 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__312_
timestamp 0
transform -1 0 330 0 1 250
box -6 -8 26 248
use FILL  FILL_3__313_
timestamp 0
transform 1 0 310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__314_
timestamp 0
transform 1 0 310 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__315_
timestamp 0
transform 1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__316_
timestamp 0
transform -1 0 850 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__317_
timestamp 0
transform 1 0 550 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__318_
timestamp 0
transform -1 0 750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__319_
timestamp 0
transform -1 0 850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__320_
timestamp 0
transform -1 0 1390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__321_
timestamp 0
transform 1 0 1530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__322_
timestamp 0
transform 1 0 1390 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__323_
timestamp 0
transform -1 0 490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__324_
timestamp 0
transform 1 0 70 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__325_
timestamp 0
transform 1 0 310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__326_
timestamp 0
transform -1 0 330 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__327_
timestamp 0
transform -1 0 90 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__328_
timestamp 0
transform 1 0 610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__329_
timestamp 0
transform 1 0 370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__330_
timestamp 0
transform 1 0 2790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__331_
timestamp 0
transform 1 0 3350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__332_
timestamp 0
transform 1 0 3050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__333_
timestamp 0
transform 1 0 2270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__334_
timestamp 0
transform 1 0 2010 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__335_
timestamp 0
transform -1 0 1990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__336_
timestamp 0
transform -1 0 90 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__337_
timestamp 0
transform 1 0 70 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__338_
timestamp 0
transform -1 0 350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__339_
timestamp 0
transform 1 0 3510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__340_
timestamp 0
transform -1 0 4030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__341_
timestamp 0
transform -1 0 4510 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__342_
timestamp 0
transform 1 0 4190 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__343_
timestamp 0
transform 1 0 3530 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__344_
timestamp 0
transform 1 0 3550 0 1 730
box -6 -8 26 248
use FILL  FILL_3__345_
timestamp 0
transform 1 0 3990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__346_
timestamp 0
transform 1 0 4070 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__347_
timestamp 0
transform -1 0 4850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__348_
timestamp 0
transform 1 0 4590 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__349_
timestamp 0
transform 1 0 2550 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__350_
timestamp 0
transform -1 0 2970 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__351_
timestamp 0
transform 1 0 2930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__352_
timestamp 0
transform -1 0 2710 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__353_
timestamp 0
transform 1 0 2330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__354_
timestamp 0
transform -1 0 3250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__355_
timestamp 0
transform -1 0 4090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__356_
timestamp 0
transform 1 0 3770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__357_
timestamp 0
transform -1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__358_
timestamp 0
transform -1 0 2830 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__359_
timestamp 0
transform 1 0 3090 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__360_
timestamp 0
transform -1 0 3390 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__361_
timestamp 0
transform -1 0 3170 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__362_
timestamp 0
transform -1 0 3110 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__363_
timestamp 0
transform 1 0 2290 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__364_
timestamp 0
transform 1 0 2150 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__365_
timestamp 0
transform 1 0 3130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__366_
timestamp 0
transform 1 0 2810 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__367_
timestamp 0
transform -1 0 2070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__368_
timestamp 0
transform 1 0 2830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__369_
timestamp 0
transform -1 0 3270 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__370_
timestamp 0
transform 1 0 4870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__371_
timestamp 0
transform 1 0 4570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__372_
timestamp 0
transform 1 0 3250 0 1 250
box -6 -8 26 248
use FILL  FILL_3__373_
timestamp 0
transform 1 0 3250 0 1 730
box -6 -8 26 248
use FILL  FILL_3__374_
timestamp 0
transform 1 0 4070 0 1 730
box -6 -8 26 248
use FILL  FILL_3__375_
timestamp 0
transform 1 0 3790 0 1 730
box -6 -8 26 248
use FILL  FILL_3__376_
timestamp 0
transform 1 0 4350 0 1 730
box -6 -8 26 248
use FILL  FILL_3__377_
timestamp 0
transform -1 0 4050 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__378_
timestamp 0
transform -1 0 4170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__379_
timestamp 0
transform -1 0 2270 0 1 250
box -6 -8 26 248
use FILL  FILL_3__380_
timestamp 0
transform 1 0 1590 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__381_
timestamp 0
transform 1 0 1290 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__382_
timestamp 0
transform -1 0 970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__383_
timestamp 0
transform 1 0 1430 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__384_
timestamp 0
transform -1 0 890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__385_
timestamp 0
transform -1 0 930 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__386_
timestamp 0
transform 1 0 990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__387_
timestamp 0
transform -1 0 810 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__388_
timestamp 0
transform -1 0 3910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__389_
timestamp 0
transform -1 0 1510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__390_
timestamp 0
transform -1 0 1210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__391_
timestamp 0
transform 1 0 890 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__392_
timestamp 0
transform -1 0 690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__393_
timestamp 0
transform 1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__394_
timestamp 0
transform 1 0 1710 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__395_
timestamp 0
transform -1 0 3670 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__396_
timestamp 0
transform 1 0 1150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__397_
timestamp 0
transform 1 0 1410 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__398_
timestamp 0
transform 1 0 1950 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__399_
timestamp 0
transform 1 0 1950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__400_
timestamp 0
transform 1 0 1690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__401_
timestamp 0
transform 1 0 1410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__402_
timestamp 0
transform 1 0 1730 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__403_
timestamp 0
transform -1 0 2810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__404_
timestamp 0
transform 1 0 2510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__405_
timestamp 0
transform -1 0 1290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__406_
timestamp 0
transform 1 0 1170 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__407_
timestamp 0
transform -1 0 1450 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__408_
timestamp 0
transform -1 0 930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__409_
timestamp 0
transform 1 0 1190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__410_
timestamp 0
transform -1 0 1110 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__411_
timestamp 0
transform -1 0 3190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__412_
timestamp 0
transform -1 0 1690 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__413_
timestamp 0
transform 1 0 1530 0 1 730
box -6 -8 26 248
use FILL  FILL_3__414_
timestamp 0
transform 1 0 1810 0 1 730
box -6 -8 26 248
use FILL  FILL_3__415_
timestamp 0
transform 1 0 2670 0 1 730
box -6 -8 26 248
use FILL  FILL_3__416_
timestamp 0
transform -1 0 2030 0 1 250
box -6 -8 26 248
use FILL  FILL_3__417_
timestamp 0
transform 1 0 2390 0 1 730
box -6 -8 26 248
use FILL  FILL_3__418_
timestamp 0
transform 1 0 2230 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__419_
timestamp 0
transform -1 0 2990 0 1 730
box -6 -8 26 248
use FILL  FILL_3__420_
timestamp 0
transform -1 0 2890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__421_
timestamp 0
transform 1 0 4550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__422_
timestamp 0
transform 1 0 4330 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__423_
timestamp 0
transform 1 0 4870 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__424_
timestamp 0
transform 1 0 4870 0 1 250
box -6 -8 26 248
use FILL  FILL_3__425_
timestamp 0
transform 1 0 4330 0 1 250
box -6 -8 26 248
use FILL  FILL_3__426_
timestamp 0
transform -1 0 4610 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__427_
timestamp 0
transform -1 0 2550 0 1 250
box -6 -8 26 248
use FILL  FILL_3__428_
timestamp 0
transform 1 0 2110 0 1 730
box -6 -8 26 248
use FILL  FILL_3__429_
timestamp 0
transform 1 0 2510 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__430_
timestamp 0
transform -1 0 1390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__431_
timestamp 0
transform 1 0 1670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__432_
timestamp 0
transform -1 0 2270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__433_
timestamp 0
transform 1 0 2530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__434_
timestamp 0
transform -1 0 4310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__435_
timestamp 0
transform 1 0 3430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__436_
timestamp 0
transform -1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__437_
timestamp 0
transform -1 0 2270 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__438_
timestamp 0
transform -1 0 2530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__439_
timestamp 0
transform 1 0 2550 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__440_
timestamp 0
transform -1 0 3110 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__441_
timestamp 0
transform 1 0 1490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__442_
timestamp 0
transform -1 0 2070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__443_
timestamp 0
transform -1 0 1690 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__444_
timestamp 0
transform -1 0 2130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__445_
timestamp 0
transform -1 0 1830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__446_
timestamp 0
transform 1 0 1970 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__447_
timestamp 0
transform -1 0 4210 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__448_
timestamp 0
transform -1 0 1770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__449_
timestamp 0
transform 1 0 2250 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__450_
timestamp 0
transform 1 0 2330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__451_
timestamp 0
transform 1 0 2510 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__452_
timestamp 0
transform -1 0 3650 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__453_
timestamp 0
transform 1 0 1410 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__454_
timestamp 0
transform -1 0 1650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__455_
timestamp 0
transform 1 0 1990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__456_
timestamp 0
transform -1 0 1930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__457_
timestamp 0
transform 1 0 1670 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__458_
timestamp 0
transform 1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__459_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__460_
timestamp 0
transform -1 0 2530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__461_
timestamp 0
transform -1 0 2070 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__462_
timestamp 0
transform 1 0 2330 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__463_
timestamp 0
transform 1 0 2630 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__464_
timestamp 0
transform -1 0 2950 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__465_
timestamp 0
transform 1 0 1210 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__466_
timestamp 0
transform -1 0 930 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__467_
timestamp 0
transform 1 0 610 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__468_
timestamp 0
transform -1 0 370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__469_
timestamp 0
transform -1 0 350 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__470_
timestamp 0
transform -1 0 650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__471_
timestamp 0
transform 1 0 650 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__472_
timestamp 0
transform -1 0 890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__473_
timestamp 0
transform 1 0 830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__474_
timestamp 0
transform 1 0 910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__475_
timestamp 0
transform -1 0 90 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__476_
timestamp 0
transform -1 0 90 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__477_
timestamp 0
transform 1 0 330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__478_
timestamp 0
transform -1 0 370 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__479_
timestamp 0
transform -1 0 3470 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__480_
timestamp 0
transform -1 0 1250 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__481_
timestamp 0
transform -1 0 90 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__482_
timestamp 0
transform -1 0 1210 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__483_
timestamp 0
transform -1 0 1490 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__484_
timestamp 0
transform 1 0 1650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__485_
timestamp 0
transform 1 0 1950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__486_
timestamp 0
transform 1 0 2230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__487_
timestamp 0
transform 1 0 2810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__488_
timestamp 0
transform 1 0 2510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__489_
timestamp 0
transform 1 0 1490 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__490_
timestamp 0
transform -1 0 1770 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__491_
timestamp 0
transform 1 0 2050 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__492_
timestamp 0
transform 1 0 2330 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__493_
timestamp 0
transform -1 0 2650 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__494_
timestamp 0
transform 1 0 1130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__495_
timestamp 0
transform 1 0 1410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__496_
timestamp 0
transform 1 0 1690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__497_
timestamp 0
transform 1 0 2070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__498_
timestamp 0
transform -1 0 2290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__499_
timestamp 0
transform -1 0 1770 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__500_
timestamp 0
transform -1 0 2310 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__501_
timestamp 0
transform -1 0 2690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__502_
timestamp 0
transform -1 0 3250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__503_
timestamp 0
transform -1 0 3330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__504_
timestamp 0
transform 1 0 4530 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__505_
timestamp 0
transform -1 0 4810 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__506_
timestamp 0
transform 1 0 4610 0 1 250
box -6 -8 26 248
use FILL  FILL_3__507_
timestamp 0
transform -1 0 4650 0 1 730
box -6 -8 26 248
use FILL  FILL_3__508_
timestamp 0
transform -1 0 2890 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__509_
timestamp 0
transform 1 0 2030 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__510_
timestamp 0
transform -1 0 2590 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__511_
timestamp 0
transform 1 0 1490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__512_
timestamp 0
transform 1 0 2370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__513_
timestamp 0
transform -1 0 3150 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__514_
timestamp 0
transform 1 0 3390 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__515_
timestamp 0
transform -1 0 3710 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__516_
timestamp 0
transform 1 0 610 0 1 250
box -6 -8 26 248
use FILL  FILL_3__517_
timestamp 0
transform 1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_3__518_
timestamp 0
transform 1 0 1450 0 1 250
box -6 -8 26 248
use FILL  FILL_3__519_
timestamp 0
transform 1 0 1730 0 1 250
box -6 -8 26 248
use FILL  FILL_3__520_
timestamp 0
transform -1 0 1590 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__521_
timestamp 0
transform -1 0 1870 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__522_
timestamp 0
transform -1 0 3530 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__523_
timestamp 0
transform -1 0 3810 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__524_
timestamp 0
transform -1 0 1150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__525_
timestamp 0
transform 1 0 1170 0 1 250
box -6 -8 26 248
use FILL  FILL_3__526_
timestamp 0
transform -1 0 870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__527_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__528_
timestamp 0
transform 1 0 3070 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__529_
timestamp 0
transform 1 0 1250 0 1 730
box -6 -8 26 248
use FILL  FILL_3__530_
timestamp 0
transform 1 0 950 0 1 730
box -6 -8 26 248
use FILL  FILL_3__531_
timestamp 0
transform -1 0 490 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__532_
timestamp 0
transform 1 0 330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__533_
timestamp 0
transform -1 0 370 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__534_
timestamp 0
transform 1 0 630 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__535_
timestamp 0
transform -1 0 2390 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__536_
timestamp 0
transform -1 0 2670 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__537_
timestamp 0
transform -1 0 2950 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__538_
timestamp 0
transform -1 0 3230 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__539_
timestamp 0
transform -1 0 90 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__540_
timestamp 0
transform -1 0 90 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__541_
timestamp 0
transform 1 0 350 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__542_
timestamp 0
transform -1 0 390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__543_
timestamp 0
transform -1 0 3450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__544_
timestamp 0
transform -1 0 3710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__545_
timestamp 0
transform -1 0 3870 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__546_
timestamp 0
transform 1 0 3550 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__547_
timestamp 0
transform 1 0 2630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__548_
timestamp 0
transform -1 0 2210 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__549_
timestamp 0
transform -1 0 3530 0 1 250
box -6 -8 26 248
use FILL  FILL_3__550_
timestamp 0
transform -1 0 3810 0 1 250
box -6 -8 26 248
use FILL  FILL_3__551_
timestamp 0
transform 1 0 950 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__552_
timestamp 0
transform 1 0 650 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__553_
timestamp 0
transform -1 0 890 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__554_
timestamp 0
transform 1 0 590 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__555_
timestamp 0
transform 1 0 370 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__556_
timestamp 0
transform -1 0 90 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__613_
timestamp 0
transform 1 0 4790 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__614_
timestamp 0
transform -1 0 4770 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__615_
timestamp 0
transform 1 0 4310 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__616_
timestamp 0
transform -1 0 4370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__617_
timestamp 0
transform 1 0 4510 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__618_
timestamp 0
transform 1 0 4830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__619_
timestamp 0
transform 1 0 4810 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__620_
timestamp 0
transform 1 0 4670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__621_
timestamp 0
transform 1 0 4810 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__622_
timestamp 0
transform 1 0 4870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__623_
timestamp 0
transform 1 0 4590 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__624_
timestamp 0
transform 1 0 4630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__625_
timestamp 0
transform 1 0 3310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert7
timestamp 0
transform 1 0 4490 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert8
timestamp 0
transform -1 0 4410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert9
timestamp 0
transform 1 0 4530 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert10
timestamp 0
transform 1 0 4550 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform -1 0 1230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 1790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform 1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform 1 0 2430 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform -1 0 610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 2810 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 1870 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform 1 0 2970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform -1 0 970 0 1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert20
timestamp 0
transform 1 0 2890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert21
timestamp 0
transform 1 0 3950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert22
timestamp 0
transform -1 0 3190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert23
timestamp 0
transform -1 0 3450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert24
timestamp 0
transform -1 0 2890 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert25
timestamp 0
transform 1 0 2810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert0
timestamp 0
transform -1 0 3610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert1
timestamp 0
transform -1 0 90 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert2
timestamp 0
transform 1 0 70 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert3
timestamp 0
transform 1 0 2490 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert4
timestamp 0
transform 1 0 4130 0 -1 730
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert5
timestamp 0
transform -1 0 330 0 1 730
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert6
timestamp 0
transform 1 0 3630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__273_
timestamp 0
transform -1 0 4350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__274_
timestamp 0
transform -1 0 4590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__275_
timestamp 0
transform -1 0 4870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__276_
timestamp 0
transform -1 0 3670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__277_
timestamp 0
transform 1 0 4890 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__278_
timestamp 0
transform 1 0 4850 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__279_
timestamp 0
transform 1 0 4490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__280_
timestamp 0
transform -1 0 4710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__281_
timestamp 0
transform -1 0 4770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__282_
timestamp 0
transform 1 0 3950 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__283_
timestamp 0
transform -1 0 3470 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__284_
timestamp 0
transform 1 0 3970 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__285_
timestamp 0
transform 1 0 3350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__286_
timestamp 0
transform -1 0 4590 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__287_
timestamp 0
transform 1 0 4550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__288_
timestamp 0
transform 1 0 3490 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__289_
timestamp 0
transform -1 0 4270 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__290_
timestamp 0
transform 1 0 4010 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__291_
timestamp 0
transform 1 0 1410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__292_
timestamp 0
transform -1 0 4010 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__293_
timestamp 0
transform -1 0 4270 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__294_
timestamp 0
transform 1 0 3850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__295_
timestamp 0
transform -1 0 4310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__296_
timestamp 0
transform 1 0 4590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__297_
timestamp 0
transform 1 0 4110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__298_
timestamp 0
transform -1 0 4030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__299_
timestamp 0
transform -1 0 4070 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__300_
timestamp 0
transform 1 0 3210 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__301_
timestamp 0
transform -1 0 3750 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__302_
timestamp 0
transform -1 0 3770 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__303_
timestamp 0
transform 1 0 3770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__304_
timestamp 0
transform -1 0 4030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__305_
timestamp 0
transform -1 0 4310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__306_
timestamp 0
transform 1 0 3850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__307_
timestamp 0
transform 1 0 4310 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__308_
timestamp 0
transform 1 0 4110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__309_
timestamp 0
transform -1 0 690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__310_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__311_
timestamp 0
transform -1 0 110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__312_
timestamp 0
transform -1 0 350 0 1 250
box -6 -8 26 248
use FILL  FILL_4__313_
timestamp 0
transform 1 0 330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__314_
timestamp 0
transform 1 0 330 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__315_
timestamp 0
transform 1 0 1510 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__316_
timestamp 0
transform -1 0 870 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__317_
timestamp 0
transform 1 0 570 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__318_
timestamp 0
transform -1 0 770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__319_
timestamp 0
transform -1 0 870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__320_
timestamp 0
transform -1 0 1410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__321_
timestamp 0
transform 1 0 1550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__322_
timestamp 0
transform 1 0 1410 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__323_
timestamp 0
transform -1 0 510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__324_
timestamp 0
transform 1 0 90 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__325_
timestamp 0
transform 1 0 330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__326_
timestamp 0
transform -1 0 350 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__327_
timestamp 0
transform -1 0 110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__328_
timestamp 0
transform 1 0 630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__329_
timestamp 0
transform 1 0 390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__330_
timestamp 0
transform 1 0 2810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__331_
timestamp 0
transform 1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__332_
timestamp 0
transform 1 0 3070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__333_
timestamp 0
transform 1 0 2290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__334_
timestamp 0
transform 1 0 2030 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__335_
timestamp 0
transform -1 0 2010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__336_
timestamp 0
transform -1 0 110 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__337_
timestamp 0
transform 1 0 90 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__338_
timestamp 0
transform -1 0 370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__339_
timestamp 0
transform 1 0 3530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__340_
timestamp 0
transform -1 0 4050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__341_
timestamp 0
transform -1 0 4530 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__342_
timestamp 0
transform 1 0 4210 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__343_
timestamp 0
transform 1 0 3550 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__344_
timestamp 0
transform 1 0 3570 0 1 730
box -6 -8 26 248
use FILL  FILL_4__345_
timestamp 0
transform 1 0 4010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__346_
timestamp 0
transform 1 0 4090 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__347_
timestamp 0
transform -1 0 4870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__348_
timestamp 0
transform 1 0 4610 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__349_
timestamp 0
transform 1 0 2570 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__350_
timestamp 0
transform -1 0 2990 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__351_
timestamp 0
transform 1 0 2950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__352_
timestamp 0
transform -1 0 2730 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__353_
timestamp 0
transform 1 0 2350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__354_
timestamp 0
transform -1 0 3270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__355_
timestamp 0
transform -1 0 4110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__356_
timestamp 0
transform 1 0 3790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__357_
timestamp 0
transform -1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__358_
timestamp 0
transform -1 0 2850 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__359_
timestamp 0
transform 1 0 3110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__360_
timestamp 0
transform -1 0 3410 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__361_
timestamp 0
transform -1 0 3190 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__362_
timestamp 0
transform -1 0 3130 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__363_
timestamp 0
transform 1 0 2310 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__364_
timestamp 0
transform 1 0 2170 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__365_
timestamp 0
transform 1 0 3150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__366_
timestamp 0
transform 1 0 2830 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__367_
timestamp 0
transform -1 0 2090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__368_
timestamp 0
transform 1 0 2850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__369_
timestamp 0
transform -1 0 3290 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__370_
timestamp 0
transform 1 0 4890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__371_
timestamp 0
transform 1 0 4590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__372_
timestamp 0
transform 1 0 3270 0 1 250
box -6 -8 26 248
use FILL  FILL_4__373_
timestamp 0
transform 1 0 3270 0 1 730
box -6 -8 26 248
use FILL  FILL_4__374_
timestamp 0
transform 1 0 4090 0 1 730
box -6 -8 26 248
use FILL  FILL_4__375_
timestamp 0
transform 1 0 3810 0 1 730
box -6 -8 26 248
use FILL  FILL_4__376_
timestamp 0
transform 1 0 4370 0 1 730
box -6 -8 26 248
use FILL  FILL_4__377_
timestamp 0
transform -1 0 4070 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__378_
timestamp 0
transform -1 0 4190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__379_
timestamp 0
transform -1 0 2290 0 1 250
box -6 -8 26 248
use FILL  FILL_4__380_
timestamp 0
transform 1 0 1610 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__381_
timestamp 0
transform 1 0 1310 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__382_
timestamp 0
transform -1 0 990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__383_
timestamp 0
transform 1 0 1450 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__384_
timestamp 0
transform -1 0 910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__385_
timestamp 0
transform -1 0 950 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__386_
timestamp 0
transform 1 0 1010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__387_
timestamp 0
transform -1 0 830 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__388_
timestamp 0
transform -1 0 3930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__389_
timestamp 0
transform -1 0 1530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__390_
timestamp 0
transform -1 0 1230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__391_
timestamp 0
transform 1 0 910 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__392_
timestamp 0
transform -1 0 710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__393_
timestamp 0
transform 1 0 1170 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__394_
timestamp 0
transform 1 0 1730 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__395_
timestamp 0
transform -1 0 3690 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__396_
timestamp 0
transform 1 0 1170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__397_
timestamp 0
transform 1 0 1430 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__398_
timestamp 0
transform 1 0 1970 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__399_
timestamp 0
transform 1 0 1970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__400_
timestamp 0
transform 1 0 1710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__401_
timestamp 0
transform 1 0 1430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__402_
timestamp 0
transform 1 0 1750 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__403_
timestamp 0
transform -1 0 2830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__404_
timestamp 0
transform 1 0 2530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__405_
timestamp 0
transform -1 0 1310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__406_
timestamp 0
transform 1 0 1190 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__407_
timestamp 0
transform -1 0 1470 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__408_
timestamp 0
transform -1 0 950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__409_
timestamp 0
transform 1 0 1210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__410_
timestamp 0
transform -1 0 1130 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__411_
timestamp 0
transform -1 0 3210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__412_
timestamp 0
transform -1 0 1710 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__413_
timestamp 0
transform 1 0 1550 0 1 730
box -6 -8 26 248
use FILL  FILL_4__414_
timestamp 0
transform 1 0 1830 0 1 730
box -6 -8 26 248
use FILL  FILL_4__415_
timestamp 0
transform 1 0 2690 0 1 730
box -6 -8 26 248
use FILL  FILL_4__416_
timestamp 0
transform -1 0 2050 0 1 250
box -6 -8 26 248
use FILL  FILL_4__417_
timestamp 0
transform 1 0 2410 0 1 730
box -6 -8 26 248
use FILL  FILL_4__418_
timestamp 0
transform 1 0 2250 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__419_
timestamp 0
transform -1 0 3010 0 1 730
box -6 -8 26 248
use FILL  FILL_4__420_
timestamp 0
transform -1 0 2910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__421_
timestamp 0
transform 1 0 4570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__422_
timestamp 0
transform 1 0 4350 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__423_
timestamp 0
transform 1 0 4890 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__424_
timestamp 0
transform 1 0 4890 0 1 250
box -6 -8 26 248
use FILL  FILL_4__425_
timestamp 0
transform 1 0 4350 0 1 250
box -6 -8 26 248
use FILL  FILL_4__426_
timestamp 0
transform -1 0 4630 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__427_
timestamp 0
transform -1 0 2570 0 1 250
box -6 -8 26 248
use FILL  FILL_4__428_
timestamp 0
transform 1 0 2130 0 1 730
box -6 -8 26 248
use FILL  FILL_4__429_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__430_
timestamp 0
transform -1 0 1410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__431_
timestamp 0
transform 1 0 1690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__432_
timestamp 0
transform -1 0 2290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__433_
timestamp 0
transform 1 0 2550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__434_
timestamp 0
transform -1 0 4330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__435_
timestamp 0
transform 1 0 3450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__436_
timestamp 0
transform -1 0 3750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__437_
timestamp 0
transform -1 0 2290 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__438_
timestamp 0
transform -1 0 2550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__439_
timestamp 0
transform 1 0 2570 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__440_
timestamp 0
transform -1 0 3130 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__441_
timestamp 0
transform 1 0 1510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__442_
timestamp 0
transform -1 0 2090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__443_
timestamp 0
transform -1 0 1710 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__444_
timestamp 0
transform -1 0 2150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__445_
timestamp 0
transform -1 0 1850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__446_
timestamp 0
transform 1 0 1990 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__447_
timestamp 0
transform -1 0 4230 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__448_
timestamp 0
transform -1 0 1790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__449_
timestamp 0
transform 1 0 2270 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__450_
timestamp 0
transform 1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__451_
timestamp 0
transform 1 0 2530 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__452_
timestamp 0
transform -1 0 3670 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__453_
timestamp 0
transform 1 0 1430 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__454_
timestamp 0
transform -1 0 1670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__455_
timestamp 0
transform 1 0 2010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__456_
timestamp 0
transform -1 0 1950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__457_
timestamp 0
transform 1 0 1690 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__458_
timestamp 0
transform 1 0 1770 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__459_
timestamp 0
transform 1 0 2230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__460_
timestamp 0
transform -1 0 2550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__461_
timestamp 0
transform -1 0 2090 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__462_
timestamp 0
transform 1 0 2350 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__463_
timestamp 0
transform 1 0 2650 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__464_
timestamp 0
transform -1 0 2970 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__465_
timestamp 0
transform 1 0 1230 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__466_
timestamp 0
transform -1 0 950 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__467_
timestamp 0
transform 1 0 630 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__468_
timestamp 0
transform -1 0 390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__469_
timestamp 0
transform -1 0 370 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__470_
timestamp 0
transform -1 0 670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__471_
timestamp 0
transform 1 0 670 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__472_
timestamp 0
transform -1 0 910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__473_
timestamp 0
transform 1 0 850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__474_
timestamp 0
transform 1 0 930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__475_
timestamp 0
transform -1 0 110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__476_
timestamp 0
transform -1 0 110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__477_
timestamp 0
transform 1 0 350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__478_
timestamp 0
transform -1 0 390 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__479_
timestamp 0
transform -1 0 3490 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__480_
timestamp 0
transform -1 0 1270 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__481_
timestamp 0
transform -1 0 110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__482_
timestamp 0
transform -1 0 1230 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__483_
timestamp 0
transform -1 0 1510 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__484_
timestamp 0
transform 1 0 1670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__485_
timestamp 0
transform 1 0 1970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__486_
timestamp 0
transform 1 0 2250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__487_
timestamp 0
transform 1 0 2830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__488_
timestamp 0
transform 1 0 2530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__489_
timestamp 0
transform 1 0 1510 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__490_
timestamp 0
transform -1 0 1790 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__491_
timestamp 0
transform 1 0 2070 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__492_
timestamp 0
transform 1 0 2350 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__493_
timestamp 0
transform -1 0 2670 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__494_
timestamp 0
transform 1 0 1150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__495_
timestamp 0
transform 1 0 1430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__496_
timestamp 0
transform 1 0 1710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__497_
timestamp 0
transform 1 0 2090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__498_
timestamp 0
transform -1 0 2310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__499_
timestamp 0
transform -1 0 1790 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__500_
timestamp 0
transform -1 0 2330 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__501_
timestamp 0
transform -1 0 2710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__502_
timestamp 0
transform -1 0 3270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__503_
timestamp 0
transform -1 0 3350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__504_
timestamp 0
transform 1 0 4550 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__505_
timestamp 0
transform -1 0 4830 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__506_
timestamp 0
transform 1 0 4630 0 1 250
box -6 -8 26 248
use FILL  FILL_4__507_
timestamp 0
transform -1 0 4670 0 1 730
box -6 -8 26 248
use FILL  FILL_4__508_
timestamp 0
transform -1 0 2910 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__509_
timestamp 0
transform 1 0 2050 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__510_
timestamp 0
transform -1 0 2610 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__511_
timestamp 0
transform 1 0 1510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__512_
timestamp 0
transform 1 0 2390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__513_
timestamp 0
transform -1 0 3170 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__514_
timestamp 0
transform 1 0 3410 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__515_
timestamp 0
transform -1 0 3730 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__516_
timestamp 0
transform 1 0 630 0 1 250
box -6 -8 26 248
use FILL  FILL_4__517_
timestamp 0
transform 1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_4__518_
timestamp 0
transform 1 0 1470 0 1 250
box -6 -8 26 248
use FILL  FILL_4__519_
timestamp 0
transform 1 0 1750 0 1 250
box -6 -8 26 248
use FILL  FILL_4__520_
timestamp 0
transform -1 0 1610 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__521_
timestamp 0
transform -1 0 1890 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__522_
timestamp 0
transform -1 0 3550 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__523_
timestamp 0
transform -1 0 3830 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__524_
timestamp 0
transform -1 0 1170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__525_
timestamp 0
transform 1 0 1190 0 1 250
box -6 -8 26 248
use FILL  FILL_4__526_
timestamp 0
transform -1 0 890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__527_
timestamp 0
transform -1 0 1030 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__528_
timestamp 0
transform 1 0 3090 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__529_
timestamp 0
transform 1 0 1270 0 1 730
box -6 -8 26 248
use FILL  FILL_4__530_
timestamp 0
transform 1 0 970 0 1 730
box -6 -8 26 248
use FILL  FILL_4__531_
timestamp 0
transform -1 0 510 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__532_
timestamp 0
transform 1 0 350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__533_
timestamp 0
transform -1 0 390 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__534_
timestamp 0
transform 1 0 650 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__535_
timestamp 0
transform -1 0 2410 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__536_
timestamp 0
transform -1 0 2690 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__537_
timestamp 0
transform -1 0 2970 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__538_
timestamp 0
transform -1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__539_
timestamp 0
transform -1 0 110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__540_
timestamp 0
transform -1 0 110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__541_
timestamp 0
transform 1 0 370 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__542_
timestamp 0
transform -1 0 410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__543_
timestamp 0
transform -1 0 3470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__544_
timestamp 0
transform -1 0 3730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__545_
timestamp 0
transform -1 0 3890 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__546_
timestamp 0
transform 1 0 3570 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__547_
timestamp 0
transform 1 0 2650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__548_
timestamp 0
transform -1 0 2230 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__549_
timestamp 0
transform -1 0 3550 0 1 250
box -6 -8 26 248
use FILL  FILL_4__550_
timestamp 0
transform -1 0 3830 0 1 250
box -6 -8 26 248
use FILL  FILL_4__551_
timestamp 0
transform 1 0 970 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__552_
timestamp 0
transform 1 0 670 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__553_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__554_
timestamp 0
transform 1 0 610 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__555_
timestamp 0
transform 1 0 390 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__556_
timestamp 0
transform -1 0 110 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__613_
timestamp 0
transform 1 0 4810 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__614_
timestamp 0
transform -1 0 4790 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__615_
timestamp 0
transform 1 0 4330 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__616_
timestamp 0
transform -1 0 4390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__617_
timestamp 0
transform 1 0 4530 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__618_
timestamp 0
transform 1 0 4850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__619_
timestamp 0
transform 1 0 4830 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__620_
timestamp 0
transform 1 0 4690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__621_
timestamp 0
transform 1 0 4830 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__622_
timestamp 0
transform 1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__623_
timestamp 0
transform 1 0 4610 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__624_
timestamp 0
transform 1 0 4650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__625_
timestamp 0
transform 1 0 3330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert7
timestamp 0
transform 1 0 4510 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert8
timestamp 0
transform -1 0 4430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert9
timestamp 0
transform 1 0 4550 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert10
timestamp 0
transform 1 0 4570 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert11
timestamp 0
transform -1 0 1250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert12
timestamp 0
transform 1 0 1810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform 1 0 1790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform 1 0 2450 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert15
timestamp 0
transform -1 0 630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert16
timestamp 0
transform 1 0 2830 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform 1 0 1890 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert18
timestamp 0
transform 1 0 2990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert19
timestamp 0
transform -1 0 990 0 1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert20
timestamp 0
transform 1 0 2910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert21
timestamp 0
transform 1 0 3970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert22
timestamp 0
transform -1 0 3210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert23
timestamp 0
transform -1 0 3470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert24
timestamp 0
transform -1 0 2910 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert25
timestamp 0
transform 1 0 2830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert0
timestamp 0
transform -1 0 3630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert1
timestamp 0
transform -1 0 110 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert2
timestamp 0
transform 1 0 90 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert3
timestamp 0
transform 1 0 2510 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert4
timestamp 0
transform 1 0 4150 0 -1 730
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert5
timestamp 0
transform -1 0 350 0 1 730
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert6
timestamp 0
transform 1 0 3650 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__273_
timestamp 0
transform -1 0 4370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__274_
timestamp 0
transform -1 0 4610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__275_
timestamp 0
transform -1 0 4890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__276_
timestamp 0
transform -1 0 3690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__277_
timestamp 0
transform 1 0 4910 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__278_
timestamp 0
transform 1 0 4870 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__279_
timestamp 0
transform 1 0 4510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__280_
timestamp 0
transform -1 0 4730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__281_
timestamp 0
transform -1 0 4790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__282_
timestamp 0
transform 1 0 3970 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__283_
timestamp 0
transform -1 0 3490 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__284_
timestamp 0
transform 1 0 3990 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__285_
timestamp 0
transform 1 0 3370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__286_
timestamp 0
transform -1 0 4610 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__287_
timestamp 0
transform 1 0 4570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__288_
timestamp 0
transform 1 0 3510 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__289_
timestamp 0
transform -1 0 4290 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__290_
timestamp 0
transform 1 0 4030 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__291_
timestamp 0
transform 1 0 1430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__292_
timestamp 0
transform -1 0 4030 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__293_
timestamp 0
transform -1 0 4290 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__294_
timestamp 0
transform 1 0 3870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__295_
timestamp 0
transform -1 0 4330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__296_
timestamp 0
transform 1 0 4610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__297_
timestamp 0
transform 1 0 4130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__298_
timestamp 0
transform -1 0 4050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__299_
timestamp 0
transform -1 0 4090 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__300_
timestamp 0
transform 1 0 3230 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__301_
timestamp 0
transform -1 0 3770 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__302_
timestamp 0
transform -1 0 3790 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__303_
timestamp 0
transform 1 0 3790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__304_
timestamp 0
transform -1 0 4050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__305_
timestamp 0
transform -1 0 4330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__306_
timestamp 0
transform 1 0 3870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__307_
timestamp 0
transform 1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__308_
timestamp 0
transform 1 0 4130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__309_
timestamp 0
transform -1 0 710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__310_
timestamp 0
transform -1 0 130 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__311_
timestamp 0
transform -1 0 130 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__312_
timestamp 0
transform -1 0 370 0 1 250
box -6 -8 26 248
use FILL  FILL_5__313_
timestamp 0
transform 1 0 350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__314_
timestamp 0
transform 1 0 350 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__315_
timestamp 0
transform 1 0 1530 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__316_
timestamp 0
transform -1 0 890 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__317_
timestamp 0
transform 1 0 590 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__318_
timestamp 0
transform -1 0 790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__319_
timestamp 0
transform -1 0 890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__320_
timestamp 0
transform -1 0 1430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__321_
timestamp 0
transform 1 0 1570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__322_
timestamp 0
transform 1 0 1430 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__323_
timestamp 0
transform -1 0 530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__324_
timestamp 0
transform 1 0 110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__325_
timestamp 0
transform 1 0 350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__326_
timestamp 0
transform -1 0 370 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__327_
timestamp 0
transform -1 0 130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__328_
timestamp 0
transform 1 0 650 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__329_
timestamp 0
transform 1 0 410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__330_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__331_
timestamp 0
transform 1 0 3390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__332_
timestamp 0
transform 1 0 3090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__333_
timestamp 0
transform 1 0 2310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__334_
timestamp 0
transform 1 0 2050 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__335_
timestamp 0
transform -1 0 2030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__336_
timestamp 0
transform -1 0 130 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__337_
timestamp 0
transform 1 0 110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__338_
timestamp 0
transform -1 0 390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__339_
timestamp 0
transform 1 0 3550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__340_
timestamp 0
transform -1 0 4070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__341_
timestamp 0
transform -1 0 4550 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__342_
timestamp 0
transform 1 0 4230 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__343_
timestamp 0
transform 1 0 3570 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__344_
timestamp 0
transform 1 0 3590 0 1 730
box -6 -8 26 248
use FILL  FILL_5__345_
timestamp 0
transform 1 0 4030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__346_
timestamp 0
transform 1 0 4110 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__347_
timestamp 0
transform -1 0 4890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__348_
timestamp 0
transform 1 0 4630 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__349_
timestamp 0
transform 1 0 2590 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__350_
timestamp 0
transform -1 0 3010 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__351_
timestamp 0
transform 1 0 2970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__352_
timestamp 0
transform -1 0 2750 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__353_
timestamp 0
transform 1 0 2370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__354_
timestamp 0
transform -1 0 3290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__355_
timestamp 0
transform -1 0 4130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__356_
timestamp 0
transform 1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__357_
timestamp 0
transform -1 0 2690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__358_
timestamp 0
transform -1 0 2870 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__359_
timestamp 0
transform 1 0 3130 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__360_
timestamp 0
transform -1 0 3430 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__361_
timestamp 0
transform -1 0 3210 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__362_
timestamp 0
transform -1 0 3150 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__363_
timestamp 0
transform 1 0 2330 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__364_
timestamp 0
transform 1 0 2190 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__365_
timestamp 0
transform 1 0 3170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__366_
timestamp 0
transform 1 0 2850 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__367_
timestamp 0
transform -1 0 2110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__368_
timestamp 0
transform 1 0 2870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__369_
timestamp 0
transform -1 0 3310 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__370_
timestamp 0
transform 1 0 4910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__371_
timestamp 0
transform 1 0 4610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__372_
timestamp 0
transform 1 0 3290 0 1 250
box -6 -8 26 248
use FILL  FILL_5__373_
timestamp 0
transform 1 0 3290 0 1 730
box -6 -8 26 248
use FILL  FILL_5__374_
timestamp 0
transform 1 0 4110 0 1 730
box -6 -8 26 248
use FILL  FILL_5__375_
timestamp 0
transform 1 0 3830 0 1 730
box -6 -8 26 248
use FILL  FILL_5__376_
timestamp 0
transform 1 0 4390 0 1 730
box -6 -8 26 248
use FILL  FILL_5__377_
timestamp 0
transform -1 0 4090 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__378_
timestamp 0
transform -1 0 4210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__379_
timestamp 0
transform -1 0 2310 0 1 250
box -6 -8 26 248
use FILL  FILL_5__380_
timestamp 0
transform 1 0 1630 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__381_
timestamp 0
transform 1 0 1330 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__382_
timestamp 0
transform -1 0 1010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__383_
timestamp 0
transform 1 0 1470 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__384_
timestamp 0
transform -1 0 930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__385_
timestamp 0
transform -1 0 970 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__386_
timestamp 0
transform 1 0 1030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__387_
timestamp 0
transform -1 0 850 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__388_
timestamp 0
transform -1 0 3950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__389_
timestamp 0
transform -1 0 1550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__390_
timestamp 0
transform -1 0 1250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__391_
timestamp 0
transform 1 0 930 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__392_
timestamp 0
transform -1 0 730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__393_
timestamp 0
transform 1 0 1190 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__394_
timestamp 0
transform 1 0 1750 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__395_
timestamp 0
transform -1 0 3710 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__396_
timestamp 0
transform 1 0 1190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__397_
timestamp 0
transform 1 0 1450 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__398_
timestamp 0
transform 1 0 1990 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__399_
timestamp 0
transform 1 0 1990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__400_
timestamp 0
transform 1 0 1730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__401_
timestamp 0
transform 1 0 1450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__402_
timestamp 0
transform 1 0 1770 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__403_
timestamp 0
transform -1 0 2850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__404_
timestamp 0
transform 1 0 2550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__405_
timestamp 0
transform -1 0 1330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__406_
timestamp 0
transform 1 0 1210 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__407_
timestamp 0
transform -1 0 1490 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__408_
timestamp 0
transform -1 0 970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__409_
timestamp 0
transform 1 0 1230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__410_
timestamp 0
transform -1 0 1150 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__411_
timestamp 0
transform -1 0 3230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__412_
timestamp 0
transform -1 0 1730 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__413_
timestamp 0
transform 1 0 1570 0 1 730
box -6 -8 26 248
use FILL  FILL_5__414_
timestamp 0
transform 1 0 1850 0 1 730
box -6 -8 26 248
use FILL  FILL_5__415_
timestamp 0
transform 1 0 2710 0 1 730
box -6 -8 26 248
use FILL  FILL_5__416_
timestamp 0
transform -1 0 2070 0 1 250
box -6 -8 26 248
use FILL  FILL_5__417_
timestamp 0
transform 1 0 2430 0 1 730
box -6 -8 26 248
use FILL  FILL_5__418_
timestamp 0
transform 1 0 2270 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__419_
timestamp 0
transform -1 0 3030 0 1 730
box -6 -8 26 248
use FILL  FILL_5__420_
timestamp 0
transform -1 0 2930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__421_
timestamp 0
transform 1 0 4590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__422_
timestamp 0
transform 1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__423_
timestamp 0
transform 1 0 4910 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__424_
timestamp 0
transform 1 0 4910 0 1 250
box -6 -8 26 248
use FILL  FILL_5__425_
timestamp 0
transform 1 0 4370 0 1 250
box -6 -8 26 248
use FILL  FILL_5__426_
timestamp 0
transform -1 0 4650 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__427_
timestamp 0
transform -1 0 2590 0 1 250
box -6 -8 26 248
use FILL  FILL_5__428_
timestamp 0
transform 1 0 2150 0 1 730
box -6 -8 26 248
use FILL  FILL_5__429_
timestamp 0
transform 1 0 2550 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__430_
timestamp 0
transform -1 0 1430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__431_
timestamp 0
transform 1 0 1710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__432_
timestamp 0
transform -1 0 2310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__433_
timestamp 0
transform 1 0 2570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__434_
timestamp 0
transform -1 0 4350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__435_
timestamp 0
transform 1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__436_
timestamp 0
transform -1 0 3770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__437_
timestamp 0
transform -1 0 2310 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__438_
timestamp 0
transform -1 0 2570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5__439_
timestamp 0
transform 1 0 2590 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__440_
timestamp 0
transform -1 0 3150 0 1 2170
box -6 -8 26 248
use FILL  FILL_5__441_
timestamp 0
transform 1 0 1530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__442_
timestamp 0
transform -1 0 2110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__443_
timestamp 0
transform -1 0 1730 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__444_
timestamp 0
transform -1 0 2170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__445_
timestamp 0
transform -1 0 1870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__446_
timestamp 0
transform 1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__447_
timestamp 0
transform -1 0 4250 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__448_
timestamp 0
transform -1 0 1810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__449_
timestamp 0
transform 1 0 2290 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__450_
timestamp 0
transform 1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5__451_
timestamp 0
transform 1 0 2550 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__452_
timestamp 0
transform -1 0 3690 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__453_
timestamp 0
transform 1 0 1450 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__454_
timestamp 0
transform -1 0 1690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__455_
timestamp 0
transform 1 0 2030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__456_
timestamp 0
transform -1 0 1970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__457_
timestamp 0
transform 1 0 1710 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__458_
timestamp 0
transform 1 0 1790 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__459_
timestamp 0
transform 1 0 2250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__460_
timestamp 0
transform -1 0 2570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__461_
timestamp 0
transform -1 0 2110 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__462_
timestamp 0
transform 1 0 2370 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__463_
timestamp 0
transform 1 0 2670 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__464_
timestamp 0
transform -1 0 2990 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__465_
timestamp 0
transform 1 0 1250 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__466_
timestamp 0
transform -1 0 970 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__467_
timestamp 0
transform 1 0 650 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__468_
timestamp 0
transform -1 0 410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__469_
timestamp 0
transform -1 0 390 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__470_
timestamp 0
transform -1 0 690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__471_
timestamp 0
transform 1 0 690 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__472_
timestamp 0
transform -1 0 930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__473_
timestamp 0
transform 1 0 870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__474_
timestamp 0
transform 1 0 950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__475_
timestamp 0
transform -1 0 130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__476_
timestamp 0
transform -1 0 130 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__477_
timestamp 0
transform 1 0 370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__478_
timestamp 0
transform -1 0 410 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__479_
timestamp 0
transform -1 0 3510 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__480_
timestamp 0
transform -1 0 1290 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__481_
timestamp 0
transform -1 0 130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__482_
timestamp 0
transform -1 0 1250 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__483_
timestamp 0
transform -1 0 1530 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__484_
timestamp 0
transform 1 0 1690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__485_
timestamp 0
transform 1 0 1990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__486_
timestamp 0
transform 1 0 2270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__487_
timestamp 0
transform 1 0 2850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__488_
timestamp 0
transform 1 0 2550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__489_
timestamp 0
transform 1 0 1530 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__490_
timestamp 0
transform -1 0 1810 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__491_
timestamp 0
transform 1 0 2090 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__492_
timestamp 0
transform 1 0 2370 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__493_
timestamp 0
transform -1 0 2690 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__494_
timestamp 0
transform 1 0 1170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__495_
timestamp 0
transform 1 0 1450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__496_
timestamp 0
transform 1 0 1730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__497_
timestamp 0
transform 1 0 2110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__498_
timestamp 0
transform -1 0 2330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__499_
timestamp 0
transform -1 0 1810 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__500_
timestamp 0
transform -1 0 2350 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__501_
timestamp 0
transform -1 0 2730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__502_
timestamp 0
transform -1 0 3290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__503_
timestamp 0
transform -1 0 3370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__504_
timestamp 0
transform 1 0 4570 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__505_
timestamp 0
transform -1 0 4850 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__506_
timestamp 0
transform 1 0 4650 0 1 250
box -6 -8 26 248
use FILL  FILL_5__507_
timestamp 0
transform -1 0 4690 0 1 730
box -6 -8 26 248
use FILL  FILL_5__508_
timestamp 0
transform -1 0 2930 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__509_
timestamp 0
transform 1 0 2070 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__510_
timestamp 0
transform -1 0 2630 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__511_
timestamp 0
transform 1 0 1530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__512_
timestamp 0
transform 1 0 2410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__513_
timestamp 0
transform -1 0 3190 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__514_
timestamp 0
transform 1 0 3430 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__515_
timestamp 0
transform -1 0 3750 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__516_
timestamp 0
transform 1 0 650 0 1 250
box -6 -8 26 248
use FILL  FILL_5__517_
timestamp 0
transform 1 0 930 0 1 250
box -6 -8 26 248
use FILL  FILL_5__518_
timestamp 0
transform 1 0 1490 0 1 250
box -6 -8 26 248
use FILL  FILL_5__519_
timestamp 0
transform 1 0 1770 0 1 250
box -6 -8 26 248
use FILL  FILL_5__520_
timestamp 0
transform -1 0 1630 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__521_
timestamp 0
transform -1 0 1910 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__522_
timestamp 0
transform -1 0 3570 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__523_
timestamp 0
transform -1 0 3850 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__524_
timestamp 0
transform -1 0 1190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__525_
timestamp 0
transform 1 0 1210 0 1 250
box -6 -8 26 248
use FILL  FILL_5__526_
timestamp 0
transform -1 0 910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__527_
timestamp 0
transform -1 0 1050 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__528_
timestamp 0
transform 1 0 3110 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__529_
timestamp 0
transform 1 0 1290 0 1 730
box -6 -8 26 248
use FILL  FILL_5__530_
timestamp 0
transform 1 0 990 0 1 730
box -6 -8 26 248
use FILL  FILL_5__531_
timestamp 0
transform -1 0 530 0 1 1210
box -6 -8 26 248
use FILL  FILL_5__532_
timestamp 0
transform 1 0 370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__533_
timestamp 0
transform -1 0 410 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__534_
timestamp 0
transform 1 0 670 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__535_
timestamp 0
transform -1 0 2430 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__536_
timestamp 0
transform -1 0 2710 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__537_
timestamp 0
transform -1 0 2990 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__538_
timestamp 0
transform -1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_5__539_
timestamp 0
transform -1 0 130 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__540_
timestamp 0
transform -1 0 130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__541_
timestamp 0
transform 1 0 390 0 1 1690
box -6 -8 26 248
use FILL  FILL_5__542_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5__543_
timestamp 0
transform -1 0 3490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__544_
timestamp 0
transform -1 0 3750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_5__545_
timestamp 0
transform -1 0 3910 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__546_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 26 248
use FILL  FILL_5__547_
timestamp 0
transform 1 0 2670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5__548_
timestamp 0
transform -1 0 2250 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__549_
timestamp 0
transform -1 0 3570 0 1 250
box -6 -8 26 248
use FILL  FILL_5__550_
timestamp 0
transform -1 0 3850 0 1 250
box -6 -8 26 248
use FILL  FILL_5__551_
timestamp 0
transform 1 0 990 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__552_
timestamp 0
transform 1 0 690 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__553_
timestamp 0
transform -1 0 930 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__554_
timestamp 0
transform 1 0 630 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__555_
timestamp 0
transform 1 0 410 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__556_
timestamp 0
transform -1 0 130 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__613_
timestamp 0
transform 1 0 4830 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__614_
timestamp 0
transform -1 0 4810 0 1 2650
box -6 -8 26 248
use FILL  FILL_5__615_
timestamp 0
transform 1 0 4350 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__616_
timestamp 0
transform -1 0 4410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__617_
timestamp 0
transform 1 0 4550 0 1 3130
box -6 -8 26 248
use FILL  FILL_5__618_
timestamp 0
transform 1 0 4870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5__619_
timestamp 0
transform 1 0 4850 0 1 3610
box -6 -8 26 248
use FILL  FILL_5__620_
timestamp 0
transform 1 0 4710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5__621_
timestamp 0
transform 1 0 4850 0 1 4090
box -6 -8 26 248
use FILL  FILL_5__622_
timestamp 0
transform 1 0 4910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5__623_
timestamp 0
transform 1 0 4630 0 1 4570
box -6 -8 26 248
use FILL  FILL_5__624_
timestamp 0
transform 1 0 4670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5__625_
timestamp 0
transform 1 0 3350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert7
timestamp 0
transform 1 0 4530 0 1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert8
timestamp 0
transform -1 0 4450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert9
timestamp 0
transform 1 0 4570 0 1 4090
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert10
timestamp 0
transform 1 0 4590 0 1 3610
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert11
timestamp 0
transform -1 0 1270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert12
timestamp 0
transform 1 0 1830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert13
timestamp 0
transform 1 0 1810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert14
timestamp 0
transform 1 0 2470 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert15
timestamp 0
transform -1 0 650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert16
timestamp 0
transform 1 0 2850 0 1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert17
timestamp 0
transform 1 0 1910 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert18
timestamp 0
transform 1 0 3010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert19
timestamp 0
transform -1 0 1010 0 1 4570
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert20
timestamp 0
transform 1 0 2930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert21
timestamp 0
transform 1 0 3990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert22
timestamp 0
transform -1 0 3230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert23
timestamp 0
transform -1 0 3490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert24
timestamp 0
transform -1 0 2930 0 1 3130
box -6 -8 26 248
use FILL  FILL_5_BUFX2_insert25
timestamp 0
transform 1 0 2850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert0
timestamp 0
transform -1 0 3650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert1
timestamp 0
transform -1 0 130 0 1 1210
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert2
timestamp 0
transform 1 0 110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert3
timestamp 0
transform 1 0 2530 0 1 3130
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert4
timestamp 0
transform 1 0 4170 0 -1 730
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert5
timestamp 0
transform -1 0 370 0 1 730
box -6 -8 26 248
use FILL  FILL_5_CLKBUF1_insert6
timestamp 0
transform 1 0 3670 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__273_
timestamp 0
transform -1 0 4390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__274_
timestamp 0
transform -1 0 4630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__275_
timestamp 0
transform -1 0 4910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__276_
timestamp 0
transform -1 0 3710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__277_
timestamp 0
transform 1 0 4930 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__278_
timestamp 0
transform 1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__279_
timestamp 0
transform 1 0 4530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__280_
timestamp 0
transform -1 0 4750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__281_
timestamp 0
transform -1 0 4810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__282_
timestamp 0
transform 1 0 3990 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__283_
timestamp 0
transform -1 0 3510 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__284_
timestamp 0
transform 1 0 4010 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__285_
timestamp 0
transform 1 0 3390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__286_
timestamp 0
transform -1 0 4630 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__287_
timestamp 0
transform 1 0 4590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__288_
timestamp 0
transform 1 0 3530 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__289_
timestamp 0
transform -1 0 4310 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__290_
timestamp 0
transform 1 0 4050 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__291_
timestamp 0
transform 1 0 1450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__292_
timestamp 0
transform -1 0 4050 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__293_
timestamp 0
transform -1 0 4310 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__294_
timestamp 0
transform 1 0 3890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__295_
timestamp 0
transform -1 0 4350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__296_
timestamp 0
transform 1 0 4630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__297_
timestamp 0
transform 1 0 4150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__298_
timestamp 0
transform -1 0 4070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__299_
timestamp 0
transform -1 0 4110 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__300_
timestamp 0
transform 1 0 3250 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__301_
timestamp 0
transform -1 0 3790 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__302_
timestamp 0
transform -1 0 3810 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__303_
timestamp 0
transform 1 0 3810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__304_
timestamp 0
transform -1 0 4070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__305_
timestamp 0
transform -1 0 4350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__306_
timestamp 0
transform 1 0 3890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__307_
timestamp 0
transform 1 0 4350 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__308_
timestamp 0
transform 1 0 4150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__309_
timestamp 0
transform -1 0 730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__310_
timestamp 0
transform -1 0 150 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__311_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__312_
timestamp 0
transform -1 0 390 0 1 250
box -6 -8 26 248
use FILL  FILL_6__313_
timestamp 0
transform 1 0 370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__314_
timestamp 0
transform 1 0 370 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__315_
timestamp 0
transform 1 0 1550 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__316_
timestamp 0
transform -1 0 910 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__317_
timestamp 0
transform 1 0 610 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__318_
timestamp 0
transform -1 0 810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__319_
timestamp 0
transform -1 0 910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__320_
timestamp 0
transform -1 0 1450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__321_
timestamp 0
transform 1 0 1590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__322_
timestamp 0
transform 1 0 1450 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__323_
timestamp 0
transform -1 0 550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__324_
timestamp 0
transform 1 0 130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__325_
timestamp 0
transform 1 0 370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__326_
timestamp 0
transform -1 0 390 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__327_
timestamp 0
transform -1 0 150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__328_
timestamp 0
transform 1 0 670 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__329_
timestamp 0
transform 1 0 430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__330_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__331_
timestamp 0
transform 1 0 3410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__332_
timestamp 0
transform 1 0 3110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__333_
timestamp 0
transform 1 0 2330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__334_
timestamp 0
transform 1 0 2070 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__335_
timestamp 0
transform -1 0 2050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__336_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__337_
timestamp 0
transform 1 0 130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__338_
timestamp 0
transform -1 0 410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__339_
timestamp 0
transform 1 0 3570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__340_
timestamp 0
transform -1 0 4090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__341_
timestamp 0
transform -1 0 4570 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__342_
timestamp 0
transform 1 0 4250 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__343_
timestamp 0
transform 1 0 3590 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__344_
timestamp 0
transform 1 0 3610 0 1 730
box -6 -8 26 248
use FILL  FILL_6__345_
timestamp 0
transform 1 0 4050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__346_
timestamp 0
transform 1 0 4130 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__347_
timestamp 0
transform -1 0 4910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__348_
timestamp 0
transform 1 0 4650 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__349_
timestamp 0
transform 1 0 2610 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__350_
timestamp 0
transform -1 0 3030 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__351_
timestamp 0
transform 1 0 2990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__352_
timestamp 0
transform -1 0 2770 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__353_
timestamp 0
transform 1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__354_
timestamp 0
transform -1 0 3310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__355_
timestamp 0
transform -1 0 4150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__356_
timestamp 0
transform 1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__357_
timestamp 0
transform -1 0 2710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__358_
timestamp 0
transform -1 0 2890 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__359_
timestamp 0
transform 1 0 3150 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__360_
timestamp 0
transform -1 0 3450 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__361_
timestamp 0
transform -1 0 3230 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__362_
timestamp 0
transform -1 0 3170 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__363_
timestamp 0
transform 1 0 2350 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__364_
timestamp 0
transform 1 0 2210 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__365_
timestamp 0
transform 1 0 3190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__366_
timestamp 0
transform 1 0 2870 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__367_
timestamp 0
transform -1 0 2130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__368_
timestamp 0
transform 1 0 2890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__369_
timestamp 0
transform -1 0 3330 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__370_
timestamp 0
transform 1 0 4930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__371_
timestamp 0
transform 1 0 4630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__372_
timestamp 0
transform 1 0 3310 0 1 250
box -6 -8 26 248
use FILL  FILL_6__373_
timestamp 0
transform 1 0 3310 0 1 730
box -6 -8 26 248
use FILL  FILL_6__374_
timestamp 0
transform 1 0 4130 0 1 730
box -6 -8 26 248
use FILL  FILL_6__375_
timestamp 0
transform 1 0 3850 0 1 730
box -6 -8 26 248
use FILL  FILL_6__376_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 26 248
use FILL  FILL_6__377_
timestamp 0
transform -1 0 4110 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__378_
timestamp 0
transform -1 0 4230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__379_
timestamp 0
transform -1 0 2330 0 1 250
box -6 -8 26 248
use FILL  FILL_6__380_
timestamp 0
transform 1 0 1650 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__381_
timestamp 0
transform 1 0 1350 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__382_
timestamp 0
transform -1 0 1030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__383_
timestamp 0
transform 1 0 1490 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__384_
timestamp 0
transform -1 0 950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__385_
timestamp 0
transform -1 0 990 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__386_
timestamp 0
transform 1 0 1050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__387_
timestamp 0
transform -1 0 870 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__388_
timestamp 0
transform -1 0 3970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__389_
timestamp 0
transform -1 0 1570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__390_
timestamp 0
transform -1 0 1270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__391_
timestamp 0
transform 1 0 950 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__392_
timestamp 0
transform -1 0 750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__393_
timestamp 0
transform 1 0 1210 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__394_
timestamp 0
transform 1 0 1770 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__395_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__396_
timestamp 0
transform 1 0 1210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__397_
timestamp 0
transform 1 0 1470 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__398_
timestamp 0
transform 1 0 2010 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__399_
timestamp 0
transform 1 0 2010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__400_
timestamp 0
transform 1 0 1750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__401_
timestamp 0
transform 1 0 1470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__402_
timestamp 0
transform 1 0 1790 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__403_
timestamp 0
transform -1 0 2870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__404_
timestamp 0
transform 1 0 2570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__405_
timestamp 0
transform -1 0 1350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__406_
timestamp 0
transform 1 0 1230 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__407_
timestamp 0
transform -1 0 1510 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__408_
timestamp 0
transform -1 0 990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__409_
timestamp 0
transform 1 0 1250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__410_
timestamp 0
transform -1 0 1170 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__411_
timestamp 0
transform -1 0 3250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__412_
timestamp 0
transform -1 0 1750 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__413_
timestamp 0
transform 1 0 1590 0 1 730
box -6 -8 26 248
use FILL  FILL_6__414_
timestamp 0
transform 1 0 1870 0 1 730
box -6 -8 26 248
use FILL  FILL_6__415_
timestamp 0
transform 1 0 2730 0 1 730
box -6 -8 26 248
use FILL  FILL_6__416_
timestamp 0
transform -1 0 2090 0 1 250
box -6 -8 26 248
use FILL  FILL_6__417_
timestamp 0
transform 1 0 2450 0 1 730
box -6 -8 26 248
use FILL  FILL_6__418_
timestamp 0
transform 1 0 2290 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__419_
timestamp 0
transform -1 0 3050 0 1 730
box -6 -8 26 248
use FILL  FILL_6__420_
timestamp 0
transform -1 0 2950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__421_
timestamp 0
transform 1 0 4610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__422_
timestamp 0
transform 1 0 4390 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__423_
timestamp 0
transform 1 0 4930 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__424_
timestamp 0
transform 1 0 4930 0 1 250
box -6 -8 26 248
use FILL  FILL_6__425_
timestamp 0
transform 1 0 4390 0 1 250
box -6 -8 26 248
use FILL  FILL_6__426_
timestamp 0
transform -1 0 4670 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__427_
timestamp 0
transform -1 0 2610 0 1 250
box -6 -8 26 248
use FILL  FILL_6__428_
timestamp 0
transform 1 0 2170 0 1 730
box -6 -8 26 248
use FILL  FILL_6__429_
timestamp 0
transform 1 0 2570 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__430_
timestamp 0
transform -1 0 1450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__431_
timestamp 0
transform 1 0 1730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__432_
timestamp 0
transform -1 0 2330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__433_
timestamp 0
transform 1 0 2590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__434_
timestamp 0
transform -1 0 4370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__435_
timestamp 0
transform 1 0 3490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__436_
timestamp 0
transform -1 0 3790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__437_
timestamp 0
transform -1 0 2330 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__438_
timestamp 0
transform -1 0 2590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6__439_
timestamp 0
transform 1 0 2610 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__440_
timestamp 0
transform -1 0 3170 0 1 2170
box -6 -8 26 248
use FILL  FILL_6__441_
timestamp 0
transform 1 0 1550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__442_
timestamp 0
transform -1 0 2130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__443_
timestamp 0
transform -1 0 1750 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__444_
timestamp 0
transform -1 0 2190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__445_
timestamp 0
transform -1 0 1890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__446_
timestamp 0
transform 1 0 2030 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__447_
timestamp 0
transform -1 0 4270 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__448_
timestamp 0
transform -1 0 1830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__449_
timestamp 0
transform 1 0 2310 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__450_
timestamp 0
transform 1 0 2390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6__451_
timestamp 0
transform 1 0 2570 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__452_
timestamp 0
transform -1 0 3710 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__453_
timestamp 0
transform 1 0 1470 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__454_
timestamp 0
transform -1 0 1710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__455_
timestamp 0
transform 1 0 2050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__456_
timestamp 0
transform -1 0 1990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__457_
timestamp 0
transform 1 0 1730 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__458_
timestamp 0
transform 1 0 1810 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__459_
timestamp 0
transform 1 0 2270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__460_
timestamp 0
transform -1 0 2590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__461_
timestamp 0
transform -1 0 2130 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__462_
timestamp 0
transform 1 0 2390 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__463_
timestamp 0
transform 1 0 2690 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__464_
timestamp 0
transform -1 0 3010 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__465_
timestamp 0
transform 1 0 1270 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__466_
timestamp 0
transform -1 0 990 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__467_
timestamp 0
transform 1 0 670 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__468_
timestamp 0
transform -1 0 430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__469_
timestamp 0
transform -1 0 410 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__470_
timestamp 0
transform -1 0 710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__471_
timestamp 0
transform 1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__472_
timestamp 0
transform -1 0 950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__473_
timestamp 0
transform 1 0 890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__474_
timestamp 0
transform 1 0 970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__475_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__476_
timestamp 0
transform -1 0 150 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__477_
timestamp 0
transform 1 0 390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__478_
timestamp 0
transform -1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__479_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__480_
timestamp 0
transform -1 0 1310 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__481_
timestamp 0
transform -1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__482_
timestamp 0
transform -1 0 1270 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__483_
timestamp 0
transform -1 0 1550 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__484_
timestamp 0
transform 1 0 1710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__485_
timestamp 0
transform 1 0 2010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__486_
timestamp 0
transform 1 0 2290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__487_
timestamp 0
transform 1 0 2870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__488_
timestamp 0
transform 1 0 2570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__489_
timestamp 0
transform 1 0 1550 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__490_
timestamp 0
transform -1 0 1830 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__491_
timestamp 0
transform 1 0 2110 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__492_
timestamp 0
transform 1 0 2390 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__493_
timestamp 0
transform -1 0 2710 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__494_
timestamp 0
transform 1 0 1190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__495_
timestamp 0
transform 1 0 1470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__496_
timestamp 0
transform 1 0 1750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__497_
timestamp 0
transform 1 0 2130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__498_
timestamp 0
transform -1 0 2350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__499_
timestamp 0
transform -1 0 1830 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__500_
timestamp 0
transform -1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__501_
timestamp 0
transform -1 0 2750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__502_
timestamp 0
transform -1 0 3310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__503_
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__504_
timestamp 0
transform 1 0 4590 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__505_
timestamp 0
transform -1 0 4870 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__506_
timestamp 0
transform 1 0 4670 0 1 250
box -6 -8 26 248
use FILL  FILL_6__507_
timestamp 0
transform -1 0 4710 0 1 730
box -6 -8 26 248
use FILL  FILL_6__508_
timestamp 0
transform -1 0 2950 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__509_
timestamp 0
transform 1 0 2090 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__510_
timestamp 0
transform -1 0 2650 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__511_
timestamp 0
transform 1 0 1550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__512_
timestamp 0
transform 1 0 2430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__513_
timestamp 0
transform -1 0 3210 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__514_
timestamp 0
transform 1 0 3450 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__515_
timestamp 0
transform -1 0 3770 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__516_
timestamp 0
transform 1 0 670 0 1 250
box -6 -8 26 248
use FILL  FILL_6__517_
timestamp 0
transform 1 0 950 0 1 250
box -6 -8 26 248
use FILL  FILL_6__518_
timestamp 0
transform 1 0 1510 0 1 250
box -6 -8 26 248
use FILL  FILL_6__519_
timestamp 0
transform 1 0 1790 0 1 250
box -6 -8 26 248
use FILL  FILL_6__520_
timestamp 0
transform -1 0 1650 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__521_
timestamp 0
transform -1 0 1930 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__522_
timestamp 0
transform -1 0 3590 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__523_
timestamp 0
transform -1 0 3870 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__524_
timestamp 0
transform -1 0 1210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__525_
timestamp 0
transform 1 0 1230 0 1 250
box -6 -8 26 248
use FILL  FILL_6__526_
timestamp 0
transform -1 0 930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__527_
timestamp 0
transform -1 0 1070 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__528_
timestamp 0
transform 1 0 3130 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__529_
timestamp 0
transform 1 0 1310 0 1 730
box -6 -8 26 248
use FILL  FILL_6__530_
timestamp 0
transform 1 0 1010 0 1 730
box -6 -8 26 248
use FILL  FILL_6__531_
timestamp 0
transform -1 0 550 0 1 1210
box -6 -8 26 248
use FILL  FILL_6__532_
timestamp 0
transform 1 0 390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__533_
timestamp 0
transform -1 0 430 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__534_
timestamp 0
transform 1 0 690 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__535_
timestamp 0
transform -1 0 2450 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__536_
timestamp 0
transform -1 0 2730 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__537_
timestamp 0
transform -1 0 3010 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__538_
timestamp 0
transform -1 0 3290 0 -1 250
box -6 -8 26 248
use FILL  FILL_6__539_
timestamp 0
transform -1 0 150 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__540_
timestamp 0
transform -1 0 150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__541_
timestamp 0
transform 1 0 410 0 1 1690
box -6 -8 26 248
use FILL  FILL_6__542_
timestamp 0
transform -1 0 450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6__543_
timestamp 0
transform -1 0 3510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__544_
timestamp 0
transform -1 0 3770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_6__545_
timestamp 0
transform -1 0 3930 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__546_
timestamp 0
transform 1 0 3610 0 -1 730
box -6 -8 26 248
use FILL  FILL_6__547_
timestamp 0
transform 1 0 2690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6__548_
timestamp 0
transform -1 0 2270 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__549_
timestamp 0
transform -1 0 3590 0 1 250
box -6 -8 26 248
use FILL  FILL_6__550_
timestamp 0
transform -1 0 3870 0 1 250
box -6 -8 26 248
use FILL  FILL_6__551_
timestamp 0
transform 1 0 1010 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__552_
timestamp 0
transform 1 0 710 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__553_
timestamp 0
transform -1 0 950 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__554_
timestamp 0
transform 1 0 650 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__555_
timestamp 0
transform 1 0 430 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__556_
timestamp 0
transform -1 0 150 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__613_
timestamp 0
transform 1 0 4850 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__614_
timestamp 0
transform -1 0 4830 0 1 2650
box -6 -8 26 248
use FILL  FILL_6__615_
timestamp 0
transform 1 0 4370 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__616_
timestamp 0
transform -1 0 4430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__617_
timestamp 0
transform 1 0 4570 0 1 3130
box -6 -8 26 248
use FILL  FILL_6__618_
timestamp 0
transform 1 0 4890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6__619_
timestamp 0
transform 1 0 4870 0 1 3610
box -6 -8 26 248
use FILL  FILL_6__620_
timestamp 0
transform 1 0 4730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6__621_
timestamp 0
transform 1 0 4870 0 1 4090
box -6 -8 26 248
use FILL  FILL_6__622_
timestamp 0
transform 1 0 4930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6__623_
timestamp 0
transform 1 0 4650 0 1 4570
box -6 -8 26 248
use FILL  FILL_6__624_
timestamp 0
transform 1 0 4690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6__625_
timestamp 0
transform 1 0 3370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert7
timestamp 0
transform 1 0 4550 0 1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert8
timestamp 0
transform -1 0 4470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert9
timestamp 0
transform 1 0 4590 0 1 4090
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert10
timestamp 0
transform 1 0 4610 0 1 3610
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert11
timestamp 0
transform -1 0 1290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert12
timestamp 0
transform 1 0 1850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert13
timestamp 0
transform 1 0 1830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert14
timestamp 0
transform 1 0 2490 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert15
timestamp 0
transform -1 0 670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert16
timestamp 0
transform 1 0 2870 0 1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert17
timestamp 0
transform 1 0 1930 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert18
timestamp 0
transform 1 0 3030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert19
timestamp 0
transform -1 0 1030 0 1 4570
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert20
timestamp 0
transform 1 0 2950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert21
timestamp 0
transform 1 0 4010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert22
timestamp 0
transform -1 0 3250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert23
timestamp 0
transform -1 0 3510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert24
timestamp 0
transform -1 0 2950 0 1 3130
box -6 -8 26 248
use FILL  FILL_6_BUFX2_insert25
timestamp 0
transform 1 0 2870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert0
timestamp 0
transform -1 0 3670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert1
timestamp 0
transform -1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert2
timestamp 0
transform 1 0 130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert3
timestamp 0
transform 1 0 2550 0 1 3130
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert4
timestamp 0
transform 1 0 4190 0 -1 730
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert5
timestamp 0
transform -1 0 390 0 1 730
box -6 -8 26 248
use FILL  FILL_6_CLKBUF1_insert6
timestamp 0
transform 1 0 3690 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__273_
timestamp 0
transform -1 0 4410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__274_
timestamp 0
transform -1 0 4650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__275_
timestamp 0
transform -1 0 4930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__276_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__277_
timestamp 0
transform 1 0 4950 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__278_
timestamp 0
transform 1 0 4910 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__279_
timestamp 0
transform 1 0 4550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__280_
timestamp 0
transform -1 0 4770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__281_
timestamp 0
transform -1 0 4830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__282_
timestamp 0
transform 1 0 4010 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__283_
timestamp 0
transform -1 0 3530 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__284_
timestamp 0
transform 1 0 4030 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__285_
timestamp 0
transform 1 0 3410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__286_
timestamp 0
transform -1 0 4650 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__287_
timestamp 0
transform 1 0 4610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__288_
timestamp 0
transform 1 0 3550 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__289_
timestamp 0
transform -1 0 4330 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__290_
timestamp 0
transform 1 0 4070 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__291_
timestamp 0
transform 1 0 1470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__292_
timestamp 0
transform -1 0 4070 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__293_
timestamp 0
transform -1 0 4330 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__294_
timestamp 0
transform 1 0 3910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__295_
timestamp 0
transform -1 0 4370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__296_
timestamp 0
transform 1 0 4650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__297_
timestamp 0
transform 1 0 4170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__298_
timestamp 0
transform -1 0 4090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__299_
timestamp 0
transform -1 0 4130 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__300_
timestamp 0
transform 1 0 3270 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__301_
timestamp 0
transform -1 0 3810 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__302_
timestamp 0
transform -1 0 3830 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__303_
timestamp 0
transform 1 0 3830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__304_
timestamp 0
transform -1 0 4090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__305_
timestamp 0
transform -1 0 4370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__306_
timestamp 0
transform 1 0 3910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__307_
timestamp 0
transform 1 0 4370 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__308_
timestamp 0
transform 1 0 4170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__309_
timestamp 0
transform -1 0 750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__310_
timestamp 0
transform -1 0 170 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__311_
timestamp 0
transform -1 0 170 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__312_
timestamp 0
transform -1 0 410 0 1 250
box -6 -8 26 248
use FILL  FILL_7__313_
timestamp 0
transform 1 0 390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__314_
timestamp 0
transform 1 0 390 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__315_
timestamp 0
transform 1 0 1570 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__316_
timestamp 0
transform -1 0 930 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__317_
timestamp 0
transform 1 0 630 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__318_
timestamp 0
transform -1 0 830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__319_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__320_
timestamp 0
transform -1 0 1470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__321_
timestamp 0
transform 1 0 1610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__322_
timestamp 0
transform 1 0 1470 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__323_
timestamp 0
transform -1 0 570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__324_
timestamp 0
transform 1 0 150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__325_
timestamp 0
transform 1 0 390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__326_
timestamp 0
transform -1 0 410 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__327_
timestamp 0
transform -1 0 170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__328_
timestamp 0
transform 1 0 690 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__329_
timestamp 0
transform 1 0 450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__330_
timestamp 0
transform 1 0 2870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__331_
timestamp 0
transform 1 0 3430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__332_
timestamp 0
transform 1 0 3130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__333_
timestamp 0
transform 1 0 2350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__334_
timestamp 0
transform 1 0 2090 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__335_
timestamp 0
transform -1 0 2070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__336_
timestamp 0
transform -1 0 170 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__337_
timestamp 0
transform 1 0 150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__338_
timestamp 0
transform -1 0 430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__339_
timestamp 0
transform 1 0 3590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__340_
timestamp 0
transform -1 0 4110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__341_
timestamp 0
transform -1 0 4590 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__342_
timestamp 0
transform 1 0 4270 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__343_
timestamp 0
transform 1 0 3610 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__344_
timestamp 0
transform 1 0 3630 0 1 730
box -6 -8 26 248
use FILL  FILL_7__345_
timestamp 0
transform 1 0 4070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__346_
timestamp 0
transform 1 0 4150 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__347_
timestamp 0
transform -1 0 4930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__348_
timestamp 0
transform 1 0 4670 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__349_
timestamp 0
transform 1 0 2630 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__350_
timestamp 0
transform -1 0 3050 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__351_
timestamp 0
transform 1 0 3010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__352_
timestamp 0
transform -1 0 2790 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__353_
timestamp 0
transform 1 0 2410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__354_
timestamp 0
transform -1 0 3330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__355_
timestamp 0
transform -1 0 4170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__356_
timestamp 0
transform 1 0 3850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__357_
timestamp 0
transform -1 0 2730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__358_
timestamp 0
transform -1 0 2910 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__359_
timestamp 0
transform 1 0 3170 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__360_
timestamp 0
transform -1 0 3470 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__361_
timestamp 0
transform -1 0 3250 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__362_
timestamp 0
transform -1 0 3190 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__363_
timestamp 0
transform 1 0 2370 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__364_
timestamp 0
transform 1 0 2230 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__365_
timestamp 0
transform 1 0 3210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__366_
timestamp 0
transform 1 0 2890 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__367_
timestamp 0
transform -1 0 2150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__368_
timestamp 0
transform 1 0 2910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__369_
timestamp 0
transform -1 0 3350 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__370_
timestamp 0
transform 1 0 4950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__371_
timestamp 0
transform 1 0 4650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__372_
timestamp 0
transform 1 0 3330 0 1 250
box -6 -8 26 248
use FILL  FILL_7__373_
timestamp 0
transform 1 0 3330 0 1 730
box -6 -8 26 248
use FILL  FILL_7__374_
timestamp 0
transform 1 0 4150 0 1 730
box -6 -8 26 248
use FILL  FILL_7__375_
timestamp 0
transform 1 0 3870 0 1 730
box -6 -8 26 248
use FILL  FILL_7__376_
timestamp 0
transform 1 0 4430 0 1 730
box -6 -8 26 248
use FILL  FILL_7__377_
timestamp 0
transform -1 0 4130 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__378_
timestamp 0
transform -1 0 4250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__379_
timestamp 0
transform -1 0 2350 0 1 250
box -6 -8 26 248
use FILL  FILL_7__380_
timestamp 0
transform 1 0 1670 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__381_
timestamp 0
transform 1 0 1370 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__382_
timestamp 0
transform -1 0 1050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__383_
timestamp 0
transform 1 0 1510 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__384_
timestamp 0
transform -1 0 970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__385_
timestamp 0
transform -1 0 1010 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__386_
timestamp 0
transform 1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__387_
timestamp 0
transform -1 0 890 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__388_
timestamp 0
transform -1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__389_
timestamp 0
transform -1 0 1590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__390_
timestamp 0
transform -1 0 1290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__391_
timestamp 0
transform 1 0 970 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__392_
timestamp 0
transform -1 0 770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__393_
timestamp 0
transform 1 0 1230 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__394_
timestamp 0
transform 1 0 1790 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__395_
timestamp 0
transform -1 0 3750 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__396_
timestamp 0
transform 1 0 1230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__397_
timestamp 0
transform 1 0 1490 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__398_
timestamp 0
transform 1 0 2030 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__399_
timestamp 0
transform 1 0 2030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__400_
timestamp 0
transform 1 0 1770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__401_
timestamp 0
transform 1 0 1490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__402_
timestamp 0
transform 1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__403_
timestamp 0
transform -1 0 2890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__404_
timestamp 0
transform 1 0 2590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__405_
timestamp 0
transform -1 0 1370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__406_
timestamp 0
transform 1 0 1250 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__407_
timestamp 0
transform -1 0 1530 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__408_
timestamp 0
transform -1 0 1010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__409_
timestamp 0
transform 1 0 1270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__410_
timestamp 0
transform -1 0 1190 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__411_
timestamp 0
transform -1 0 3270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__412_
timestamp 0
transform -1 0 1770 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__413_
timestamp 0
transform 1 0 1610 0 1 730
box -6 -8 26 248
use FILL  FILL_7__414_
timestamp 0
transform 1 0 1890 0 1 730
box -6 -8 26 248
use FILL  FILL_7__415_
timestamp 0
transform 1 0 2750 0 1 730
box -6 -8 26 248
use FILL  FILL_7__416_
timestamp 0
transform -1 0 2110 0 1 250
box -6 -8 26 248
use FILL  FILL_7__417_
timestamp 0
transform 1 0 2470 0 1 730
box -6 -8 26 248
use FILL  FILL_7__418_
timestamp 0
transform 1 0 2310 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__419_
timestamp 0
transform -1 0 3070 0 1 730
box -6 -8 26 248
use FILL  FILL_7__420_
timestamp 0
transform -1 0 2970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__421_
timestamp 0
transform 1 0 4630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__422_
timestamp 0
transform 1 0 4410 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__423_
timestamp 0
transform 1 0 4950 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__424_
timestamp 0
transform 1 0 4950 0 1 250
box -6 -8 26 248
use FILL  FILL_7__425_
timestamp 0
transform 1 0 4410 0 1 250
box -6 -8 26 248
use FILL  FILL_7__426_
timestamp 0
transform -1 0 4690 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__427_
timestamp 0
transform -1 0 2630 0 1 250
box -6 -8 26 248
use FILL  FILL_7__428_
timestamp 0
transform 1 0 2190 0 1 730
box -6 -8 26 248
use FILL  FILL_7__429_
timestamp 0
transform 1 0 2590 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__430_
timestamp 0
transform -1 0 1470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__431_
timestamp 0
transform 1 0 1750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__432_
timestamp 0
transform -1 0 2350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__433_
timestamp 0
transform 1 0 2610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__434_
timestamp 0
transform -1 0 4390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__435_
timestamp 0
transform 1 0 3510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__436_
timestamp 0
transform -1 0 3810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__437_
timestamp 0
transform -1 0 2350 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__438_
timestamp 0
transform -1 0 2610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7__439_
timestamp 0
transform 1 0 2630 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__440_
timestamp 0
transform -1 0 3190 0 1 2170
box -6 -8 26 248
use FILL  FILL_7__441_
timestamp 0
transform 1 0 1570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__442_
timestamp 0
transform -1 0 2150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__443_
timestamp 0
transform -1 0 1770 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__444_
timestamp 0
transform -1 0 2210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__445_
timestamp 0
transform -1 0 1910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__446_
timestamp 0
transform 1 0 2050 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__447_
timestamp 0
transform -1 0 4290 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__448_
timestamp 0
transform -1 0 1850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__449_
timestamp 0
transform 1 0 2330 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__450_
timestamp 0
transform 1 0 2410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7__451_
timestamp 0
transform 1 0 2590 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__452_
timestamp 0
transform -1 0 3730 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__453_
timestamp 0
transform 1 0 1490 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__454_
timestamp 0
transform -1 0 1730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__455_
timestamp 0
transform 1 0 2070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__456_
timestamp 0
transform -1 0 2010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__457_
timestamp 0
transform 1 0 1750 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__458_
timestamp 0
transform 1 0 1830 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__459_
timestamp 0
transform 1 0 2290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__460_
timestamp 0
transform -1 0 2610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__461_
timestamp 0
transform -1 0 2150 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__462_
timestamp 0
transform 1 0 2410 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__463_
timestamp 0
transform 1 0 2710 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__464_
timestamp 0
transform -1 0 3030 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__465_
timestamp 0
transform 1 0 1290 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__466_
timestamp 0
transform -1 0 1010 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__467_
timestamp 0
transform 1 0 690 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__468_
timestamp 0
transform -1 0 450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__469_
timestamp 0
transform -1 0 430 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__470_
timestamp 0
transform -1 0 730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__471_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__472_
timestamp 0
transform -1 0 970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__473_
timestamp 0
transform 1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__474_
timestamp 0
transform 1 0 990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__475_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__476_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__477_
timestamp 0
transform 1 0 410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__478_
timestamp 0
transform -1 0 450 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__479_
timestamp 0
transform -1 0 3550 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__480_
timestamp 0
transform -1 0 1330 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__481_
timestamp 0
transform -1 0 170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__482_
timestamp 0
transform -1 0 1290 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__483_
timestamp 0
transform -1 0 1570 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__484_
timestamp 0
transform 1 0 1730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__485_
timestamp 0
transform 1 0 2030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__486_
timestamp 0
transform 1 0 2310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__487_
timestamp 0
transform 1 0 2890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__488_
timestamp 0
transform 1 0 2590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__489_
timestamp 0
transform 1 0 1570 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__490_
timestamp 0
transform -1 0 1850 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__491_
timestamp 0
transform 1 0 2130 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__492_
timestamp 0
transform 1 0 2410 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__493_
timestamp 0
transform -1 0 2730 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__494_
timestamp 0
transform 1 0 1210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__495_
timestamp 0
transform 1 0 1490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__496_
timestamp 0
transform 1 0 1770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__497_
timestamp 0
transform 1 0 2150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__498_
timestamp 0
transform -1 0 2370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__499_
timestamp 0
transform -1 0 1850 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__500_
timestamp 0
transform -1 0 2390 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__501_
timestamp 0
transform -1 0 2770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__502_
timestamp 0
transform -1 0 3330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__503_
timestamp 0
transform -1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__504_
timestamp 0
transform 1 0 4610 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__505_
timestamp 0
transform -1 0 4890 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__506_
timestamp 0
transform 1 0 4690 0 1 250
box -6 -8 26 248
use FILL  FILL_7__507_
timestamp 0
transform -1 0 4730 0 1 730
box -6 -8 26 248
use FILL  FILL_7__508_
timestamp 0
transform -1 0 2970 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__509_
timestamp 0
transform 1 0 2110 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__510_
timestamp 0
transform -1 0 2670 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__511_
timestamp 0
transform 1 0 1570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__512_
timestamp 0
transform 1 0 2450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__513_
timestamp 0
transform -1 0 3230 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__514_
timestamp 0
transform 1 0 3470 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__515_
timestamp 0
transform -1 0 3790 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__516_
timestamp 0
transform 1 0 690 0 1 250
box -6 -8 26 248
use FILL  FILL_7__517_
timestamp 0
transform 1 0 970 0 1 250
box -6 -8 26 248
use FILL  FILL_7__518_
timestamp 0
transform 1 0 1530 0 1 250
box -6 -8 26 248
use FILL  FILL_7__519_
timestamp 0
transform 1 0 1810 0 1 250
box -6 -8 26 248
use FILL  FILL_7__520_
timestamp 0
transform -1 0 1670 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__521_
timestamp 0
transform -1 0 1950 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__522_
timestamp 0
transform -1 0 3610 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__523_
timestamp 0
transform -1 0 3890 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__524_
timestamp 0
transform -1 0 1230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__525_
timestamp 0
transform 1 0 1250 0 1 250
box -6 -8 26 248
use FILL  FILL_7__526_
timestamp 0
transform -1 0 950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__527_
timestamp 0
transform -1 0 1090 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__528_
timestamp 0
transform 1 0 3150 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__529_
timestamp 0
transform 1 0 1330 0 1 730
box -6 -8 26 248
use FILL  FILL_7__530_
timestamp 0
transform 1 0 1030 0 1 730
box -6 -8 26 248
use FILL  FILL_7__531_
timestamp 0
transform -1 0 570 0 1 1210
box -6 -8 26 248
use FILL  FILL_7__532_
timestamp 0
transform 1 0 410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__533_
timestamp 0
transform -1 0 450 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__534_
timestamp 0
transform 1 0 710 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__535_
timestamp 0
transform -1 0 2470 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__536_
timestamp 0
transform -1 0 2750 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__537_
timestamp 0
transform -1 0 3030 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__538_
timestamp 0
transform -1 0 3310 0 -1 250
box -6 -8 26 248
use FILL  FILL_7__539_
timestamp 0
transform -1 0 170 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__540_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__541_
timestamp 0
transform 1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_7__542_
timestamp 0
transform -1 0 470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7__543_
timestamp 0
transform -1 0 3530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__544_
timestamp 0
transform -1 0 3790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_7__545_
timestamp 0
transform -1 0 3950 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__546_
timestamp 0
transform 1 0 3630 0 -1 730
box -6 -8 26 248
use FILL  FILL_7__547_
timestamp 0
transform 1 0 2710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7__548_
timestamp 0
transform -1 0 2290 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__549_
timestamp 0
transform -1 0 3610 0 1 250
box -6 -8 26 248
use FILL  FILL_7__550_
timestamp 0
transform -1 0 3890 0 1 250
box -6 -8 26 248
use FILL  FILL_7__551_
timestamp 0
transform 1 0 1030 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__552_
timestamp 0
transform 1 0 730 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__553_
timestamp 0
transform -1 0 970 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__554_
timestamp 0
transform 1 0 670 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__555_
timestamp 0
transform 1 0 450 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__556_
timestamp 0
transform -1 0 170 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__613_
timestamp 0
transform 1 0 4870 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__614_
timestamp 0
transform -1 0 4850 0 1 2650
box -6 -8 26 248
use FILL  FILL_7__615_
timestamp 0
transform 1 0 4390 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__616_
timestamp 0
transform -1 0 4450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__617_
timestamp 0
transform 1 0 4590 0 1 3130
box -6 -8 26 248
use FILL  FILL_7__618_
timestamp 0
transform 1 0 4910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7__619_
timestamp 0
transform 1 0 4890 0 1 3610
box -6 -8 26 248
use FILL  FILL_7__620_
timestamp 0
transform 1 0 4750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7__621_
timestamp 0
transform 1 0 4890 0 1 4090
box -6 -8 26 248
use FILL  FILL_7__622_
timestamp 0
transform 1 0 4950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7__623_
timestamp 0
transform 1 0 4670 0 1 4570
box -6 -8 26 248
use FILL  FILL_7__624_
timestamp 0
transform 1 0 4710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7__625_
timestamp 0
transform 1 0 3390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert7
timestamp 0
transform 1 0 4570 0 1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert8
timestamp 0
transform -1 0 4490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert9
timestamp 0
transform 1 0 4610 0 1 4090
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert10
timestamp 0
transform 1 0 4630 0 1 3610
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert11
timestamp 0
transform -1 0 1310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert12
timestamp 0
transform 1 0 1870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert13
timestamp 0
transform 1 0 1850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert14
timestamp 0
transform 1 0 2510 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert15
timestamp 0
transform -1 0 690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert16
timestamp 0
transform 1 0 2890 0 1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert17
timestamp 0
transform 1 0 1950 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert18
timestamp 0
transform 1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert19
timestamp 0
transform -1 0 1050 0 1 4570
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert20
timestamp 0
transform 1 0 2970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert21
timestamp 0
transform 1 0 4030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert22
timestamp 0
transform -1 0 3270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert23
timestamp 0
transform -1 0 3530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert24
timestamp 0
transform -1 0 2970 0 1 3130
box -6 -8 26 248
use FILL  FILL_7_BUFX2_insert25
timestamp 0
transform 1 0 2890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert0
timestamp 0
transform -1 0 3690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert1
timestamp 0
transform -1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert2
timestamp 0
transform 1 0 150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert3
timestamp 0
transform 1 0 2570 0 1 3130
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert4
timestamp 0
transform 1 0 4210 0 -1 730
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert5
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_7_CLKBUF1_insert6
timestamp 0
transform 1 0 3710 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__273_
timestamp 0
transform -1 0 4430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__274_
timestamp 0
transform -1 0 4670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__275_
timestamp 0
transform -1 0 4950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__276_
timestamp 0
transform -1 0 3750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__277_
timestamp 0
transform 1 0 4970 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__278_
timestamp 0
transform 1 0 4930 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__279_
timestamp 0
transform 1 0 4570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__280_
timestamp 0
transform -1 0 4790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__281_
timestamp 0
transform -1 0 4850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__282_
timestamp 0
transform 1 0 4030 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__283_
timestamp 0
transform -1 0 3550 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__284_
timestamp 0
transform 1 0 4050 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__285_
timestamp 0
transform 1 0 3430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__286_
timestamp 0
transform -1 0 4670 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__287_
timestamp 0
transform 1 0 4630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__288_
timestamp 0
transform 1 0 3570 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__289_
timestamp 0
transform -1 0 4350 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__290_
timestamp 0
transform 1 0 4090 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__291_
timestamp 0
transform 1 0 1490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__292_
timestamp 0
transform -1 0 4090 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__293_
timestamp 0
transform -1 0 4350 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__294_
timestamp 0
transform 1 0 3930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__295_
timestamp 0
transform -1 0 4390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__296_
timestamp 0
transform 1 0 4670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__297_
timestamp 0
transform 1 0 4190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__298_
timestamp 0
transform -1 0 4110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__299_
timestamp 0
transform -1 0 4150 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__300_
timestamp 0
transform 1 0 3290 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__301_
timestamp 0
transform -1 0 3830 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__302_
timestamp 0
transform -1 0 3850 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__303_
timestamp 0
transform 1 0 3850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__304_
timestamp 0
transform -1 0 4110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__305_
timestamp 0
transform -1 0 4390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__306_
timestamp 0
transform 1 0 3930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__307_
timestamp 0
transform 1 0 4390 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__308_
timestamp 0
transform 1 0 4190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__309_
timestamp 0
transform -1 0 770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__310_
timestamp 0
transform -1 0 190 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__311_
timestamp 0
transform -1 0 190 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__312_
timestamp 0
transform -1 0 430 0 1 250
box -6 -8 26 248
use FILL  FILL_8__313_
timestamp 0
transform 1 0 410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__314_
timestamp 0
transform 1 0 410 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__315_
timestamp 0
transform 1 0 1590 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__316_
timestamp 0
transform -1 0 950 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__317_
timestamp 0
transform 1 0 650 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__318_
timestamp 0
transform -1 0 850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__319_
timestamp 0
transform -1 0 950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__320_
timestamp 0
transform -1 0 1490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__321_
timestamp 0
transform 1 0 1630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__322_
timestamp 0
transform 1 0 1490 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__323_
timestamp 0
transform -1 0 590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__324_
timestamp 0
transform 1 0 170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__325_
timestamp 0
transform 1 0 410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__326_
timestamp 0
transform -1 0 430 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__327_
timestamp 0
transform -1 0 190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__328_
timestamp 0
transform 1 0 710 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__329_
timestamp 0
transform 1 0 470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__330_
timestamp 0
transform 1 0 2890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__331_
timestamp 0
transform 1 0 3450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__332_
timestamp 0
transform 1 0 3150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__333_
timestamp 0
transform 1 0 2370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__334_
timestamp 0
transform 1 0 2110 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__335_
timestamp 0
transform -1 0 2090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__336_
timestamp 0
transform -1 0 190 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__337_
timestamp 0
transform 1 0 170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__338_
timestamp 0
transform -1 0 450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__339_
timestamp 0
transform 1 0 3610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__340_
timestamp 0
transform -1 0 4130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__341_
timestamp 0
transform -1 0 4610 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__342_
timestamp 0
transform 1 0 4290 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__343_
timestamp 0
transform 1 0 3630 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__344_
timestamp 0
transform 1 0 3650 0 1 730
box -6 -8 26 248
use FILL  FILL_8__345_
timestamp 0
transform 1 0 4090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__346_
timestamp 0
transform 1 0 4170 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__347_
timestamp 0
transform -1 0 4950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__348_
timestamp 0
transform 1 0 4690 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__349_
timestamp 0
transform 1 0 2650 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__350_
timestamp 0
transform -1 0 3070 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__351_
timestamp 0
transform 1 0 3030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__352_
timestamp 0
transform -1 0 2810 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__353_
timestamp 0
transform 1 0 2430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__354_
timestamp 0
transform -1 0 3350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__355_
timestamp 0
transform -1 0 4190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__356_
timestamp 0
transform 1 0 3870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__357_
timestamp 0
transform -1 0 2750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__358_
timestamp 0
transform -1 0 2930 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__359_
timestamp 0
transform 1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__360_
timestamp 0
transform -1 0 3490 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__361_
timestamp 0
transform -1 0 3270 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__362_
timestamp 0
transform -1 0 3210 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__363_
timestamp 0
transform 1 0 2390 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__364_
timestamp 0
transform 1 0 2250 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__365_
timestamp 0
transform 1 0 3230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__366_
timestamp 0
transform 1 0 2910 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__367_
timestamp 0
transform -1 0 2170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__368_
timestamp 0
transform 1 0 2930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__369_
timestamp 0
transform -1 0 3370 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__370_
timestamp 0
transform 1 0 4970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__371_
timestamp 0
transform 1 0 4670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__372_
timestamp 0
transform 1 0 3350 0 1 250
box -6 -8 26 248
use FILL  FILL_8__373_
timestamp 0
transform 1 0 3350 0 1 730
box -6 -8 26 248
use FILL  FILL_8__374_
timestamp 0
transform 1 0 4170 0 1 730
box -6 -8 26 248
use FILL  FILL_8__375_
timestamp 0
transform 1 0 3890 0 1 730
box -6 -8 26 248
use FILL  FILL_8__376_
timestamp 0
transform 1 0 4450 0 1 730
box -6 -8 26 248
use FILL  FILL_8__377_
timestamp 0
transform -1 0 4150 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__378_
timestamp 0
transform -1 0 4270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__379_
timestamp 0
transform -1 0 2370 0 1 250
box -6 -8 26 248
use FILL  FILL_8__380_
timestamp 0
transform 1 0 1690 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__381_
timestamp 0
transform 1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__382_
timestamp 0
transform -1 0 1070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__383_
timestamp 0
transform 1 0 1530 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__384_
timestamp 0
transform -1 0 990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__385_
timestamp 0
transform -1 0 1030 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__386_
timestamp 0
transform 1 0 1090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__387_
timestamp 0
transform -1 0 910 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__388_
timestamp 0
transform -1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__389_
timestamp 0
transform -1 0 1610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__390_
timestamp 0
transform -1 0 1310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__391_
timestamp 0
transform 1 0 990 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__392_
timestamp 0
transform -1 0 790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__393_
timestamp 0
transform 1 0 1250 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__394_
timestamp 0
transform 1 0 1810 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__395_
timestamp 0
transform -1 0 3770 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__396_
timestamp 0
transform 1 0 1250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__397_
timestamp 0
transform 1 0 1510 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__398_
timestamp 0
transform 1 0 2050 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__399_
timestamp 0
transform 1 0 2050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__400_
timestamp 0
transform 1 0 1790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__401_
timestamp 0
transform 1 0 1510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__402_
timestamp 0
transform 1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__403_
timestamp 0
transform -1 0 2910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__404_
timestamp 0
transform 1 0 2610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__405_
timestamp 0
transform -1 0 1390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__406_
timestamp 0
transform 1 0 1270 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__407_
timestamp 0
transform -1 0 1550 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__408_
timestamp 0
transform -1 0 1030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__409_
timestamp 0
transform 1 0 1290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__410_
timestamp 0
transform -1 0 1210 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__411_
timestamp 0
transform -1 0 3290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__412_
timestamp 0
transform -1 0 1790 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__413_
timestamp 0
transform 1 0 1630 0 1 730
box -6 -8 26 248
use FILL  FILL_8__414_
timestamp 0
transform 1 0 1910 0 1 730
box -6 -8 26 248
use FILL  FILL_8__415_
timestamp 0
transform 1 0 2770 0 1 730
box -6 -8 26 248
use FILL  FILL_8__416_
timestamp 0
transform -1 0 2130 0 1 250
box -6 -8 26 248
use FILL  FILL_8__417_
timestamp 0
transform 1 0 2490 0 1 730
box -6 -8 26 248
use FILL  FILL_8__418_
timestamp 0
transform 1 0 2330 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__419_
timestamp 0
transform -1 0 3090 0 1 730
box -6 -8 26 248
use FILL  FILL_8__420_
timestamp 0
transform -1 0 2990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__421_
timestamp 0
transform 1 0 4650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__422_
timestamp 0
transform 1 0 4430 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__423_
timestamp 0
transform 1 0 4970 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__424_
timestamp 0
transform 1 0 4970 0 1 250
box -6 -8 26 248
use FILL  FILL_8__425_
timestamp 0
transform 1 0 4430 0 1 250
box -6 -8 26 248
use FILL  FILL_8__426_
timestamp 0
transform -1 0 4710 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__427_
timestamp 0
transform -1 0 2650 0 1 250
box -6 -8 26 248
use FILL  FILL_8__428_
timestamp 0
transform 1 0 2210 0 1 730
box -6 -8 26 248
use FILL  FILL_8__429_
timestamp 0
transform 1 0 2610 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__430_
timestamp 0
transform -1 0 1490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__431_
timestamp 0
transform 1 0 1770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__432_
timestamp 0
transform -1 0 2370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__433_
timestamp 0
transform 1 0 2630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__434_
timestamp 0
transform -1 0 4410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__435_
timestamp 0
transform 1 0 3530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__436_
timestamp 0
transform -1 0 3830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__437_
timestamp 0
transform -1 0 2370 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__438_
timestamp 0
transform -1 0 2630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8__439_
timestamp 0
transform 1 0 2650 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__440_
timestamp 0
transform -1 0 3210 0 1 2170
box -6 -8 26 248
use FILL  FILL_8__441_
timestamp 0
transform 1 0 1590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__442_
timestamp 0
transform -1 0 2170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__443_
timestamp 0
transform -1 0 1790 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__444_
timestamp 0
transform -1 0 2230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__445_
timestamp 0
transform -1 0 1930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__446_
timestamp 0
transform 1 0 2070 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__447_
timestamp 0
transform -1 0 4310 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__448_
timestamp 0
transform -1 0 1870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__449_
timestamp 0
transform 1 0 2350 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__450_
timestamp 0
transform 1 0 2430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8__451_
timestamp 0
transform 1 0 2610 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__452_
timestamp 0
transform -1 0 3750 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__453_
timestamp 0
transform 1 0 1510 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__454_
timestamp 0
transform -1 0 1750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__455_
timestamp 0
transform 1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__456_
timestamp 0
transform -1 0 2030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__457_
timestamp 0
transform 1 0 1770 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__458_
timestamp 0
transform 1 0 1850 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__459_
timestamp 0
transform 1 0 2310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__460_
timestamp 0
transform -1 0 2630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__461_
timestamp 0
transform -1 0 2170 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__462_
timestamp 0
transform 1 0 2430 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__463_
timestamp 0
transform 1 0 2730 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__464_
timestamp 0
transform -1 0 3050 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__465_
timestamp 0
transform 1 0 1310 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__466_
timestamp 0
transform -1 0 1030 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__467_
timestamp 0
transform 1 0 710 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__468_
timestamp 0
transform -1 0 470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__469_
timestamp 0
transform -1 0 450 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__470_
timestamp 0
transform -1 0 750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__471_
timestamp 0
transform 1 0 750 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__472_
timestamp 0
transform -1 0 990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__473_
timestamp 0
transform 1 0 930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__474_
timestamp 0
transform 1 0 1010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__475_
timestamp 0
transform -1 0 190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__476_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__477_
timestamp 0
transform 1 0 430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__478_
timestamp 0
transform -1 0 470 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__479_
timestamp 0
transform -1 0 3570 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__480_
timestamp 0
transform -1 0 1350 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__481_
timestamp 0
transform -1 0 190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__482_
timestamp 0
transform -1 0 1310 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__483_
timestamp 0
transform -1 0 1590 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__484_
timestamp 0
transform 1 0 1750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__485_
timestamp 0
transform 1 0 2050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__486_
timestamp 0
transform 1 0 2330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__487_
timestamp 0
transform 1 0 2910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__488_
timestamp 0
transform 1 0 2610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__489_
timestamp 0
transform 1 0 1590 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__490_
timestamp 0
transform -1 0 1870 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__491_
timestamp 0
transform 1 0 2150 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__492_
timestamp 0
transform 1 0 2430 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__493_
timestamp 0
transform -1 0 2750 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__494_
timestamp 0
transform 1 0 1230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__495_
timestamp 0
transform 1 0 1510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__496_
timestamp 0
transform 1 0 1790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__497_
timestamp 0
transform 1 0 2170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__498_
timestamp 0
transform -1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__499_
timestamp 0
transform -1 0 1870 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__500_
timestamp 0
transform -1 0 2410 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__501_
timestamp 0
transform -1 0 2790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__502_
timestamp 0
transform -1 0 3350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__503_
timestamp 0
transform -1 0 3430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__504_
timestamp 0
transform 1 0 4630 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__505_
timestamp 0
transform -1 0 4910 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__506_
timestamp 0
transform 1 0 4710 0 1 250
box -6 -8 26 248
use FILL  FILL_8__507_
timestamp 0
transform -1 0 4750 0 1 730
box -6 -8 26 248
use FILL  FILL_8__508_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__509_
timestamp 0
transform 1 0 2130 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__510_
timestamp 0
transform -1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__511_
timestamp 0
transform 1 0 1590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__512_
timestamp 0
transform 1 0 2470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__513_
timestamp 0
transform -1 0 3250 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__514_
timestamp 0
transform 1 0 3490 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__515_
timestamp 0
transform -1 0 3810 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__516_
timestamp 0
transform 1 0 710 0 1 250
box -6 -8 26 248
use FILL  FILL_8__517_
timestamp 0
transform 1 0 990 0 1 250
box -6 -8 26 248
use FILL  FILL_8__518_
timestamp 0
transform 1 0 1550 0 1 250
box -6 -8 26 248
use FILL  FILL_8__519_
timestamp 0
transform 1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_8__520_
timestamp 0
transform -1 0 1690 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__521_
timestamp 0
transform -1 0 1970 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__522_
timestamp 0
transform -1 0 3630 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__523_
timestamp 0
transform -1 0 3910 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__524_
timestamp 0
transform -1 0 1250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__525_
timestamp 0
transform 1 0 1270 0 1 250
box -6 -8 26 248
use FILL  FILL_8__526_
timestamp 0
transform -1 0 970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__527_
timestamp 0
transform -1 0 1110 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__528_
timestamp 0
transform 1 0 3170 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__529_
timestamp 0
transform 1 0 1350 0 1 730
box -6 -8 26 248
use FILL  FILL_8__530_
timestamp 0
transform 1 0 1050 0 1 730
box -6 -8 26 248
use FILL  FILL_8__531_
timestamp 0
transform -1 0 590 0 1 1210
box -6 -8 26 248
use FILL  FILL_8__532_
timestamp 0
transform 1 0 430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__533_
timestamp 0
transform -1 0 470 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__534_
timestamp 0
transform 1 0 730 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__535_
timestamp 0
transform -1 0 2490 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__536_
timestamp 0
transform -1 0 2770 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__537_
timestamp 0
transform -1 0 3050 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__538_
timestamp 0
transform -1 0 3330 0 -1 250
box -6 -8 26 248
use FILL  FILL_8__539_
timestamp 0
transform -1 0 190 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__540_
timestamp 0
transform -1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__541_
timestamp 0
transform 1 0 450 0 1 1690
box -6 -8 26 248
use FILL  FILL_8__542_
timestamp 0
transform -1 0 490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8__543_
timestamp 0
transform -1 0 3550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__544_
timestamp 0
transform -1 0 3810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_8__545_
timestamp 0
transform -1 0 3970 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__546_
timestamp 0
transform 1 0 3650 0 -1 730
box -6 -8 26 248
use FILL  FILL_8__547_
timestamp 0
transform 1 0 2730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8__548_
timestamp 0
transform -1 0 2310 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__549_
timestamp 0
transform -1 0 3630 0 1 250
box -6 -8 26 248
use FILL  FILL_8__550_
timestamp 0
transform -1 0 3910 0 1 250
box -6 -8 26 248
use FILL  FILL_8__551_
timestamp 0
transform 1 0 1050 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__552_
timestamp 0
transform 1 0 750 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__553_
timestamp 0
transform -1 0 990 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__554_
timestamp 0
transform 1 0 690 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__555_
timestamp 0
transform 1 0 470 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__556_
timestamp 0
transform -1 0 190 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__613_
timestamp 0
transform 1 0 4890 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__614_
timestamp 0
transform -1 0 4870 0 1 2650
box -6 -8 26 248
use FILL  FILL_8__615_
timestamp 0
transform 1 0 4410 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__616_
timestamp 0
transform -1 0 4470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__617_
timestamp 0
transform 1 0 4610 0 1 3130
box -6 -8 26 248
use FILL  FILL_8__618_
timestamp 0
transform 1 0 4930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8__619_
timestamp 0
transform 1 0 4910 0 1 3610
box -6 -8 26 248
use FILL  FILL_8__620_
timestamp 0
transform 1 0 4770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8__621_
timestamp 0
transform 1 0 4910 0 1 4090
box -6 -8 26 248
use FILL  FILL_8__622_
timestamp 0
transform 1 0 4970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8__623_
timestamp 0
transform 1 0 4690 0 1 4570
box -6 -8 26 248
use FILL  FILL_8__624_
timestamp 0
transform 1 0 4730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8__625_
timestamp 0
transform 1 0 3410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert7
timestamp 0
transform 1 0 4590 0 1 2650
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert8
timestamp 0
transform -1 0 4510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert9
timestamp 0
transform 1 0 4630 0 1 4090
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert10
timestamp 0
transform 1 0 4650 0 1 3610
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert11
timestamp 0
transform -1 0 1330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert12
timestamp 0
transform 1 0 1890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert13
timestamp 0
transform 1 0 1870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert14
timestamp 0
transform 1 0 2530 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert15
timestamp 0
transform -1 0 710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert16
timestamp 0
transform 1 0 2910 0 1 2650
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert17
timestamp 0
transform 1 0 1970 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert18
timestamp 0
transform 1 0 3070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert19
timestamp 0
transform -1 0 1070 0 1 4570
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert20
timestamp 0
transform 1 0 2990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert21
timestamp 0
transform 1 0 4050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert22
timestamp 0
transform -1 0 3290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert23
timestamp 0
transform -1 0 3550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert24
timestamp 0
transform -1 0 2990 0 1 3130
box -6 -8 26 248
use FILL  FILL_8_BUFX2_insert25
timestamp 0
transform 1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert0
timestamp 0
transform -1 0 3710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert1
timestamp 0
transform -1 0 190 0 1 1210
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert2
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert3
timestamp 0
transform 1 0 2590 0 1 3130
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert4
timestamp 0
transform 1 0 4230 0 -1 730
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert5
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 26 248
use FILL  FILL_8_CLKBUF1_insert6
timestamp 0
transform 1 0 3730 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__274_
timestamp 0
transform -1 0 4690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__275_
timestamp 0
transform -1 0 4970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__276_
timestamp 0
transform -1 0 3770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__278_
timestamp 0
transform 1 0 4950 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__279_
timestamp 0
transform 1 0 4590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__281_
timestamp 0
transform -1 0 4870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__282_
timestamp 0
transform 1 0 4050 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__283_
timestamp 0
transform -1 0 3570 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__285_
timestamp 0
transform 1 0 3450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__286_
timestamp 0
transform -1 0 4690 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__287_
timestamp 0
transform 1 0 4650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__289_
timestamp 0
transform -1 0 4370 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__290_
timestamp 0
transform 1 0 4110 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__291_
timestamp 0
transform 1 0 1510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__293_
timestamp 0
transform -1 0 4370 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__294_
timestamp 0
transform 1 0 3950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__296_
timestamp 0
transform 1 0 4690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__297_
timestamp 0
transform 1 0 4210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__298_
timestamp 0
transform -1 0 4130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__300_
timestamp 0
transform 1 0 3310 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__301_
timestamp 0
transform -1 0 3850 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__302_
timestamp 0
transform -1 0 3870 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__304_
timestamp 0
transform -1 0 4130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__305_
timestamp 0
transform -1 0 4410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__306_
timestamp 0
transform 1 0 3950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__308_
timestamp 0
transform 1 0 4210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__309_
timestamp 0
transform -1 0 790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__311_
timestamp 0
transform -1 0 210 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__312_
timestamp 0
transform -1 0 450 0 1 250
box -6 -8 26 248
use FILL  FILL_9__313_
timestamp 0
transform 1 0 430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__315_
timestamp 0
transform 1 0 1610 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__316_
timestamp 0
transform -1 0 970 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__317_
timestamp 0
transform 1 0 670 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__319_
timestamp 0
transform -1 0 970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__320_
timestamp 0
transform -1 0 1510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__321_
timestamp 0
transform 1 0 1650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__323_
timestamp 0
transform -1 0 610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__324_
timestamp 0
transform 1 0 190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__326_
timestamp 0
transform -1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__327_
timestamp 0
transform -1 0 210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__328_
timestamp 0
transform 1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__330_
timestamp 0
transform 1 0 2910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__331_
timestamp 0
transform 1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__332_
timestamp 0
transform 1 0 3170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__334_
timestamp 0
transform 1 0 2130 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__335_
timestamp 0
transform -1 0 2110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__336_
timestamp 0
transform -1 0 210 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__338_
timestamp 0
transform -1 0 470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__339_
timestamp 0
transform 1 0 3630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__341_
timestamp 0
transform -1 0 4630 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__342_
timestamp 0
transform 1 0 4310 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__343_
timestamp 0
transform 1 0 3650 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__345_
timestamp 0
transform 1 0 4110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__346_
timestamp 0
transform 1 0 4190 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__347_
timestamp 0
transform -1 0 4970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__349_
timestamp 0
transform 1 0 2670 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__350_
timestamp 0
transform -1 0 3090 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__351_
timestamp 0
transform 1 0 3050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__353_
timestamp 0
transform 1 0 2450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__354_
timestamp 0
transform -1 0 3370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__356_
timestamp 0
transform 1 0 3890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__357_
timestamp 0
transform -1 0 2770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__358_
timestamp 0
transform -1 0 2950 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__360_
timestamp 0
transform -1 0 3510 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__361_
timestamp 0
transform -1 0 3290 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__362_
timestamp 0
transform -1 0 3230 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__364_
timestamp 0
transform 1 0 2270 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__365_
timestamp 0
transform 1 0 3250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__366_
timestamp 0
transform 1 0 2930 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__368_
timestamp 0
transform 1 0 2950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__369_
timestamp 0
transform -1 0 3390 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__371_
timestamp 0
transform 1 0 4690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__372_
timestamp 0
transform 1 0 3370 0 1 250
box -6 -8 26 248
use FILL  FILL_9__373_
timestamp 0
transform 1 0 3370 0 1 730
box -6 -8 26 248
use FILL  FILL_9__375_
timestamp 0
transform 1 0 3910 0 1 730
box -6 -8 26 248
use FILL  FILL_9__376_
timestamp 0
transform 1 0 4470 0 1 730
box -6 -8 26 248
use FILL  FILL_9__377_
timestamp 0
transform -1 0 4170 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__379_
timestamp 0
transform -1 0 2390 0 1 250
box -6 -8 26 248
use FILL  FILL_9__380_
timestamp 0
transform 1 0 1710 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__381_
timestamp 0
transform 1 0 1410 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__383_
timestamp 0
transform 1 0 1550 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__384_
timestamp 0
transform -1 0 1010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__386_
timestamp 0
transform 1 0 1110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__387_
timestamp 0
transform -1 0 930 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__388_
timestamp 0
transform -1 0 4030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__390_
timestamp 0
transform -1 0 1330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__391_
timestamp 0
transform 1 0 1010 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__392_
timestamp 0
transform -1 0 810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__394_
timestamp 0
transform 1 0 1830 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__395_
timestamp 0
transform -1 0 3790 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__396_
timestamp 0
transform 1 0 1270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__398_
timestamp 0
transform 1 0 2070 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__399_
timestamp 0
transform 1 0 2070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__401_
timestamp 0
transform 1 0 1530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9__402_
timestamp 0
transform 1 0 1850 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__403_
timestamp 0
transform -1 0 2930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__405_
timestamp 0
transform -1 0 1410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__406_
timestamp 0
transform 1 0 1290 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__407_
timestamp 0
transform -1 0 1570 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__409_
timestamp 0
transform 1 0 1310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__410_
timestamp 0
transform -1 0 1230 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__411_
timestamp 0
transform -1 0 3310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__413_
timestamp 0
transform 1 0 1650 0 1 730
box -6 -8 26 248
use FILL  FILL_9__414_
timestamp 0
transform 1 0 1930 0 1 730
box -6 -8 26 248
use FILL  FILL_9__415_
timestamp 0
transform 1 0 2790 0 1 730
box -6 -8 26 248
use FILL  FILL_9__417_
timestamp 0
transform 1 0 2510 0 1 730
box -6 -8 26 248
use FILL  FILL_9__418_
timestamp 0
transform 1 0 2350 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__420_
timestamp 0
transform -1 0 3010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__421_
timestamp 0
transform 1 0 4670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__422_
timestamp 0
transform 1 0 4450 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__424_
timestamp 0
transform 1 0 4990 0 1 250
box -6 -8 26 248
use FILL  FILL_9__425_
timestamp 0
transform 1 0 4450 0 1 250
box -6 -8 26 248
use FILL  FILL_9__426_
timestamp 0
transform -1 0 4730 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__428_
timestamp 0
transform 1 0 2230 0 1 730
box -6 -8 26 248
use FILL  FILL_9__429_
timestamp 0
transform 1 0 2630 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__430_
timestamp 0
transform -1 0 1510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__432_
timestamp 0
transform -1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__433_
timestamp 0
transform 1 0 2650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__435_
timestamp 0
transform 1 0 3550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__436_
timestamp 0
transform -1 0 3850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__437_
timestamp 0
transform -1 0 2390 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__439_
timestamp 0
transform 1 0 2670 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__440_
timestamp 0
transform -1 0 3230 0 1 2170
box -6 -8 26 248
use FILL  FILL_9__441_
timestamp 0
transform 1 0 1610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__443_
timestamp 0
transform -1 0 1810 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__444_
timestamp 0
transform -1 0 2250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__445_
timestamp 0
transform -1 0 1950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9__447_
timestamp 0
transform -1 0 4330 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__448_
timestamp 0
transform -1 0 1890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__450_
timestamp 0
transform 1 0 2450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9__451_
timestamp 0
transform 1 0 2630 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__452_
timestamp 0
transform -1 0 3770 0 1 2650
box -6 -8 26 248
use FILL  FILL_9__454_
timestamp 0
transform -1 0 1770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__455_
timestamp 0
transform 1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__456_
timestamp 0
transform -1 0 2050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__458_
timestamp 0
transform 1 0 1870 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__459_
timestamp 0
transform 1 0 2330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__460_
timestamp 0
transform -1 0 2650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9__462_
timestamp 0
transform 1 0 2450 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__463_
timestamp 0
transform 1 0 2750 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__465_
timestamp 0
transform 1 0 1330 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__466_
timestamp 0
transform -1 0 1050 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__467_
timestamp 0
transform 1 0 730 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__469_
timestamp 0
transform -1 0 470 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__470_
timestamp 0
transform -1 0 770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__471_
timestamp 0
transform 1 0 770 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__473_
timestamp 0
transform 1 0 950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__474_
timestamp 0
transform 1 0 1030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__475_
timestamp 0
transform -1 0 210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__477_
timestamp 0
transform 1 0 450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__478_
timestamp 0
transform -1 0 490 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__480_
timestamp 0
transform -1 0 1370 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__481_
timestamp 0
transform -1 0 210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__482_
timestamp 0
transform -1 0 1330 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__484_
timestamp 0
transform 1 0 1770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__485_
timestamp 0
transform 1 0 2070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__486_
timestamp 0
transform 1 0 2350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__488_
timestamp 0
transform 1 0 2630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__489_
timestamp 0
transform 1 0 1610 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__490_
timestamp 0
transform -1 0 1890 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__492_
timestamp 0
transform 1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__493_
timestamp 0
transform -1 0 2770 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__495_
timestamp 0
transform 1 0 1530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__496_
timestamp 0
transform 1 0 1810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__497_
timestamp 0
transform 1 0 2190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__499_
timestamp 0
transform -1 0 1890 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__500_
timestamp 0
transform -1 0 2430 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__501_
timestamp 0
transform -1 0 2810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__503_
timestamp 0
transform -1 0 3450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__504_
timestamp 0
transform 1 0 4650 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__505_
timestamp 0
transform -1 0 4930 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__507_
timestamp 0
transform -1 0 4770 0 1 730
box -6 -8 26 248
use FILL  FILL_9__508_
timestamp 0
transform -1 0 3010 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__510_
timestamp 0
transform -1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__511_
timestamp 0
transform 1 0 1610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__512_
timestamp 0
transform 1 0 2490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9__514_
timestamp 0
transform 1 0 3510 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__515_
timestamp 0
transform -1 0 3830 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__516_
timestamp 0
transform 1 0 730 0 1 250
box -6 -8 26 248
use FILL  FILL_9__518_
timestamp 0
transform 1 0 1570 0 1 250
box -6 -8 26 248
use FILL  FILL_9__519_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_9__520_
timestamp 0
transform -1 0 1710 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__522_
timestamp 0
transform -1 0 3650 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__523_
timestamp 0
transform -1 0 3930 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__525_
timestamp 0
transform 1 0 1290 0 1 250
box -6 -8 26 248
use FILL  FILL_9__526_
timestamp 0
transform -1 0 990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__527_
timestamp 0
transform -1 0 1130 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__529_
timestamp 0
transform 1 0 1370 0 1 730
box -6 -8 26 248
use FILL  FILL_9__530_
timestamp 0
transform 1 0 1070 0 1 730
box -6 -8 26 248
use FILL  FILL_9__531_
timestamp 0
transform -1 0 610 0 1 1210
box -6 -8 26 248
use FILL  FILL_9__533_
timestamp 0
transform -1 0 490 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__534_
timestamp 0
transform 1 0 750 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__535_
timestamp 0
transform -1 0 2510 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__537_
timestamp 0
transform -1 0 3070 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__538_
timestamp 0
transform -1 0 3350 0 -1 250
box -6 -8 26 248
use FILL  FILL_9__540_
timestamp 0
transform -1 0 210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__541_
timestamp 0
transform 1 0 470 0 1 1690
box -6 -8 26 248
use FILL  FILL_9__542_
timestamp 0
transform -1 0 510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9__544_
timestamp 0
transform -1 0 3830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_9__545_
timestamp 0
transform -1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__546_
timestamp 0
transform 1 0 3670 0 -1 730
box -6 -8 26 248
use FILL  FILL_9__548_
timestamp 0
transform -1 0 2330 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__549_
timestamp 0
transform -1 0 3650 0 1 250
box -6 -8 26 248
use FILL  FILL_9__550_
timestamp 0
transform -1 0 3930 0 1 250
box -6 -8 26 248
use FILL  FILL_9__552_
timestamp 0
transform 1 0 770 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__553_
timestamp 0
transform -1 0 1010 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__555_
timestamp 0
transform 1 0 490 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__556_
timestamp 0
transform -1 0 210 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__613_
timestamp 0
transform 1 0 4910 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__615_
timestamp 0
transform 1 0 4430 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__616_
timestamp 0
transform -1 0 4490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__617_
timestamp 0
transform 1 0 4630 0 1 3130
box -6 -8 26 248
use FILL  FILL_9__619_
timestamp 0
transform 1 0 4930 0 1 3610
box -6 -8 26 248
use FILL  FILL_9__620_
timestamp 0
transform 1 0 4790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9__621_
timestamp 0
transform 1 0 4930 0 1 4090
box -6 -8 26 248
use FILL  FILL_9__623_
timestamp 0
transform 1 0 4710 0 1 4570
box -6 -8 26 248
use FILL  FILL_9__624_
timestamp 0
transform 1 0 4750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9__625_
timestamp 0
transform 1 0 3430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert8
timestamp 0
transform -1 0 4530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert9
timestamp 0
transform 1 0 4650 0 1 4090
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert11
timestamp 0
transform -1 0 1350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert12
timestamp 0
transform 1 0 1910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert13
timestamp 0
transform 1 0 1890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert15
timestamp 0
transform -1 0 730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert16
timestamp 0
transform 1 0 2930 0 1 2650
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert17
timestamp 0
transform 1 0 1990 0 1 1210
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert19
timestamp 0
transform -1 0 1090 0 1 4570
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert20
timestamp 0
transform 1 0 3010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert21
timestamp 0
transform 1 0 4070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert23
timestamp 0
transform -1 0 3570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert24
timestamp 0
transform -1 0 3010 0 1 3130
box -6 -8 26 248
use FILL  FILL_9_BUFX2_insert25
timestamp 0
transform 1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert0
timestamp 0
transform -1 0 3730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert1
timestamp 0
transform -1 0 210 0 1 1210
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert2
timestamp 0
transform 1 0 190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert4
timestamp 0
transform 1 0 4250 0 -1 730
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert5
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_9_CLKBUF1_insert6
timestamp 0
transform 1 0 3750 0 1 2170
box -6 -8 26 248
<< labels >>
flabel metal1 s 5082 2 5142 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 4417 5097 4423 5103 3 FreeSans 16 90 0 0 Dout[11]
port 2 nsew
flabel metal2 s 4477 5097 4483 5103 3 FreeSans 16 90 0 0 Dout[10]
port 3 nsew
flabel metal2 s 4717 5097 4723 5103 3 FreeSans 16 90 0 0 Dout[9]
port 4 nsew
flabel metal2 s 4757 5097 4763 5103 3 FreeSans 16 90 0 0 Dout[8]
port 5 nsew
flabel metal2 s 5037 5097 5043 5103 3 FreeSans 16 90 0 0 Dout[7]
port 6 nsew
flabel metal3 s 5116 4196 5124 4204 3 FreeSans 16 0 0 0 Dout[6]
port 7 nsew
flabel metal3 s 5116 3956 5124 3964 3 FreeSans 16 0 0 0 Dout[5]
port 8 nsew
flabel metal3 s 5116 3716 5124 3724 3 FreeSans 16 0 0 0 Dout[4]
port 9 nsew
flabel metal3 s 5116 3476 5124 3484 3 FreeSans 16 0 0 0 Dout[3]
port 10 nsew
flabel metal3 s 5116 3296 5124 3304 3 FreeSans 16 0 0 0 Dout[2]
port 11 nsew
flabel metal3 s 5116 3256 5124 3264 3 FreeSans 16 0 0 0 Dout[1]
port 12 nsew
flabel metal3 s 5116 3216 5124 3224 3 FreeSans 16 0 0 0 Dout[0]
port 13 nsew
flabel metal3 s -24 4916 -16 4924 7 FreeSans 16 0 0 0 ISin
port 14 nsew
flabel metal3 s -24 3056 -16 3064 7 FreeSans 16 0 0 0 Rdy
port 15 nsew
flabel metal2 s 3477 5097 3483 5103 3 FreeSans 16 90 0 0 Vld
port 16 nsew
flabel metal2 s 3037 -23 3043 -17 7 FreeSans 16 270 0 0 Xin[1]
port 17 nsew
flabel metal2 s 3077 -23 3083 -17 7 FreeSans 16 270 0 0 Xin[0]
port 18 nsew
flabel metal2 s 3557 -23 3563 -17 7 FreeSans 16 270 0 0 Yin[1]
port 19 nsew
flabel metal2 s 3597 -23 3603 -17 7 FreeSans 16 270 0 0 Yin[0]
port 20 nsew
flabel metal3 s -24 3016 -16 3024 7 FreeSans 16 0 0 0 clk
port 21 nsew
flabel metal2 s 4957 -23 4963 -17 7 FreeSans 16 270 0 0 selSign
port 22 nsew
flabel metal2 s 4637 -23 4643 -17 7 FreeSans 16 270 0 0 selXY
port 23 nsew
<< properties >>
string FIXED_BBOX -40 -40 5120 5100
<< error_p >>
rect 2753 1593 2767 1607
<< end >>