/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module output_terminal(
    inout vdd,
    inout gnd,
    output [11:0] Dout,
    input ISin,
    input Rdy,
    output Vld,
    input [1:0] Xin,
    input [1:0] Yin,
    input clk,
    input selSign,
    input selXY
);

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire [6:0] LoadCtl ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire ISin ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _256_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _48_ ;
wire _121_ ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire _118_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire _212_ ;
wire _250_ ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire ISreg_bF$buf0 ;
wire ISreg_bF$buf1 ;
wire ISreg_bF$buf2 ;
wire ISreg_bF$buf3 ;
wire ISreg_bF$buf4 ;
wire _80_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _147_ ;
wire _185_ ;
wire selXY ;
wire selSign ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire [11:0] Ycalc ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _96__bF$buf0 ;
wire _96__bF$buf1 ;
wire _96__bF$buf2 ;
wire _96__bF$buf3 ;
wire _96__bF$buf4 ;
wire _138_ ;
wire _30_ ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire ISreg ;
wire _264_ ;
wire [11:0] Dout ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire [11:4] Xin12b ;
wire [1:0] Yin ;
wire _255_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire [11:0] Xcalc ;
wire [1:0] Yin0 ;
wire [1:0] Yin1 ;
wire _214_ ;
wire _252_ ;
wire _117_ ;
wire _155_ ;
wire _193_ ;
wire _249_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire [1:0] Xin0 ;
wire [1:0] Xin1 ;
wire _114_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire _146_ ;
wire _184_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire [11:0] _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire LoadCtl_6_bF$buf0 ;
wire LoadCtl_6_bF$buf1 ;
wire LoadCtl_6_bF$buf2 ;
wire LoadCtl_6_bF$buf3 ;
wire LoadCtl_6_bF$buf4 ;
wire _119_ ;
wire _11_ ;
wire [11:4] Yin12b ;
wire _157_ ;
wire _195_ ;
wire _5_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _116_ ;
wire _154_ ;
wire _192_ ;
wire _248_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire [1:0] Xin ;
wire _245_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

FILL FILL_2__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _588_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_39_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[4])
);

FILL FILL_1__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[6]),
    .B(Xin12b[7]),
    .Y(_145_)
);

FILL FILL_5__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_242_),
    .C(_219_),
    .Y(_245_)
);

FILL FILL_4__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .B(_80_),
    .Y(_83_)
);

FILL FILL_7__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_251_),
    .C(_268_),
    .Y(_46_)
);

FILL FILL_5__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _606_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Rdy),
    .CLK(clk_bF$buf5),
    .Q(LoadCtl[0])
);

FILL FILL_4__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf1),
    .B(Xin12b[10]),
    .C(_160_),
    .Y(_161_)
);

FILL FILL_4__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[0]),
    .B(Yin1[1]),
    .Y(_193_)
);

FILL FILL_4__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf3),
    .B(Yin12b[10]),
    .Y(_242_)
);

FILL FILL_4__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .B(_80_),
    .Y(_81_)
);

FILL FILL_1__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

FILL FILL_5__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .B(_251_),
    .Y(_267_)
);

FILL FILL_1__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf2),
    .B(_108_),
    .C(_109_),
    .Y(_11_)
);

FILL FILL_4__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _585_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .CLK(clk_bF$buf1),
    .Q(Xin12b[9])
);

FILL FILL_2__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf3),
    .B(_139_),
    .C(_142_),
    .Y(_143_)
);

FILL FILL_5__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf0),
    .B(_222_),
    .C(_223_),
    .Y(_29_)
);

FILL FILL_2__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[8]),
    .Y(_65_)
);

FILL FILL_2__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _603_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf5),
    .Q(Yin1[1])
);

FILL FILL_4__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_145_),
    .Y(_158_)
);

FILL FILL_4__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(Yin1[1]),
    .Y(_191_)
);

FILL FILL_5__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[11]),
    .B(_169_),
    .Y(_239_)
);

FILL FILL_4__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[4]),
    .Y(_78_)
);

FILL FILL_7__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_95_),
    .C(_265_),
    .Y(_43_)
);

FILL FILL_4__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_106_),
    .C(_103_),
    .Y(_107_)
);

FILL FILL_4__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_153_),
    .C(_96__bF$buf3),
    .Y(_156_)
);

FILL FILL_1__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _582_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[10])
);

FILL FILL_2__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[7]),
    .Y(_140_)
);

FILL FILL_5__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_53_),
    .B(LoadCtl_6_bF$buf4),
    .C(_188_),
    .Y(_23_)
);

FILL FILL_4__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_219_),
    .Y(_221_)
);

FILL FILL_2__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[7]),
    .Y(_63_)
);

FILL FILL_2__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _579_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[9])
);

FILL FILL_1__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[7]),
    .Y(_137_)
);

FILL FILL_3__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _600_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[4])
);

FILL FILL_8__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[11]),
    .B(_96__bF$buf1),
    .Y(_236_)
);

FILL FILL_4__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(LoadCtl[3]),
    .C(_75_),
    .Y(_76_)
);

FILL FILL_7__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[1]),
    .Y(_264_)
);

FILL FILL_5__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73050x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin0[0]),
    .B(Xin0[1]),
    .C(ISreg_bF$buf1),
    .Y(_104_)
);

FILL FILL_5__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[9]),
    .Y(_153_)
);

FILL FILL_4__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .B(Yin0[1]),
    .Y(_186_)
);

FILL FILL_4__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .Y(_73_)
);

FILL FILL_3_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_217_),
    .Y(_218_)
);

FILL FILL_2__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_80_),
    .C(_262_),
    .Y(_40_)
);

FILL FILL_1__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[6]),
    .Y(_61_)
);

FILL FILL_6__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[1]),
    .B(_96__bF$buf4),
    .Y(_102_)
);

FILL FILL_1__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _576_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .CLK(clk_bF$buf4),
    .Q(Ycalc[6])
);

FILL FILL_1__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(_134_),
    .Y(_135_)
);

FILL FILL_2__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_63_),
    .B(LoadCtl_6_bF$buf2),
    .C(_215_),
    .Y(_28_)
);

FILL FILL_2__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[5]),
    .Y(_59_)
);

FILL FILL_1__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_233_),
    .Y(_234_)
);

FILL FILL_1__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[8]),
    .B(_96__bF$buf1),
    .Y(_151_)
);

FILL FILL_4__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[0]),
    .Y(_183_)
);

FILL FILL_5__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[11]),
    .Y(_71_)
);

FILL FILL_1__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(_80_),
    .Y(_261_)
);

FILL FILL_4__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin0[1]),
    .Y(_99_)
);

FILL FILL_5__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _573_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf0),
    .Q(Ycalc[3])
);

FILL FILL_5__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[6]),
    .Y(_132_)
);

FILL FILL_2__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_93_),
    .C(_91_),
    .Y(_181_)
);

FILL FILL_4__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf4),
    .B(Yin12b[6]),
    .Y(_213_)
);

FILL FILL_5__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[4]),
    .Y(_57_)
);

FILL FILL_2__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[4]),
    .B(Xin12b[5]),
    .Y(_129_)
);

FILL FILL_2__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_144_),
    .Y(_148_)
);

FILL FILL_7__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[10]),
    .Y(_69_)
);

FILL FILL_7__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_76_),
    .C(_259_),
    .Y(_37_)
);

FILL FILL_4__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[0]),
    .B(_96__bF$buf4),
    .Y(_97_)
);

FILL FILL_5__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _570_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf3),
    .Q(Ycalc[0])
);

FILL FILL_5__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .B(LoadCtl_6_bF$buf0),
    .Y(_179_)
);

FILL FILL_4__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73050x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_203_),
    .C(_197_),
    .Y(_210_)
);

FILL FILL_5__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[9]),
    .B(_255_),
    .Y(_258_)
);

FILL FILL_1__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[3]),
    .Y(_55_)
);

FILL FILL_2__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf1),
    .B(_93_),
    .C(_94_),
    .Y(_8_)
);

FILL FILL_1__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _567_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[9])
);

FILL FILL_1__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_125_),
    .Y(_127_)
);

FILL FILL_2__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[2]),
    .Y(_53_)
);

FILL FILL_1__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[9]),
    .Y(_67_)
);

FILL FILL_7__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[8]),
    .Y(Dout[8])
);

FILL FILL_4__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_176_),
    .Y(_177_)
);

FILL FILL_4__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_207_),
    .Y(_208_)
);

FILL FILL_5__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[8]),
    .B(_255_),
    .Y(_256_)
);

FILL FILL_1__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_91_),
    .C(_92_),
    .Y(_7_)
);

FILL FILL_8__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _564_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf5),
    .Q(Xcalc[6])
);

FILL FILL75750x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[4]),
    .B(_116_),
    .C(ISreg_bF$buf1),
    .Y(_124_)
);

FILL FILL_5__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_173_),
    .C(_163_),
    .Y(_174_)
);

FILL FILL_4__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf4),
    .B(Yin12b[6]),
    .C(_204_),
    .Y(_205_)
);

FILL FILL_4__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[1]),
    .Y(_51_)
);

FILL FILL_1__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _599_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[7])
);

FILL FILL_1__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[5]),
    .Y(Dout[5])
);

FILL FILL_2__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_251_),
    .C(_253_),
    .Y(_34_)
);

FILL FILL_4__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_89_),
    .C(_90_),
    .Y(_6_)
);

FILL FILL_8__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _561_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[3])
);

FILL FILL_5__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[2]),
    .Y(Dout[2])
);

FILL FILL_1__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[4]),
    .B(_96__bF$buf4),
    .Y(_122_)
);

FILL FILL_5__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_170_),
    .Y(_171_)
);

FILL FILL_4__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_96__bF$buf1),
    .C(_201_),
    .D(_202_),
    .Y(_26_)
);

FILL FILL_4__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[0]),
    .Y(_49_)
);

FILL FILL_2__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_86_),
    .C(_88_),
    .Y(_5_)
);

FILL FILL_1__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _558_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[0])
);

FILL FILL_1__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .B(_115_),
    .Y(_119_)
);

FILL FILL_4__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _596_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_47_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[8])
);

FILL FILL_1__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf1)
);

FILL FILL_4__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf3),
    .B(_230_),
    .Y(_233_)
);

FILL FILL_1__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(_251_),
    .Y(_252_)
);

FILL FILL_8__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[1]),
    .Y(Dout[1])
);

FILL FILL_4__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .B(_167_),
    .Y(_168_)
);

FILL FILL_4__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_78_),
    .C(_195_),
    .Y(_200_)
);

FILL FILL_5__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_248_),
    .Y(_249_)
);

FILL FILL_1__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[0]),
    .Y(_87_)
);

FILL FILL_4_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[6]),
    .B(_76_),
    .Y(_271_)
);

FILL FILL_4__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .B(_115_),
    .Y(_116_)
);

FILL FILL_4__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _593_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_44_),
    .CLK(clk_bF$buf2),
    .Q(Xin0[1])
);

FILL FILL_2__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_197_),
    .C(_78_),
    .Y(_198_)
);

FILL FILL_4__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_197_),
    .C(_228_),
    .Y(_230_)
);

FILL FILL_1__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_146_),
    .C(ISreg_bF$buf2),
    .Y(_147_)
);

FILL FILL_2__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _611_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[4]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[5])
);

FILL FILL_8__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(LoadCtl_6_bF$buf4),
    .C(_165_),
    .Y(_19_)
);

FILL FILL_7__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf2),
    .B(_246_),
    .C(_243_),
    .Y(_247_)
);

FILL FILL_4__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .Y(_84_)
);

FILL FILL_7__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_255_),
    .C(_269_),
    .Y(_47_)
);

FILL FILL_4__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _608_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[1]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[2])
);

FILL FILL_4__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[3]),
    .B(_96__bF$buf1),
    .Y(_114_)
);

FILL FILL_5__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf2),
    .B(_160_),
    .Y(_163_)
);

FILL FILL_1__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _590_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_41_),
    .CLK(clk_bF$buf5),
    .Q(Xin1[0])
);

FILL FILL_5__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf3),
    .B(_194_),
    .Y(_195_)
);

FILL FILL_4__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .B(_96__bF$buf0),
    .C(_226_),
    .D(_227_),
    .Y(_30_)
);

FILL FILL_2__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .B(_251_),
    .Y(_268_)
);

FILL FILL_1__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin1[1]),
    .B(_110_),
    .Y(_111_)
);

FILL FILL_4__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _587_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .CLK(clk_bF$buf1),
    .Q(Xin12b[7])
);

FILL FILL74850x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73350x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[8]),
    .Y(_144_)
);

FILL FILL_5__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_65_),
    .C(_66_),
    .Y(_272_[8])
);

FILL FILL_2__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .C(ISreg_bF$buf4),
    .Y(_244_)
);

FILL FILL_8__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[5]),
    .Y(_82_)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_96__bF$buf4)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_96__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_96__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_96__bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_96__bF$buf0)
);

FILL FILL_7__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _605_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf3),
    .Q(Yin0[1])
);

FILL FILL_4__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_119_),
    .C(_158_),
    .Y(_160_)
);

FILL FILL_4__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(LoadCtl_6_bF$buf4),
    .C(_192_),
    .Y(_24_)
);

FILL FILL_4__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .Y(_241_)
);

FILL FILL_4__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(_79_),
    .Y(_80_)
);

FILL FILL_1__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_216_),
    .C(_219_),
    .Y(_225_)
);

FILL FILL_5__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_99_),
    .C(_266_),
    .Y(_44_)
);

FILL FILL_1__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[2]),
    .B(_96__bF$buf2),
    .Y(_109_)
);

FILL FILL_4__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _584_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .CLK(clk_bF$buf5),
    .Q(Xin12b[8])
);

FILL FILL_2__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_141_),
    .C(_133_),
    .Y(_142_)
);

FILL FILL_5__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[1]),
    .B(_189_),
    .Y(_190_)
);

FILL FILL_4__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Ycalc[8]),
    .B(_96__bF$buf0),
    .Y(_223_)
);

FILL FILL_2__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_63_),
    .C(_64_),
    .Y(_272_[7])
);

FILL FILL_2__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _602_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf5),
    .Q(Yin1[0])
);

FILL FILL_4__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[10]),
    .Y(_157_)
);

FILL FILL_7__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .B(_237_),
    .Y(_238_)
);

FILL FILL_4__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_76_),
    .C(_77_),
    .Y(_1_)
);

FILL FILL_7__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(Xin[0]),
    .Y(_265_)
);

FILL FILL_4__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin0[0]),
    .B(Xin0[1]),
    .Y(_106_)
);

FILL FILL_4__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_153_),
    .Y(_155_)
);

FILL FILL_4__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _581_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[11])
);

FILL FILL_5__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf0),
    .B(Xin12b[7]),
    .C(_138_),
    .Y(_139_)
);

FILL FILL_5__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf0),
    .B(_187_),
    .C(_185_),
    .Y(_188_)
);

FILL FILL_4__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_216_),
    .Y(_220_)
);

FILL FILL_2__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_61_),
    .C(_62_),
    .Y(_272_[6])
);

FILL FILL_2__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin1[0]),
    .Y(_103_)
);

FILL FILL_1__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _578_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[8])
);

FILL FILL_1__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf3),
    .B(_135_),
    .C(_136_),
    .Y(_15_)
);

FILL FILL_2__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(LoadCtl_6_bF$buf2),
    .C(_235_),
    .Y(_31_)
);

FILL FILL_4__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(LoadCtl[1]),
    .Y(_75_)
);

FILL FILL75150x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_86_),
    .C(_263_),
    .Y(_41_)
);

FILL FILL_5__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[9]),
    .Y(_152_)
);

FILL FILL_4__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_183_),
    .Y(_185_)
);

FILL FILL_4__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_71_),
    .C(_72_),
    .Y(_272_[11])
);

FILL FILL_1__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[6]),
    .B(Yin12b[7]),
    .Y(_217_)
);

FILL FILL_5__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(_80_),
    .Y(_262_)
);

FILL FILL75450x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(_59_),
    .C(_60_),
    .Y(_272_[5])
);

FILL FILL_6__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_100_),
    .Y(_101_)
);

FILL FILL_1__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _575_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[5])
);

FILL FILL_5__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_133_),
    .Y(_134_)
);

FILL FILL_2__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf1),
    .B(_211_),
    .C(_214_),
    .Y(_215_)
);

FILL FILL_3__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(_57_),
    .C(_58_),
    .Y(_272_[4])
);

FILL FILL_1__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_148_),
    .Y(_150_)
);

FILL FILL_4__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .B(LoadCtl_6_bF$buf4),
    .C(_182_),
    .Y(_22_)
);

FILL FILL_5__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_69_),
    .C(_70_),
    .Y(_272_[10])
);

FILL FILL_7__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_76_),
    .C(_260_),
    .Y(_38_)
);

FILL FILL_4__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf1),
    .B(Xin0[0]),
    .C(Xin0[1]),
    .Y(_98_)
);

FILL FILL_5__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _572_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf0),
    .Q(Ycalc[2])
);

FILL FILL73950x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf0),
    .B(Xin12b[6]),
    .C(_130_),
    .Y(_131_)
);

FILL FILL_5__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf2),
    .Y(_180_)
);

FILL FILL_4__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[7]),
    .Y(_212_)
);

FILL FILL_5__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(_55_),
    .C(_56_),
    .Y(_272_[3])
);

FILL FILL_2__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _569_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf2),
    .Q(Xcalc[11])
);

FILL FILL_1__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf2),
    .B(_127_),
    .C(_128_),
    .Y(_14_)
);

FILL FILL_2__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(_67_),
    .C(_68_),
    .Y(_272_[9])
);

FILL FILL_7__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[6]),
    .B(_76_),
    .Y(_259_)
);

FILL FILL_8__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf4),
    .Y(_96_)
);

FILL FILL_5__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf2),
    .Y(Vld)
);

FILL FILL_4__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_178_),
    .Y(_20_)
);

FILL FILL_4__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(LoadCtl_6_bF$buf1),
    .C(_209_),
    .Y(_27_)
);

FILL FILL_5__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .Y(_257_)
);

FILL FILL_1__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_53_),
    .C(_54_),
    .Y(_272_[2])
);

FILL FILL_8__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISin),
    .B(LoadCtl_6_bF$buf1),
    .Y(_94_)
);

FILL FILL_1__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _566_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf6),
    .Q(Xcalc[8])
);

FILL FILL_1__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_124_),
    .Y(_126_)
);

FILL FILL_2__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf4),
    .B(_204_),
    .Y(_207_)
);

FILL FILL_4__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_51_),
    .C(_52_),
    .Y(_272_[1])
);

FILL FILL_1__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[7]),
    .Y(Dout[7])
);

FILL FILL_4__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_173_),
    .C(_147_),
    .Y(_176_)
);

FILL FILL_1__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .B(_249_),
    .Y(_255_)
);

FILL FILL_4__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(Yin[1]),
    .Y(_92_)
);

FILL FILL_8__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _563_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[5])
);

FILL FILL_4__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[4]),
    .Y(Dout[4])
);

FILL FILL_1__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[5]),
    .Y(_123_)
);

FILL FILL_5__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf2),
    .B(Xin12b[10]),
    .Y(_173_)
);

FILL FILL_4__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_197_),
    .Y(_204_)
);

FILL FILL_2_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(_49_),
    .C(_50_),
    .Y(_272_[0])
);

FILL FILL_2__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73050x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_120_),
    .Y(_121_)
);

FILL FILL_4__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _598_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[6])
);

FILL FILL_1__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(_251_),
    .Y(_253_)
);

FILL FILL_4__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(Yin[0]),
    .Y(_90_)
);

FILL FILL_1__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _560_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[2])
);

FILL FILL_5__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[11]),
    .Y(Dout[11])
);

FILL FILL_1__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[11]),
    .B(_169_),
    .Y(_170_)
);

FILL FILL_4__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_82_),
    .C(_96__bF$buf1),
    .Y(_202_)
);

FILL FILL_4__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .B(_250_),
    .Y(_251_)
);

FILL FILL_1__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Yin1[1]),
    .Y(_88_)
);

FILL FILL_1__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _557_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf4),
    .Q(ISreg)
);

FILL FILL_1__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[4]),
    .Y(_118_)
);

FILL FILL_4__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _595_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_46_),
    .CLK(clk_bF$buf2),
    .Q(Yin12b[11])
);

FILL FILL_2__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[10]),
    .Y(_232_)
);

FILL FILL_1__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73350x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[0]),
    .Y(Dout[0])
);

FILL FILL_4__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[11]),
    .Y(_167_)
);

FILL FILL_4__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(LoadCtl_6_bF$buf0),
    .C(_199_),
    .Y(_25_)
);

FILL FILL_5__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(LoadCtl[3]),
    .Y(_248_)
);

FILL FILL_1__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(LoadCtl[0]),
    .Y(_86_)
);

FILL FILL_4_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_255_),
    .C(_270_),
    .Y(_48_)
);

FILL FILL_4__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin1[0]),
    .B(Xin1[1]),
    .Y(_115_)
);

FILL FILL_4__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf3),
    .B(_161_),
    .C(_164_),
    .Y(_165_)
);

FILL FILL_1__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _592_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_43_),
    .CLK(clk_bF$buf2),
    .Q(Xin0[0])
);

FILL FILL_2__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_193_),
    .Y(_197_)
);

FILL FILL_4__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[8]),
    .B(Yin12b[9]),
    .Y(_229_)
);

FILL FILL_2__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _589_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_40_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[5])
);

FILL FILL_1__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_145_),
    .Y(_146_)
);

FILL FILL_3__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _610_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[3]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[4])
);

FILL FILL_8__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_245_),
    .Y(_246_)
);

FILL FILL_4__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_80_),
    .C(_83_),
    .Y(_3_)
);

FILL FILL_7__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[8]),
    .B(_255_),
    .Y(_269_)
);

FILL FILL_5__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _607_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[0]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[1])
);

FILL FILL_4__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_112_),
    .Y(_113_)
);

FILL FILL_5__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[10]),
    .Y(_162_)
);

FILL FILL_1__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_193_),
    .Y(_194_)
);

FILL FILL_4__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_80_),
    .C(_81_),
    .Y(_2_)
);

FILL FILL_1__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_224_),
    .C(_96__bF$buf0),
    .Y(_227_)
);

FILL FILL_2__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_251_),
    .C(_267_),
    .Y(_45_)
);

FILL FILL_1__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_103_),
    .C(_104_),
    .Y(_110_)
);

FILL FILL_4__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _586_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .CLK(clk_bF$buf5),
    .Q(Xin12b[6])
);

FILL FILL_1__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(LoadCtl_6_bF$buf3),
    .C(_143_),
    .Y(_16_)
);

FILL FILL_5__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[9]),
    .Y(_224_)
);

FILL FILL_1__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(Xcalc[8]),
    .Y(_66_)
);

FILL FILL_2__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_242_),
    .C(_233_),
    .Y(_243_)
);

FILL FILL_8__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg),
    .Y(ISreg_bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg),
    .Y(ISreg_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg),
    .Y(ISreg_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg),
    .Y(ISreg_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg),
    .Y(ISreg_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf4)
);

FILL FILL_7__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[6]),
    .Y(LoadCtl_6_bF$buf1)
);

FILL FILL_1__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _604_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf3),
    .Q(Yin0[0])
);

FILL FILL_4__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .Y(_159_)
);

FILL FILL_4__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf0),
    .B(_190_),
    .C(_191_),
    .Y(_192_)
);

FILL FILL_5__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_239_),
    .Y(_240_)
);

FILL FILL_4__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .Y(_79_)
);

FILL FILL_1__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(Xin[1]),
    .Y(_266_)
);

FILL FILL73650x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_105_),
    .Y(_108_)
);

FILL FILL_4__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _583_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .CLK(clk_bF$buf2),
    .Q(Xin12b[11])
);

FILL FILL_2__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf0),
    .B(Xin12b[6]),
    .Y(_141_)
);

FILL FILL_5__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_183_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_4__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_220_),
    .Y(_222_)
);

FILL FILL_2__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(Xcalc[7]),
    .Y(_64_)
);

FILL FILL_2__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_129_),
    .C(_119_),
    .Y(_138_)
);

FILL FILL_2__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _601_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[5])
);

FILL FILL_8__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_96__bF$buf3),
    .C(_155_),
    .D(_156_),
    .Y(_18_)
);

FILL FILL_7__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[11]),
    .Y(_237_)
);

FILL FILL_4__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[7]),
    .B(_76_),
    .Y(_77_)
);

FILL FILL_7__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_86_),
    .C(_264_),
    .Y(_42_)
);

FILL FILL_4__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_103_),
    .Y(_105_)
);

FILL FILL_5__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_144_),
    .C(_147_),
    .Y(_154_)
);

FILL FILL_4__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _580_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[10])
);

FILL FILL_5__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_186_),
    .C(_183_),
    .Y(_187_)
);

FILL FILL_4__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_218_),
    .C(ISreg_bF$buf3),
    .Y(_219_)
);

FILL FILL_2__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .B(_85_),
    .C(Xin1[0]),
    .Y(_263_)
);

FILL FILL_1__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf1),
    .B(Xcalc[6]),
    .Y(_62_)
);

FILL FILL_2__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf4),
    .B(_101_),
    .C(_102_),
    .Y(_10_)
);

FILL FILL_1__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _577_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[7])
);

FILL FILL_1__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[6]),
    .B(_96__bF$buf3),
    .Y(_136_)
);

FILL FILL_2__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL72750x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(Xcalc[5]),
    .Y(_60_)
);

FILL FILL_1__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf2),
    .B(_231_),
    .C(_234_),
    .Y(_235_)
);

FILL FILL_1__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .Y(_74_)
);

FILL FILL_7__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf0),
    .B(_150_),
    .C(_151_),
    .Y(_17_)
);

FILL FILL_4__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .B(Yin0[1]),
    .C(ISreg_bF$buf2),
    .Y(_184_)
);

FILL FILL_4__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(Xcalc[11]),
    .Y(_72_)
);

FILL FILL_1__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[8]),
    .Y(_216_)
);

FILL FILL_5__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_80_),
    .C(_261_),
    .Y(_39_)
);

FILL FILL_1__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_95_),
    .C(_99_),
    .Y(_100_)
);

FILL FILL_4__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _574_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf6),
    .Q(Ycalc[4])
);

FILL FILL_5__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf0),
    .B(_130_),
    .Y(_133_)
);

FILL FILL_2__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf3),
    .B(_180_),
    .C(_181_),
    .Y(_182_)
);

FILL FILL_4__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_213_),
    .C(_207_),
    .Y(_214_)
);

FILL FILL75450x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(Xcalc[4]),
    .Y(_58_)
);

FILL FILL_1__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_147_),
    .Y(_149_)
);

FILL FILL_7__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf2),
    .B(Xcalc[10]),
    .Y(_70_)
);

FILL FILL_7__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[7]),
    .B(_76_),
    .Y(_260_)
);

FILL FILL_4__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_96__bF$buf2),
    .C(_97_),
    .Y(_9_)
);

FILL FILL_5__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _571_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf3),
    .Q(Ycalc[1])
);

FILL FILL_5__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_119_),
    .Y(_130_)
);

FILL FILL_5__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf4),
    .B(_49_),
    .C(_179_),
    .Y(_21_)
);

FILL FILL_4__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf4),
    .B(Yin12b[7]),
    .C(_210_),
    .Y(_211_)
);

FILL FILL_5__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(Xcalc[3]),
    .Y(_56_)
);

FILL FILL_2__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin0[0]),
    .Y(_95_)
);

FILL FILL_1__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _568_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf3),
    .Q(Xcalc[10])
);

FILL FILL_1__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[5]),
    .B(_96__bF$buf2),
    .Y(_128_)
);

FILL FILL_2__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf0),
    .B(Xcalc[9]),
    .Y(_68_)
);

FILL FILL_7__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_255_),
    .C(_258_),
    .Y(_36_)
);

FILL FILL_8__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL72750x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[9]),
    .Y(Dout[9])
);

FILL FILL73350x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf3),
    .B(_177_),
    .C(_174_),
    .Y(_178_)
);

FILL FILL_4__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf1),
    .B(_205_),
    .C(_208_),
    .Y(_209_)
);

FILL FILL_5__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_255_),
    .C(_256_),
    .Y(_35_)
);

FILL FILL_1__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(Xcalc[2]),
    .Y(_54_)
);

FILL FILL_8__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf4),
    .Y(_93_)
);

FILL FILL_1__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _565_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[7])
);

FILL FILL_4__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_123_),
    .Y(_125_)
);

FILL FILL_5__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[6]),
    .Y(_206_)
);

FILL FILL_4__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selXY_bF$buf3),
    .B(Xcalc[1]),
    .Y(_52_)
);

FILL FILL73950x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[6]),
    .Y(Dout[6])
);

FILL FILL_7__273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin12b[8]),
    .B(Xin12b[9]),
    .C(ISreg_bF$buf0),
    .Y(_175_)
);

FILL FILL_1__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .Y(_254_)
);

FILL FILL_4__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[1]),
    .Y(_91_)
);

FILL FILL_8__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _562_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[4])
);

FILL FILL_4__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[3]),
    .Y(Dout[3])
);

FILL FILL_1__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf4),
    .B(_121_),
    .C(_122_),
    .Y(_13_)
);

FILL FILL_5__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .Y(_172_)
);

FILL FILL_4__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[4]),
    .B(Yin12b[5]),
    .Y(_203_)
);

FILL FILL_4__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[0]),
    .B(selXY_bF$buf0),
    .Y(_50_)
);

FILL FILL_2__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _559_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf0),
    .Q(Xcalc[1])
);

FILL FILL_1__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_119_),
    .C(_118_),
    .Y(_120_)
);

FILL FILL_4__296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _597_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_48_),
    .CLK(clk_bF$buf4),
    .Q(Yin12b[9])
);

FILL FILL75450x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_251_),
    .C(_252_),
    .Y(_33_)
);

FILL FILL_8__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .Y(_89_)
);

FILL FILL_1__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_[10]),
    .Y(Dout[10])
);

FILL FILL_4__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__289_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(selSign),
    .Y(_169_)
);

FILL FILL_4__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_82_),
    .Y(_201_)
);

FILL FILL_2_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[5]),
    .B(_249_),
    .Y(_250_)
);

FILL FILL73350x72150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_86_),
    .C(_87_),
    .Y(_4_)
);

FILL FILL_1__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__277_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_76_),
    .C(_271_),
    .Y(_0_)
);

FILL FILL_1__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf1),
    .B(Xin12b[4]),
    .C(_116_),
    .Y(_117_)
);

FILL FILL_4__293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _594_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_45_),
    .CLK(clk_bF$buf3),
    .Q(Yin12b[10])
);

FILL FILL_2__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_6_bF$buf0),
    .B(_198_),
    .C(_196_),
    .Y(_199_)
);

FILL FILL_4__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ISreg_bF$buf3),
    .B(Yin12b[10]),
    .C(_230_),
    .Y(_231_)
);

FILL FILL_1__281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__298_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_7__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _612_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[5]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[6])
);

FILL FILL_4__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xcalc[11]),
    .B(_96__bF$buf4),
    .Y(_166_)
);

FILL FILL74550x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_247_),
    .Y(_32_)
);

FILL FILL_4__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[1]),
    .Y(_85_)
);

FILL FILL_7__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__308_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin12b[9]),
    .B(_255_),
    .Y(_270_)
);

FILL FILL_4__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _609_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[2]),
    .CLK(clk_bF$buf1),
    .Q(LoadCtl[3])
);

FILL FILL_4__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96__bF$buf3),
    .B(_113_),
    .C(_114_),
    .Y(_12_)
);

FILL FILL_4__290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_163_),
    .Y(_164_)
);

FILL FILL_1__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _591_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_42_),
    .CLK(clk_bF$buf5),
    .Q(Xin1[1])
);

FILL FILL_5__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_78_),
    .Y(_196_)
);

FILL FILL_4__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_217_),
    .Y(_228_)
);

FILL FILL_2__312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(Xin1[1]),
    .Y(_112_)
);

FILL FILL_4__287_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule
