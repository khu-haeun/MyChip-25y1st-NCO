magic
tech scmos
magscale 1 3
timestamp 1569533753
<< checkpaint >>
rect -64 -64 64 64
<< gv2 >>
rect -4 -4 4 4
<< end >>
