magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect 8700 8700 29300 29320
<< metal1 >>
rect 11840 28719 26820 28720
rect 9961 28696 26820 28719
rect 9961 28680 9980 28696
rect 9996 28680 10012 28696
rect 10028 28680 10044 28696
rect 10060 28680 10076 28696
rect 10092 28680 10108 28696
rect 10124 28680 10140 28696
rect 10156 28680 10172 28696
rect 10188 28680 10204 28696
rect 10220 28680 10236 28696
rect 10252 28680 10268 28696
rect 10284 28680 10300 28696
rect 10316 28680 10332 28696
rect 10348 28680 10364 28696
rect 10380 28680 10396 28696
rect 10412 28680 10428 28696
rect 10444 28680 10460 28696
rect 10476 28680 10492 28696
rect 10508 28680 10524 28696
rect 10540 28680 10556 28696
rect 10572 28680 10588 28696
rect 10604 28680 10620 28696
rect 10636 28680 10652 28696
rect 10668 28680 10684 28696
rect 10700 28680 10716 28696
rect 10732 28680 10748 28696
rect 10764 28680 10780 28696
rect 10796 28680 10812 28696
rect 10828 28680 10844 28696
rect 10860 28680 10876 28696
rect 10892 28680 10908 28696
rect 10924 28680 10940 28696
rect 10956 28680 10972 28696
rect 10988 28680 11004 28696
rect 11020 28680 11036 28696
rect 11052 28680 11068 28696
rect 11084 28680 11100 28696
rect 11116 28680 11132 28696
rect 11148 28680 11164 28696
rect 11180 28680 11196 28696
rect 11212 28680 11228 28696
rect 11244 28680 11260 28696
rect 11276 28680 11292 28696
rect 11308 28680 11324 28696
rect 11340 28680 11356 28696
rect 11372 28680 11388 28696
rect 11404 28680 11420 28696
rect 11436 28680 11452 28696
rect 11468 28680 11484 28696
rect 11500 28680 11516 28696
rect 11532 28680 11548 28696
rect 11564 28680 11580 28696
rect 11596 28680 11612 28696
rect 11628 28680 11644 28696
rect 11660 28680 11676 28696
rect 11692 28680 11708 28696
rect 11724 28680 11740 28696
rect 11756 28680 11772 28696
rect 11788 28680 11804 28696
rect 11820 28680 26820 28696
rect 9961 28664 26820 28680
rect 9961 28648 9980 28664
rect 9996 28648 10012 28664
rect 10028 28648 10044 28664
rect 10060 28648 10076 28664
rect 10092 28648 10108 28664
rect 10124 28648 10140 28664
rect 10156 28648 10172 28664
rect 10188 28648 10204 28664
rect 10220 28648 10236 28664
rect 10252 28648 10268 28664
rect 10284 28648 10300 28664
rect 10316 28648 10332 28664
rect 10348 28648 10364 28664
rect 10380 28648 10396 28664
rect 10412 28648 10428 28664
rect 10444 28648 10460 28664
rect 10476 28648 10492 28664
rect 10508 28648 10524 28664
rect 10540 28648 10556 28664
rect 10572 28648 10588 28664
rect 10604 28648 10620 28664
rect 10636 28648 10652 28664
rect 10668 28648 10684 28664
rect 10700 28648 10716 28664
rect 10732 28648 10748 28664
rect 10764 28648 10780 28664
rect 10796 28648 10812 28664
rect 10828 28648 10844 28664
rect 10860 28648 10876 28664
rect 10892 28648 10908 28664
rect 10924 28648 10940 28664
rect 10956 28648 10972 28664
rect 10988 28648 11004 28664
rect 11020 28648 11036 28664
rect 11052 28648 11068 28664
rect 11084 28648 11100 28664
rect 11116 28648 11132 28664
rect 11148 28648 11164 28664
rect 11180 28648 11196 28664
rect 11212 28648 11228 28664
rect 11244 28648 11260 28664
rect 11276 28648 11292 28664
rect 11308 28648 11324 28664
rect 11340 28648 11356 28664
rect 11372 28648 11388 28664
rect 11404 28648 11420 28664
rect 11436 28648 11452 28664
rect 11468 28648 11484 28664
rect 11500 28648 11516 28664
rect 11532 28648 11548 28664
rect 11564 28648 11580 28664
rect 11596 28648 11612 28664
rect 11628 28648 11644 28664
rect 11660 28648 11676 28664
rect 11692 28648 11708 28664
rect 11724 28648 11740 28664
rect 11756 28648 11772 28664
rect 11788 28648 11804 28664
rect 11820 28648 26820 28664
rect 9961 28632 26820 28648
rect 9961 28616 9980 28632
rect 9996 28616 10012 28632
rect 10028 28616 10044 28632
rect 10060 28616 10076 28632
rect 10092 28616 10108 28632
rect 10124 28616 10140 28632
rect 10156 28616 10172 28632
rect 10188 28616 10204 28632
rect 10220 28616 10236 28632
rect 10252 28616 10268 28632
rect 10284 28616 10300 28632
rect 10316 28616 10332 28632
rect 10348 28616 10364 28632
rect 10380 28616 10396 28632
rect 10412 28616 10428 28632
rect 10444 28616 10460 28632
rect 10476 28616 10492 28632
rect 10508 28616 10524 28632
rect 10540 28616 10556 28632
rect 10572 28616 10588 28632
rect 10604 28616 10620 28632
rect 10636 28616 10652 28632
rect 10668 28616 10684 28632
rect 10700 28616 10716 28632
rect 10732 28616 10748 28632
rect 10764 28616 10780 28632
rect 10796 28616 10812 28632
rect 10828 28616 10844 28632
rect 10860 28616 10876 28632
rect 10892 28616 10908 28632
rect 10924 28616 10940 28632
rect 10956 28616 10972 28632
rect 10988 28616 11004 28632
rect 11020 28616 11036 28632
rect 11052 28616 11068 28632
rect 11084 28616 11100 28632
rect 11116 28616 11132 28632
rect 11148 28616 11164 28632
rect 11180 28616 11196 28632
rect 11212 28616 11228 28632
rect 11244 28616 11260 28632
rect 11276 28616 11292 28632
rect 11308 28616 11324 28632
rect 11340 28616 11356 28632
rect 11372 28616 11388 28632
rect 11404 28616 11420 28632
rect 11436 28616 11452 28632
rect 11468 28616 11484 28632
rect 11500 28616 11516 28632
rect 11532 28616 11548 28632
rect 11564 28616 11580 28632
rect 11596 28616 11612 28632
rect 11628 28616 11644 28632
rect 11660 28616 11676 28632
rect 11692 28616 11708 28632
rect 11724 28616 11740 28632
rect 11756 28616 11772 28632
rect 11788 28616 11804 28632
rect 11820 28616 26820 28632
rect 9961 28600 26820 28616
rect 9961 28584 9980 28600
rect 9996 28584 10012 28600
rect 10028 28584 10044 28600
rect 10060 28584 10076 28600
rect 10092 28584 10108 28600
rect 10124 28584 10140 28600
rect 10156 28584 10172 28600
rect 10188 28584 10204 28600
rect 10220 28584 10236 28600
rect 10252 28584 10268 28600
rect 10284 28584 10300 28600
rect 10316 28584 10332 28600
rect 10348 28584 10364 28600
rect 10380 28584 10396 28600
rect 10412 28584 10428 28600
rect 10444 28584 10460 28600
rect 10476 28584 10492 28600
rect 10508 28584 10524 28600
rect 10540 28584 10556 28600
rect 10572 28584 10588 28600
rect 10604 28584 10620 28600
rect 10636 28584 10652 28600
rect 10668 28584 10684 28600
rect 10700 28584 10716 28600
rect 10732 28584 10748 28600
rect 10764 28584 10780 28600
rect 10796 28584 10812 28600
rect 10828 28584 10844 28600
rect 10860 28584 10876 28600
rect 10892 28584 10908 28600
rect 10924 28584 10940 28600
rect 10956 28584 10972 28600
rect 10988 28584 11004 28600
rect 11020 28584 11036 28600
rect 11052 28584 11068 28600
rect 11084 28584 11100 28600
rect 11116 28584 11132 28600
rect 11148 28584 11164 28600
rect 11180 28584 11196 28600
rect 11212 28584 11228 28600
rect 11244 28584 11260 28600
rect 11276 28584 11292 28600
rect 11308 28584 11324 28600
rect 11340 28584 11356 28600
rect 11372 28584 11388 28600
rect 11404 28584 11420 28600
rect 11436 28584 11452 28600
rect 11468 28584 11484 28600
rect 11500 28584 11516 28600
rect 11532 28584 11548 28600
rect 11564 28584 11580 28600
rect 11596 28584 11612 28600
rect 11628 28584 11644 28600
rect 11660 28584 11676 28600
rect 11692 28584 11708 28600
rect 11724 28584 11740 28600
rect 11756 28584 11772 28600
rect 11788 28584 11804 28600
rect 11820 28584 26820 28600
rect 9961 28568 26820 28584
rect 9961 28552 9980 28568
rect 9996 28552 10012 28568
rect 10028 28552 10044 28568
rect 10060 28552 10076 28568
rect 10092 28552 10108 28568
rect 10124 28552 10140 28568
rect 10156 28552 10172 28568
rect 10188 28552 10204 28568
rect 10220 28552 10236 28568
rect 10252 28552 10268 28568
rect 10284 28552 10300 28568
rect 10316 28552 10332 28568
rect 10348 28552 10364 28568
rect 10380 28552 10396 28568
rect 10412 28552 10428 28568
rect 10444 28552 10460 28568
rect 10476 28552 10492 28568
rect 10508 28552 10524 28568
rect 10540 28552 10556 28568
rect 10572 28552 10588 28568
rect 10604 28552 10620 28568
rect 10636 28552 10652 28568
rect 10668 28552 10684 28568
rect 10700 28552 10716 28568
rect 10732 28552 10748 28568
rect 10764 28552 10780 28568
rect 10796 28552 10812 28568
rect 10828 28552 10844 28568
rect 10860 28552 10876 28568
rect 10892 28552 10908 28568
rect 10924 28552 10940 28568
rect 10956 28552 10972 28568
rect 10988 28552 11004 28568
rect 11020 28552 11036 28568
rect 11052 28552 11068 28568
rect 11084 28552 11100 28568
rect 11116 28552 11132 28568
rect 11148 28552 11164 28568
rect 11180 28552 11196 28568
rect 11212 28552 11228 28568
rect 11244 28552 11260 28568
rect 11276 28552 11292 28568
rect 11308 28552 11324 28568
rect 11340 28552 11356 28568
rect 11372 28552 11388 28568
rect 11404 28552 11420 28568
rect 11436 28552 11452 28568
rect 11468 28552 11484 28568
rect 11500 28552 11516 28568
rect 11532 28552 11548 28568
rect 11564 28552 11580 28568
rect 11596 28552 11612 28568
rect 11628 28552 11644 28568
rect 11660 28552 11676 28568
rect 11692 28552 11708 28568
rect 11724 28552 11740 28568
rect 11756 28552 11772 28568
rect 11788 28552 11804 28568
rect 11820 28552 26820 28568
rect 9961 28536 26820 28552
rect 9961 28520 9980 28536
rect 9996 28520 10012 28536
rect 10028 28520 10044 28536
rect 10060 28520 10076 28536
rect 10092 28520 10108 28536
rect 10124 28520 10140 28536
rect 10156 28520 10172 28536
rect 10188 28520 10204 28536
rect 10220 28520 10236 28536
rect 10252 28520 10268 28536
rect 10284 28520 10300 28536
rect 10316 28520 10332 28536
rect 10348 28520 10364 28536
rect 10380 28520 10396 28536
rect 10412 28520 10428 28536
rect 10444 28520 10460 28536
rect 10476 28520 10492 28536
rect 10508 28520 10524 28536
rect 10540 28520 10556 28536
rect 10572 28520 10588 28536
rect 10604 28520 10620 28536
rect 10636 28520 10652 28536
rect 10668 28520 10684 28536
rect 10700 28520 10716 28536
rect 10732 28520 10748 28536
rect 10764 28520 10780 28536
rect 10796 28520 10812 28536
rect 10828 28520 10844 28536
rect 10860 28520 10876 28536
rect 10892 28520 10908 28536
rect 10924 28520 10940 28536
rect 10956 28520 10972 28536
rect 10988 28520 11004 28536
rect 11020 28520 11036 28536
rect 11052 28520 11068 28536
rect 11084 28520 11100 28536
rect 11116 28520 11132 28536
rect 11148 28520 11164 28536
rect 11180 28520 11196 28536
rect 11212 28520 11228 28536
rect 11244 28520 11260 28536
rect 11276 28520 11292 28536
rect 11308 28520 11324 28536
rect 11340 28520 11356 28536
rect 11372 28520 11388 28536
rect 11404 28520 11420 28536
rect 11436 28520 11452 28536
rect 11468 28520 11484 28536
rect 11500 28520 11516 28536
rect 11532 28520 11548 28536
rect 11564 28520 11580 28536
rect 11596 28520 11612 28536
rect 11628 28520 11644 28536
rect 11660 28520 11676 28536
rect 11692 28520 11708 28536
rect 11724 28520 11740 28536
rect 11756 28520 11772 28536
rect 11788 28520 11804 28536
rect 11820 28520 26820 28536
rect 9961 28504 26820 28520
rect 9961 28488 9980 28504
rect 9996 28488 10012 28504
rect 10028 28488 10044 28504
rect 10060 28488 10076 28504
rect 10092 28488 10108 28504
rect 10124 28488 10140 28504
rect 10156 28488 10172 28504
rect 10188 28488 10204 28504
rect 10220 28488 10236 28504
rect 10252 28488 10268 28504
rect 10284 28488 10300 28504
rect 10316 28488 10332 28504
rect 10348 28488 10364 28504
rect 10380 28488 10396 28504
rect 10412 28488 10428 28504
rect 10444 28488 10460 28504
rect 10476 28488 10492 28504
rect 10508 28488 10524 28504
rect 10540 28488 10556 28504
rect 10572 28488 10588 28504
rect 10604 28488 10620 28504
rect 10636 28488 10652 28504
rect 10668 28488 10684 28504
rect 10700 28488 10716 28504
rect 10732 28488 10748 28504
rect 10764 28488 10780 28504
rect 10796 28488 10812 28504
rect 10828 28488 10844 28504
rect 10860 28488 10876 28504
rect 10892 28488 10908 28504
rect 10924 28488 10940 28504
rect 10956 28488 10972 28504
rect 10988 28488 11004 28504
rect 11020 28488 11036 28504
rect 11052 28488 11068 28504
rect 11084 28488 11100 28504
rect 11116 28488 11132 28504
rect 11148 28488 11164 28504
rect 11180 28488 11196 28504
rect 11212 28488 11228 28504
rect 11244 28488 11260 28504
rect 11276 28488 11292 28504
rect 11308 28488 11324 28504
rect 11340 28488 11356 28504
rect 11372 28488 11388 28504
rect 11404 28488 11420 28504
rect 11436 28488 11452 28504
rect 11468 28488 11484 28504
rect 11500 28488 11516 28504
rect 11532 28488 11548 28504
rect 11564 28488 11580 28504
rect 11596 28488 11612 28504
rect 11628 28488 11644 28504
rect 11660 28488 11676 28504
rect 11692 28488 11708 28504
rect 11724 28488 11740 28504
rect 11756 28488 11772 28504
rect 11788 28488 11804 28504
rect 11820 28488 26820 28504
rect 9961 28472 26820 28488
rect 9961 28456 9980 28472
rect 9996 28456 10012 28472
rect 10028 28456 10044 28472
rect 10060 28456 10076 28472
rect 10092 28456 10108 28472
rect 10124 28456 10140 28472
rect 10156 28456 10172 28472
rect 10188 28456 10204 28472
rect 10220 28456 10236 28472
rect 10252 28456 10268 28472
rect 10284 28456 10300 28472
rect 10316 28456 10332 28472
rect 10348 28456 10364 28472
rect 10380 28456 10396 28472
rect 10412 28456 10428 28472
rect 10444 28456 10460 28472
rect 10476 28456 10492 28472
rect 10508 28456 10524 28472
rect 10540 28456 10556 28472
rect 10572 28456 10588 28472
rect 10604 28456 10620 28472
rect 10636 28456 10652 28472
rect 10668 28456 10684 28472
rect 10700 28456 10716 28472
rect 10732 28456 10748 28472
rect 10764 28456 10780 28472
rect 10796 28456 10812 28472
rect 10828 28456 10844 28472
rect 10860 28456 10876 28472
rect 10892 28456 10908 28472
rect 10924 28456 10940 28472
rect 10956 28456 10972 28472
rect 10988 28456 11004 28472
rect 11020 28456 11036 28472
rect 11052 28456 11068 28472
rect 11084 28456 11100 28472
rect 11116 28456 11132 28472
rect 11148 28456 11164 28472
rect 11180 28456 11196 28472
rect 11212 28456 11228 28472
rect 11244 28456 11260 28472
rect 11276 28456 11292 28472
rect 11308 28456 11324 28472
rect 11340 28456 11356 28472
rect 11372 28456 11388 28472
rect 11404 28456 11420 28472
rect 11436 28456 11452 28472
rect 11468 28456 11484 28472
rect 11500 28456 11516 28472
rect 11532 28456 11548 28472
rect 11564 28456 11580 28472
rect 11596 28456 11612 28472
rect 11628 28456 11644 28472
rect 11660 28456 11676 28472
rect 11692 28456 11708 28472
rect 11724 28456 11740 28472
rect 11756 28456 11772 28472
rect 11788 28456 11804 28472
rect 11820 28456 26820 28472
rect 9961 28440 26820 28456
rect 9961 28424 9980 28440
rect 9996 28424 10012 28440
rect 10028 28424 10044 28440
rect 10060 28424 10076 28440
rect 10092 28424 10108 28440
rect 10124 28424 10140 28440
rect 10156 28424 10172 28440
rect 10188 28424 10204 28440
rect 10220 28424 10236 28440
rect 10252 28424 10268 28440
rect 10284 28424 10300 28440
rect 10316 28424 10332 28440
rect 10348 28424 10364 28440
rect 10380 28424 10396 28440
rect 10412 28424 10428 28440
rect 10444 28424 10460 28440
rect 10476 28424 10492 28440
rect 10508 28424 10524 28440
rect 10540 28424 10556 28440
rect 10572 28424 10588 28440
rect 10604 28424 10620 28440
rect 10636 28424 10652 28440
rect 10668 28424 10684 28440
rect 10700 28424 10716 28440
rect 10732 28424 10748 28440
rect 10764 28424 10780 28440
rect 10796 28424 10812 28440
rect 10828 28424 10844 28440
rect 10860 28424 10876 28440
rect 10892 28424 10908 28440
rect 10924 28424 10940 28440
rect 10956 28424 10972 28440
rect 10988 28424 11004 28440
rect 11020 28424 11036 28440
rect 11052 28424 11068 28440
rect 11084 28424 11100 28440
rect 11116 28424 11132 28440
rect 11148 28424 11164 28440
rect 11180 28424 11196 28440
rect 11212 28424 11228 28440
rect 11244 28424 11260 28440
rect 11276 28424 11292 28440
rect 11308 28424 11324 28440
rect 11340 28424 11356 28440
rect 11372 28424 11388 28440
rect 11404 28424 11420 28440
rect 11436 28424 11452 28440
rect 11468 28424 11484 28440
rect 11500 28424 11516 28440
rect 11532 28424 11548 28440
rect 11564 28424 11580 28440
rect 11596 28424 11612 28440
rect 11628 28424 11644 28440
rect 11660 28424 11676 28440
rect 11692 28424 11708 28440
rect 11724 28424 11740 28440
rect 11756 28424 11772 28440
rect 11788 28424 11804 28440
rect 11820 28424 26820 28440
rect 9961 28408 26820 28424
rect 9961 28392 9980 28408
rect 9996 28392 10012 28408
rect 10028 28392 10044 28408
rect 10060 28392 10076 28408
rect 10092 28392 10108 28408
rect 10124 28392 10140 28408
rect 10156 28392 10172 28408
rect 10188 28392 10204 28408
rect 10220 28392 10236 28408
rect 10252 28392 10268 28408
rect 10284 28392 10300 28408
rect 10316 28392 10332 28408
rect 10348 28392 10364 28408
rect 10380 28392 10396 28408
rect 10412 28392 10428 28408
rect 10444 28392 10460 28408
rect 10476 28392 10492 28408
rect 10508 28392 10524 28408
rect 10540 28392 10556 28408
rect 10572 28392 10588 28408
rect 10604 28392 10620 28408
rect 10636 28392 10652 28408
rect 10668 28392 10684 28408
rect 10700 28392 10716 28408
rect 10732 28392 10748 28408
rect 10764 28392 10780 28408
rect 10796 28392 10812 28408
rect 10828 28392 10844 28408
rect 10860 28392 10876 28408
rect 10892 28392 10908 28408
rect 10924 28392 10940 28408
rect 10956 28392 10972 28408
rect 10988 28392 11004 28408
rect 11020 28392 11036 28408
rect 11052 28392 11068 28408
rect 11084 28392 11100 28408
rect 11116 28392 11132 28408
rect 11148 28392 11164 28408
rect 11180 28392 11196 28408
rect 11212 28392 11228 28408
rect 11244 28392 11260 28408
rect 11276 28392 11292 28408
rect 11308 28392 11324 28408
rect 11340 28392 11356 28408
rect 11372 28392 11388 28408
rect 11404 28392 11420 28408
rect 11436 28392 11452 28408
rect 11468 28392 11484 28408
rect 11500 28392 11516 28408
rect 11532 28392 11548 28408
rect 11564 28392 11580 28408
rect 11596 28392 11612 28408
rect 11628 28392 11644 28408
rect 11660 28392 11676 28408
rect 11692 28392 11708 28408
rect 11724 28392 11740 28408
rect 11756 28392 11772 28408
rect 11788 28392 11804 28408
rect 11820 28392 26820 28408
rect 9961 28376 26820 28392
rect 9961 28360 9980 28376
rect 9996 28360 10012 28376
rect 10028 28360 10044 28376
rect 10060 28360 10076 28376
rect 10092 28360 10108 28376
rect 10124 28360 10140 28376
rect 10156 28360 10172 28376
rect 10188 28360 10204 28376
rect 10220 28360 10236 28376
rect 10252 28360 10268 28376
rect 10284 28360 10300 28376
rect 10316 28360 10332 28376
rect 10348 28360 10364 28376
rect 10380 28360 10396 28376
rect 10412 28360 10428 28376
rect 10444 28360 10460 28376
rect 10476 28360 10492 28376
rect 10508 28360 10524 28376
rect 10540 28360 10556 28376
rect 10572 28360 10588 28376
rect 10604 28360 10620 28376
rect 10636 28360 10652 28376
rect 10668 28360 10684 28376
rect 10700 28360 10716 28376
rect 10732 28360 10748 28376
rect 10764 28360 10780 28376
rect 10796 28360 10812 28376
rect 10828 28360 10844 28376
rect 10860 28360 10876 28376
rect 10892 28360 10908 28376
rect 10924 28360 10940 28376
rect 10956 28360 10972 28376
rect 10988 28360 11004 28376
rect 11020 28360 11036 28376
rect 11052 28360 11068 28376
rect 11084 28360 11100 28376
rect 11116 28360 11132 28376
rect 11148 28360 11164 28376
rect 11180 28360 11196 28376
rect 11212 28360 11228 28376
rect 11244 28360 11260 28376
rect 11276 28360 11292 28376
rect 11308 28360 11324 28376
rect 11340 28360 11356 28376
rect 11372 28360 11388 28376
rect 11404 28360 11420 28376
rect 11436 28360 11452 28376
rect 11468 28360 11484 28376
rect 11500 28360 11516 28376
rect 11532 28360 11548 28376
rect 11564 28360 11580 28376
rect 11596 28360 11612 28376
rect 11628 28360 11644 28376
rect 11660 28360 11676 28376
rect 11692 28360 11708 28376
rect 11724 28360 11740 28376
rect 11756 28360 11772 28376
rect 11788 28360 11804 28376
rect 11820 28360 26820 28376
rect 9961 28344 26820 28360
rect 9961 28328 9980 28344
rect 9996 28328 10012 28344
rect 10028 28328 10044 28344
rect 10060 28328 10076 28344
rect 10092 28328 10108 28344
rect 10124 28328 10140 28344
rect 10156 28328 10172 28344
rect 10188 28328 10204 28344
rect 10220 28328 10236 28344
rect 10252 28328 10268 28344
rect 10284 28328 10300 28344
rect 10316 28328 10332 28344
rect 10348 28328 10364 28344
rect 10380 28328 10396 28344
rect 10412 28328 10428 28344
rect 10444 28328 10460 28344
rect 10476 28328 10492 28344
rect 10508 28328 10524 28344
rect 10540 28328 10556 28344
rect 10572 28328 10588 28344
rect 10604 28328 10620 28344
rect 10636 28328 10652 28344
rect 10668 28328 10684 28344
rect 10700 28328 10716 28344
rect 10732 28328 10748 28344
rect 10764 28328 10780 28344
rect 10796 28328 10812 28344
rect 10828 28328 10844 28344
rect 10860 28328 10876 28344
rect 10892 28328 10908 28344
rect 10924 28328 10940 28344
rect 10956 28328 10972 28344
rect 10988 28328 11004 28344
rect 11020 28328 11036 28344
rect 11052 28328 11068 28344
rect 11084 28328 11100 28344
rect 11116 28328 11132 28344
rect 11148 28328 11164 28344
rect 11180 28328 11196 28344
rect 11212 28328 11228 28344
rect 11244 28328 11260 28344
rect 11276 28328 11292 28344
rect 11308 28328 11324 28344
rect 11340 28328 11356 28344
rect 11372 28328 11388 28344
rect 11404 28328 11420 28344
rect 11436 28328 11452 28344
rect 11468 28328 11484 28344
rect 11500 28328 11516 28344
rect 11532 28328 11548 28344
rect 11564 28328 11580 28344
rect 11596 28328 11612 28344
rect 11628 28328 11644 28344
rect 11660 28328 11676 28344
rect 11692 28328 11708 28344
rect 11724 28328 11740 28344
rect 11756 28328 11772 28344
rect 11788 28328 11804 28344
rect 11820 28328 26820 28344
rect 9961 28312 26820 28328
rect 9961 28296 9980 28312
rect 9996 28296 10012 28312
rect 10028 28296 10044 28312
rect 10060 28296 10076 28312
rect 10092 28296 10108 28312
rect 10124 28296 10140 28312
rect 10156 28296 10172 28312
rect 10188 28296 10204 28312
rect 10220 28296 10236 28312
rect 10252 28296 10268 28312
rect 10284 28296 10300 28312
rect 10316 28296 10332 28312
rect 10348 28296 10364 28312
rect 10380 28296 10396 28312
rect 10412 28296 10428 28312
rect 10444 28296 10460 28312
rect 10476 28296 10492 28312
rect 10508 28296 10524 28312
rect 10540 28296 10556 28312
rect 10572 28296 10588 28312
rect 10604 28296 10620 28312
rect 10636 28296 10652 28312
rect 10668 28296 10684 28312
rect 10700 28296 10716 28312
rect 10732 28296 10748 28312
rect 10764 28296 10780 28312
rect 10796 28296 10812 28312
rect 10828 28296 10844 28312
rect 10860 28296 10876 28312
rect 10892 28296 10908 28312
rect 10924 28296 10940 28312
rect 10956 28296 10972 28312
rect 10988 28296 11004 28312
rect 11020 28296 11036 28312
rect 11052 28296 11068 28312
rect 11084 28296 11100 28312
rect 11116 28296 11132 28312
rect 11148 28296 11164 28312
rect 11180 28296 11196 28312
rect 11212 28296 11228 28312
rect 11244 28296 11260 28312
rect 11276 28296 11292 28312
rect 11308 28296 11324 28312
rect 11340 28296 11356 28312
rect 11372 28296 11388 28312
rect 11404 28296 11420 28312
rect 11436 28296 11452 28312
rect 11468 28296 11484 28312
rect 11500 28296 11516 28312
rect 11532 28296 11548 28312
rect 11564 28296 11580 28312
rect 11596 28296 11612 28312
rect 11628 28296 11644 28312
rect 11660 28296 11676 28312
rect 11692 28296 11708 28312
rect 11724 28296 11740 28312
rect 11756 28296 11772 28312
rect 11788 28296 11804 28312
rect 11820 28296 26820 28312
rect 9961 28280 26820 28296
rect 9961 28264 9980 28280
rect 9996 28264 10012 28280
rect 10028 28264 10044 28280
rect 10060 28264 10076 28280
rect 10092 28264 10108 28280
rect 10124 28264 10140 28280
rect 10156 28264 10172 28280
rect 10188 28264 10204 28280
rect 10220 28264 10236 28280
rect 10252 28264 10268 28280
rect 10284 28264 10300 28280
rect 10316 28264 10332 28280
rect 10348 28264 10364 28280
rect 10380 28264 10396 28280
rect 10412 28264 10428 28280
rect 10444 28264 10460 28280
rect 10476 28264 10492 28280
rect 10508 28264 10524 28280
rect 10540 28264 10556 28280
rect 10572 28264 10588 28280
rect 10604 28264 10620 28280
rect 10636 28264 10652 28280
rect 10668 28264 10684 28280
rect 10700 28264 10716 28280
rect 10732 28264 10748 28280
rect 10764 28264 10780 28280
rect 10796 28264 10812 28280
rect 10828 28264 10844 28280
rect 10860 28264 10876 28280
rect 10892 28264 10908 28280
rect 10924 28264 10940 28280
rect 10956 28264 10972 28280
rect 10988 28264 11004 28280
rect 11020 28264 11036 28280
rect 11052 28264 11068 28280
rect 11084 28264 11100 28280
rect 11116 28264 11132 28280
rect 11148 28264 11164 28280
rect 11180 28264 11196 28280
rect 11212 28264 11228 28280
rect 11244 28264 11260 28280
rect 11276 28264 11292 28280
rect 11308 28264 11324 28280
rect 11340 28264 11356 28280
rect 11372 28264 11388 28280
rect 11404 28264 11420 28280
rect 11436 28264 11452 28280
rect 11468 28264 11484 28280
rect 11500 28264 11516 28280
rect 11532 28264 11548 28280
rect 11564 28264 11580 28280
rect 11596 28264 11612 28280
rect 11628 28264 11644 28280
rect 11660 28264 11676 28280
rect 11692 28264 11708 28280
rect 11724 28264 11740 28280
rect 11756 28264 11772 28280
rect 11788 28264 11804 28280
rect 11820 28264 26820 28280
rect 9961 28241 26820 28264
rect 11840 28240 26820 28241
rect 9820 27779 10200 27780
rect 9321 27764 10200 27779
rect 9321 27748 9338 27764
rect 9354 27748 9370 27764
rect 9386 27748 9402 27764
rect 9418 27748 9434 27764
rect 9450 27748 9466 27764
rect 9482 27748 9498 27764
rect 9514 27748 9530 27764
rect 9546 27748 9562 27764
rect 9578 27748 9594 27764
rect 9610 27748 9626 27764
rect 9642 27748 9658 27764
rect 9674 27748 9690 27764
rect 9706 27748 9722 27764
rect 9738 27748 9754 27764
rect 9770 27748 9786 27764
rect 9802 27748 10200 27764
rect 9321 27740 10200 27748
rect 9321 27732 10240 27740
rect 9321 27716 9338 27732
rect 9354 27716 9370 27732
rect 9386 27716 9402 27732
rect 9418 27716 9434 27732
rect 9450 27716 9466 27732
rect 9482 27716 9498 27732
rect 9514 27716 9530 27732
rect 9546 27716 9562 27732
rect 9578 27716 9594 27732
rect 9610 27716 9626 27732
rect 9642 27716 9658 27732
rect 9674 27716 9690 27732
rect 9706 27716 9722 27732
rect 9738 27716 9754 27732
rect 9770 27716 9786 27732
rect 9802 27720 10240 27732
rect 9802 27716 10280 27720
rect 9321 27700 10280 27716
rect 9321 27684 9338 27700
rect 9354 27684 9370 27700
rect 9386 27684 9402 27700
rect 9418 27684 9434 27700
rect 9450 27684 9466 27700
rect 9482 27684 9498 27700
rect 9514 27684 9530 27700
rect 9546 27684 9562 27700
rect 9578 27684 9594 27700
rect 9610 27684 9626 27700
rect 9642 27684 9658 27700
rect 9674 27684 9690 27700
rect 9706 27684 9722 27700
rect 9738 27684 9754 27700
rect 9770 27684 9786 27700
rect 9802 27684 10280 27700
rect 9321 27680 10280 27684
rect 9321 27668 10320 27680
rect 9321 27652 9338 27668
rect 9354 27652 9370 27668
rect 9386 27652 9402 27668
rect 9418 27652 9434 27668
rect 9450 27652 9466 27668
rect 9482 27652 9498 27668
rect 9514 27652 9530 27668
rect 9546 27652 9562 27668
rect 9578 27652 9594 27668
rect 9610 27652 9626 27668
rect 9642 27652 9658 27668
rect 9674 27652 9690 27668
rect 9706 27652 9722 27668
rect 9738 27652 9754 27668
rect 9770 27652 9786 27668
rect 9802 27652 10320 27668
rect 9321 27640 10320 27652
rect 9321 27636 10360 27640
rect 9321 27620 9338 27636
rect 9354 27620 9370 27636
rect 9386 27620 9402 27636
rect 9418 27620 9434 27636
rect 9450 27620 9466 27636
rect 9482 27620 9498 27636
rect 9514 27620 9530 27636
rect 9546 27620 9562 27636
rect 9578 27620 9594 27636
rect 9610 27620 9626 27636
rect 9642 27620 9658 27636
rect 9674 27620 9690 27636
rect 9706 27620 9722 27636
rect 9738 27620 9754 27636
rect 9770 27620 9786 27636
rect 9802 27620 10360 27636
rect 9321 27604 10360 27620
rect 9321 27588 9338 27604
rect 9354 27588 9370 27604
rect 9386 27588 9402 27604
rect 9418 27588 9434 27604
rect 9450 27588 9466 27604
rect 9482 27588 9498 27604
rect 9514 27588 9530 27604
rect 9546 27588 9562 27604
rect 9578 27588 9594 27604
rect 9610 27588 9626 27604
rect 9642 27588 9658 27604
rect 9674 27588 9690 27604
rect 9706 27588 9722 27604
rect 9738 27588 9754 27604
rect 9770 27588 9786 27604
rect 9802 27600 10360 27604
rect 9802 27588 10400 27600
rect 9321 27572 10400 27588
rect 9321 27556 9338 27572
rect 9354 27556 9370 27572
rect 9386 27556 9402 27572
rect 9418 27556 9434 27572
rect 9450 27556 9466 27572
rect 9482 27556 9498 27572
rect 9514 27556 9530 27572
rect 9546 27556 9562 27572
rect 9578 27556 9594 27572
rect 9610 27556 9626 27572
rect 9642 27556 9658 27572
rect 9674 27556 9690 27572
rect 9706 27556 9722 27572
rect 9738 27556 9754 27572
rect 9770 27556 9786 27572
rect 9802 27560 10400 27572
rect 9802 27556 10440 27560
rect 9321 27540 10440 27556
rect 9321 27524 9338 27540
rect 9354 27524 9370 27540
rect 9386 27524 9402 27540
rect 9418 27524 9434 27540
rect 9450 27524 9466 27540
rect 9482 27524 9498 27540
rect 9514 27524 9530 27540
rect 9546 27524 9562 27540
rect 9578 27524 9594 27540
rect 9610 27524 9626 27540
rect 9642 27524 9658 27540
rect 9674 27524 9690 27540
rect 9706 27524 9722 27540
rect 9738 27524 9754 27540
rect 9770 27524 9786 27540
rect 9802 27524 10440 27540
rect 9321 27520 10440 27524
rect 9321 27508 10480 27520
rect 9321 27492 9338 27508
rect 9354 27492 9370 27508
rect 9386 27492 9402 27508
rect 9418 27492 9434 27508
rect 9450 27492 9466 27508
rect 9482 27492 9498 27508
rect 9514 27492 9530 27508
rect 9546 27492 9562 27508
rect 9578 27492 9594 27508
rect 9610 27492 9626 27508
rect 9642 27492 9658 27508
rect 9674 27492 9690 27508
rect 9706 27492 9722 27508
rect 9738 27492 9754 27508
rect 9770 27492 9786 27508
rect 9802 27492 10480 27508
rect 9321 27480 10480 27492
rect 9321 27476 10520 27480
rect 9321 27460 9338 27476
rect 9354 27460 9370 27476
rect 9386 27460 9402 27476
rect 9418 27460 9434 27476
rect 9450 27460 9466 27476
rect 9482 27460 9498 27476
rect 9514 27460 9530 27476
rect 9546 27460 9562 27476
rect 9578 27460 9594 27476
rect 9610 27460 9626 27476
rect 9642 27460 9658 27476
rect 9674 27460 9690 27476
rect 9706 27460 9722 27476
rect 9738 27460 9754 27476
rect 9770 27460 9786 27476
rect 9802 27460 10520 27476
rect 9321 27444 10520 27460
rect 9321 27428 9338 27444
rect 9354 27428 9370 27444
rect 9386 27428 9402 27444
rect 9418 27428 9434 27444
rect 9450 27428 9466 27444
rect 9482 27428 9498 27444
rect 9514 27428 9530 27444
rect 9546 27428 9562 27444
rect 9578 27428 9594 27444
rect 9610 27428 9626 27444
rect 9642 27428 9658 27444
rect 9674 27428 9690 27444
rect 9706 27428 9722 27444
rect 9738 27428 9754 27444
rect 9770 27428 9786 27444
rect 9802 27440 10520 27444
rect 9802 27428 10560 27440
rect 9321 27412 10560 27428
rect 9321 27396 9338 27412
rect 9354 27396 9370 27412
rect 9386 27396 9402 27412
rect 9418 27396 9434 27412
rect 9450 27396 9466 27412
rect 9482 27396 9498 27412
rect 9514 27396 9530 27412
rect 9546 27396 9562 27412
rect 9578 27396 9594 27412
rect 9610 27396 9626 27412
rect 9642 27396 9658 27412
rect 9674 27396 9690 27412
rect 9706 27396 9722 27412
rect 9738 27396 9754 27412
rect 9770 27396 9786 27412
rect 9802 27400 10560 27412
rect 9802 27396 10600 27400
rect 9321 27380 10600 27396
rect 9321 27364 9338 27380
rect 9354 27364 9370 27380
rect 9386 27364 9402 27380
rect 9418 27364 9434 27380
rect 9450 27364 9466 27380
rect 9482 27364 9498 27380
rect 9514 27364 9530 27380
rect 9546 27364 9562 27380
rect 9578 27364 9594 27380
rect 9610 27364 9626 27380
rect 9642 27364 9658 27380
rect 9674 27364 9690 27380
rect 9706 27364 9722 27380
rect 9738 27364 9754 27380
rect 9770 27364 9786 27380
rect 9802 27364 10600 27380
rect 9321 27360 10600 27364
rect 9321 27348 10640 27360
rect 9321 27332 9338 27348
rect 9354 27332 9370 27348
rect 9386 27332 9402 27348
rect 9418 27332 9434 27348
rect 9450 27332 9466 27348
rect 9482 27332 9498 27348
rect 9514 27332 9530 27348
rect 9546 27332 9562 27348
rect 9578 27332 9594 27348
rect 9610 27332 9626 27348
rect 9642 27332 9658 27348
rect 9674 27332 9690 27348
rect 9706 27332 9722 27348
rect 9738 27332 9754 27348
rect 9770 27332 9786 27348
rect 9802 27332 10640 27348
rect 9321 27320 10640 27332
rect 9321 27316 10680 27320
rect 9321 27300 9338 27316
rect 9354 27300 9370 27316
rect 9386 27300 9402 27316
rect 9418 27300 9434 27316
rect 9450 27300 9466 27316
rect 9482 27300 9498 27316
rect 9514 27300 9530 27316
rect 9546 27300 9562 27316
rect 9578 27300 9594 27316
rect 9610 27300 9626 27316
rect 9642 27300 9658 27316
rect 9674 27300 9690 27316
rect 9706 27300 9722 27316
rect 9738 27300 9754 27316
rect 9770 27300 9786 27316
rect 9802 27300 10680 27316
rect 9321 27284 10680 27300
rect 9321 27268 9338 27284
rect 9354 27268 9370 27284
rect 9386 27268 9402 27284
rect 9418 27268 9434 27284
rect 9450 27268 9466 27284
rect 9482 27268 9498 27284
rect 9514 27268 9530 27284
rect 9546 27268 9562 27284
rect 9578 27268 9594 27284
rect 9610 27268 9626 27284
rect 9642 27268 9658 27284
rect 9674 27268 9690 27284
rect 9706 27268 9722 27284
rect 9738 27268 9754 27284
rect 9770 27268 9786 27284
rect 9802 27280 10680 27284
rect 9802 27268 10720 27280
rect 9321 27252 10720 27268
rect 9321 27236 9338 27252
rect 9354 27236 9370 27252
rect 9386 27236 9402 27252
rect 9418 27236 9434 27252
rect 9450 27236 9466 27252
rect 9482 27236 9498 27252
rect 9514 27236 9530 27252
rect 9546 27236 9562 27252
rect 9578 27236 9594 27252
rect 9610 27236 9626 27252
rect 9642 27236 9658 27252
rect 9674 27236 9690 27252
rect 9706 27236 9722 27252
rect 9738 27236 9754 27252
rect 9770 27236 9786 27252
rect 9802 27240 10720 27252
rect 9802 27236 10760 27240
rect 9321 27220 10760 27236
rect 9321 27204 9338 27220
rect 9354 27204 9370 27220
rect 9386 27204 9402 27220
rect 9418 27204 9434 27220
rect 9450 27204 9466 27220
rect 9482 27204 9498 27220
rect 9514 27204 9530 27220
rect 9546 27204 9562 27220
rect 9578 27204 9594 27220
rect 9610 27204 9626 27220
rect 9642 27204 9658 27220
rect 9674 27204 9690 27220
rect 9706 27204 9722 27220
rect 9738 27204 9754 27220
rect 9770 27204 9786 27220
rect 9802 27204 10760 27220
rect 9321 27200 10760 27204
rect 9321 27188 10800 27200
rect 9321 27172 9338 27188
rect 9354 27172 9370 27188
rect 9386 27172 9402 27188
rect 9418 27172 9434 27188
rect 9450 27172 9466 27188
rect 9482 27172 9498 27188
rect 9514 27172 9530 27188
rect 9546 27172 9562 27188
rect 9578 27172 9594 27188
rect 9610 27172 9626 27188
rect 9642 27172 9658 27188
rect 9674 27172 9690 27188
rect 9706 27172 9722 27188
rect 9738 27172 9754 27188
rect 9770 27172 9786 27188
rect 9802 27172 10800 27188
rect 9321 27160 10800 27172
rect 9321 27156 10840 27160
rect 9321 27140 9338 27156
rect 9354 27140 9370 27156
rect 9386 27140 9402 27156
rect 9418 27140 9434 27156
rect 9450 27140 9466 27156
rect 9482 27140 9498 27156
rect 9514 27140 9530 27156
rect 9546 27140 9562 27156
rect 9578 27140 9594 27156
rect 9610 27140 9626 27156
rect 9642 27140 9658 27156
rect 9674 27140 9690 27156
rect 9706 27140 9722 27156
rect 9738 27140 9754 27156
rect 9770 27140 9786 27156
rect 9802 27140 10840 27156
rect 9321 27124 10840 27140
rect 9321 27108 9338 27124
rect 9354 27108 9370 27124
rect 9386 27108 9402 27124
rect 9418 27108 9434 27124
rect 9450 27108 9466 27124
rect 9482 27108 9498 27124
rect 9514 27108 9530 27124
rect 9546 27108 9562 27124
rect 9578 27108 9594 27124
rect 9610 27108 9626 27124
rect 9642 27108 9658 27124
rect 9674 27108 9690 27124
rect 9706 27108 9722 27124
rect 9738 27108 9754 27124
rect 9770 27108 9786 27124
rect 9802 27120 10840 27124
rect 9802 27108 10880 27120
rect 9321 27092 10880 27108
rect 9321 27076 9338 27092
rect 9354 27076 9370 27092
rect 9386 27076 9402 27092
rect 9418 27076 9434 27092
rect 9450 27076 9466 27092
rect 9482 27076 9498 27092
rect 9514 27076 9530 27092
rect 9546 27076 9562 27092
rect 9578 27076 9594 27092
rect 9610 27076 9626 27092
rect 9642 27076 9658 27092
rect 9674 27076 9690 27092
rect 9706 27076 9722 27092
rect 9738 27076 9754 27092
rect 9770 27076 9786 27092
rect 9802 27080 10880 27092
rect 9802 27076 10920 27080
rect 9321 27060 10920 27076
rect 9321 27044 9338 27060
rect 9354 27044 9370 27060
rect 9386 27044 9402 27060
rect 9418 27044 9434 27060
rect 9450 27044 9466 27060
rect 9482 27044 9498 27060
rect 9514 27044 9530 27060
rect 9546 27044 9562 27060
rect 9578 27044 9594 27060
rect 9610 27044 9626 27060
rect 9642 27044 9658 27060
rect 9674 27044 9690 27060
rect 9706 27044 9722 27060
rect 9738 27044 9754 27060
rect 9770 27044 9786 27060
rect 9802 27044 10920 27060
rect 9321 27040 10920 27044
rect 9321 27028 10960 27040
rect 9321 27012 9338 27028
rect 9354 27012 9370 27028
rect 9386 27012 9402 27028
rect 9418 27012 9434 27028
rect 9450 27012 9466 27028
rect 9482 27012 9498 27028
rect 9514 27012 9530 27028
rect 9546 27012 9562 27028
rect 9578 27012 9594 27028
rect 9610 27012 9626 27028
rect 9642 27012 9658 27028
rect 9674 27012 9690 27028
rect 9706 27012 9722 27028
rect 9738 27012 9754 27028
rect 9770 27012 9786 27028
rect 9802 27012 10960 27028
rect 9321 27000 10960 27012
rect 9321 26996 11000 27000
rect 9321 26980 9338 26996
rect 9354 26980 9370 26996
rect 9386 26980 9402 26996
rect 9418 26980 9434 26996
rect 9450 26980 9466 26996
rect 9482 26980 9498 26996
rect 9514 26980 9530 26996
rect 9546 26980 9562 26996
rect 9578 26980 9594 26996
rect 9610 26980 9626 26996
rect 9642 26980 9658 26996
rect 9674 26980 9690 26996
rect 9706 26980 9722 26996
rect 9738 26980 9754 26996
rect 9770 26980 9786 26996
rect 9802 26980 11000 26996
rect 9321 26964 11000 26980
rect 9321 26948 9338 26964
rect 9354 26948 9370 26964
rect 9386 26948 9402 26964
rect 9418 26948 9434 26964
rect 9450 26948 9466 26964
rect 9482 26948 9498 26964
rect 9514 26948 9530 26964
rect 9546 26948 9562 26964
rect 9578 26948 9594 26964
rect 9610 26948 9626 26964
rect 9642 26948 9658 26964
rect 9674 26948 9690 26964
rect 9706 26948 9722 26964
rect 9738 26948 9754 26964
rect 9770 26948 9786 26964
rect 9802 26960 11000 26964
rect 9802 26948 11040 26960
rect 9321 26932 11040 26948
rect 9321 26916 9338 26932
rect 9354 26916 9370 26932
rect 9386 26916 9402 26932
rect 9418 26916 9434 26932
rect 9450 26916 9466 26932
rect 9482 26916 9498 26932
rect 9514 26916 9530 26932
rect 9546 26916 9562 26932
rect 9578 26916 9594 26932
rect 9610 26916 9626 26932
rect 9642 26916 9658 26932
rect 9674 26916 9690 26932
rect 9706 26916 9722 26932
rect 9738 26916 9754 26932
rect 9770 26916 9786 26932
rect 9802 26920 11040 26932
rect 9802 26916 11080 26920
rect 9321 26900 11080 26916
rect 9321 26884 9338 26900
rect 9354 26884 9370 26900
rect 9386 26884 9402 26900
rect 9418 26884 9434 26900
rect 9450 26884 9466 26900
rect 9482 26884 9498 26900
rect 9514 26884 9530 26900
rect 9546 26884 9562 26900
rect 9578 26884 9594 26900
rect 9610 26884 9626 26900
rect 9642 26884 9658 26900
rect 9674 26884 9690 26900
rect 9706 26884 9722 26900
rect 9738 26884 9754 26900
rect 9770 26884 9786 26900
rect 9802 26884 11120 26900
rect 9321 26868 11120 26884
rect 9321 26852 9338 26868
rect 9354 26852 9370 26868
rect 9386 26852 9402 26868
rect 9418 26852 9434 26868
rect 9450 26852 9466 26868
rect 9482 26852 9498 26868
rect 9514 26852 9530 26868
rect 9546 26852 9562 26868
rect 9578 26852 9594 26868
rect 9610 26852 9626 26868
rect 9642 26852 9658 26868
rect 9674 26852 9690 26868
rect 9706 26852 9722 26868
rect 9738 26852 9754 26868
rect 9770 26852 9786 26868
rect 9802 26860 11120 26868
rect 9802 26852 11160 26860
rect 9321 26836 11160 26852
rect 9321 26820 9338 26836
rect 9354 26820 9370 26836
rect 9386 26820 9402 26836
rect 9418 26820 9434 26836
rect 9450 26820 9466 26836
rect 9482 26820 9498 26836
rect 9514 26820 9530 26836
rect 9546 26820 9562 26836
rect 9578 26820 9594 26836
rect 9610 26820 9626 26836
rect 9642 26820 9658 26836
rect 9674 26820 9690 26836
rect 9706 26820 9722 26836
rect 9738 26820 9754 26836
rect 9770 26820 9786 26836
rect 9802 26820 11160 26836
rect 9321 26804 11200 26820
rect 9321 26788 9338 26804
rect 9354 26788 9370 26804
rect 9386 26788 9402 26804
rect 9418 26788 9434 26804
rect 9450 26788 9466 26804
rect 9482 26788 9498 26804
rect 9514 26788 9530 26804
rect 9546 26788 9562 26804
rect 9578 26788 9594 26804
rect 9610 26788 9626 26804
rect 9642 26788 9658 26804
rect 9674 26788 9690 26804
rect 9706 26788 9722 26804
rect 9738 26788 9754 26804
rect 9770 26788 9786 26804
rect 9802 26788 11200 26804
rect 9321 26780 11200 26788
rect 9321 26772 11240 26780
rect 9321 26756 9338 26772
rect 9354 26756 9370 26772
rect 9386 26756 9402 26772
rect 9418 26756 9434 26772
rect 9450 26756 9466 26772
rect 9482 26756 9498 26772
rect 9514 26756 9530 26772
rect 9546 26756 9562 26772
rect 9578 26756 9594 26772
rect 9610 26756 9626 26772
rect 9642 26756 9658 26772
rect 9674 26756 9690 26772
rect 9706 26756 9722 26772
rect 9738 26756 9754 26772
rect 9770 26756 9786 26772
rect 9802 26756 11240 26772
rect 9321 26740 11240 26756
rect 9321 26724 9338 26740
rect 9354 26724 9370 26740
rect 9386 26724 9402 26740
rect 9418 26724 9434 26740
rect 9450 26724 9466 26740
rect 9482 26724 9498 26740
rect 9514 26724 9530 26740
rect 9546 26724 9562 26740
rect 9578 26724 9594 26740
rect 9610 26724 9626 26740
rect 9642 26724 9658 26740
rect 9674 26724 9690 26740
rect 9706 26724 9722 26740
rect 9738 26724 9754 26740
rect 9770 26724 9786 26740
rect 9802 26724 11280 26740
rect 9321 26708 11280 26724
rect 9321 26692 9338 26708
rect 9354 26692 9370 26708
rect 9386 26692 9402 26708
rect 9418 26692 9434 26708
rect 9450 26692 9466 26708
rect 9482 26692 9498 26708
rect 9514 26692 9530 26708
rect 9546 26692 9562 26708
rect 9578 26692 9594 26708
rect 9610 26692 9626 26708
rect 9642 26692 9658 26708
rect 9674 26692 9690 26708
rect 9706 26692 9722 26708
rect 9738 26692 9754 26708
rect 9770 26692 9786 26708
rect 9802 26700 11280 26708
rect 9802 26692 11320 26700
rect 9321 26676 11320 26692
rect 9321 26660 9338 26676
rect 9354 26660 9370 26676
rect 9386 26660 9402 26676
rect 9418 26660 9434 26676
rect 9450 26660 9466 26676
rect 9482 26660 9498 26676
rect 9514 26660 9530 26676
rect 9546 26660 9562 26676
rect 9578 26660 9594 26676
rect 9610 26660 9626 26676
rect 9642 26660 9658 26676
rect 9674 26660 9690 26676
rect 9706 26660 9722 26676
rect 9738 26660 9754 26676
rect 9770 26660 9786 26676
rect 9802 26660 11320 26676
rect 9321 26644 11320 26660
rect 9321 26628 9338 26644
rect 9354 26628 9370 26644
rect 9386 26628 9402 26644
rect 9418 26628 9434 26644
rect 9450 26628 9466 26644
rect 9482 26628 9498 26644
rect 9514 26628 9530 26644
rect 9546 26628 9562 26644
rect 9578 26628 9594 26644
rect 9610 26628 9626 26644
rect 9642 26628 9658 26644
rect 9674 26628 9690 26644
rect 9706 26628 9722 26644
rect 9738 26628 9754 26644
rect 9770 26628 9786 26644
rect 9802 26628 11320 26644
rect 9321 26612 11320 26628
rect 9321 26596 9338 26612
rect 9354 26596 9370 26612
rect 9386 26596 9402 26612
rect 9418 26596 9434 26612
rect 9450 26596 9466 26612
rect 9482 26596 9498 26612
rect 9514 26596 9530 26612
rect 9546 26596 9562 26612
rect 9578 26596 9594 26612
rect 9610 26596 9626 26612
rect 9642 26596 9658 26612
rect 9674 26596 9690 26612
rect 9706 26596 9722 26612
rect 9738 26596 9754 26612
rect 9770 26596 9786 26612
rect 9802 26596 11320 26612
rect 9321 26580 11320 26596
rect 9321 26564 9338 26580
rect 9354 26564 9370 26580
rect 9386 26564 9402 26580
rect 9418 26564 9434 26580
rect 9450 26564 9466 26580
rect 9482 26564 9498 26580
rect 9514 26564 9530 26580
rect 9546 26564 9562 26580
rect 9578 26564 9594 26580
rect 9610 26564 9626 26580
rect 9642 26564 9658 26580
rect 9674 26564 9690 26580
rect 9706 26564 9722 26580
rect 9738 26564 9754 26580
rect 9770 26564 9786 26580
rect 9802 26564 11320 26580
rect 9321 26548 11320 26564
rect 9321 26532 9338 26548
rect 9354 26532 9370 26548
rect 9386 26532 9402 26548
rect 9418 26532 9434 26548
rect 9450 26532 9466 26548
rect 9482 26532 9498 26548
rect 9514 26532 9530 26548
rect 9546 26532 9562 26548
rect 9578 26532 9594 26548
rect 9610 26532 9626 26548
rect 9642 26532 9658 26548
rect 9674 26532 9690 26548
rect 9706 26532 9722 26548
rect 9738 26532 9754 26548
rect 9770 26532 9786 26548
rect 9802 26532 11320 26548
rect 9321 26516 11320 26532
rect 26640 26520 26820 28240
rect 9321 26500 9338 26516
rect 9354 26500 9370 26516
rect 9386 26500 9402 26516
rect 9418 26500 9434 26516
rect 9450 26500 9466 26516
rect 9482 26500 9498 26516
rect 9514 26500 9530 26516
rect 9546 26500 9562 26516
rect 9578 26500 9594 26516
rect 9610 26500 9626 26516
rect 9642 26500 9658 26516
rect 9674 26500 9690 26516
rect 9706 26500 9722 26516
rect 9738 26500 9754 26516
rect 9770 26500 9786 26516
rect 9802 26500 11320 26516
rect 9321 26484 11320 26500
rect 9321 26468 9338 26484
rect 9354 26468 9370 26484
rect 9386 26468 9402 26484
rect 9418 26468 9434 26484
rect 9450 26468 9466 26484
rect 9482 26468 9498 26484
rect 9514 26468 9530 26484
rect 9546 26468 9562 26484
rect 9578 26468 9594 26484
rect 9610 26468 9626 26484
rect 9642 26468 9658 26484
rect 9674 26468 9690 26484
rect 9706 26468 9722 26484
rect 9738 26468 9754 26484
rect 9770 26468 9786 26484
rect 9802 26468 11320 26484
rect 9321 26452 11320 26468
rect 9321 26436 9338 26452
rect 9354 26436 9370 26452
rect 9386 26436 9402 26452
rect 9418 26436 9434 26452
rect 9450 26436 9466 26452
rect 9482 26436 9498 26452
rect 9514 26436 9530 26452
rect 9546 26436 9562 26452
rect 9578 26436 9594 26452
rect 9610 26436 9626 26452
rect 9642 26436 9658 26452
rect 9674 26436 9690 26452
rect 9706 26436 9722 26452
rect 9738 26436 9754 26452
rect 9770 26436 9786 26452
rect 9802 26436 11320 26452
rect 9321 26421 11320 26436
rect 9820 26420 11320 26421
<< m2contact >>
rect 9980 28680 9996 28696
rect 10012 28680 10028 28696
rect 10044 28680 10060 28696
rect 10076 28680 10092 28696
rect 10108 28680 10124 28696
rect 10140 28680 10156 28696
rect 10172 28680 10188 28696
rect 10204 28680 10220 28696
rect 10236 28680 10252 28696
rect 10268 28680 10284 28696
rect 10300 28680 10316 28696
rect 10332 28680 10348 28696
rect 10364 28680 10380 28696
rect 10396 28680 10412 28696
rect 10428 28680 10444 28696
rect 10460 28680 10476 28696
rect 10492 28680 10508 28696
rect 10524 28680 10540 28696
rect 10556 28680 10572 28696
rect 10588 28680 10604 28696
rect 10620 28680 10636 28696
rect 10652 28680 10668 28696
rect 10684 28680 10700 28696
rect 10716 28680 10732 28696
rect 10748 28680 10764 28696
rect 10780 28680 10796 28696
rect 10812 28680 10828 28696
rect 10844 28680 10860 28696
rect 10876 28680 10892 28696
rect 10908 28680 10924 28696
rect 10940 28680 10956 28696
rect 10972 28680 10988 28696
rect 11004 28680 11020 28696
rect 11036 28680 11052 28696
rect 11068 28680 11084 28696
rect 11100 28680 11116 28696
rect 11132 28680 11148 28696
rect 11164 28680 11180 28696
rect 11196 28680 11212 28696
rect 11228 28680 11244 28696
rect 11260 28680 11276 28696
rect 11292 28680 11308 28696
rect 11324 28680 11340 28696
rect 11356 28680 11372 28696
rect 11388 28680 11404 28696
rect 11420 28680 11436 28696
rect 11452 28680 11468 28696
rect 11484 28680 11500 28696
rect 11516 28680 11532 28696
rect 11548 28680 11564 28696
rect 11580 28680 11596 28696
rect 11612 28680 11628 28696
rect 11644 28680 11660 28696
rect 11676 28680 11692 28696
rect 11708 28680 11724 28696
rect 11740 28680 11756 28696
rect 11772 28680 11788 28696
rect 11804 28680 11820 28696
rect 9980 28648 9996 28664
rect 10012 28648 10028 28664
rect 10044 28648 10060 28664
rect 10076 28648 10092 28664
rect 10108 28648 10124 28664
rect 10140 28648 10156 28664
rect 10172 28648 10188 28664
rect 10204 28648 10220 28664
rect 10236 28648 10252 28664
rect 10268 28648 10284 28664
rect 10300 28648 10316 28664
rect 10332 28648 10348 28664
rect 10364 28648 10380 28664
rect 10396 28648 10412 28664
rect 10428 28648 10444 28664
rect 10460 28648 10476 28664
rect 10492 28648 10508 28664
rect 10524 28648 10540 28664
rect 10556 28648 10572 28664
rect 10588 28648 10604 28664
rect 10620 28648 10636 28664
rect 10652 28648 10668 28664
rect 10684 28648 10700 28664
rect 10716 28648 10732 28664
rect 10748 28648 10764 28664
rect 10780 28648 10796 28664
rect 10812 28648 10828 28664
rect 10844 28648 10860 28664
rect 10876 28648 10892 28664
rect 10908 28648 10924 28664
rect 10940 28648 10956 28664
rect 10972 28648 10988 28664
rect 11004 28648 11020 28664
rect 11036 28648 11052 28664
rect 11068 28648 11084 28664
rect 11100 28648 11116 28664
rect 11132 28648 11148 28664
rect 11164 28648 11180 28664
rect 11196 28648 11212 28664
rect 11228 28648 11244 28664
rect 11260 28648 11276 28664
rect 11292 28648 11308 28664
rect 11324 28648 11340 28664
rect 11356 28648 11372 28664
rect 11388 28648 11404 28664
rect 11420 28648 11436 28664
rect 11452 28648 11468 28664
rect 11484 28648 11500 28664
rect 11516 28648 11532 28664
rect 11548 28648 11564 28664
rect 11580 28648 11596 28664
rect 11612 28648 11628 28664
rect 11644 28648 11660 28664
rect 11676 28648 11692 28664
rect 11708 28648 11724 28664
rect 11740 28648 11756 28664
rect 11772 28648 11788 28664
rect 11804 28648 11820 28664
rect 9980 28616 9996 28632
rect 10012 28616 10028 28632
rect 10044 28616 10060 28632
rect 10076 28616 10092 28632
rect 10108 28616 10124 28632
rect 10140 28616 10156 28632
rect 10172 28616 10188 28632
rect 10204 28616 10220 28632
rect 10236 28616 10252 28632
rect 10268 28616 10284 28632
rect 10300 28616 10316 28632
rect 10332 28616 10348 28632
rect 10364 28616 10380 28632
rect 10396 28616 10412 28632
rect 10428 28616 10444 28632
rect 10460 28616 10476 28632
rect 10492 28616 10508 28632
rect 10524 28616 10540 28632
rect 10556 28616 10572 28632
rect 10588 28616 10604 28632
rect 10620 28616 10636 28632
rect 10652 28616 10668 28632
rect 10684 28616 10700 28632
rect 10716 28616 10732 28632
rect 10748 28616 10764 28632
rect 10780 28616 10796 28632
rect 10812 28616 10828 28632
rect 10844 28616 10860 28632
rect 10876 28616 10892 28632
rect 10908 28616 10924 28632
rect 10940 28616 10956 28632
rect 10972 28616 10988 28632
rect 11004 28616 11020 28632
rect 11036 28616 11052 28632
rect 11068 28616 11084 28632
rect 11100 28616 11116 28632
rect 11132 28616 11148 28632
rect 11164 28616 11180 28632
rect 11196 28616 11212 28632
rect 11228 28616 11244 28632
rect 11260 28616 11276 28632
rect 11292 28616 11308 28632
rect 11324 28616 11340 28632
rect 11356 28616 11372 28632
rect 11388 28616 11404 28632
rect 11420 28616 11436 28632
rect 11452 28616 11468 28632
rect 11484 28616 11500 28632
rect 11516 28616 11532 28632
rect 11548 28616 11564 28632
rect 11580 28616 11596 28632
rect 11612 28616 11628 28632
rect 11644 28616 11660 28632
rect 11676 28616 11692 28632
rect 11708 28616 11724 28632
rect 11740 28616 11756 28632
rect 11772 28616 11788 28632
rect 11804 28616 11820 28632
rect 9980 28584 9996 28600
rect 10012 28584 10028 28600
rect 10044 28584 10060 28600
rect 10076 28584 10092 28600
rect 10108 28584 10124 28600
rect 10140 28584 10156 28600
rect 10172 28584 10188 28600
rect 10204 28584 10220 28600
rect 10236 28584 10252 28600
rect 10268 28584 10284 28600
rect 10300 28584 10316 28600
rect 10332 28584 10348 28600
rect 10364 28584 10380 28600
rect 10396 28584 10412 28600
rect 10428 28584 10444 28600
rect 10460 28584 10476 28600
rect 10492 28584 10508 28600
rect 10524 28584 10540 28600
rect 10556 28584 10572 28600
rect 10588 28584 10604 28600
rect 10620 28584 10636 28600
rect 10652 28584 10668 28600
rect 10684 28584 10700 28600
rect 10716 28584 10732 28600
rect 10748 28584 10764 28600
rect 10780 28584 10796 28600
rect 10812 28584 10828 28600
rect 10844 28584 10860 28600
rect 10876 28584 10892 28600
rect 10908 28584 10924 28600
rect 10940 28584 10956 28600
rect 10972 28584 10988 28600
rect 11004 28584 11020 28600
rect 11036 28584 11052 28600
rect 11068 28584 11084 28600
rect 11100 28584 11116 28600
rect 11132 28584 11148 28600
rect 11164 28584 11180 28600
rect 11196 28584 11212 28600
rect 11228 28584 11244 28600
rect 11260 28584 11276 28600
rect 11292 28584 11308 28600
rect 11324 28584 11340 28600
rect 11356 28584 11372 28600
rect 11388 28584 11404 28600
rect 11420 28584 11436 28600
rect 11452 28584 11468 28600
rect 11484 28584 11500 28600
rect 11516 28584 11532 28600
rect 11548 28584 11564 28600
rect 11580 28584 11596 28600
rect 11612 28584 11628 28600
rect 11644 28584 11660 28600
rect 11676 28584 11692 28600
rect 11708 28584 11724 28600
rect 11740 28584 11756 28600
rect 11772 28584 11788 28600
rect 11804 28584 11820 28600
rect 9980 28552 9996 28568
rect 10012 28552 10028 28568
rect 10044 28552 10060 28568
rect 10076 28552 10092 28568
rect 10108 28552 10124 28568
rect 10140 28552 10156 28568
rect 10172 28552 10188 28568
rect 10204 28552 10220 28568
rect 10236 28552 10252 28568
rect 10268 28552 10284 28568
rect 10300 28552 10316 28568
rect 10332 28552 10348 28568
rect 10364 28552 10380 28568
rect 10396 28552 10412 28568
rect 10428 28552 10444 28568
rect 10460 28552 10476 28568
rect 10492 28552 10508 28568
rect 10524 28552 10540 28568
rect 10556 28552 10572 28568
rect 10588 28552 10604 28568
rect 10620 28552 10636 28568
rect 10652 28552 10668 28568
rect 10684 28552 10700 28568
rect 10716 28552 10732 28568
rect 10748 28552 10764 28568
rect 10780 28552 10796 28568
rect 10812 28552 10828 28568
rect 10844 28552 10860 28568
rect 10876 28552 10892 28568
rect 10908 28552 10924 28568
rect 10940 28552 10956 28568
rect 10972 28552 10988 28568
rect 11004 28552 11020 28568
rect 11036 28552 11052 28568
rect 11068 28552 11084 28568
rect 11100 28552 11116 28568
rect 11132 28552 11148 28568
rect 11164 28552 11180 28568
rect 11196 28552 11212 28568
rect 11228 28552 11244 28568
rect 11260 28552 11276 28568
rect 11292 28552 11308 28568
rect 11324 28552 11340 28568
rect 11356 28552 11372 28568
rect 11388 28552 11404 28568
rect 11420 28552 11436 28568
rect 11452 28552 11468 28568
rect 11484 28552 11500 28568
rect 11516 28552 11532 28568
rect 11548 28552 11564 28568
rect 11580 28552 11596 28568
rect 11612 28552 11628 28568
rect 11644 28552 11660 28568
rect 11676 28552 11692 28568
rect 11708 28552 11724 28568
rect 11740 28552 11756 28568
rect 11772 28552 11788 28568
rect 11804 28552 11820 28568
rect 9980 28520 9996 28536
rect 10012 28520 10028 28536
rect 10044 28520 10060 28536
rect 10076 28520 10092 28536
rect 10108 28520 10124 28536
rect 10140 28520 10156 28536
rect 10172 28520 10188 28536
rect 10204 28520 10220 28536
rect 10236 28520 10252 28536
rect 10268 28520 10284 28536
rect 10300 28520 10316 28536
rect 10332 28520 10348 28536
rect 10364 28520 10380 28536
rect 10396 28520 10412 28536
rect 10428 28520 10444 28536
rect 10460 28520 10476 28536
rect 10492 28520 10508 28536
rect 10524 28520 10540 28536
rect 10556 28520 10572 28536
rect 10588 28520 10604 28536
rect 10620 28520 10636 28536
rect 10652 28520 10668 28536
rect 10684 28520 10700 28536
rect 10716 28520 10732 28536
rect 10748 28520 10764 28536
rect 10780 28520 10796 28536
rect 10812 28520 10828 28536
rect 10844 28520 10860 28536
rect 10876 28520 10892 28536
rect 10908 28520 10924 28536
rect 10940 28520 10956 28536
rect 10972 28520 10988 28536
rect 11004 28520 11020 28536
rect 11036 28520 11052 28536
rect 11068 28520 11084 28536
rect 11100 28520 11116 28536
rect 11132 28520 11148 28536
rect 11164 28520 11180 28536
rect 11196 28520 11212 28536
rect 11228 28520 11244 28536
rect 11260 28520 11276 28536
rect 11292 28520 11308 28536
rect 11324 28520 11340 28536
rect 11356 28520 11372 28536
rect 11388 28520 11404 28536
rect 11420 28520 11436 28536
rect 11452 28520 11468 28536
rect 11484 28520 11500 28536
rect 11516 28520 11532 28536
rect 11548 28520 11564 28536
rect 11580 28520 11596 28536
rect 11612 28520 11628 28536
rect 11644 28520 11660 28536
rect 11676 28520 11692 28536
rect 11708 28520 11724 28536
rect 11740 28520 11756 28536
rect 11772 28520 11788 28536
rect 11804 28520 11820 28536
rect 9980 28488 9996 28504
rect 10012 28488 10028 28504
rect 10044 28488 10060 28504
rect 10076 28488 10092 28504
rect 10108 28488 10124 28504
rect 10140 28488 10156 28504
rect 10172 28488 10188 28504
rect 10204 28488 10220 28504
rect 10236 28488 10252 28504
rect 10268 28488 10284 28504
rect 10300 28488 10316 28504
rect 10332 28488 10348 28504
rect 10364 28488 10380 28504
rect 10396 28488 10412 28504
rect 10428 28488 10444 28504
rect 10460 28488 10476 28504
rect 10492 28488 10508 28504
rect 10524 28488 10540 28504
rect 10556 28488 10572 28504
rect 10588 28488 10604 28504
rect 10620 28488 10636 28504
rect 10652 28488 10668 28504
rect 10684 28488 10700 28504
rect 10716 28488 10732 28504
rect 10748 28488 10764 28504
rect 10780 28488 10796 28504
rect 10812 28488 10828 28504
rect 10844 28488 10860 28504
rect 10876 28488 10892 28504
rect 10908 28488 10924 28504
rect 10940 28488 10956 28504
rect 10972 28488 10988 28504
rect 11004 28488 11020 28504
rect 11036 28488 11052 28504
rect 11068 28488 11084 28504
rect 11100 28488 11116 28504
rect 11132 28488 11148 28504
rect 11164 28488 11180 28504
rect 11196 28488 11212 28504
rect 11228 28488 11244 28504
rect 11260 28488 11276 28504
rect 11292 28488 11308 28504
rect 11324 28488 11340 28504
rect 11356 28488 11372 28504
rect 11388 28488 11404 28504
rect 11420 28488 11436 28504
rect 11452 28488 11468 28504
rect 11484 28488 11500 28504
rect 11516 28488 11532 28504
rect 11548 28488 11564 28504
rect 11580 28488 11596 28504
rect 11612 28488 11628 28504
rect 11644 28488 11660 28504
rect 11676 28488 11692 28504
rect 11708 28488 11724 28504
rect 11740 28488 11756 28504
rect 11772 28488 11788 28504
rect 11804 28488 11820 28504
rect 9980 28456 9996 28472
rect 10012 28456 10028 28472
rect 10044 28456 10060 28472
rect 10076 28456 10092 28472
rect 10108 28456 10124 28472
rect 10140 28456 10156 28472
rect 10172 28456 10188 28472
rect 10204 28456 10220 28472
rect 10236 28456 10252 28472
rect 10268 28456 10284 28472
rect 10300 28456 10316 28472
rect 10332 28456 10348 28472
rect 10364 28456 10380 28472
rect 10396 28456 10412 28472
rect 10428 28456 10444 28472
rect 10460 28456 10476 28472
rect 10492 28456 10508 28472
rect 10524 28456 10540 28472
rect 10556 28456 10572 28472
rect 10588 28456 10604 28472
rect 10620 28456 10636 28472
rect 10652 28456 10668 28472
rect 10684 28456 10700 28472
rect 10716 28456 10732 28472
rect 10748 28456 10764 28472
rect 10780 28456 10796 28472
rect 10812 28456 10828 28472
rect 10844 28456 10860 28472
rect 10876 28456 10892 28472
rect 10908 28456 10924 28472
rect 10940 28456 10956 28472
rect 10972 28456 10988 28472
rect 11004 28456 11020 28472
rect 11036 28456 11052 28472
rect 11068 28456 11084 28472
rect 11100 28456 11116 28472
rect 11132 28456 11148 28472
rect 11164 28456 11180 28472
rect 11196 28456 11212 28472
rect 11228 28456 11244 28472
rect 11260 28456 11276 28472
rect 11292 28456 11308 28472
rect 11324 28456 11340 28472
rect 11356 28456 11372 28472
rect 11388 28456 11404 28472
rect 11420 28456 11436 28472
rect 11452 28456 11468 28472
rect 11484 28456 11500 28472
rect 11516 28456 11532 28472
rect 11548 28456 11564 28472
rect 11580 28456 11596 28472
rect 11612 28456 11628 28472
rect 11644 28456 11660 28472
rect 11676 28456 11692 28472
rect 11708 28456 11724 28472
rect 11740 28456 11756 28472
rect 11772 28456 11788 28472
rect 11804 28456 11820 28472
rect 9980 28424 9996 28440
rect 10012 28424 10028 28440
rect 10044 28424 10060 28440
rect 10076 28424 10092 28440
rect 10108 28424 10124 28440
rect 10140 28424 10156 28440
rect 10172 28424 10188 28440
rect 10204 28424 10220 28440
rect 10236 28424 10252 28440
rect 10268 28424 10284 28440
rect 10300 28424 10316 28440
rect 10332 28424 10348 28440
rect 10364 28424 10380 28440
rect 10396 28424 10412 28440
rect 10428 28424 10444 28440
rect 10460 28424 10476 28440
rect 10492 28424 10508 28440
rect 10524 28424 10540 28440
rect 10556 28424 10572 28440
rect 10588 28424 10604 28440
rect 10620 28424 10636 28440
rect 10652 28424 10668 28440
rect 10684 28424 10700 28440
rect 10716 28424 10732 28440
rect 10748 28424 10764 28440
rect 10780 28424 10796 28440
rect 10812 28424 10828 28440
rect 10844 28424 10860 28440
rect 10876 28424 10892 28440
rect 10908 28424 10924 28440
rect 10940 28424 10956 28440
rect 10972 28424 10988 28440
rect 11004 28424 11020 28440
rect 11036 28424 11052 28440
rect 11068 28424 11084 28440
rect 11100 28424 11116 28440
rect 11132 28424 11148 28440
rect 11164 28424 11180 28440
rect 11196 28424 11212 28440
rect 11228 28424 11244 28440
rect 11260 28424 11276 28440
rect 11292 28424 11308 28440
rect 11324 28424 11340 28440
rect 11356 28424 11372 28440
rect 11388 28424 11404 28440
rect 11420 28424 11436 28440
rect 11452 28424 11468 28440
rect 11484 28424 11500 28440
rect 11516 28424 11532 28440
rect 11548 28424 11564 28440
rect 11580 28424 11596 28440
rect 11612 28424 11628 28440
rect 11644 28424 11660 28440
rect 11676 28424 11692 28440
rect 11708 28424 11724 28440
rect 11740 28424 11756 28440
rect 11772 28424 11788 28440
rect 11804 28424 11820 28440
rect 9980 28392 9996 28408
rect 10012 28392 10028 28408
rect 10044 28392 10060 28408
rect 10076 28392 10092 28408
rect 10108 28392 10124 28408
rect 10140 28392 10156 28408
rect 10172 28392 10188 28408
rect 10204 28392 10220 28408
rect 10236 28392 10252 28408
rect 10268 28392 10284 28408
rect 10300 28392 10316 28408
rect 10332 28392 10348 28408
rect 10364 28392 10380 28408
rect 10396 28392 10412 28408
rect 10428 28392 10444 28408
rect 10460 28392 10476 28408
rect 10492 28392 10508 28408
rect 10524 28392 10540 28408
rect 10556 28392 10572 28408
rect 10588 28392 10604 28408
rect 10620 28392 10636 28408
rect 10652 28392 10668 28408
rect 10684 28392 10700 28408
rect 10716 28392 10732 28408
rect 10748 28392 10764 28408
rect 10780 28392 10796 28408
rect 10812 28392 10828 28408
rect 10844 28392 10860 28408
rect 10876 28392 10892 28408
rect 10908 28392 10924 28408
rect 10940 28392 10956 28408
rect 10972 28392 10988 28408
rect 11004 28392 11020 28408
rect 11036 28392 11052 28408
rect 11068 28392 11084 28408
rect 11100 28392 11116 28408
rect 11132 28392 11148 28408
rect 11164 28392 11180 28408
rect 11196 28392 11212 28408
rect 11228 28392 11244 28408
rect 11260 28392 11276 28408
rect 11292 28392 11308 28408
rect 11324 28392 11340 28408
rect 11356 28392 11372 28408
rect 11388 28392 11404 28408
rect 11420 28392 11436 28408
rect 11452 28392 11468 28408
rect 11484 28392 11500 28408
rect 11516 28392 11532 28408
rect 11548 28392 11564 28408
rect 11580 28392 11596 28408
rect 11612 28392 11628 28408
rect 11644 28392 11660 28408
rect 11676 28392 11692 28408
rect 11708 28392 11724 28408
rect 11740 28392 11756 28408
rect 11772 28392 11788 28408
rect 11804 28392 11820 28408
rect 9980 28360 9996 28376
rect 10012 28360 10028 28376
rect 10044 28360 10060 28376
rect 10076 28360 10092 28376
rect 10108 28360 10124 28376
rect 10140 28360 10156 28376
rect 10172 28360 10188 28376
rect 10204 28360 10220 28376
rect 10236 28360 10252 28376
rect 10268 28360 10284 28376
rect 10300 28360 10316 28376
rect 10332 28360 10348 28376
rect 10364 28360 10380 28376
rect 10396 28360 10412 28376
rect 10428 28360 10444 28376
rect 10460 28360 10476 28376
rect 10492 28360 10508 28376
rect 10524 28360 10540 28376
rect 10556 28360 10572 28376
rect 10588 28360 10604 28376
rect 10620 28360 10636 28376
rect 10652 28360 10668 28376
rect 10684 28360 10700 28376
rect 10716 28360 10732 28376
rect 10748 28360 10764 28376
rect 10780 28360 10796 28376
rect 10812 28360 10828 28376
rect 10844 28360 10860 28376
rect 10876 28360 10892 28376
rect 10908 28360 10924 28376
rect 10940 28360 10956 28376
rect 10972 28360 10988 28376
rect 11004 28360 11020 28376
rect 11036 28360 11052 28376
rect 11068 28360 11084 28376
rect 11100 28360 11116 28376
rect 11132 28360 11148 28376
rect 11164 28360 11180 28376
rect 11196 28360 11212 28376
rect 11228 28360 11244 28376
rect 11260 28360 11276 28376
rect 11292 28360 11308 28376
rect 11324 28360 11340 28376
rect 11356 28360 11372 28376
rect 11388 28360 11404 28376
rect 11420 28360 11436 28376
rect 11452 28360 11468 28376
rect 11484 28360 11500 28376
rect 11516 28360 11532 28376
rect 11548 28360 11564 28376
rect 11580 28360 11596 28376
rect 11612 28360 11628 28376
rect 11644 28360 11660 28376
rect 11676 28360 11692 28376
rect 11708 28360 11724 28376
rect 11740 28360 11756 28376
rect 11772 28360 11788 28376
rect 11804 28360 11820 28376
rect 9980 28328 9996 28344
rect 10012 28328 10028 28344
rect 10044 28328 10060 28344
rect 10076 28328 10092 28344
rect 10108 28328 10124 28344
rect 10140 28328 10156 28344
rect 10172 28328 10188 28344
rect 10204 28328 10220 28344
rect 10236 28328 10252 28344
rect 10268 28328 10284 28344
rect 10300 28328 10316 28344
rect 10332 28328 10348 28344
rect 10364 28328 10380 28344
rect 10396 28328 10412 28344
rect 10428 28328 10444 28344
rect 10460 28328 10476 28344
rect 10492 28328 10508 28344
rect 10524 28328 10540 28344
rect 10556 28328 10572 28344
rect 10588 28328 10604 28344
rect 10620 28328 10636 28344
rect 10652 28328 10668 28344
rect 10684 28328 10700 28344
rect 10716 28328 10732 28344
rect 10748 28328 10764 28344
rect 10780 28328 10796 28344
rect 10812 28328 10828 28344
rect 10844 28328 10860 28344
rect 10876 28328 10892 28344
rect 10908 28328 10924 28344
rect 10940 28328 10956 28344
rect 10972 28328 10988 28344
rect 11004 28328 11020 28344
rect 11036 28328 11052 28344
rect 11068 28328 11084 28344
rect 11100 28328 11116 28344
rect 11132 28328 11148 28344
rect 11164 28328 11180 28344
rect 11196 28328 11212 28344
rect 11228 28328 11244 28344
rect 11260 28328 11276 28344
rect 11292 28328 11308 28344
rect 11324 28328 11340 28344
rect 11356 28328 11372 28344
rect 11388 28328 11404 28344
rect 11420 28328 11436 28344
rect 11452 28328 11468 28344
rect 11484 28328 11500 28344
rect 11516 28328 11532 28344
rect 11548 28328 11564 28344
rect 11580 28328 11596 28344
rect 11612 28328 11628 28344
rect 11644 28328 11660 28344
rect 11676 28328 11692 28344
rect 11708 28328 11724 28344
rect 11740 28328 11756 28344
rect 11772 28328 11788 28344
rect 11804 28328 11820 28344
rect 9980 28296 9996 28312
rect 10012 28296 10028 28312
rect 10044 28296 10060 28312
rect 10076 28296 10092 28312
rect 10108 28296 10124 28312
rect 10140 28296 10156 28312
rect 10172 28296 10188 28312
rect 10204 28296 10220 28312
rect 10236 28296 10252 28312
rect 10268 28296 10284 28312
rect 10300 28296 10316 28312
rect 10332 28296 10348 28312
rect 10364 28296 10380 28312
rect 10396 28296 10412 28312
rect 10428 28296 10444 28312
rect 10460 28296 10476 28312
rect 10492 28296 10508 28312
rect 10524 28296 10540 28312
rect 10556 28296 10572 28312
rect 10588 28296 10604 28312
rect 10620 28296 10636 28312
rect 10652 28296 10668 28312
rect 10684 28296 10700 28312
rect 10716 28296 10732 28312
rect 10748 28296 10764 28312
rect 10780 28296 10796 28312
rect 10812 28296 10828 28312
rect 10844 28296 10860 28312
rect 10876 28296 10892 28312
rect 10908 28296 10924 28312
rect 10940 28296 10956 28312
rect 10972 28296 10988 28312
rect 11004 28296 11020 28312
rect 11036 28296 11052 28312
rect 11068 28296 11084 28312
rect 11100 28296 11116 28312
rect 11132 28296 11148 28312
rect 11164 28296 11180 28312
rect 11196 28296 11212 28312
rect 11228 28296 11244 28312
rect 11260 28296 11276 28312
rect 11292 28296 11308 28312
rect 11324 28296 11340 28312
rect 11356 28296 11372 28312
rect 11388 28296 11404 28312
rect 11420 28296 11436 28312
rect 11452 28296 11468 28312
rect 11484 28296 11500 28312
rect 11516 28296 11532 28312
rect 11548 28296 11564 28312
rect 11580 28296 11596 28312
rect 11612 28296 11628 28312
rect 11644 28296 11660 28312
rect 11676 28296 11692 28312
rect 11708 28296 11724 28312
rect 11740 28296 11756 28312
rect 11772 28296 11788 28312
rect 11804 28296 11820 28312
rect 9980 28264 9996 28280
rect 10012 28264 10028 28280
rect 10044 28264 10060 28280
rect 10076 28264 10092 28280
rect 10108 28264 10124 28280
rect 10140 28264 10156 28280
rect 10172 28264 10188 28280
rect 10204 28264 10220 28280
rect 10236 28264 10252 28280
rect 10268 28264 10284 28280
rect 10300 28264 10316 28280
rect 10332 28264 10348 28280
rect 10364 28264 10380 28280
rect 10396 28264 10412 28280
rect 10428 28264 10444 28280
rect 10460 28264 10476 28280
rect 10492 28264 10508 28280
rect 10524 28264 10540 28280
rect 10556 28264 10572 28280
rect 10588 28264 10604 28280
rect 10620 28264 10636 28280
rect 10652 28264 10668 28280
rect 10684 28264 10700 28280
rect 10716 28264 10732 28280
rect 10748 28264 10764 28280
rect 10780 28264 10796 28280
rect 10812 28264 10828 28280
rect 10844 28264 10860 28280
rect 10876 28264 10892 28280
rect 10908 28264 10924 28280
rect 10940 28264 10956 28280
rect 10972 28264 10988 28280
rect 11004 28264 11020 28280
rect 11036 28264 11052 28280
rect 11068 28264 11084 28280
rect 11100 28264 11116 28280
rect 11132 28264 11148 28280
rect 11164 28264 11180 28280
rect 11196 28264 11212 28280
rect 11228 28264 11244 28280
rect 11260 28264 11276 28280
rect 11292 28264 11308 28280
rect 11324 28264 11340 28280
rect 11356 28264 11372 28280
rect 11388 28264 11404 28280
rect 11420 28264 11436 28280
rect 11452 28264 11468 28280
rect 11484 28264 11500 28280
rect 11516 28264 11532 28280
rect 11548 28264 11564 28280
rect 11580 28264 11596 28280
rect 11612 28264 11628 28280
rect 11644 28264 11660 28280
rect 11676 28264 11692 28280
rect 11708 28264 11724 28280
rect 11740 28264 11756 28280
rect 11772 28264 11788 28280
rect 11804 28264 11820 28280
rect 9338 27748 9354 27764
rect 9370 27748 9386 27764
rect 9402 27748 9418 27764
rect 9434 27748 9450 27764
rect 9466 27748 9482 27764
rect 9498 27748 9514 27764
rect 9530 27748 9546 27764
rect 9562 27748 9578 27764
rect 9594 27748 9610 27764
rect 9626 27748 9642 27764
rect 9658 27748 9674 27764
rect 9690 27748 9706 27764
rect 9722 27748 9738 27764
rect 9754 27748 9770 27764
rect 9786 27748 9802 27764
rect 9338 27716 9354 27732
rect 9370 27716 9386 27732
rect 9402 27716 9418 27732
rect 9434 27716 9450 27732
rect 9466 27716 9482 27732
rect 9498 27716 9514 27732
rect 9530 27716 9546 27732
rect 9562 27716 9578 27732
rect 9594 27716 9610 27732
rect 9626 27716 9642 27732
rect 9658 27716 9674 27732
rect 9690 27716 9706 27732
rect 9722 27716 9738 27732
rect 9754 27716 9770 27732
rect 9786 27716 9802 27732
rect 9338 27684 9354 27700
rect 9370 27684 9386 27700
rect 9402 27684 9418 27700
rect 9434 27684 9450 27700
rect 9466 27684 9482 27700
rect 9498 27684 9514 27700
rect 9530 27684 9546 27700
rect 9562 27684 9578 27700
rect 9594 27684 9610 27700
rect 9626 27684 9642 27700
rect 9658 27684 9674 27700
rect 9690 27684 9706 27700
rect 9722 27684 9738 27700
rect 9754 27684 9770 27700
rect 9786 27684 9802 27700
rect 9338 27652 9354 27668
rect 9370 27652 9386 27668
rect 9402 27652 9418 27668
rect 9434 27652 9450 27668
rect 9466 27652 9482 27668
rect 9498 27652 9514 27668
rect 9530 27652 9546 27668
rect 9562 27652 9578 27668
rect 9594 27652 9610 27668
rect 9626 27652 9642 27668
rect 9658 27652 9674 27668
rect 9690 27652 9706 27668
rect 9722 27652 9738 27668
rect 9754 27652 9770 27668
rect 9786 27652 9802 27668
rect 9338 27620 9354 27636
rect 9370 27620 9386 27636
rect 9402 27620 9418 27636
rect 9434 27620 9450 27636
rect 9466 27620 9482 27636
rect 9498 27620 9514 27636
rect 9530 27620 9546 27636
rect 9562 27620 9578 27636
rect 9594 27620 9610 27636
rect 9626 27620 9642 27636
rect 9658 27620 9674 27636
rect 9690 27620 9706 27636
rect 9722 27620 9738 27636
rect 9754 27620 9770 27636
rect 9786 27620 9802 27636
rect 9338 27588 9354 27604
rect 9370 27588 9386 27604
rect 9402 27588 9418 27604
rect 9434 27588 9450 27604
rect 9466 27588 9482 27604
rect 9498 27588 9514 27604
rect 9530 27588 9546 27604
rect 9562 27588 9578 27604
rect 9594 27588 9610 27604
rect 9626 27588 9642 27604
rect 9658 27588 9674 27604
rect 9690 27588 9706 27604
rect 9722 27588 9738 27604
rect 9754 27588 9770 27604
rect 9786 27588 9802 27604
rect 9338 27556 9354 27572
rect 9370 27556 9386 27572
rect 9402 27556 9418 27572
rect 9434 27556 9450 27572
rect 9466 27556 9482 27572
rect 9498 27556 9514 27572
rect 9530 27556 9546 27572
rect 9562 27556 9578 27572
rect 9594 27556 9610 27572
rect 9626 27556 9642 27572
rect 9658 27556 9674 27572
rect 9690 27556 9706 27572
rect 9722 27556 9738 27572
rect 9754 27556 9770 27572
rect 9786 27556 9802 27572
rect 9338 27524 9354 27540
rect 9370 27524 9386 27540
rect 9402 27524 9418 27540
rect 9434 27524 9450 27540
rect 9466 27524 9482 27540
rect 9498 27524 9514 27540
rect 9530 27524 9546 27540
rect 9562 27524 9578 27540
rect 9594 27524 9610 27540
rect 9626 27524 9642 27540
rect 9658 27524 9674 27540
rect 9690 27524 9706 27540
rect 9722 27524 9738 27540
rect 9754 27524 9770 27540
rect 9786 27524 9802 27540
rect 9338 27492 9354 27508
rect 9370 27492 9386 27508
rect 9402 27492 9418 27508
rect 9434 27492 9450 27508
rect 9466 27492 9482 27508
rect 9498 27492 9514 27508
rect 9530 27492 9546 27508
rect 9562 27492 9578 27508
rect 9594 27492 9610 27508
rect 9626 27492 9642 27508
rect 9658 27492 9674 27508
rect 9690 27492 9706 27508
rect 9722 27492 9738 27508
rect 9754 27492 9770 27508
rect 9786 27492 9802 27508
rect 9338 27460 9354 27476
rect 9370 27460 9386 27476
rect 9402 27460 9418 27476
rect 9434 27460 9450 27476
rect 9466 27460 9482 27476
rect 9498 27460 9514 27476
rect 9530 27460 9546 27476
rect 9562 27460 9578 27476
rect 9594 27460 9610 27476
rect 9626 27460 9642 27476
rect 9658 27460 9674 27476
rect 9690 27460 9706 27476
rect 9722 27460 9738 27476
rect 9754 27460 9770 27476
rect 9786 27460 9802 27476
rect 9338 27428 9354 27444
rect 9370 27428 9386 27444
rect 9402 27428 9418 27444
rect 9434 27428 9450 27444
rect 9466 27428 9482 27444
rect 9498 27428 9514 27444
rect 9530 27428 9546 27444
rect 9562 27428 9578 27444
rect 9594 27428 9610 27444
rect 9626 27428 9642 27444
rect 9658 27428 9674 27444
rect 9690 27428 9706 27444
rect 9722 27428 9738 27444
rect 9754 27428 9770 27444
rect 9786 27428 9802 27444
rect 9338 27396 9354 27412
rect 9370 27396 9386 27412
rect 9402 27396 9418 27412
rect 9434 27396 9450 27412
rect 9466 27396 9482 27412
rect 9498 27396 9514 27412
rect 9530 27396 9546 27412
rect 9562 27396 9578 27412
rect 9594 27396 9610 27412
rect 9626 27396 9642 27412
rect 9658 27396 9674 27412
rect 9690 27396 9706 27412
rect 9722 27396 9738 27412
rect 9754 27396 9770 27412
rect 9786 27396 9802 27412
rect 9338 27364 9354 27380
rect 9370 27364 9386 27380
rect 9402 27364 9418 27380
rect 9434 27364 9450 27380
rect 9466 27364 9482 27380
rect 9498 27364 9514 27380
rect 9530 27364 9546 27380
rect 9562 27364 9578 27380
rect 9594 27364 9610 27380
rect 9626 27364 9642 27380
rect 9658 27364 9674 27380
rect 9690 27364 9706 27380
rect 9722 27364 9738 27380
rect 9754 27364 9770 27380
rect 9786 27364 9802 27380
rect 9338 27332 9354 27348
rect 9370 27332 9386 27348
rect 9402 27332 9418 27348
rect 9434 27332 9450 27348
rect 9466 27332 9482 27348
rect 9498 27332 9514 27348
rect 9530 27332 9546 27348
rect 9562 27332 9578 27348
rect 9594 27332 9610 27348
rect 9626 27332 9642 27348
rect 9658 27332 9674 27348
rect 9690 27332 9706 27348
rect 9722 27332 9738 27348
rect 9754 27332 9770 27348
rect 9786 27332 9802 27348
rect 9338 27300 9354 27316
rect 9370 27300 9386 27316
rect 9402 27300 9418 27316
rect 9434 27300 9450 27316
rect 9466 27300 9482 27316
rect 9498 27300 9514 27316
rect 9530 27300 9546 27316
rect 9562 27300 9578 27316
rect 9594 27300 9610 27316
rect 9626 27300 9642 27316
rect 9658 27300 9674 27316
rect 9690 27300 9706 27316
rect 9722 27300 9738 27316
rect 9754 27300 9770 27316
rect 9786 27300 9802 27316
rect 9338 27268 9354 27284
rect 9370 27268 9386 27284
rect 9402 27268 9418 27284
rect 9434 27268 9450 27284
rect 9466 27268 9482 27284
rect 9498 27268 9514 27284
rect 9530 27268 9546 27284
rect 9562 27268 9578 27284
rect 9594 27268 9610 27284
rect 9626 27268 9642 27284
rect 9658 27268 9674 27284
rect 9690 27268 9706 27284
rect 9722 27268 9738 27284
rect 9754 27268 9770 27284
rect 9786 27268 9802 27284
rect 9338 27236 9354 27252
rect 9370 27236 9386 27252
rect 9402 27236 9418 27252
rect 9434 27236 9450 27252
rect 9466 27236 9482 27252
rect 9498 27236 9514 27252
rect 9530 27236 9546 27252
rect 9562 27236 9578 27252
rect 9594 27236 9610 27252
rect 9626 27236 9642 27252
rect 9658 27236 9674 27252
rect 9690 27236 9706 27252
rect 9722 27236 9738 27252
rect 9754 27236 9770 27252
rect 9786 27236 9802 27252
rect 9338 27204 9354 27220
rect 9370 27204 9386 27220
rect 9402 27204 9418 27220
rect 9434 27204 9450 27220
rect 9466 27204 9482 27220
rect 9498 27204 9514 27220
rect 9530 27204 9546 27220
rect 9562 27204 9578 27220
rect 9594 27204 9610 27220
rect 9626 27204 9642 27220
rect 9658 27204 9674 27220
rect 9690 27204 9706 27220
rect 9722 27204 9738 27220
rect 9754 27204 9770 27220
rect 9786 27204 9802 27220
rect 9338 27172 9354 27188
rect 9370 27172 9386 27188
rect 9402 27172 9418 27188
rect 9434 27172 9450 27188
rect 9466 27172 9482 27188
rect 9498 27172 9514 27188
rect 9530 27172 9546 27188
rect 9562 27172 9578 27188
rect 9594 27172 9610 27188
rect 9626 27172 9642 27188
rect 9658 27172 9674 27188
rect 9690 27172 9706 27188
rect 9722 27172 9738 27188
rect 9754 27172 9770 27188
rect 9786 27172 9802 27188
rect 9338 27140 9354 27156
rect 9370 27140 9386 27156
rect 9402 27140 9418 27156
rect 9434 27140 9450 27156
rect 9466 27140 9482 27156
rect 9498 27140 9514 27156
rect 9530 27140 9546 27156
rect 9562 27140 9578 27156
rect 9594 27140 9610 27156
rect 9626 27140 9642 27156
rect 9658 27140 9674 27156
rect 9690 27140 9706 27156
rect 9722 27140 9738 27156
rect 9754 27140 9770 27156
rect 9786 27140 9802 27156
rect 9338 27108 9354 27124
rect 9370 27108 9386 27124
rect 9402 27108 9418 27124
rect 9434 27108 9450 27124
rect 9466 27108 9482 27124
rect 9498 27108 9514 27124
rect 9530 27108 9546 27124
rect 9562 27108 9578 27124
rect 9594 27108 9610 27124
rect 9626 27108 9642 27124
rect 9658 27108 9674 27124
rect 9690 27108 9706 27124
rect 9722 27108 9738 27124
rect 9754 27108 9770 27124
rect 9786 27108 9802 27124
rect 9338 27076 9354 27092
rect 9370 27076 9386 27092
rect 9402 27076 9418 27092
rect 9434 27076 9450 27092
rect 9466 27076 9482 27092
rect 9498 27076 9514 27092
rect 9530 27076 9546 27092
rect 9562 27076 9578 27092
rect 9594 27076 9610 27092
rect 9626 27076 9642 27092
rect 9658 27076 9674 27092
rect 9690 27076 9706 27092
rect 9722 27076 9738 27092
rect 9754 27076 9770 27092
rect 9786 27076 9802 27092
rect 9338 27044 9354 27060
rect 9370 27044 9386 27060
rect 9402 27044 9418 27060
rect 9434 27044 9450 27060
rect 9466 27044 9482 27060
rect 9498 27044 9514 27060
rect 9530 27044 9546 27060
rect 9562 27044 9578 27060
rect 9594 27044 9610 27060
rect 9626 27044 9642 27060
rect 9658 27044 9674 27060
rect 9690 27044 9706 27060
rect 9722 27044 9738 27060
rect 9754 27044 9770 27060
rect 9786 27044 9802 27060
rect 9338 27012 9354 27028
rect 9370 27012 9386 27028
rect 9402 27012 9418 27028
rect 9434 27012 9450 27028
rect 9466 27012 9482 27028
rect 9498 27012 9514 27028
rect 9530 27012 9546 27028
rect 9562 27012 9578 27028
rect 9594 27012 9610 27028
rect 9626 27012 9642 27028
rect 9658 27012 9674 27028
rect 9690 27012 9706 27028
rect 9722 27012 9738 27028
rect 9754 27012 9770 27028
rect 9786 27012 9802 27028
rect 9338 26980 9354 26996
rect 9370 26980 9386 26996
rect 9402 26980 9418 26996
rect 9434 26980 9450 26996
rect 9466 26980 9482 26996
rect 9498 26980 9514 26996
rect 9530 26980 9546 26996
rect 9562 26980 9578 26996
rect 9594 26980 9610 26996
rect 9626 26980 9642 26996
rect 9658 26980 9674 26996
rect 9690 26980 9706 26996
rect 9722 26980 9738 26996
rect 9754 26980 9770 26996
rect 9786 26980 9802 26996
rect 9338 26948 9354 26964
rect 9370 26948 9386 26964
rect 9402 26948 9418 26964
rect 9434 26948 9450 26964
rect 9466 26948 9482 26964
rect 9498 26948 9514 26964
rect 9530 26948 9546 26964
rect 9562 26948 9578 26964
rect 9594 26948 9610 26964
rect 9626 26948 9642 26964
rect 9658 26948 9674 26964
rect 9690 26948 9706 26964
rect 9722 26948 9738 26964
rect 9754 26948 9770 26964
rect 9786 26948 9802 26964
rect 9338 26916 9354 26932
rect 9370 26916 9386 26932
rect 9402 26916 9418 26932
rect 9434 26916 9450 26932
rect 9466 26916 9482 26932
rect 9498 26916 9514 26932
rect 9530 26916 9546 26932
rect 9562 26916 9578 26932
rect 9594 26916 9610 26932
rect 9626 26916 9642 26932
rect 9658 26916 9674 26932
rect 9690 26916 9706 26932
rect 9722 26916 9738 26932
rect 9754 26916 9770 26932
rect 9786 26916 9802 26932
rect 9338 26884 9354 26900
rect 9370 26884 9386 26900
rect 9402 26884 9418 26900
rect 9434 26884 9450 26900
rect 9466 26884 9482 26900
rect 9498 26884 9514 26900
rect 9530 26884 9546 26900
rect 9562 26884 9578 26900
rect 9594 26884 9610 26900
rect 9626 26884 9642 26900
rect 9658 26884 9674 26900
rect 9690 26884 9706 26900
rect 9722 26884 9738 26900
rect 9754 26884 9770 26900
rect 9786 26884 9802 26900
rect 9338 26852 9354 26868
rect 9370 26852 9386 26868
rect 9402 26852 9418 26868
rect 9434 26852 9450 26868
rect 9466 26852 9482 26868
rect 9498 26852 9514 26868
rect 9530 26852 9546 26868
rect 9562 26852 9578 26868
rect 9594 26852 9610 26868
rect 9626 26852 9642 26868
rect 9658 26852 9674 26868
rect 9690 26852 9706 26868
rect 9722 26852 9738 26868
rect 9754 26852 9770 26868
rect 9786 26852 9802 26868
rect 9338 26820 9354 26836
rect 9370 26820 9386 26836
rect 9402 26820 9418 26836
rect 9434 26820 9450 26836
rect 9466 26820 9482 26836
rect 9498 26820 9514 26836
rect 9530 26820 9546 26836
rect 9562 26820 9578 26836
rect 9594 26820 9610 26836
rect 9626 26820 9642 26836
rect 9658 26820 9674 26836
rect 9690 26820 9706 26836
rect 9722 26820 9738 26836
rect 9754 26820 9770 26836
rect 9786 26820 9802 26836
rect 9338 26788 9354 26804
rect 9370 26788 9386 26804
rect 9402 26788 9418 26804
rect 9434 26788 9450 26804
rect 9466 26788 9482 26804
rect 9498 26788 9514 26804
rect 9530 26788 9546 26804
rect 9562 26788 9578 26804
rect 9594 26788 9610 26804
rect 9626 26788 9642 26804
rect 9658 26788 9674 26804
rect 9690 26788 9706 26804
rect 9722 26788 9738 26804
rect 9754 26788 9770 26804
rect 9786 26788 9802 26804
rect 9338 26756 9354 26772
rect 9370 26756 9386 26772
rect 9402 26756 9418 26772
rect 9434 26756 9450 26772
rect 9466 26756 9482 26772
rect 9498 26756 9514 26772
rect 9530 26756 9546 26772
rect 9562 26756 9578 26772
rect 9594 26756 9610 26772
rect 9626 26756 9642 26772
rect 9658 26756 9674 26772
rect 9690 26756 9706 26772
rect 9722 26756 9738 26772
rect 9754 26756 9770 26772
rect 9786 26756 9802 26772
rect 9338 26724 9354 26740
rect 9370 26724 9386 26740
rect 9402 26724 9418 26740
rect 9434 26724 9450 26740
rect 9466 26724 9482 26740
rect 9498 26724 9514 26740
rect 9530 26724 9546 26740
rect 9562 26724 9578 26740
rect 9594 26724 9610 26740
rect 9626 26724 9642 26740
rect 9658 26724 9674 26740
rect 9690 26724 9706 26740
rect 9722 26724 9738 26740
rect 9754 26724 9770 26740
rect 9786 26724 9802 26740
rect 9338 26692 9354 26708
rect 9370 26692 9386 26708
rect 9402 26692 9418 26708
rect 9434 26692 9450 26708
rect 9466 26692 9482 26708
rect 9498 26692 9514 26708
rect 9530 26692 9546 26708
rect 9562 26692 9578 26708
rect 9594 26692 9610 26708
rect 9626 26692 9642 26708
rect 9658 26692 9674 26708
rect 9690 26692 9706 26708
rect 9722 26692 9738 26708
rect 9754 26692 9770 26708
rect 9786 26692 9802 26708
rect 9338 26660 9354 26676
rect 9370 26660 9386 26676
rect 9402 26660 9418 26676
rect 9434 26660 9450 26676
rect 9466 26660 9482 26676
rect 9498 26660 9514 26676
rect 9530 26660 9546 26676
rect 9562 26660 9578 26676
rect 9594 26660 9610 26676
rect 9626 26660 9642 26676
rect 9658 26660 9674 26676
rect 9690 26660 9706 26676
rect 9722 26660 9738 26676
rect 9754 26660 9770 26676
rect 9786 26660 9802 26676
rect 9338 26628 9354 26644
rect 9370 26628 9386 26644
rect 9402 26628 9418 26644
rect 9434 26628 9450 26644
rect 9466 26628 9482 26644
rect 9498 26628 9514 26644
rect 9530 26628 9546 26644
rect 9562 26628 9578 26644
rect 9594 26628 9610 26644
rect 9626 26628 9642 26644
rect 9658 26628 9674 26644
rect 9690 26628 9706 26644
rect 9722 26628 9738 26644
rect 9754 26628 9770 26644
rect 9786 26628 9802 26644
rect 9338 26596 9354 26612
rect 9370 26596 9386 26612
rect 9402 26596 9418 26612
rect 9434 26596 9450 26612
rect 9466 26596 9482 26612
rect 9498 26596 9514 26612
rect 9530 26596 9546 26612
rect 9562 26596 9578 26612
rect 9594 26596 9610 26612
rect 9626 26596 9642 26612
rect 9658 26596 9674 26612
rect 9690 26596 9706 26612
rect 9722 26596 9738 26612
rect 9754 26596 9770 26612
rect 9786 26596 9802 26612
rect 9338 26564 9354 26580
rect 9370 26564 9386 26580
rect 9402 26564 9418 26580
rect 9434 26564 9450 26580
rect 9466 26564 9482 26580
rect 9498 26564 9514 26580
rect 9530 26564 9546 26580
rect 9562 26564 9578 26580
rect 9594 26564 9610 26580
rect 9626 26564 9642 26580
rect 9658 26564 9674 26580
rect 9690 26564 9706 26580
rect 9722 26564 9738 26580
rect 9754 26564 9770 26580
rect 9786 26564 9802 26580
rect 9338 26532 9354 26548
rect 9370 26532 9386 26548
rect 9402 26532 9418 26548
rect 9434 26532 9450 26548
rect 9466 26532 9482 26548
rect 9498 26532 9514 26548
rect 9530 26532 9546 26548
rect 9562 26532 9578 26548
rect 9594 26532 9610 26548
rect 9626 26532 9642 26548
rect 9658 26532 9674 26548
rect 9690 26532 9706 26548
rect 9722 26532 9738 26548
rect 9754 26532 9770 26548
rect 9786 26532 9802 26548
rect 9338 26500 9354 26516
rect 9370 26500 9386 26516
rect 9402 26500 9418 26516
rect 9434 26500 9450 26516
rect 9466 26500 9482 26516
rect 9498 26500 9514 26516
rect 9530 26500 9546 26516
rect 9562 26500 9578 26516
rect 9594 26500 9610 26516
rect 9626 26500 9642 26516
rect 9658 26500 9674 26516
rect 9690 26500 9706 26516
rect 9722 26500 9738 26516
rect 9754 26500 9770 26516
rect 9786 26500 9802 26516
rect 9338 26468 9354 26484
rect 9370 26468 9386 26484
rect 9402 26468 9418 26484
rect 9434 26468 9450 26484
rect 9466 26468 9482 26484
rect 9498 26468 9514 26484
rect 9530 26468 9546 26484
rect 9562 26468 9578 26484
rect 9594 26468 9610 26484
rect 9626 26468 9642 26484
rect 9658 26468 9674 26484
rect 9690 26468 9706 26484
rect 9722 26468 9738 26484
rect 9754 26468 9770 26484
rect 9786 26468 9802 26484
rect 9338 26436 9354 26452
rect 9370 26436 9386 26452
rect 9402 26436 9418 26452
rect 9434 26436 9450 26452
rect 9466 26436 9482 26452
rect 9498 26436 9514 26452
rect 9530 26436 9546 26452
rect 9562 26436 9578 26452
rect 9594 26436 9610 26452
rect 9626 26436 9642 26452
rect 9658 26436 9674 26452
rect 9690 26436 9706 26452
rect 9722 26436 9738 26452
rect 9754 26436 9770 26452
rect 9786 26436 9802 26452
<< metal2 >>
rect 9960 28720 11840 29200
rect 9961 28696 11839 28720
rect 9961 28680 9980 28696
rect 9996 28680 10012 28696
rect 10028 28680 10044 28696
rect 10060 28680 10076 28696
rect 10092 28680 10108 28696
rect 10124 28680 10140 28696
rect 10156 28680 10172 28696
rect 10188 28680 10204 28696
rect 10220 28680 10236 28696
rect 10252 28680 10268 28696
rect 10284 28680 10300 28696
rect 10316 28680 10332 28696
rect 10348 28680 10364 28696
rect 10380 28680 10396 28696
rect 10412 28680 10428 28696
rect 10444 28680 10460 28696
rect 10476 28680 10492 28696
rect 10508 28680 10524 28696
rect 10540 28680 10556 28696
rect 10572 28680 10588 28696
rect 10604 28680 10620 28696
rect 10636 28680 10652 28696
rect 10668 28680 10684 28696
rect 10700 28680 10716 28696
rect 10732 28680 10748 28696
rect 10764 28680 10780 28696
rect 10796 28680 10812 28696
rect 10828 28680 10844 28696
rect 10860 28680 10876 28696
rect 10892 28680 10908 28696
rect 10924 28680 10940 28696
rect 10956 28680 10972 28696
rect 10988 28680 11004 28696
rect 11020 28680 11036 28696
rect 11052 28680 11068 28696
rect 11084 28680 11100 28696
rect 11116 28680 11132 28696
rect 11148 28680 11164 28696
rect 11180 28680 11196 28696
rect 11212 28680 11228 28696
rect 11244 28680 11260 28696
rect 11276 28680 11292 28696
rect 11308 28680 11324 28696
rect 11340 28680 11356 28696
rect 11372 28680 11388 28696
rect 11404 28680 11420 28696
rect 11436 28680 11452 28696
rect 11468 28680 11484 28696
rect 11500 28680 11516 28696
rect 11532 28680 11548 28696
rect 11564 28680 11580 28696
rect 11596 28680 11612 28696
rect 11628 28680 11644 28696
rect 11660 28680 11676 28696
rect 11692 28680 11708 28696
rect 11724 28680 11740 28696
rect 11756 28680 11772 28696
rect 11788 28680 11804 28696
rect 11820 28680 11839 28696
rect 9961 28664 11839 28680
rect 9961 28648 9980 28664
rect 9996 28648 10012 28664
rect 10028 28648 10044 28664
rect 10060 28648 10076 28664
rect 10092 28648 10108 28664
rect 10124 28648 10140 28664
rect 10156 28648 10172 28664
rect 10188 28648 10204 28664
rect 10220 28648 10236 28664
rect 10252 28648 10268 28664
rect 10284 28648 10300 28664
rect 10316 28648 10332 28664
rect 10348 28648 10364 28664
rect 10380 28648 10396 28664
rect 10412 28648 10428 28664
rect 10444 28648 10460 28664
rect 10476 28648 10492 28664
rect 10508 28648 10524 28664
rect 10540 28648 10556 28664
rect 10572 28648 10588 28664
rect 10604 28648 10620 28664
rect 10636 28648 10652 28664
rect 10668 28648 10684 28664
rect 10700 28648 10716 28664
rect 10732 28648 10748 28664
rect 10764 28648 10780 28664
rect 10796 28648 10812 28664
rect 10828 28648 10844 28664
rect 10860 28648 10876 28664
rect 10892 28648 10908 28664
rect 10924 28648 10940 28664
rect 10956 28648 10972 28664
rect 10988 28648 11004 28664
rect 11020 28648 11036 28664
rect 11052 28648 11068 28664
rect 11084 28648 11100 28664
rect 11116 28648 11132 28664
rect 11148 28648 11164 28664
rect 11180 28648 11196 28664
rect 11212 28648 11228 28664
rect 11244 28648 11260 28664
rect 11276 28648 11292 28664
rect 11308 28648 11324 28664
rect 11340 28648 11356 28664
rect 11372 28648 11388 28664
rect 11404 28648 11420 28664
rect 11436 28648 11452 28664
rect 11468 28648 11484 28664
rect 11500 28648 11516 28664
rect 11532 28648 11548 28664
rect 11564 28648 11580 28664
rect 11596 28648 11612 28664
rect 11628 28648 11644 28664
rect 11660 28648 11676 28664
rect 11692 28648 11708 28664
rect 11724 28648 11740 28664
rect 11756 28648 11772 28664
rect 11788 28648 11804 28664
rect 11820 28648 11839 28664
rect 9961 28632 11839 28648
rect 9961 28616 9980 28632
rect 9996 28616 10012 28632
rect 10028 28616 10044 28632
rect 10060 28616 10076 28632
rect 10092 28616 10108 28632
rect 10124 28616 10140 28632
rect 10156 28616 10172 28632
rect 10188 28616 10204 28632
rect 10220 28616 10236 28632
rect 10252 28616 10268 28632
rect 10284 28616 10300 28632
rect 10316 28616 10332 28632
rect 10348 28616 10364 28632
rect 10380 28616 10396 28632
rect 10412 28616 10428 28632
rect 10444 28616 10460 28632
rect 10476 28616 10492 28632
rect 10508 28616 10524 28632
rect 10540 28616 10556 28632
rect 10572 28616 10588 28632
rect 10604 28616 10620 28632
rect 10636 28616 10652 28632
rect 10668 28616 10684 28632
rect 10700 28616 10716 28632
rect 10732 28616 10748 28632
rect 10764 28616 10780 28632
rect 10796 28616 10812 28632
rect 10828 28616 10844 28632
rect 10860 28616 10876 28632
rect 10892 28616 10908 28632
rect 10924 28616 10940 28632
rect 10956 28616 10972 28632
rect 10988 28616 11004 28632
rect 11020 28616 11036 28632
rect 11052 28616 11068 28632
rect 11084 28616 11100 28632
rect 11116 28616 11132 28632
rect 11148 28616 11164 28632
rect 11180 28616 11196 28632
rect 11212 28616 11228 28632
rect 11244 28616 11260 28632
rect 11276 28616 11292 28632
rect 11308 28616 11324 28632
rect 11340 28616 11356 28632
rect 11372 28616 11388 28632
rect 11404 28616 11420 28632
rect 11436 28616 11452 28632
rect 11468 28616 11484 28632
rect 11500 28616 11516 28632
rect 11532 28616 11548 28632
rect 11564 28616 11580 28632
rect 11596 28616 11612 28632
rect 11628 28616 11644 28632
rect 11660 28616 11676 28632
rect 11692 28616 11708 28632
rect 11724 28616 11740 28632
rect 11756 28616 11772 28632
rect 11788 28616 11804 28632
rect 11820 28616 11839 28632
rect 9961 28600 11839 28616
rect 9961 28584 9980 28600
rect 9996 28584 10012 28600
rect 10028 28584 10044 28600
rect 10060 28584 10076 28600
rect 10092 28584 10108 28600
rect 10124 28584 10140 28600
rect 10156 28584 10172 28600
rect 10188 28584 10204 28600
rect 10220 28584 10236 28600
rect 10252 28584 10268 28600
rect 10284 28584 10300 28600
rect 10316 28584 10332 28600
rect 10348 28584 10364 28600
rect 10380 28584 10396 28600
rect 10412 28584 10428 28600
rect 10444 28584 10460 28600
rect 10476 28584 10492 28600
rect 10508 28584 10524 28600
rect 10540 28584 10556 28600
rect 10572 28584 10588 28600
rect 10604 28584 10620 28600
rect 10636 28584 10652 28600
rect 10668 28584 10684 28600
rect 10700 28584 10716 28600
rect 10732 28584 10748 28600
rect 10764 28584 10780 28600
rect 10796 28584 10812 28600
rect 10828 28584 10844 28600
rect 10860 28584 10876 28600
rect 10892 28584 10908 28600
rect 10924 28584 10940 28600
rect 10956 28584 10972 28600
rect 10988 28584 11004 28600
rect 11020 28584 11036 28600
rect 11052 28584 11068 28600
rect 11084 28584 11100 28600
rect 11116 28584 11132 28600
rect 11148 28584 11164 28600
rect 11180 28584 11196 28600
rect 11212 28584 11228 28600
rect 11244 28584 11260 28600
rect 11276 28584 11292 28600
rect 11308 28584 11324 28600
rect 11340 28584 11356 28600
rect 11372 28584 11388 28600
rect 11404 28584 11420 28600
rect 11436 28584 11452 28600
rect 11468 28584 11484 28600
rect 11500 28584 11516 28600
rect 11532 28584 11548 28600
rect 11564 28584 11580 28600
rect 11596 28584 11612 28600
rect 11628 28584 11644 28600
rect 11660 28584 11676 28600
rect 11692 28584 11708 28600
rect 11724 28584 11740 28600
rect 11756 28584 11772 28600
rect 11788 28584 11804 28600
rect 11820 28584 11839 28600
rect 9961 28568 11839 28584
rect 9961 28552 9980 28568
rect 9996 28552 10012 28568
rect 10028 28552 10044 28568
rect 10060 28552 10076 28568
rect 10092 28552 10108 28568
rect 10124 28552 10140 28568
rect 10156 28552 10172 28568
rect 10188 28552 10204 28568
rect 10220 28552 10236 28568
rect 10252 28552 10268 28568
rect 10284 28552 10300 28568
rect 10316 28552 10332 28568
rect 10348 28552 10364 28568
rect 10380 28552 10396 28568
rect 10412 28552 10428 28568
rect 10444 28552 10460 28568
rect 10476 28552 10492 28568
rect 10508 28552 10524 28568
rect 10540 28552 10556 28568
rect 10572 28552 10588 28568
rect 10604 28552 10620 28568
rect 10636 28552 10652 28568
rect 10668 28552 10684 28568
rect 10700 28552 10716 28568
rect 10732 28552 10748 28568
rect 10764 28552 10780 28568
rect 10796 28552 10812 28568
rect 10828 28552 10844 28568
rect 10860 28552 10876 28568
rect 10892 28552 10908 28568
rect 10924 28552 10940 28568
rect 10956 28552 10972 28568
rect 10988 28552 11004 28568
rect 11020 28552 11036 28568
rect 11052 28552 11068 28568
rect 11084 28552 11100 28568
rect 11116 28552 11132 28568
rect 11148 28552 11164 28568
rect 11180 28552 11196 28568
rect 11212 28552 11228 28568
rect 11244 28552 11260 28568
rect 11276 28552 11292 28568
rect 11308 28552 11324 28568
rect 11340 28552 11356 28568
rect 11372 28552 11388 28568
rect 11404 28552 11420 28568
rect 11436 28552 11452 28568
rect 11468 28552 11484 28568
rect 11500 28552 11516 28568
rect 11532 28552 11548 28568
rect 11564 28552 11580 28568
rect 11596 28552 11612 28568
rect 11628 28552 11644 28568
rect 11660 28552 11676 28568
rect 11692 28552 11708 28568
rect 11724 28552 11740 28568
rect 11756 28552 11772 28568
rect 11788 28552 11804 28568
rect 11820 28552 11839 28568
rect 9961 28536 11839 28552
rect 9961 28520 9980 28536
rect 9996 28520 10012 28536
rect 10028 28520 10044 28536
rect 10060 28520 10076 28536
rect 10092 28520 10108 28536
rect 10124 28520 10140 28536
rect 10156 28520 10172 28536
rect 10188 28520 10204 28536
rect 10220 28520 10236 28536
rect 10252 28520 10268 28536
rect 10284 28520 10300 28536
rect 10316 28520 10332 28536
rect 10348 28520 10364 28536
rect 10380 28520 10396 28536
rect 10412 28520 10428 28536
rect 10444 28520 10460 28536
rect 10476 28520 10492 28536
rect 10508 28520 10524 28536
rect 10540 28520 10556 28536
rect 10572 28520 10588 28536
rect 10604 28520 10620 28536
rect 10636 28520 10652 28536
rect 10668 28520 10684 28536
rect 10700 28520 10716 28536
rect 10732 28520 10748 28536
rect 10764 28520 10780 28536
rect 10796 28520 10812 28536
rect 10828 28520 10844 28536
rect 10860 28520 10876 28536
rect 10892 28520 10908 28536
rect 10924 28520 10940 28536
rect 10956 28520 10972 28536
rect 10988 28520 11004 28536
rect 11020 28520 11036 28536
rect 11052 28520 11068 28536
rect 11084 28520 11100 28536
rect 11116 28520 11132 28536
rect 11148 28520 11164 28536
rect 11180 28520 11196 28536
rect 11212 28520 11228 28536
rect 11244 28520 11260 28536
rect 11276 28520 11292 28536
rect 11308 28520 11324 28536
rect 11340 28520 11356 28536
rect 11372 28520 11388 28536
rect 11404 28520 11420 28536
rect 11436 28520 11452 28536
rect 11468 28520 11484 28536
rect 11500 28520 11516 28536
rect 11532 28520 11548 28536
rect 11564 28520 11580 28536
rect 11596 28520 11612 28536
rect 11628 28520 11644 28536
rect 11660 28520 11676 28536
rect 11692 28520 11708 28536
rect 11724 28520 11740 28536
rect 11756 28520 11772 28536
rect 11788 28520 11804 28536
rect 11820 28520 11839 28536
rect 9961 28504 11839 28520
rect 9961 28488 9980 28504
rect 9996 28488 10012 28504
rect 10028 28488 10044 28504
rect 10060 28488 10076 28504
rect 10092 28488 10108 28504
rect 10124 28488 10140 28504
rect 10156 28488 10172 28504
rect 10188 28488 10204 28504
rect 10220 28488 10236 28504
rect 10252 28488 10268 28504
rect 10284 28488 10300 28504
rect 10316 28488 10332 28504
rect 10348 28488 10364 28504
rect 10380 28488 10396 28504
rect 10412 28488 10428 28504
rect 10444 28488 10460 28504
rect 10476 28488 10492 28504
rect 10508 28488 10524 28504
rect 10540 28488 10556 28504
rect 10572 28488 10588 28504
rect 10604 28488 10620 28504
rect 10636 28488 10652 28504
rect 10668 28488 10684 28504
rect 10700 28488 10716 28504
rect 10732 28488 10748 28504
rect 10764 28488 10780 28504
rect 10796 28488 10812 28504
rect 10828 28488 10844 28504
rect 10860 28488 10876 28504
rect 10892 28488 10908 28504
rect 10924 28488 10940 28504
rect 10956 28488 10972 28504
rect 10988 28488 11004 28504
rect 11020 28488 11036 28504
rect 11052 28488 11068 28504
rect 11084 28488 11100 28504
rect 11116 28488 11132 28504
rect 11148 28488 11164 28504
rect 11180 28488 11196 28504
rect 11212 28488 11228 28504
rect 11244 28488 11260 28504
rect 11276 28488 11292 28504
rect 11308 28488 11324 28504
rect 11340 28488 11356 28504
rect 11372 28488 11388 28504
rect 11404 28488 11420 28504
rect 11436 28488 11452 28504
rect 11468 28488 11484 28504
rect 11500 28488 11516 28504
rect 11532 28488 11548 28504
rect 11564 28488 11580 28504
rect 11596 28488 11612 28504
rect 11628 28488 11644 28504
rect 11660 28488 11676 28504
rect 11692 28488 11708 28504
rect 11724 28488 11740 28504
rect 11756 28488 11772 28504
rect 11788 28488 11804 28504
rect 11820 28488 11839 28504
rect 9961 28472 11839 28488
rect 9961 28456 9980 28472
rect 9996 28456 10012 28472
rect 10028 28456 10044 28472
rect 10060 28456 10076 28472
rect 10092 28456 10108 28472
rect 10124 28456 10140 28472
rect 10156 28456 10172 28472
rect 10188 28456 10204 28472
rect 10220 28456 10236 28472
rect 10252 28456 10268 28472
rect 10284 28456 10300 28472
rect 10316 28456 10332 28472
rect 10348 28456 10364 28472
rect 10380 28456 10396 28472
rect 10412 28456 10428 28472
rect 10444 28456 10460 28472
rect 10476 28456 10492 28472
rect 10508 28456 10524 28472
rect 10540 28456 10556 28472
rect 10572 28456 10588 28472
rect 10604 28456 10620 28472
rect 10636 28456 10652 28472
rect 10668 28456 10684 28472
rect 10700 28456 10716 28472
rect 10732 28456 10748 28472
rect 10764 28456 10780 28472
rect 10796 28456 10812 28472
rect 10828 28456 10844 28472
rect 10860 28456 10876 28472
rect 10892 28456 10908 28472
rect 10924 28456 10940 28472
rect 10956 28456 10972 28472
rect 10988 28456 11004 28472
rect 11020 28456 11036 28472
rect 11052 28456 11068 28472
rect 11084 28456 11100 28472
rect 11116 28456 11132 28472
rect 11148 28456 11164 28472
rect 11180 28456 11196 28472
rect 11212 28456 11228 28472
rect 11244 28456 11260 28472
rect 11276 28456 11292 28472
rect 11308 28456 11324 28472
rect 11340 28456 11356 28472
rect 11372 28456 11388 28472
rect 11404 28456 11420 28472
rect 11436 28456 11452 28472
rect 11468 28456 11484 28472
rect 11500 28456 11516 28472
rect 11532 28456 11548 28472
rect 11564 28456 11580 28472
rect 11596 28456 11612 28472
rect 11628 28456 11644 28472
rect 11660 28456 11676 28472
rect 11692 28456 11708 28472
rect 11724 28456 11740 28472
rect 11756 28456 11772 28472
rect 11788 28456 11804 28472
rect 11820 28456 11839 28472
rect 9961 28440 11839 28456
rect 9961 28424 9980 28440
rect 9996 28424 10012 28440
rect 10028 28424 10044 28440
rect 10060 28424 10076 28440
rect 10092 28424 10108 28440
rect 10124 28424 10140 28440
rect 10156 28424 10172 28440
rect 10188 28424 10204 28440
rect 10220 28424 10236 28440
rect 10252 28424 10268 28440
rect 10284 28424 10300 28440
rect 10316 28424 10332 28440
rect 10348 28424 10364 28440
rect 10380 28424 10396 28440
rect 10412 28424 10428 28440
rect 10444 28424 10460 28440
rect 10476 28424 10492 28440
rect 10508 28424 10524 28440
rect 10540 28424 10556 28440
rect 10572 28424 10588 28440
rect 10604 28424 10620 28440
rect 10636 28424 10652 28440
rect 10668 28424 10684 28440
rect 10700 28424 10716 28440
rect 10732 28424 10748 28440
rect 10764 28424 10780 28440
rect 10796 28424 10812 28440
rect 10828 28424 10844 28440
rect 10860 28424 10876 28440
rect 10892 28424 10908 28440
rect 10924 28424 10940 28440
rect 10956 28424 10972 28440
rect 10988 28424 11004 28440
rect 11020 28424 11036 28440
rect 11052 28424 11068 28440
rect 11084 28424 11100 28440
rect 11116 28424 11132 28440
rect 11148 28424 11164 28440
rect 11180 28424 11196 28440
rect 11212 28424 11228 28440
rect 11244 28424 11260 28440
rect 11276 28424 11292 28440
rect 11308 28424 11324 28440
rect 11340 28424 11356 28440
rect 11372 28424 11388 28440
rect 11404 28424 11420 28440
rect 11436 28424 11452 28440
rect 11468 28424 11484 28440
rect 11500 28424 11516 28440
rect 11532 28424 11548 28440
rect 11564 28424 11580 28440
rect 11596 28424 11612 28440
rect 11628 28424 11644 28440
rect 11660 28424 11676 28440
rect 11692 28424 11708 28440
rect 11724 28424 11740 28440
rect 11756 28424 11772 28440
rect 11788 28424 11804 28440
rect 11820 28424 11839 28440
rect 9961 28408 11839 28424
rect 9961 28392 9980 28408
rect 9996 28392 10012 28408
rect 10028 28392 10044 28408
rect 10060 28392 10076 28408
rect 10092 28392 10108 28408
rect 10124 28392 10140 28408
rect 10156 28392 10172 28408
rect 10188 28392 10204 28408
rect 10220 28392 10236 28408
rect 10252 28392 10268 28408
rect 10284 28392 10300 28408
rect 10316 28392 10332 28408
rect 10348 28392 10364 28408
rect 10380 28392 10396 28408
rect 10412 28392 10428 28408
rect 10444 28392 10460 28408
rect 10476 28392 10492 28408
rect 10508 28392 10524 28408
rect 10540 28392 10556 28408
rect 10572 28392 10588 28408
rect 10604 28392 10620 28408
rect 10636 28392 10652 28408
rect 10668 28392 10684 28408
rect 10700 28392 10716 28408
rect 10732 28392 10748 28408
rect 10764 28392 10780 28408
rect 10796 28392 10812 28408
rect 10828 28392 10844 28408
rect 10860 28392 10876 28408
rect 10892 28392 10908 28408
rect 10924 28392 10940 28408
rect 10956 28392 10972 28408
rect 10988 28392 11004 28408
rect 11020 28392 11036 28408
rect 11052 28392 11068 28408
rect 11084 28392 11100 28408
rect 11116 28392 11132 28408
rect 11148 28392 11164 28408
rect 11180 28392 11196 28408
rect 11212 28392 11228 28408
rect 11244 28392 11260 28408
rect 11276 28392 11292 28408
rect 11308 28392 11324 28408
rect 11340 28392 11356 28408
rect 11372 28392 11388 28408
rect 11404 28392 11420 28408
rect 11436 28392 11452 28408
rect 11468 28392 11484 28408
rect 11500 28392 11516 28408
rect 11532 28392 11548 28408
rect 11564 28392 11580 28408
rect 11596 28392 11612 28408
rect 11628 28392 11644 28408
rect 11660 28392 11676 28408
rect 11692 28392 11708 28408
rect 11724 28392 11740 28408
rect 11756 28392 11772 28408
rect 11788 28392 11804 28408
rect 11820 28392 11839 28408
rect 9961 28376 11839 28392
rect 9961 28360 9980 28376
rect 9996 28360 10012 28376
rect 10028 28360 10044 28376
rect 10060 28360 10076 28376
rect 10092 28360 10108 28376
rect 10124 28360 10140 28376
rect 10156 28360 10172 28376
rect 10188 28360 10204 28376
rect 10220 28360 10236 28376
rect 10252 28360 10268 28376
rect 10284 28360 10300 28376
rect 10316 28360 10332 28376
rect 10348 28360 10364 28376
rect 10380 28360 10396 28376
rect 10412 28360 10428 28376
rect 10444 28360 10460 28376
rect 10476 28360 10492 28376
rect 10508 28360 10524 28376
rect 10540 28360 10556 28376
rect 10572 28360 10588 28376
rect 10604 28360 10620 28376
rect 10636 28360 10652 28376
rect 10668 28360 10684 28376
rect 10700 28360 10716 28376
rect 10732 28360 10748 28376
rect 10764 28360 10780 28376
rect 10796 28360 10812 28376
rect 10828 28360 10844 28376
rect 10860 28360 10876 28376
rect 10892 28360 10908 28376
rect 10924 28360 10940 28376
rect 10956 28360 10972 28376
rect 10988 28360 11004 28376
rect 11020 28360 11036 28376
rect 11052 28360 11068 28376
rect 11084 28360 11100 28376
rect 11116 28360 11132 28376
rect 11148 28360 11164 28376
rect 11180 28360 11196 28376
rect 11212 28360 11228 28376
rect 11244 28360 11260 28376
rect 11276 28360 11292 28376
rect 11308 28360 11324 28376
rect 11340 28360 11356 28376
rect 11372 28360 11388 28376
rect 11404 28360 11420 28376
rect 11436 28360 11452 28376
rect 11468 28360 11484 28376
rect 11500 28360 11516 28376
rect 11532 28360 11548 28376
rect 11564 28360 11580 28376
rect 11596 28360 11612 28376
rect 11628 28360 11644 28376
rect 11660 28360 11676 28376
rect 11692 28360 11708 28376
rect 11724 28360 11740 28376
rect 11756 28360 11772 28376
rect 11788 28360 11804 28376
rect 11820 28360 11839 28376
rect 9961 28344 11839 28360
rect 9961 28328 9980 28344
rect 9996 28328 10012 28344
rect 10028 28328 10044 28344
rect 10060 28328 10076 28344
rect 10092 28328 10108 28344
rect 10124 28328 10140 28344
rect 10156 28328 10172 28344
rect 10188 28328 10204 28344
rect 10220 28328 10236 28344
rect 10252 28328 10268 28344
rect 10284 28328 10300 28344
rect 10316 28328 10332 28344
rect 10348 28328 10364 28344
rect 10380 28328 10396 28344
rect 10412 28328 10428 28344
rect 10444 28328 10460 28344
rect 10476 28328 10492 28344
rect 10508 28328 10524 28344
rect 10540 28328 10556 28344
rect 10572 28328 10588 28344
rect 10604 28328 10620 28344
rect 10636 28328 10652 28344
rect 10668 28328 10684 28344
rect 10700 28328 10716 28344
rect 10732 28328 10748 28344
rect 10764 28328 10780 28344
rect 10796 28328 10812 28344
rect 10828 28328 10844 28344
rect 10860 28328 10876 28344
rect 10892 28328 10908 28344
rect 10924 28328 10940 28344
rect 10956 28328 10972 28344
rect 10988 28328 11004 28344
rect 11020 28328 11036 28344
rect 11052 28328 11068 28344
rect 11084 28328 11100 28344
rect 11116 28328 11132 28344
rect 11148 28328 11164 28344
rect 11180 28328 11196 28344
rect 11212 28328 11228 28344
rect 11244 28328 11260 28344
rect 11276 28328 11292 28344
rect 11308 28328 11324 28344
rect 11340 28328 11356 28344
rect 11372 28328 11388 28344
rect 11404 28328 11420 28344
rect 11436 28328 11452 28344
rect 11468 28328 11484 28344
rect 11500 28328 11516 28344
rect 11532 28328 11548 28344
rect 11564 28328 11580 28344
rect 11596 28328 11612 28344
rect 11628 28328 11644 28344
rect 11660 28328 11676 28344
rect 11692 28328 11708 28344
rect 11724 28328 11740 28344
rect 11756 28328 11772 28344
rect 11788 28328 11804 28344
rect 11820 28328 11839 28344
rect 9961 28312 11839 28328
rect 9961 28296 9980 28312
rect 9996 28296 10012 28312
rect 10028 28296 10044 28312
rect 10060 28296 10076 28312
rect 10092 28296 10108 28312
rect 10124 28296 10140 28312
rect 10156 28296 10172 28312
rect 10188 28296 10204 28312
rect 10220 28296 10236 28312
rect 10252 28296 10268 28312
rect 10284 28296 10300 28312
rect 10316 28296 10332 28312
rect 10348 28296 10364 28312
rect 10380 28296 10396 28312
rect 10412 28296 10428 28312
rect 10444 28296 10460 28312
rect 10476 28296 10492 28312
rect 10508 28296 10524 28312
rect 10540 28296 10556 28312
rect 10572 28296 10588 28312
rect 10604 28296 10620 28312
rect 10636 28296 10652 28312
rect 10668 28296 10684 28312
rect 10700 28296 10716 28312
rect 10732 28296 10748 28312
rect 10764 28296 10780 28312
rect 10796 28296 10812 28312
rect 10828 28296 10844 28312
rect 10860 28296 10876 28312
rect 10892 28296 10908 28312
rect 10924 28296 10940 28312
rect 10956 28296 10972 28312
rect 10988 28296 11004 28312
rect 11020 28296 11036 28312
rect 11052 28296 11068 28312
rect 11084 28296 11100 28312
rect 11116 28296 11132 28312
rect 11148 28296 11164 28312
rect 11180 28296 11196 28312
rect 11212 28296 11228 28312
rect 11244 28296 11260 28312
rect 11276 28296 11292 28312
rect 11308 28296 11324 28312
rect 11340 28296 11356 28312
rect 11372 28296 11388 28312
rect 11404 28296 11420 28312
rect 11436 28296 11452 28312
rect 11468 28296 11484 28312
rect 11500 28296 11516 28312
rect 11532 28296 11548 28312
rect 11564 28296 11580 28312
rect 11596 28296 11612 28312
rect 11628 28296 11644 28312
rect 11660 28296 11676 28312
rect 11692 28296 11708 28312
rect 11724 28296 11740 28312
rect 11756 28296 11772 28312
rect 11788 28296 11804 28312
rect 11820 28296 11839 28312
rect 9961 28280 11839 28296
rect 9961 28264 9980 28280
rect 9996 28264 10012 28280
rect 10028 28264 10044 28280
rect 10060 28264 10076 28280
rect 10092 28264 10108 28280
rect 10124 28264 10140 28280
rect 10156 28264 10172 28280
rect 10188 28264 10204 28280
rect 10220 28264 10236 28280
rect 10252 28264 10268 28280
rect 10284 28264 10300 28280
rect 10316 28264 10332 28280
rect 10348 28264 10364 28280
rect 10380 28264 10396 28280
rect 10412 28264 10428 28280
rect 10444 28264 10460 28280
rect 10476 28264 10492 28280
rect 10508 28264 10524 28280
rect 10540 28264 10556 28280
rect 10572 28264 10588 28280
rect 10604 28264 10620 28280
rect 10636 28264 10652 28280
rect 10668 28264 10684 28280
rect 10700 28264 10716 28280
rect 10732 28264 10748 28280
rect 10764 28264 10780 28280
rect 10796 28264 10812 28280
rect 10828 28264 10844 28280
rect 10860 28264 10876 28280
rect 10892 28264 10908 28280
rect 10924 28264 10940 28280
rect 10956 28264 10972 28280
rect 10988 28264 11004 28280
rect 11020 28264 11036 28280
rect 11052 28264 11068 28280
rect 11084 28264 11100 28280
rect 11116 28264 11132 28280
rect 11148 28264 11164 28280
rect 11180 28264 11196 28280
rect 11212 28264 11228 28280
rect 11244 28264 11260 28280
rect 11276 28264 11292 28280
rect 11308 28264 11324 28280
rect 11340 28264 11356 28280
rect 11372 28264 11388 28280
rect 11404 28264 11420 28280
rect 11436 28264 11452 28280
rect 11468 28264 11484 28280
rect 11500 28264 11516 28280
rect 11532 28264 11548 28280
rect 11564 28264 11580 28280
rect 11596 28264 11612 28280
rect 11628 28264 11644 28280
rect 11660 28264 11676 28280
rect 11692 28264 11708 28280
rect 11724 28264 11740 28280
rect 11756 28264 11772 28280
rect 11788 28264 11804 28280
rect 11820 28264 11839 28280
rect 9961 28241 11839 28264
rect 8820 27779 9320 27780
rect 8820 27764 9819 27779
rect 8820 27748 9338 27764
rect 9354 27748 9370 27764
rect 9386 27748 9402 27764
rect 9418 27748 9434 27764
rect 9450 27748 9466 27764
rect 9482 27748 9498 27764
rect 9514 27748 9530 27764
rect 9546 27748 9562 27764
rect 9578 27748 9594 27764
rect 9610 27748 9626 27764
rect 9642 27748 9658 27764
rect 9674 27748 9690 27764
rect 9706 27748 9722 27764
rect 9738 27748 9754 27764
rect 9770 27748 9786 27764
rect 9802 27748 9819 27764
rect 8820 27732 9819 27748
rect 8820 27716 9338 27732
rect 9354 27716 9370 27732
rect 9386 27716 9402 27732
rect 9418 27716 9434 27732
rect 9450 27716 9466 27732
rect 9482 27716 9498 27732
rect 9514 27716 9530 27732
rect 9546 27716 9562 27732
rect 9578 27716 9594 27732
rect 9610 27716 9626 27732
rect 9642 27716 9658 27732
rect 9674 27716 9690 27732
rect 9706 27716 9722 27732
rect 9738 27716 9754 27732
rect 9770 27716 9786 27732
rect 9802 27716 9819 27732
rect 8820 27700 9819 27716
rect 8820 27684 9338 27700
rect 9354 27684 9370 27700
rect 9386 27684 9402 27700
rect 9418 27684 9434 27700
rect 9450 27684 9466 27700
rect 9482 27684 9498 27700
rect 9514 27684 9530 27700
rect 9546 27684 9562 27700
rect 9578 27684 9594 27700
rect 9610 27684 9626 27700
rect 9642 27684 9658 27700
rect 9674 27684 9690 27700
rect 9706 27684 9722 27700
rect 9738 27684 9754 27700
rect 9770 27684 9786 27700
rect 9802 27684 9819 27700
rect 8820 27668 9819 27684
rect 8820 27652 9338 27668
rect 9354 27652 9370 27668
rect 9386 27652 9402 27668
rect 9418 27652 9434 27668
rect 9450 27652 9466 27668
rect 9482 27652 9498 27668
rect 9514 27652 9530 27668
rect 9546 27652 9562 27668
rect 9578 27652 9594 27668
rect 9610 27652 9626 27668
rect 9642 27652 9658 27668
rect 9674 27652 9690 27668
rect 9706 27652 9722 27668
rect 9738 27652 9754 27668
rect 9770 27652 9786 27668
rect 9802 27652 9819 27668
rect 8820 27636 9819 27652
rect 8820 27620 9338 27636
rect 9354 27620 9370 27636
rect 9386 27620 9402 27636
rect 9418 27620 9434 27636
rect 9450 27620 9466 27636
rect 9482 27620 9498 27636
rect 9514 27620 9530 27636
rect 9546 27620 9562 27636
rect 9578 27620 9594 27636
rect 9610 27620 9626 27636
rect 9642 27620 9658 27636
rect 9674 27620 9690 27636
rect 9706 27620 9722 27636
rect 9738 27620 9754 27636
rect 9770 27620 9786 27636
rect 9802 27620 9819 27636
rect 8820 27604 9819 27620
rect 8820 27588 9338 27604
rect 9354 27588 9370 27604
rect 9386 27588 9402 27604
rect 9418 27588 9434 27604
rect 9450 27588 9466 27604
rect 9482 27588 9498 27604
rect 9514 27588 9530 27604
rect 9546 27588 9562 27604
rect 9578 27588 9594 27604
rect 9610 27588 9626 27604
rect 9642 27588 9658 27604
rect 9674 27588 9690 27604
rect 9706 27588 9722 27604
rect 9738 27588 9754 27604
rect 9770 27588 9786 27604
rect 9802 27588 9819 27604
rect 8820 27572 9819 27588
rect 8820 27556 9338 27572
rect 9354 27556 9370 27572
rect 9386 27556 9402 27572
rect 9418 27556 9434 27572
rect 9450 27556 9466 27572
rect 9482 27556 9498 27572
rect 9514 27556 9530 27572
rect 9546 27556 9562 27572
rect 9578 27556 9594 27572
rect 9610 27556 9626 27572
rect 9642 27556 9658 27572
rect 9674 27556 9690 27572
rect 9706 27556 9722 27572
rect 9738 27556 9754 27572
rect 9770 27556 9786 27572
rect 9802 27556 9819 27572
rect 8820 27540 9819 27556
rect 8820 27524 9338 27540
rect 9354 27524 9370 27540
rect 9386 27524 9402 27540
rect 9418 27524 9434 27540
rect 9450 27524 9466 27540
rect 9482 27524 9498 27540
rect 9514 27524 9530 27540
rect 9546 27524 9562 27540
rect 9578 27524 9594 27540
rect 9610 27524 9626 27540
rect 9642 27524 9658 27540
rect 9674 27524 9690 27540
rect 9706 27524 9722 27540
rect 9738 27524 9754 27540
rect 9770 27524 9786 27540
rect 9802 27524 9819 27540
rect 8820 27508 9819 27524
rect 8820 27492 9338 27508
rect 9354 27492 9370 27508
rect 9386 27492 9402 27508
rect 9418 27492 9434 27508
rect 9450 27492 9466 27508
rect 9482 27492 9498 27508
rect 9514 27492 9530 27508
rect 9546 27492 9562 27508
rect 9578 27492 9594 27508
rect 9610 27492 9626 27508
rect 9642 27492 9658 27508
rect 9674 27492 9690 27508
rect 9706 27492 9722 27508
rect 9738 27492 9754 27508
rect 9770 27492 9786 27508
rect 9802 27492 9819 27508
rect 8820 27476 9819 27492
rect 8820 27460 9338 27476
rect 9354 27460 9370 27476
rect 9386 27460 9402 27476
rect 9418 27460 9434 27476
rect 9450 27460 9466 27476
rect 9482 27460 9498 27476
rect 9514 27460 9530 27476
rect 9546 27460 9562 27476
rect 9578 27460 9594 27476
rect 9610 27460 9626 27476
rect 9642 27460 9658 27476
rect 9674 27460 9690 27476
rect 9706 27460 9722 27476
rect 9738 27460 9754 27476
rect 9770 27460 9786 27476
rect 9802 27460 9819 27476
rect 8820 27444 9819 27460
rect 8820 27428 9338 27444
rect 9354 27428 9370 27444
rect 9386 27428 9402 27444
rect 9418 27428 9434 27444
rect 9450 27428 9466 27444
rect 9482 27428 9498 27444
rect 9514 27428 9530 27444
rect 9546 27428 9562 27444
rect 9578 27428 9594 27444
rect 9610 27428 9626 27444
rect 9642 27428 9658 27444
rect 9674 27428 9690 27444
rect 9706 27428 9722 27444
rect 9738 27428 9754 27444
rect 9770 27428 9786 27444
rect 9802 27428 9819 27444
rect 8820 27412 9819 27428
rect 8820 27396 9338 27412
rect 9354 27396 9370 27412
rect 9386 27396 9402 27412
rect 9418 27396 9434 27412
rect 9450 27396 9466 27412
rect 9482 27396 9498 27412
rect 9514 27396 9530 27412
rect 9546 27396 9562 27412
rect 9578 27396 9594 27412
rect 9610 27396 9626 27412
rect 9642 27396 9658 27412
rect 9674 27396 9690 27412
rect 9706 27396 9722 27412
rect 9738 27396 9754 27412
rect 9770 27396 9786 27412
rect 9802 27396 9819 27412
rect 8820 27380 9819 27396
rect 8820 27364 9338 27380
rect 9354 27364 9370 27380
rect 9386 27364 9402 27380
rect 9418 27364 9434 27380
rect 9450 27364 9466 27380
rect 9482 27364 9498 27380
rect 9514 27364 9530 27380
rect 9546 27364 9562 27380
rect 9578 27364 9594 27380
rect 9610 27364 9626 27380
rect 9642 27364 9658 27380
rect 9674 27364 9690 27380
rect 9706 27364 9722 27380
rect 9738 27364 9754 27380
rect 9770 27364 9786 27380
rect 9802 27364 9819 27380
rect 8820 27348 9819 27364
rect 8820 27332 9338 27348
rect 9354 27332 9370 27348
rect 9386 27332 9402 27348
rect 9418 27332 9434 27348
rect 9450 27332 9466 27348
rect 9482 27332 9498 27348
rect 9514 27332 9530 27348
rect 9546 27332 9562 27348
rect 9578 27332 9594 27348
rect 9610 27332 9626 27348
rect 9642 27332 9658 27348
rect 9674 27332 9690 27348
rect 9706 27332 9722 27348
rect 9738 27332 9754 27348
rect 9770 27332 9786 27348
rect 9802 27332 9819 27348
rect 8820 27316 9819 27332
rect 8820 27300 9338 27316
rect 9354 27300 9370 27316
rect 9386 27300 9402 27316
rect 9418 27300 9434 27316
rect 9450 27300 9466 27316
rect 9482 27300 9498 27316
rect 9514 27300 9530 27316
rect 9546 27300 9562 27316
rect 9578 27300 9594 27316
rect 9610 27300 9626 27316
rect 9642 27300 9658 27316
rect 9674 27300 9690 27316
rect 9706 27300 9722 27316
rect 9738 27300 9754 27316
rect 9770 27300 9786 27316
rect 9802 27300 9819 27316
rect 8820 27284 9819 27300
rect 8820 27268 9338 27284
rect 9354 27268 9370 27284
rect 9386 27268 9402 27284
rect 9418 27268 9434 27284
rect 9450 27268 9466 27284
rect 9482 27268 9498 27284
rect 9514 27268 9530 27284
rect 9546 27268 9562 27284
rect 9578 27268 9594 27284
rect 9610 27268 9626 27284
rect 9642 27268 9658 27284
rect 9674 27268 9690 27284
rect 9706 27268 9722 27284
rect 9738 27268 9754 27284
rect 9770 27268 9786 27284
rect 9802 27268 9819 27284
rect 8820 27252 9819 27268
rect 8820 27236 9338 27252
rect 9354 27236 9370 27252
rect 9386 27236 9402 27252
rect 9418 27236 9434 27252
rect 9450 27236 9466 27252
rect 9482 27236 9498 27252
rect 9514 27236 9530 27252
rect 9546 27236 9562 27252
rect 9578 27236 9594 27252
rect 9610 27236 9626 27252
rect 9642 27236 9658 27252
rect 9674 27236 9690 27252
rect 9706 27236 9722 27252
rect 9738 27236 9754 27252
rect 9770 27236 9786 27252
rect 9802 27236 9819 27252
rect 8820 27220 9819 27236
rect 8820 27204 9338 27220
rect 9354 27204 9370 27220
rect 9386 27204 9402 27220
rect 9418 27204 9434 27220
rect 9450 27204 9466 27220
rect 9482 27204 9498 27220
rect 9514 27204 9530 27220
rect 9546 27204 9562 27220
rect 9578 27204 9594 27220
rect 9610 27204 9626 27220
rect 9642 27204 9658 27220
rect 9674 27204 9690 27220
rect 9706 27204 9722 27220
rect 9738 27204 9754 27220
rect 9770 27204 9786 27220
rect 9802 27204 9819 27220
rect 8820 27188 9819 27204
rect 8820 27172 9338 27188
rect 9354 27172 9370 27188
rect 9386 27172 9402 27188
rect 9418 27172 9434 27188
rect 9450 27172 9466 27188
rect 9482 27172 9498 27188
rect 9514 27172 9530 27188
rect 9546 27172 9562 27188
rect 9578 27172 9594 27188
rect 9610 27172 9626 27188
rect 9642 27172 9658 27188
rect 9674 27172 9690 27188
rect 9706 27172 9722 27188
rect 9738 27172 9754 27188
rect 9770 27172 9786 27188
rect 9802 27172 9819 27188
rect 8820 27156 9819 27172
rect 8820 27140 9338 27156
rect 9354 27140 9370 27156
rect 9386 27140 9402 27156
rect 9418 27140 9434 27156
rect 9450 27140 9466 27156
rect 9482 27140 9498 27156
rect 9514 27140 9530 27156
rect 9546 27140 9562 27156
rect 9578 27140 9594 27156
rect 9610 27140 9626 27156
rect 9642 27140 9658 27156
rect 9674 27140 9690 27156
rect 9706 27140 9722 27156
rect 9738 27140 9754 27156
rect 9770 27140 9786 27156
rect 9802 27140 9819 27156
rect 8820 27124 9819 27140
rect 8820 27108 9338 27124
rect 9354 27108 9370 27124
rect 9386 27108 9402 27124
rect 9418 27108 9434 27124
rect 9450 27108 9466 27124
rect 9482 27108 9498 27124
rect 9514 27108 9530 27124
rect 9546 27108 9562 27124
rect 9578 27108 9594 27124
rect 9610 27108 9626 27124
rect 9642 27108 9658 27124
rect 9674 27108 9690 27124
rect 9706 27108 9722 27124
rect 9738 27108 9754 27124
rect 9770 27108 9786 27124
rect 9802 27108 9819 27124
rect 8820 27092 9819 27108
rect 8820 27076 9338 27092
rect 9354 27076 9370 27092
rect 9386 27076 9402 27092
rect 9418 27076 9434 27092
rect 9450 27076 9466 27092
rect 9482 27076 9498 27092
rect 9514 27076 9530 27092
rect 9546 27076 9562 27092
rect 9578 27076 9594 27092
rect 9610 27076 9626 27092
rect 9642 27076 9658 27092
rect 9674 27076 9690 27092
rect 9706 27076 9722 27092
rect 9738 27076 9754 27092
rect 9770 27076 9786 27092
rect 9802 27076 9819 27092
rect 8820 27060 9819 27076
rect 8820 27044 9338 27060
rect 9354 27044 9370 27060
rect 9386 27044 9402 27060
rect 9418 27044 9434 27060
rect 9450 27044 9466 27060
rect 9482 27044 9498 27060
rect 9514 27044 9530 27060
rect 9546 27044 9562 27060
rect 9578 27044 9594 27060
rect 9610 27044 9626 27060
rect 9642 27044 9658 27060
rect 9674 27044 9690 27060
rect 9706 27044 9722 27060
rect 9738 27044 9754 27060
rect 9770 27044 9786 27060
rect 9802 27044 9819 27060
rect 8820 27028 9819 27044
rect 8820 27012 9338 27028
rect 9354 27012 9370 27028
rect 9386 27012 9402 27028
rect 9418 27012 9434 27028
rect 9450 27012 9466 27028
rect 9482 27012 9498 27028
rect 9514 27012 9530 27028
rect 9546 27012 9562 27028
rect 9578 27012 9594 27028
rect 9610 27012 9626 27028
rect 9642 27012 9658 27028
rect 9674 27012 9690 27028
rect 9706 27012 9722 27028
rect 9738 27012 9754 27028
rect 9770 27012 9786 27028
rect 9802 27012 9819 27028
rect 8820 26996 9819 27012
rect 8820 26980 9338 26996
rect 9354 26980 9370 26996
rect 9386 26980 9402 26996
rect 9418 26980 9434 26996
rect 9450 26980 9466 26996
rect 9482 26980 9498 26996
rect 9514 26980 9530 26996
rect 9546 26980 9562 26996
rect 9578 26980 9594 26996
rect 9610 26980 9626 26996
rect 9642 26980 9658 26996
rect 9674 26980 9690 26996
rect 9706 26980 9722 26996
rect 9738 26980 9754 26996
rect 9770 26980 9786 26996
rect 9802 26980 9819 26996
rect 8820 26964 9819 26980
rect 8820 26948 9338 26964
rect 9354 26948 9370 26964
rect 9386 26948 9402 26964
rect 9418 26948 9434 26964
rect 9450 26948 9466 26964
rect 9482 26948 9498 26964
rect 9514 26948 9530 26964
rect 9546 26948 9562 26964
rect 9578 26948 9594 26964
rect 9610 26948 9626 26964
rect 9642 26948 9658 26964
rect 9674 26948 9690 26964
rect 9706 26948 9722 26964
rect 9738 26948 9754 26964
rect 9770 26948 9786 26964
rect 9802 26948 9819 26964
rect 8820 26932 9819 26948
rect 8820 26916 9338 26932
rect 9354 26916 9370 26932
rect 9386 26916 9402 26932
rect 9418 26916 9434 26932
rect 9450 26916 9466 26932
rect 9482 26916 9498 26932
rect 9514 26916 9530 26932
rect 9546 26916 9562 26932
rect 9578 26916 9594 26932
rect 9610 26916 9626 26932
rect 9642 26916 9658 26932
rect 9674 26916 9690 26932
rect 9706 26916 9722 26932
rect 9738 26916 9754 26932
rect 9770 26916 9786 26932
rect 9802 26916 9819 26932
rect 8820 26900 9819 26916
rect 8820 26884 9338 26900
rect 9354 26884 9370 26900
rect 9386 26884 9402 26900
rect 9418 26884 9434 26900
rect 9450 26884 9466 26900
rect 9482 26884 9498 26900
rect 9514 26884 9530 26900
rect 9546 26884 9562 26900
rect 9578 26884 9594 26900
rect 9610 26884 9626 26900
rect 9642 26884 9658 26900
rect 9674 26884 9690 26900
rect 9706 26884 9722 26900
rect 9738 26884 9754 26900
rect 9770 26884 9786 26900
rect 9802 26884 9819 26900
rect 8820 26868 9819 26884
rect 8820 26852 9338 26868
rect 9354 26852 9370 26868
rect 9386 26852 9402 26868
rect 9418 26852 9434 26868
rect 9450 26852 9466 26868
rect 9482 26852 9498 26868
rect 9514 26852 9530 26868
rect 9546 26852 9562 26868
rect 9578 26852 9594 26868
rect 9610 26852 9626 26868
rect 9642 26852 9658 26868
rect 9674 26852 9690 26868
rect 9706 26852 9722 26868
rect 9738 26852 9754 26868
rect 9770 26852 9786 26868
rect 9802 26852 9819 26868
rect 8820 26836 9819 26852
rect 8820 26820 9338 26836
rect 9354 26820 9370 26836
rect 9386 26820 9402 26836
rect 9418 26820 9434 26836
rect 9450 26820 9466 26836
rect 9482 26820 9498 26836
rect 9514 26820 9530 26836
rect 9546 26820 9562 26836
rect 9578 26820 9594 26836
rect 9610 26820 9626 26836
rect 9642 26820 9658 26836
rect 9674 26820 9690 26836
rect 9706 26820 9722 26836
rect 9738 26820 9754 26836
rect 9770 26820 9786 26836
rect 9802 26820 9819 26836
rect 8820 26804 9819 26820
rect 8820 26788 9338 26804
rect 9354 26788 9370 26804
rect 9386 26788 9402 26804
rect 9418 26788 9434 26804
rect 9450 26788 9466 26804
rect 9482 26788 9498 26804
rect 9514 26788 9530 26804
rect 9546 26788 9562 26804
rect 9578 26788 9594 26804
rect 9610 26788 9626 26804
rect 9642 26788 9658 26804
rect 9674 26788 9690 26804
rect 9706 26788 9722 26804
rect 9738 26788 9754 26804
rect 9770 26788 9786 26804
rect 9802 26788 9819 26804
rect 8820 26772 9819 26788
rect 8820 26756 9338 26772
rect 9354 26756 9370 26772
rect 9386 26756 9402 26772
rect 9418 26756 9434 26772
rect 9450 26756 9466 26772
rect 9482 26756 9498 26772
rect 9514 26756 9530 26772
rect 9546 26756 9562 26772
rect 9578 26756 9594 26772
rect 9610 26756 9626 26772
rect 9642 26756 9658 26772
rect 9674 26756 9690 26772
rect 9706 26756 9722 26772
rect 9738 26756 9754 26772
rect 9770 26756 9786 26772
rect 9802 26756 9819 26772
rect 12480 26860 12580 29180
rect 15180 27060 15280 29180
rect 17880 27260 17980 29180
rect 20580 27460 20680 29180
rect 23280 27660 23380 29180
rect 25980 27860 26080 29180
rect 25980 27760 26500 27860
rect 23280 27560 25760 27660
rect 20580 27360 25560 27460
rect 17880 27160 24860 27260
rect 15180 26960 24660 27060
rect 12480 26760 21920 26860
rect 8820 26740 9819 26756
rect 24560 26740 24660 26960
rect 24760 26740 24860 27160
rect 25460 26740 25560 27360
rect 25660 26740 25760 27560
rect 26400 26740 26500 27760
rect 8820 26724 9338 26740
rect 9354 26724 9370 26740
rect 9386 26724 9402 26740
rect 9418 26724 9434 26740
rect 9450 26724 9466 26740
rect 9482 26724 9498 26740
rect 9514 26724 9530 26740
rect 9546 26724 9562 26740
rect 9578 26724 9594 26740
rect 9610 26724 9626 26740
rect 9642 26724 9658 26740
rect 9674 26724 9690 26740
rect 9706 26724 9722 26740
rect 9738 26724 9754 26740
rect 9770 26724 9786 26740
rect 9802 26724 9819 26740
rect 8820 26708 9819 26724
rect 8820 26692 9338 26708
rect 9354 26692 9370 26708
rect 9386 26692 9402 26708
rect 9418 26692 9434 26708
rect 9450 26692 9466 26708
rect 9482 26692 9498 26708
rect 9514 26692 9530 26708
rect 9546 26692 9562 26708
rect 9578 26692 9594 26708
rect 9610 26692 9626 26708
rect 9642 26692 9658 26708
rect 9674 26692 9690 26708
rect 9706 26692 9722 26708
rect 9738 26692 9754 26708
rect 9770 26692 9786 26708
rect 9802 26692 9819 26708
rect 8820 26676 9819 26692
rect 8820 26660 9338 26676
rect 9354 26660 9370 26676
rect 9386 26660 9402 26676
rect 9418 26660 9434 26676
rect 9450 26660 9466 26676
rect 9482 26660 9498 26676
rect 9514 26660 9530 26676
rect 9546 26660 9562 26676
rect 9578 26660 9594 26676
rect 9610 26660 9626 26676
rect 9642 26660 9658 26676
rect 9674 26660 9690 26676
rect 9706 26660 9722 26676
rect 9738 26660 9754 26676
rect 9770 26660 9786 26676
rect 9802 26660 9819 26676
rect 8820 26644 9819 26660
rect 8820 26628 9338 26644
rect 9354 26628 9370 26644
rect 9386 26628 9402 26644
rect 9418 26628 9434 26644
rect 9450 26628 9466 26644
rect 9482 26628 9498 26644
rect 9514 26628 9530 26644
rect 9546 26628 9562 26644
rect 9578 26628 9594 26644
rect 9610 26628 9626 26644
rect 9642 26628 9658 26644
rect 9674 26628 9690 26644
rect 9706 26628 9722 26644
rect 9738 26628 9754 26644
rect 9770 26628 9786 26644
rect 9802 26628 9819 26644
rect 8820 26612 9819 26628
rect 8820 26596 9338 26612
rect 9354 26596 9370 26612
rect 9386 26596 9402 26612
rect 9418 26596 9434 26612
rect 9450 26596 9466 26612
rect 9482 26596 9498 26612
rect 9514 26596 9530 26612
rect 9546 26596 9562 26612
rect 9578 26596 9594 26612
rect 9610 26596 9626 26612
rect 9642 26596 9658 26612
rect 9674 26596 9690 26612
rect 9706 26596 9722 26612
rect 9738 26596 9754 26612
rect 9770 26596 9786 26612
rect 9802 26596 9819 26612
rect 8820 26580 9819 26596
rect 8820 26564 9338 26580
rect 9354 26564 9370 26580
rect 9386 26564 9402 26580
rect 9418 26564 9434 26580
rect 9450 26564 9466 26580
rect 9482 26564 9498 26580
rect 9514 26564 9530 26580
rect 9546 26564 9562 26580
rect 9578 26564 9594 26580
rect 9610 26564 9626 26580
rect 9642 26564 9658 26580
rect 9674 26564 9690 26580
rect 9706 26564 9722 26580
rect 9738 26564 9754 26580
rect 9770 26564 9786 26580
rect 9802 26564 9819 26580
rect 8820 26548 9819 26564
rect 8820 26532 9338 26548
rect 9354 26532 9370 26548
rect 9386 26532 9402 26548
rect 9418 26532 9434 26548
rect 9450 26532 9466 26548
rect 9482 26532 9498 26548
rect 9514 26532 9530 26548
rect 9546 26532 9562 26548
rect 9578 26532 9594 26548
rect 9610 26532 9626 26548
rect 9642 26532 9658 26548
rect 9674 26532 9690 26548
rect 9706 26532 9722 26548
rect 9738 26532 9754 26548
rect 9770 26532 9786 26548
rect 9802 26532 9819 26548
rect 8820 26516 9819 26532
rect 8820 26500 9338 26516
rect 9354 26500 9370 26516
rect 9386 26500 9402 26516
rect 9418 26500 9434 26516
rect 9450 26500 9466 26516
rect 9482 26500 9498 26516
rect 9514 26500 9530 26516
rect 9546 26500 9562 26516
rect 9578 26500 9594 26516
rect 9610 26500 9626 26516
rect 9642 26500 9658 26516
rect 9674 26500 9690 26516
rect 9706 26500 9722 26516
rect 9738 26500 9754 26516
rect 9770 26500 9786 26516
rect 9802 26500 9819 26516
rect 8820 26484 9819 26500
rect 8820 26468 9338 26484
rect 9354 26468 9370 26484
rect 9386 26468 9402 26484
rect 9418 26468 9434 26484
rect 9450 26468 9466 26484
rect 9482 26468 9498 26484
rect 9514 26468 9530 26484
rect 9546 26468 9562 26484
rect 9578 26468 9594 26484
rect 9610 26468 9626 26484
rect 9642 26468 9658 26484
rect 9674 26468 9690 26484
rect 9706 26468 9722 26484
rect 9738 26468 9754 26484
rect 9770 26468 9786 26484
rect 9802 26468 9819 26484
rect 8820 26452 9819 26468
rect 8820 26436 9338 26452
rect 9354 26436 9370 26452
rect 9386 26436 9402 26452
rect 9418 26436 9434 26452
rect 9450 26436 9466 26452
rect 9482 26436 9498 26452
rect 9514 26436 9530 26452
rect 9546 26436 9562 26452
rect 9578 26436 9594 26452
rect 9610 26436 9626 26452
rect 9642 26436 9658 26452
rect 9674 26436 9690 26452
rect 9706 26436 9722 26452
rect 9738 26436 9754 26452
rect 9770 26436 9786 26452
rect 9802 26436 9819 26452
rect 8820 26421 9819 26436
rect 8820 26420 9320 26421
rect 29080 26079 29180 26080
rect 28781 26054 29180 26079
rect 28781 26038 28794 26054
rect 28810 26038 28826 26054
rect 28842 26038 28858 26054
rect 28874 26038 28890 26054
rect 28906 26038 28922 26054
rect 28938 26038 28954 26054
rect 28970 26038 28986 26054
rect 29002 26038 29018 26054
rect 29034 26038 29050 26054
rect 29066 26038 29180 26054
rect 28781 26022 29180 26038
rect 28781 26006 28794 26022
rect 28810 26006 28826 26022
rect 28842 26006 28858 26022
rect 28874 26006 28890 26022
rect 28906 26006 28922 26022
rect 28938 26006 28954 26022
rect 28970 26006 28986 26022
rect 29002 26006 29018 26022
rect 29034 26006 29050 26022
rect 29066 26006 29180 26022
rect 28781 25981 29180 26006
rect 29080 25980 29180 25981
rect 29080 23379 29180 23380
rect 8820 23359 10620 23360
rect 8820 23334 10919 23359
rect 8820 23318 10634 23334
rect 10650 23318 10666 23334
rect 10682 23318 10698 23334
rect 10714 23318 10730 23334
rect 10746 23318 10762 23334
rect 10778 23318 10794 23334
rect 10810 23318 10826 23334
rect 10842 23318 10858 23334
rect 10874 23318 10890 23334
rect 10906 23318 10919 23334
rect 8820 23302 10919 23318
rect 8820 23286 10634 23302
rect 10650 23286 10666 23302
rect 10682 23286 10698 23302
rect 10714 23286 10730 23302
rect 10746 23286 10762 23302
rect 10778 23286 10794 23302
rect 10810 23286 10826 23302
rect 10842 23286 10858 23302
rect 10874 23286 10890 23302
rect 10906 23286 10919 23302
rect 8820 23261 10919 23286
rect 28781 23354 29180 23379
rect 28781 23338 28794 23354
rect 28810 23338 28826 23354
rect 28842 23338 28858 23354
rect 28874 23338 28890 23354
rect 28906 23338 28922 23354
rect 28938 23338 28954 23354
rect 28970 23338 28986 23354
rect 29002 23338 29018 23354
rect 29034 23338 29050 23354
rect 29066 23338 29180 23354
rect 28781 23322 29180 23338
rect 28781 23306 28794 23322
rect 28810 23306 28826 23322
rect 28842 23306 28858 23322
rect 28874 23306 28890 23322
rect 28906 23306 28922 23322
rect 28938 23306 28954 23322
rect 28970 23306 28986 23322
rect 29002 23306 29018 23322
rect 29034 23306 29050 23322
rect 29066 23306 29180 23322
rect 28781 23281 29180 23306
rect 29080 23280 29180 23281
rect 8820 23260 10620 23261
rect 29080 20679 29180 20680
rect 8820 20659 8920 20660
rect 8820 20634 9219 20659
rect 8820 20618 8934 20634
rect 8950 20618 8966 20634
rect 8982 20618 8998 20634
rect 9014 20618 9030 20634
rect 9046 20618 9062 20634
rect 9078 20618 9094 20634
rect 9110 20618 9126 20634
rect 9142 20618 9158 20634
rect 9174 20618 9190 20634
rect 9206 20618 9219 20634
rect 8820 20602 9219 20618
rect 8820 20586 8934 20602
rect 8950 20586 8966 20602
rect 8982 20586 8998 20602
rect 9014 20586 9030 20602
rect 9046 20586 9062 20602
rect 9078 20586 9094 20602
rect 9110 20586 9126 20602
rect 9142 20586 9158 20602
rect 9174 20586 9190 20602
rect 9206 20586 9219 20602
rect 8820 20561 9219 20586
rect 28781 20654 29180 20679
rect 28781 20638 28794 20654
rect 28810 20638 28826 20654
rect 28842 20638 28858 20654
rect 28874 20638 28890 20654
rect 28906 20638 28922 20654
rect 28938 20638 28954 20654
rect 28970 20638 28986 20654
rect 29002 20638 29018 20654
rect 29034 20638 29050 20654
rect 29066 20638 29180 20654
rect 28781 20622 29180 20638
rect 28781 20606 28794 20622
rect 28810 20606 28826 20622
rect 28842 20606 28858 20622
rect 28874 20606 28890 20622
rect 28906 20606 28922 20622
rect 28938 20606 28954 20622
rect 28970 20606 28986 20622
rect 29002 20606 29018 20622
rect 29034 20606 29050 20622
rect 29066 20606 29180 20622
rect 28781 20581 29180 20606
rect 29080 20580 29180 20581
rect 8820 20560 8920 20561
rect 29080 17979 29180 17980
rect 28781 17954 29180 17979
rect 28781 17938 28794 17954
rect 28810 17938 28826 17954
rect 28842 17938 28858 17954
rect 28874 17938 28890 17954
rect 28906 17938 28922 17954
rect 28938 17938 28954 17954
rect 28970 17938 28986 17954
rect 29002 17938 29018 17954
rect 29034 17938 29050 17954
rect 29066 17938 29180 17954
rect 28781 17922 29180 17938
rect 28781 17906 28794 17922
rect 28810 17906 28826 17922
rect 28842 17906 28858 17922
rect 28874 17906 28890 17922
rect 28906 17906 28922 17922
rect 28938 17906 28954 17922
rect 28970 17906 28986 17922
rect 29002 17906 29018 17922
rect 29034 17906 29050 17922
rect 29066 17906 29180 17922
rect 28781 17881 29180 17906
rect 29080 17880 29180 17881
rect 29080 15279 29180 15280
rect 28781 15254 29180 15279
rect 28781 15238 28794 15254
rect 28810 15238 28826 15254
rect 28842 15238 28858 15254
rect 28874 15238 28890 15254
rect 28906 15238 28922 15254
rect 28938 15238 28954 15254
rect 28970 15238 28986 15254
rect 29002 15238 29018 15254
rect 29034 15238 29050 15254
rect 29066 15238 29180 15254
rect 28781 15222 29180 15238
rect 28781 15206 28794 15222
rect 28810 15206 28826 15222
rect 28842 15206 28858 15222
rect 28874 15206 28890 15222
rect 28906 15206 28922 15222
rect 28938 15206 28954 15222
rect 28970 15206 28986 15222
rect 29002 15206 29018 15222
rect 29034 15206 29050 15222
rect 29066 15206 29180 15222
rect 28781 15181 29180 15206
rect 29080 15180 29180 15181
rect 29080 12579 29180 12580
rect 28781 12554 29180 12579
rect 28781 12538 28794 12554
rect 28810 12538 28826 12554
rect 28842 12538 28858 12554
rect 28874 12538 28890 12554
rect 28906 12538 28922 12554
rect 28938 12538 28954 12554
rect 28970 12538 28986 12554
rect 29002 12538 29018 12554
rect 29034 12538 29050 12554
rect 29066 12538 29180 12554
rect 28781 12522 29180 12538
rect 28781 12506 28794 12522
rect 28810 12506 28826 12522
rect 28842 12506 28858 12522
rect 28874 12506 28890 12522
rect 28906 12506 28922 12522
rect 28938 12506 28954 12522
rect 28970 12506 28986 12522
rect 29002 12506 29018 12522
rect 29034 12506 29050 12522
rect 29066 12506 29180 12522
rect 28781 12481 29180 12506
rect 29080 12480 29180 12481
rect 20420 10080 20520 11440
rect 11940 9980 20520 10080
rect 8820 9899 9000 9900
rect 8820 9882 9719 9899
rect 8820 9866 9016 9882
rect 9032 9866 9048 9882
rect 9064 9866 9080 9882
rect 9096 9866 9112 9882
rect 9128 9866 9144 9882
rect 9160 9866 9176 9882
rect 9192 9866 9208 9882
rect 9224 9866 9240 9882
rect 9256 9866 9272 9882
rect 9288 9866 9304 9882
rect 9320 9866 9336 9882
rect 9352 9866 9368 9882
rect 9384 9866 9400 9882
rect 9416 9866 9432 9882
rect 9448 9866 9464 9882
rect 9480 9866 9496 9882
rect 9512 9866 9528 9882
rect 9544 9866 9560 9882
rect 9576 9866 9592 9882
rect 9608 9866 9624 9882
rect 9640 9866 9656 9882
rect 9672 9866 9688 9882
rect 9704 9866 9719 9882
rect 8820 9850 9719 9866
rect 8820 9834 9016 9850
rect 9032 9834 9048 9850
rect 9064 9834 9080 9850
rect 9096 9834 9112 9850
rect 9128 9834 9144 9850
rect 9160 9834 9176 9850
rect 9192 9834 9208 9850
rect 9224 9834 9240 9850
rect 9256 9834 9272 9850
rect 9288 9834 9304 9850
rect 9320 9834 9336 9850
rect 9352 9834 9368 9850
rect 9384 9834 9400 9850
rect 9416 9834 9432 9850
rect 9448 9834 9464 9850
rect 9480 9834 9496 9850
rect 9512 9834 9528 9850
rect 9544 9834 9560 9850
rect 9576 9834 9592 9850
rect 9608 9834 9624 9850
rect 9640 9834 9656 9850
rect 9672 9834 9688 9850
rect 9704 9834 9719 9850
rect 8820 9818 9719 9834
rect 8820 9802 9016 9818
rect 9032 9802 9048 9818
rect 9064 9802 9080 9818
rect 9096 9802 9112 9818
rect 9128 9802 9144 9818
rect 9160 9802 9176 9818
rect 9192 9802 9208 9818
rect 9224 9802 9240 9818
rect 9256 9802 9272 9818
rect 9288 9802 9304 9818
rect 9320 9802 9336 9818
rect 9352 9802 9368 9818
rect 9384 9802 9400 9818
rect 9416 9802 9432 9818
rect 9448 9802 9464 9818
rect 9480 9802 9496 9818
rect 9512 9802 9528 9818
rect 9544 9802 9560 9818
rect 9576 9802 9592 9818
rect 9608 9802 9624 9818
rect 9640 9802 9656 9818
rect 9672 9802 9688 9818
rect 9704 9802 9719 9818
rect 8820 9786 9719 9802
rect 8820 9770 9016 9786
rect 9032 9770 9048 9786
rect 9064 9770 9080 9786
rect 9096 9770 9112 9786
rect 9128 9770 9144 9786
rect 9160 9770 9176 9786
rect 9192 9770 9208 9786
rect 9224 9770 9240 9786
rect 9256 9770 9272 9786
rect 9288 9770 9304 9786
rect 9320 9770 9336 9786
rect 9352 9770 9368 9786
rect 9384 9770 9400 9786
rect 9416 9770 9432 9786
rect 9448 9770 9464 9786
rect 9480 9770 9496 9786
rect 9512 9770 9528 9786
rect 9544 9770 9560 9786
rect 9576 9770 9592 9786
rect 9608 9770 9624 9786
rect 9640 9770 9656 9786
rect 9672 9770 9688 9786
rect 9704 9770 9719 9786
rect 8820 9754 9719 9770
rect 8820 9738 9016 9754
rect 9032 9738 9048 9754
rect 9064 9738 9080 9754
rect 9096 9738 9112 9754
rect 9128 9738 9144 9754
rect 9160 9738 9176 9754
rect 9192 9738 9208 9754
rect 9224 9738 9240 9754
rect 9256 9738 9272 9754
rect 9288 9738 9304 9754
rect 9320 9738 9336 9754
rect 9352 9738 9368 9754
rect 9384 9738 9400 9754
rect 9416 9738 9432 9754
rect 9448 9738 9464 9754
rect 9480 9738 9496 9754
rect 9512 9738 9528 9754
rect 9544 9738 9560 9754
rect 9576 9738 9592 9754
rect 9608 9738 9624 9754
rect 9640 9738 9656 9754
rect 9672 9738 9688 9754
rect 9704 9738 9719 9754
rect 8820 9721 9719 9738
rect 8820 9720 9000 9721
rect 11940 8820 12040 9980
rect 20600 9880 20700 11440
rect 14640 9780 20700 9880
rect 14640 8820 14740 9780
rect 21980 9680 22080 11440
rect 17340 9580 22080 9680
rect 17340 8820 17440 9580
rect 22160 9480 22260 11440
rect 20040 9380 22260 9480
rect 20040 8820 20140 9380
rect 25260 9280 25360 11420
rect 22740 9180 25360 9280
rect 22740 8820 22840 9180
rect 26200 9080 26300 11420
rect 29080 9879 29180 9880
rect 28781 9854 29180 9879
rect 28781 9838 28794 9854
rect 28810 9838 28826 9854
rect 28842 9838 28858 9854
rect 28874 9838 28890 9854
rect 28906 9838 28922 9854
rect 28938 9838 28954 9854
rect 28970 9838 28986 9854
rect 29002 9838 29018 9854
rect 29034 9838 29050 9854
rect 29066 9838 29180 9854
rect 28781 9822 29180 9838
rect 28781 9806 28794 9822
rect 28810 9806 28826 9822
rect 28842 9806 28858 9822
rect 28874 9806 28890 9822
rect 28906 9806 28922 9822
rect 28938 9806 28954 9822
rect 28970 9806 28986 9822
rect 29002 9806 29018 9822
rect 29034 9806 29050 9822
rect 29066 9806 29180 9822
rect 28781 9781 29180 9806
rect 29080 9780 29180 9781
rect 25440 8980 26300 9080
rect 25440 8820 25540 8980
<< m3contact >>
rect 28794 26038 28810 26054
rect 28826 26038 28842 26054
rect 28858 26038 28874 26054
rect 28890 26038 28906 26054
rect 28922 26038 28938 26054
rect 28954 26038 28970 26054
rect 28986 26038 29002 26054
rect 29018 26038 29034 26054
rect 29050 26038 29066 26054
rect 28794 26006 28810 26022
rect 28826 26006 28842 26022
rect 28858 26006 28874 26022
rect 28890 26006 28906 26022
rect 28922 26006 28938 26022
rect 28954 26006 28970 26022
rect 28986 26006 29002 26022
rect 29018 26006 29034 26022
rect 29050 26006 29066 26022
rect 10634 23318 10650 23334
rect 10666 23318 10682 23334
rect 10698 23318 10714 23334
rect 10730 23318 10746 23334
rect 10762 23318 10778 23334
rect 10794 23318 10810 23334
rect 10826 23318 10842 23334
rect 10858 23318 10874 23334
rect 10890 23318 10906 23334
rect 10634 23286 10650 23302
rect 10666 23286 10682 23302
rect 10698 23286 10714 23302
rect 10730 23286 10746 23302
rect 10762 23286 10778 23302
rect 10794 23286 10810 23302
rect 10826 23286 10842 23302
rect 10858 23286 10874 23302
rect 10890 23286 10906 23302
rect 28794 23338 28810 23354
rect 28826 23338 28842 23354
rect 28858 23338 28874 23354
rect 28890 23338 28906 23354
rect 28922 23338 28938 23354
rect 28954 23338 28970 23354
rect 28986 23338 29002 23354
rect 29018 23338 29034 23354
rect 29050 23338 29066 23354
rect 28794 23306 28810 23322
rect 28826 23306 28842 23322
rect 28858 23306 28874 23322
rect 28890 23306 28906 23322
rect 28922 23306 28938 23322
rect 28954 23306 28970 23322
rect 28986 23306 29002 23322
rect 29018 23306 29034 23322
rect 29050 23306 29066 23322
rect 8934 20618 8950 20634
rect 8966 20618 8982 20634
rect 8998 20618 9014 20634
rect 9030 20618 9046 20634
rect 9062 20618 9078 20634
rect 9094 20618 9110 20634
rect 9126 20618 9142 20634
rect 9158 20618 9174 20634
rect 9190 20618 9206 20634
rect 8934 20586 8950 20602
rect 8966 20586 8982 20602
rect 8998 20586 9014 20602
rect 9030 20586 9046 20602
rect 9062 20586 9078 20602
rect 9094 20586 9110 20602
rect 9126 20586 9142 20602
rect 9158 20586 9174 20602
rect 9190 20586 9206 20602
rect 28794 20638 28810 20654
rect 28826 20638 28842 20654
rect 28858 20638 28874 20654
rect 28890 20638 28906 20654
rect 28922 20638 28938 20654
rect 28954 20638 28970 20654
rect 28986 20638 29002 20654
rect 29018 20638 29034 20654
rect 29050 20638 29066 20654
rect 28794 20606 28810 20622
rect 28826 20606 28842 20622
rect 28858 20606 28874 20622
rect 28890 20606 28906 20622
rect 28922 20606 28938 20622
rect 28954 20606 28970 20622
rect 28986 20606 29002 20622
rect 29018 20606 29034 20622
rect 29050 20606 29066 20622
rect 28794 17938 28810 17954
rect 28826 17938 28842 17954
rect 28858 17938 28874 17954
rect 28890 17938 28906 17954
rect 28922 17938 28938 17954
rect 28954 17938 28970 17954
rect 28986 17938 29002 17954
rect 29018 17938 29034 17954
rect 29050 17938 29066 17954
rect 28794 17906 28810 17922
rect 28826 17906 28842 17922
rect 28858 17906 28874 17922
rect 28890 17906 28906 17922
rect 28922 17906 28938 17922
rect 28954 17906 28970 17922
rect 28986 17906 29002 17922
rect 29018 17906 29034 17922
rect 29050 17906 29066 17922
rect 28794 15238 28810 15254
rect 28826 15238 28842 15254
rect 28858 15238 28874 15254
rect 28890 15238 28906 15254
rect 28922 15238 28938 15254
rect 28954 15238 28970 15254
rect 28986 15238 29002 15254
rect 29018 15238 29034 15254
rect 29050 15238 29066 15254
rect 28794 15206 28810 15222
rect 28826 15206 28842 15222
rect 28858 15206 28874 15222
rect 28890 15206 28906 15222
rect 28922 15206 28938 15222
rect 28954 15206 28970 15222
rect 28986 15206 29002 15222
rect 29018 15206 29034 15222
rect 29050 15206 29066 15222
rect 28794 12538 28810 12554
rect 28826 12538 28842 12554
rect 28858 12538 28874 12554
rect 28890 12538 28906 12554
rect 28922 12538 28938 12554
rect 28954 12538 28970 12554
rect 28986 12538 29002 12554
rect 29018 12538 29034 12554
rect 29050 12538 29066 12554
rect 28794 12506 28810 12522
rect 28826 12506 28842 12522
rect 28858 12506 28874 12522
rect 28890 12506 28906 12522
rect 28922 12506 28938 12522
rect 28954 12506 28970 12522
rect 28986 12506 29002 12522
rect 29018 12506 29034 12522
rect 29050 12506 29066 12522
rect 9016 9866 9032 9882
rect 9048 9866 9064 9882
rect 9080 9866 9096 9882
rect 9112 9866 9128 9882
rect 9144 9866 9160 9882
rect 9176 9866 9192 9882
rect 9208 9866 9224 9882
rect 9240 9866 9256 9882
rect 9272 9866 9288 9882
rect 9304 9866 9320 9882
rect 9336 9866 9352 9882
rect 9368 9866 9384 9882
rect 9400 9866 9416 9882
rect 9432 9866 9448 9882
rect 9464 9866 9480 9882
rect 9496 9866 9512 9882
rect 9528 9866 9544 9882
rect 9560 9866 9576 9882
rect 9592 9866 9608 9882
rect 9624 9866 9640 9882
rect 9656 9866 9672 9882
rect 9688 9866 9704 9882
rect 9016 9834 9032 9850
rect 9048 9834 9064 9850
rect 9080 9834 9096 9850
rect 9112 9834 9128 9850
rect 9144 9834 9160 9850
rect 9176 9834 9192 9850
rect 9208 9834 9224 9850
rect 9240 9834 9256 9850
rect 9272 9834 9288 9850
rect 9304 9834 9320 9850
rect 9336 9834 9352 9850
rect 9368 9834 9384 9850
rect 9400 9834 9416 9850
rect 9432 9834 9448 9850
rect 9464 9834 9480 9850
rect 9496 9834 9512 9850
rect 9528 9834 9544 9850
rect 9560 9834 9576 9850
rect 9592 9834 9608 9850
rect 9624 9834 9640 9850
rect 9656 9834 9672 9850
rect 9688 9834 9704 9850
rect 9016 9802 9032 9818
rect 9048 9802 9064 9818
rect 9080 9802 9096 9818
rect 9112 9802 9128 9818
rect 9144 9802 9160 9818
rect 9176 9802 9192 9818
rect 9208 9802 9224 9818
rect 9240 9802 9256 9818
rect 9272 9802 9288 9818
rect 9304 9802 9320 9818
rect 9336 9802 9352 9818
rect 9368 9802 9384 9818
rect 9400 9802 9416 9818
rect 9432 9802 9448 9818
rect 9464 9802 9480 9818
rect 9496 9802 9512 9818
rect 9528 9802 9544 9818
rect 9560 9802 9576 9818
rect 9592 9802 9608 9818
rect 9624 9802 9640 9818
rect 9656 9802 9672 9818
rect 9688 9802 9704 9818
rect 9016 9770 9032 9786
rect 9048 9770 9064 9786
rect 9080 9770 9096 9786
rect 9112 9770 9128 9786
rect 9144 9770 9160 9786
rect 9176 9770 9192 9786
rect 9208 9770 9224 9786
rect 9240 9770 9256 9786
rect 9272 9770 9288 9786
rect 9304 9770 9320 9786
rect 9336 9770 9352 9786
rect 9368 9770 9384 9786
rect 9400 9770 9416 9786
rect 9432 9770 9448 9786
rect 9464 9770 9480 9786
rect 9496 9770 9512 9786
rect 9528 9770 9544 9786
rect 9560 9770 9576 9786
rect 9592 9770 9608 9786
rect 9624 9770 9640 9786
rect 9656 9770 9672 9786
rect 9688 9770 9704 9786
rect 9016 9738 9032 9754
rect 9048 9738 9064 9754
rect 9080 9738 9096 9754
rect 9112 9738 9128 9754
rect 9144 9738 9160 9754
rect 9176 9738 9192 9754
rect 9208 9738 9224 9754
rect 9240 9738 9256 9754
rect 9272 9738 9288 9754
rect 9304 9738 9320 9754
rect 9336 9738 9352 9754
rect 9368 9738 9384 9754
rect 9400 9738 9416 9754
rect 9432 9738 9448 9754
rect 9464 9738 9480 9754
rect 9496 9738 9512 9754
rect 9528 9738 9544 9754
rect 9560 9738 9576 9754
rect 9592 9738 9608 9754
rect 9624 9738 9640 9754
rect 9656 9738 9672 9754
rect 9688 9738 9704 9754
rect 28794 9838 28810 9854
rect 28826 9838 28842 9854
rect 28858 9838 28874 9854
rect 28890 9838 28906 9854
rect 28922 9838 28938 9854
rect 28954 9838 28970 9854
rect 28986 9838 29002 9854
rect 29018 9838 29034 9854
rect 29050 9838 29066 9854
rect 28794 9806 28810 9822
rect 28826 9806 28842 9822
rect 28858 9806 28874 9822
rect 28890 9806 28906 9822
rect 28922 9806 28938 9822
rect 28954 9806 28970 9822
rect 28986 9806 29002 9822
rect 29018 9806 29034 9822
rect 29050 9806 29066 9822
<< metal3 >>
rect 9120 26180 11320 26280
rect 9120 20660 9220 26180
rect 28781 26054 29079 26079
rect 28781 26038 28794 26054
rect 28810 26038 28826 26054
rect 28842 26038 28858 26054
rect 28874 26038 28890 26054
rect 28906 26038 28922 26054
rect 28938 26038 28954 26054
rect 28970 26038 28986 26054
rect 29002 26038 29018 26054
rect 29034 26038 29050 26054
rect 29066 26038 29079 26054
rect 28781 26022 29079 26038
rect 28781 26006 28794 26022
rect 28810 26006 28826 26022
rect 28842 26006 28858 26022
rect 28874 26006 28890 26022
rect 28906 26006 28922 26022
rect 28938 26006 28954 26022
rect 28970 26006 28986 26022
rect 29002 26006 29018 26022
rect 29034 26006 29050 26022
rect 29066 26006 29079 26022
rect 28781 25980 29079 26006
rect 28780 24100 28880 25980
rect 26720 24000 28880 24100
rect 26720 23380 28020 23400
rect 26720 23379 28780 23380
rect 10621 23334 10919 23359
rect 10621 23318 10634 23334
rect 10650 23318 10666 23334
rect 10682 23318 10698 23334
rect 10714 23318 10730 23334
rect 10746 23318 10762 23334
rect 10778 23318 10794 23334
rect 10810 23318 10826 23334
rect 10842 23318 10858 23334
rect 10874 23318 10890 23334
rect 10906 23318 10919 23334
rect 10621 23302 10919 23318
rect 10621 23286 10634 23302
rect 10650 23286 10666 23302
rect 10682 23286 10698 23302
rect 10714 23286 10730 23302
rect 10746 23286 10762 23302
rect 10778 23286 10794 23302
rect 10810 23286 10826 23302
rect 10842 23286 10858 23302
rect 10874 23286 10890 23302
rect 10906 23286 10919 23302
rect 26720 23354 29079 23379
rect 26720 23338 28794 23354
rect 28810 23338 28826 23354
rect 28842 23338 28858 23354
rect 28874 23338 28890 23354
rect 28906 23338 28922 23354
rect 28938 23338 28954 23354
rect 28970 23338 28986 23354
rect 29002 23338 29018 23354
rect 29034 23338 29050 23354
rect 29066 23338 29079 23354
rect 26720 23322 29079 23338
rect 26720 23306 28794 23322
rect 28810 23306 28826 23322
rect 28842 23306 28858 23322
rect 28874 23306 28890 23322
rect 28906 23306 28922 23322
rect 28938 23306 28954 23322
rect 28970 23306 28986 23322
rect 29002 23306 29018 23322
rect 29034 23306 29050 23322
rect 29066 23306 29079 23322
rect 26720 23300 29079 23306
rect 10621 23260 10919 23286
rect 27920 23281 29079 23300
rect 27920 23280 28780 23281
rect 10820 20800 10920 23260
rect 26720 22560 27820 22660
rect 26720 21860 27620 21960
rect 26680 21380 27420 21460
rect 26680 21220 27220 21300
rect 26680 21060 27020 21140
rect 10820 20700 11360 20800
rect 11300 20660 11360 20700
rect 8921 20634 9219 20660
rect 8921 20618 8934 20634
rect 8950 20618 8966 20634
rect 8982 20618 8998 20634
rect 9014 20618 9030 20634
rect 9046 20618 9062 20634
rect 9078 20618 9094 20634
rect 9110 20618 9126 20634
rect 9142 20618 9158 20634
rect 9174 20618 9190 20634
rect 9206 20618 9219 20634
rect 8921 20602 9219 20618
rect 8921 20586 8934 20602
rect 8950 20586 8966 20602
rect 8982 20586 8998 20602
rect 9014 20586 9030 20602
rect 9046 20586 9062 20602
rect 9078 20586 9094 20602
rect 9110 20586 9126 20602
rect 9142 20586 9158 20602
rect 9174 20586 9190 20602
rect 9206 20586 9219 20602
rect 8921 20561 9219 20586
rect 9540 20480 11340 20560
rect 9540 20340 11060 20480
rect 9540 9900 9720 20340
rect 9001 9882 9719 9900
rect 9001 9866 9016 9882
rect 9032 9866 9048 9882
rect 9064 9866 9080 9882
rect 9096 9866 9112 9882
rect 9128 9866 9144 9882
rect 9160 9866 9176 9882
rect 9192 9866 9208 9882
rect 9224 9866 9240 9882
rect 9256 9866 9272 9882
rect 9288 9866 9304 9882
rect 9320 9866 9336 9882
rect 9352 9866 9368 9882
rect 9384 9866 9400 9882
rect 9416 9866 9432 9882
rect 9448 9866 9464 9882
rect 9480 9866 9496 9882
rect 9512 9866 9528 9882
rect 9544 9866 9560 9882
rect 9576 9866 9592 9882
rect 9608 9866 9624 9882
rect 9640 9866 9656 9882
rect 9672 9866 9688 9882
rect 9704 9866 9719 9882
rect 9001 9850 9719 9866
rect 9001 9834 9016 9850
rect 9032 9834 9048 9850
rect 9064 9834 9080 9850
rect 9096 9834 9112 9850
rect 9128 9834 9144 9850
rect 9160 9834 9176 9850
rect 9192 9834 9208 9850
rect 9224 9834 9240 9850
rect 9256 9834 9272 9850
rect 9288 9834 9304 9850
rect 9320 9834 9336 9850
rect 9352 9834 9368 9850
rect 9384 9834 9400 9850
rect 9416 9834 9432 9850
rect 9448 9834 9464 9850
rect 9480 9834 9496 9850
rect 9512 9834 9528 9850
rect 9544 9834 9560 9850
rect 9576 9834 9592 9850
rect 9608 9834 9624 9850
rect 9640 9834 9656 9850
rect 9672 9834 9688 9850
rect 9704 9834 9719 9850
rect 9001 9818 9719 9834
rect 9001 9802 9016 9818
rect 9032 9802 9048 9818
rect 9064 9802 9080 9818
rect 9096 9802 9112 9818
rect 9128 9802 9144 9818
rect 9160 9802 9176 9818
rect 9192 9802 9208 9818
rect 9224 9802 9240 9818
rect 9256 9802 9272 9818
rect 9288 9802 9304 9818
rect 9320 9802 9336 9818
rect 9352 9802 9368 9818
rect 9384 9802 9400 9818
rect 9416 9802 9432 9818
rect 9448 9802 9464 9818
rect 9480 9802 9496 9818
rect 9512 9802 9528 9818
rect 9544 9802 9560 9818
rect 9576 9802 9592 9818
rect 9608 9802 9624 9818
rect 9640 9802 9656 9818
rect 9672 9802 9688 9818
rect 9704 9802 9719 9818
rect 9001 9786 9719 9802
rect 9001 9770 9016 9786
rect 9032 9770 9048 9786
rect 9064 9770 9080 9786
rect 9096 9770 9112 9786
rect 9128 9770 9144 9786
rect 9160 9770 9176 9786
rect 9192 9770 9208 9786
rect 9224 9770 9240 9786
rect 9256 9770 9272 9786
rect 9288 9770 9304 9786
rect 9320 9770 9336 9786
rect 9352 9770 9368 9786
rect 9384 9770 9400 9786
rect 9416 9770 9432 9786
rect 9448 9770 9464 9786
rect 9480 9770 9496 9786
rect 9512 9770 9528 9786
rect 9544 9770 9560 9786
rect 9576 9770 9592 9786
rect 9608 9770 9624 9786
rect 9640 9770 9656 9786
rect 9672 9770 9688 9786
rect 9704 9770 9719 9786
rect 26920 9880 27020 21060
rect 27120 12580 27220 21220
rect 27320 15280 27420 21380
rect 27520 17980 27620 21860
rect 27720 20680 27820 22560
rect 27720 20679 28780 20680
rect 27720 20654 29079 20679
rect 27720 20638 28794 20654
rect 28810 20638 28826 20654
rect 28842 20638 28858 20654
rect 28874 20638 28890 20654
rect 28906 20638 28922 20654
rect 28938 20638 28954 20654
rect 28970 20638 28986 20654
rect 29002 20638 29018 20654
rect 29034 20638 29050 20654
rect 29066 20638 29079 20654
rect 27720 20622 29079 20638
rect 27720 20606 28794 20622
rect 28810 20606 28826 20622
rect 28842 20606 28858 20622
rect 28874 20606 28890 20622
rect 28906 20606 28922 20622
rect 28938 20606 28954 20622
rect 28970 20606 28986 20622
rect 29002 20606 29018 20622
rect 29034 20606 29050 20622
rect 29066 20606 29079 20622
rect 27720 20581 29079 20606
rect 27720 20580 28780 20581
rect 27520 17979 28780 17980
rect 27520 17954 29079 17979
rect 27520 17938 28794 17954
rect 28810 17938 28826 17954
rect 28842 17938 28858 17954
rect 28874 17938 28890 17954
rect 28906 17938 28922 17954
rect 28938 17938 28954 17954
rect 28970 17938 28986 17954
rect 29002 17938 29018 17954
rect 29034 17938 29050 17954
rect 29066 17938 29079 17954
rect 27520 17922 29079 17938
rect 27520 17906 28794 17922
rect 28810 17906 28826 17922
rect 28842 17906 28858 17922
rect 28874 17906 28890 17922
rect 28906 17906 28922 17922
rect 28938 17906 28954 17922
rect 28970 17906 28986 17922
rect 29002 17906 29018 17922
rect 29034 17906 29050 17922
rect 29066 17906 29079 17922
rect 27520 17881 29079 17906
rect 27520 17880 28780 17881
rect 27320 15279 28780 15280
rect 27320 15254 29079 15279
rect 27320 15238 28794 15254
rect 28810 15238 28826 15254
rect 28842 15238 28858 15254
rect 28874 15238 28890 15254
rect 28906 15238 28922 15254
rect 28938 15238 28954 15254
rect 28970 15238 28986 15254
rect 29002 15238 29018 15254
rect 29034 15238 29050 15254
rect 29066 15238 29079 15254
rect 27320 15222 29079 15238
rect 27320 15206 28794 15222
rect 28810 15206 28826 15222
rect 28842 15206 28858 15222
rect 28874 15206 28890 15222
rect 28906 15206 28922 15222
rect 28938 15206 28954 15222
rect 28970 15206 28986 15222
rect 29002 15206 29018 15222
rect 29034 15206 29050 15222
rect 29066 15206 29079 15222
rect 27320 15181 29079 15206
rect 27320 15180 28780 15181
rect 27120 12579 28780 12580
rect 27120 12554 29079 12579
rect 27120 12538 28794 12554
rect 28810 12538 28826 12554
rect 28842 12538 28858 12554
rect 28874 12538 28890 12554
rect 28906 12538 28922 12554
rect 28938 12538 28954 12554
rect 28970 12538 28986 12554
rect 29002 12538 29018 12554
rect 29034 12538 29050 12554
rect 29066 12538 29079 12554
rect 27120 12522 29079 12538
rect 27120 12506 28794 12522
rect 28810 12506 28826 12522
rect 28842 12506 28858 12522
rect 28874 12506 28890 12522
rect 28906 12506 28922 12522
rect 28938 12506 28954 12522
rect 28970 12506 28986 12522
rect 29002 12506 29018 12522
rect 29034 12506 29050 12522
rect 29066 12506 29079 12522
rect 27120 12481 29079 12506
rect 27120 12480 28780 12481
rect 26920 9879 28780 9880
rect 26920 9854 29079 9879
rect 26920 9838 28794 9854
rect 28810 9838 28826 9854
rect 28842 9838 28858 9854
rect 28874 9838 28890 9854
rect 28906 9838 28922 9854
rect 28938 9838 28954 9854
rect 28970 9838 28986 9854
rect 29002 9838 29018 9854
rect 29034 9838 29050 9854
rect 29066 9838 29079 9854
rect 26920 9822 29079 9838
rect 26920 9806 28794 9822
rect 28810 9806 28826 9822
rect 28842 9806 28858 9822
rect 28874 9806 28890 9822
rect 28906 9806 28922 9822
rect 28938 9806 28954 9822
rect 28970 9806 28986 9822
rect 29002 9806 29018 9822
rect 29034 9806 29050 9822
rect 29066 9806 29079 9822
rect 26920 9781 29079 9806
rect 26920 9780 28780 9781
rect 9001 9754 9719 9770
rect 9001 9738 9016 9754
rect 9032 9738 9048 9754
rect 9064 9738 9080 9754
rect 9096 9738 9112 9754
rect 9128 9738 9144 9754
rect 9160 9738 9176 9754
rect 9192 9738 9208 9754
rect 9224 9738 9240 9754
rect 9256 9738 9272 9754
rect 9288 9738 9304 9754
rect 9320 9738 9336 9754
rect 9352 9738 9368 9754
rect 9384 9738 9400 9754
rect 9416 9738 9432 9754
rect 9448 9738 9464 9754
rect 9480 9738 9496 9754
rect 9512 9738 9528 9754
rect 9544 9738 9560 9754
rect 9576 9738 9592 9754
rect 9608 9738 9624 9754
rect 9640 9738 9656 9754
rect 9672 9738 9688 9754
rect 9704 9738 9719 9754
rect 9001 9721 9719 9738
<< end >>
