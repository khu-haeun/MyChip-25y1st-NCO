/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module phase_accumulator(
    output [1:0] Aout,
    input En,
    input [19:0] FCW,
    output ISout,
    output Vld,
    input clk
);

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _73__bF$buf0 ;
wire _73__bF$buf1 ;
wire _73__bF$buf2 ;
wire _73__bF$buf3 ;
wire _73__bF$buf4 ;
wire _218_ ;
wire _256_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _197_ ;
wire _7_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire ISout ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire [11:0] Atmp ;
wire _309_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _288_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire [19:0] acc_reg ;
wire _212_ ;
wire _250_ ;
wire _306_ ;
wire En_bF$buf0 ;
wire En_bF$buf1 ;
wire En_bF$buf2 ;
wire En_bF$buf3 ;
wire En_bF$buf4 ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire _282_ ;
wire _147_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _273_ ;
wire _138_ ;
wire _30_ ;
wire En ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _264_ ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _299_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _255_ ;
wire _293_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire [1:0] _311_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire _214_ ;
wire _252_ ;
wire _308_ ;
wire _117_ ;
wire _290_ ;
wire _155_ ;
wire [1:0] Aout ;
wire _193_ ;
wire _249_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire _305_ ;
wire _114_ ;
wire [19:0] FCW ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _284_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire RdyCtl_6_bF$buf0 ;
wire RdyCtl_6_bF$buf1 ;
wire RdyCtl_6_bF$buf2 ;
wire RdyCtl_6_bF$buf3 ;
wire RdyCtl_6_bF$buf4 ;
wire _281_ ;
wire _146_ ;
wire _184_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _275_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire [6:0] RdyCtl ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _298_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _157_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _310_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _307_ ;
wire _116_ ;
wire _154_ ;
wire _192_ ;
wire _248_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _245_ ;
wire _283_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _301_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _280_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

BUFX2 BUFX2_insert20 (
    .A(_73_),
    .Y(_73__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(_73_),
    .Y(_73__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(_73_),
    .Y(_73__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(_73_),
    .Y(_73__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .A(_73_),
    .Y(_73__bF$buf4)
);

BUFX2 BUFX2_insert15 (
    .A(En),
    .Y(En_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(En),
    .Y(En_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(En),
    .Y(En_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(En),
    .Y(En_bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(En),
    .Y(En_bF$buf4)
);

BUFX2 BUFX2_insert10 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert6 (
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf4)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf5)
);

OAI21X1 _313_ (
    .A(_129_),
    .B(_147_),
    .C(_139_),
    .Y(_153_)
);

INVX1 _314_ (
    .A(_153_),
    .Y(_154_)
);

OAI21X1 _315_ (
    .A(_152_),
    .B(_149_),
    .C(_154_),
    .Y(_155_)
);

AOI21X1 _316_ (
    .A(_150_),
    .B(_111_),
    .C(_155_),
    .Y(_156_)
);

NAND2X1 _317_ (
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_157_)
);

OR2X2 _318_ (
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_158_)
);

NAND2X1 _319_ (
    .A(_157_),
    .B(_158_),
    .Y(_159_)
);

OR2X2 _320_ (
    .A(_156_),
    .B(_159_),
    .Y(_160_)
);

NAND2X1 _321_ (
    .A(_159_),
    .B(_156_),
    .Y(_161_)
);

NAND2X1 _322_ (
    .A(_161_),
    .B(_160_),
    .Y(_162_)
);

OAI21X1 _323_ (
    .A(acc_reg[8]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf4),
    .Y(_163_)
);

AOI21X1 _324_ (
    .A(_162_),
    .B(RdyCtl_6_bF$buf3),
    .C(_163_),
    .Y(_15_)
);

OAI21X1 _325_ (
    .A(_159_),
    .B(_156_),
    .C(_157_),
    .Y(_164_)
);

NAND2X1 _326_ (
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_165_)
);

INVX1 _327_ (
    .A(acc_reg[9]),
    .Y(_166_)
);

INVX1 _328_ (
    .A(FCW[9]),
    .Y(_167_)
);

NAND2X1 _329_ (
    .A(_166_),
    .B(_167_),
    .Y(_168_)
);

NAND2X1 _330_ (
    .A(_165_),
    .B(_168_),
    .Y(_169_)
);

NAND2X1 _331_ (
    .A(_169_),
    .B(_164_),
    .Y(_170_)
);

NOR2X1 _332_ (
    .A(_169_),
    .B(_164_),
    .Y(_171_)
);

NOR2X1 _333_ (
    .A(_73__bF$buf4),
    .B(_171_),
    .Y(_172_)
);

OAI21X1 _334_ (
    .A(acc_reg[9]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf3),
    .Y(_173_)
);

AOI21X1 _335_ (
    .A(_172_),
    .B(_170_),
    .C(_173_),
    .Y(_16_)
);

NOR2X1 _336_ (
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_174_)
);

OAI21X1 _337_ (
    .A(_157_),
    .B(_174_),
    .C(_165_),
    .Y(_175_)
);

INVX1 _338_ (
    .A(_175_),
    .Y(_176_)
);

OR2X2 _339_ (
    .A(_169_),
    .B(_159_),
    .Y(_177_)
);

OAI21X1 _340_ (
    .A(_177_),
    .B(_156_),
    .C(_176_),
    .Y(_178_)
);

AND2X2 _341_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_179_)
);

NOR2X1 _342_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_180_)
);

NOR2X1 _343_ (
    .A(_180_),
    .B(_179_),
    .Y(_181_)
);

NAND2X1 _344_ (
    .A(_181_),
    .B(_178_),
    .Y(_182_)
);

OR2X2 _345_ (
    .A(_178_),
    .B(_181_),
    .Y(_183_)
);

NAND2X1 _346_ (
    .A(_182_),
    .B(_183_),
    .Y(_184_)
);

OAI21X1 _347_ (
    .A(acc_reg[10]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf2),
    .Y(_185_)
);

AOI21X1 _348_ (
    .A(_184_),
    .B(RdyCtl_6_bF$buf0),
    .C(_185_),
    .Y(_17_)
);

NAND2X1 _349_ (
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_186_)
);

NAND2X1 _350_ (
    .A(_186_),
    .B(_182_),
    .Y(_187_)
);

AND2X2 _351_ (
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_188_)
);

NOR2X1 _352_ (
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_189_)
);

NOR2X1 _353_ (
    .A(_189_),
    .B(_188_),
    .Y(_190_)
);

INVX1 _354_ (
    .A(_190_),
    .Y(_191_)
);

OR2X2 _355_ (
    .A(_187_),
    .B(_191_),
    .Y(_192_)
);

AOI21X1 _356_ (
    .A(_187_),
    .B(_191_),
    .C(_73__bF$buf3),
    .Y(_193_)
);

OAI21X1 _357_ (
    .A(acc_reg[11]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_194_)
);

AOI21X1 _358_ (
    .A(_192_),
    .B(_193_),
    .C(_194_),
    .Y(_18_)
);

NAND2X1 _359_ (
    .A(acc_reg[12]),
    .B(_73__bF$buf2),
    .Y(_195_)
);

NOR2X1 _360_ (
    .A(_159_),
    .B(_169_),
    .Y(_196_)
);

NAND3X1 _361_ (
    .A(_181_),
    .B(_190_),
    .C(_196_),
    .Y(_197_)
);

NAND3X1 _362_ (
    .A(_175_),
    .B(_181_),
    .C(_190_),
    .Y(_198_)
);

INVX1 _363_ (
    .A(_189_),
    .Y(_199_)
);

AOI21X1 _364_ (
    .A(_199_),
    .B(_179_),
    .C(_188_),
    .Y(_200_)
);

AND2X2 _365_ (
    .A(_198_),
    .B(_200_),
    .Y(_201_)
);

OAI21X1 _366_ (
    .A(_197_),
    .B(_156_),
    .C(_201_),
    .Y(_202_)
);

NAND2X1 _367_ (
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_203_)
);

OR2X2 _368_ (
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_204_)
);

NAND2X1 _369_ (
    .A(_203_),
    .B(_204_),
    .Y(_205_)
);

NOR2X1 _370_ (
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

AND2X2 _371_ (
    .A(_202_),
    .B(_205_),
    .Y(_207_)
);

OAI21X1 _372_ (
    .A(_206_),
    .B(_207_),
    .C(RdyCtl_6_bF$buf3),
    .Y(_208_)
);

AOI21X1 _373_ (
    .A(_208_),
    .B(_195_),
    .C(_74_),
    .Y(_19_)
);

INVX1 _374_ (
    .A(_202_),
    .Y(_209_)
);

OAI21X1 _375_ (
    .A(_205_),
    .B(_209_),
    .C(_203_),
    .Y(_210_)
);

NAND2X1 _376_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_211_)
);

OR2X2 _377_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_212_)
);

NAND2X1 _378_ (
    .A(_211_),
    .B(_212_),
    .Y(_213_)
);

OR2X2 _379_ (
    .A(_210_),
    .B(_213_),
    .Y(_214_)
);

AOI21X1 _380_ (
    .A(_210_),
    .B(_213_),
    .C(_73__bF$buf1),
    .Y(_215_)
);

OAI21X1 _381_ (
    .A(acc_reg[13]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf0),
    .Y(_216_)
);

AOI21X1 _382_ (
    .A(_214_),
    .B(_215_),
    .C(_216_),
    .Y(_20_)
);

NOR2X1 _383_ (
    .A(_205_),
    .B(_213_),
    .Y(_217_)
);

NOR2X1 _384_ (
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_218_)
);

OAI21X1 _385_ (
    .A(_203_),
    .B(_218_),
    .C(_211_),
    .Y(_219_)
);

AOI21X1 _386_ (
    .A(_202_),
    .B(_217_),
    .C(_219_),
    .Y(_220_)
);

AND2X2 _387_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_221_)
);

NOR2X1 _388_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_222_)
);

OR2X2 _389_ (
    .A(_221_),
    .B(_222_),
    .Y(_223_)
);

OR2X2 _390_ (
    .A(_220_),
    .B(_223_),
    .Y(_224_)
);

OAI21X1 _391_ (
    .A(_221_),
    .B(_222_),
    .C(_220_),
    .Y(_225_)
);

NAND2X1 _392_ (
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

OAI21X1 _393_ (
    .A(acc_reg[14]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf4),
    .Y(_227_)
);

AOI21X1 _394_ (
    .A(_226_),
    .B(RdyCtl_6_bF$buf0),
    .C(_227_),
    .Y(_21_)
);

NAND2X1 _395_ (
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_228_)
);

NAND2X1 _396_ (
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_229_)
);

INVX1 _397_ (
    .A(_229_),
    .Y(_230_)
);

NOR2X1 _398_ (
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_231_)
);

NOR2X1 _399_ (
    .A(_231_),
    .B(_230_),
    .Y(_232_)
);

NAND3X1 _400_ (
    .A(_228_),
    .B(_232_),
    .C(_224_),
    .Y(_233_)
);

OAI21X1 _401_ (
    .A(_223_),
    .B(_220_),
    .C(_228_),
    .Y(_234_)
);

INVX1 _402_ (
    .A(_231_),
    .Y(_235_)
);

NAND2X1 _403_ (
    .A(_229_),
    .B(_235_),
    .Y(_236_)
);

AOI21X1 _404_ (
    .A(_234_),
    .B(_236_),
    .C(_73__bF$buf0),
    .Y(_237_)
);

OAI21X1 _405_ (
    .A(acc_reg[15]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf3),
    .Y(_238_)
);

AOI21X1 _406_ (
    .A(_233_),
    .B(_237_),
    .C(_238_),
    .Y(_22_)
);

NOR2X1 _407_ (
    .A(_222_),
    .B(_221_),
    .Y(_239_)
);

NAND3X1 _408_ (
    .A(_239_),
    .B(_232_),
    .C(_217_),
    .Y(_240_)
);

OR2X2 _409_ (
    .A(_197_),
    .B(_240_),
    .Y(_241_)
);

NAND2X1 _410_ (
    .A(_200_),
    .B(_198_),
    .Y(_242_)
);

NOR2X1 _411_ (
    .A(_223_),
    .B(_236_),
    .Y(_243_)
);

AND2X2 _412_ (
    .A(_243_),
    .B(_217_),
    .Y(_244_)
);

NAND3X1 _413_ (
    .A(_219_),
    .B(_239_),
    .C(_232_),
    .Y(_245_)
);

AOI21X1 _414_ (
    .A(_235_),
    .B(_221_),
    .C(_230_),
    .Y(_246_)
);

NAND2X1 _415_ (
    .A(_246_),
    .B(_245_),
    .Y(_247_)
);

AOI21X1 _416_ (
    .A(_244_),
    .B(_242_),
    .C(_247_),
    .Y(_248_)
);

OAI21X1 _417_ (
    .A(_156_),
    .B(_241_),
    .C(_248_),
    .Y(_249_)
);

AND2X2 _418_ (
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_250_)
);

NOR2X1 _419_ (
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_251_)
);

NOR2X1 _420_ (
    .A(_251_),
    .B(_250_),
    .Y(_252_)
);

NAND2X1 _421_ (
    .A(_252_),
    .B(_249_),
    .Y(_253_)
);

NOR2X1 _422_ (
    .A(_141_),
    .B(_131_),
    .Y(_254_)
);

NAND2X1 _423_ (
    .A(_254_),
    .B(_127_),
    .Y(_255_)
);

AOI21X1 _424_ (
    .A(_254_),
    .B(_126_),
    .C(_153_),
    .Y(_256_)
);

OAI21X1 _425_ (
    .A(_255_),
    .B(_107_),
    .C(_256_),
    .Y(_257_)
);

NOR2X1 _426_ (
    .A(_197_),
    .B(_240_),
    .Y(_258_)
);

AND2X2 _427_ (
    .A(_245_),
    .B(_246_),
    .Y(_259_)
);

OAI21X1 _428_ (
    .A(_240_),
    .B(_201_),
    .C(_259_),
    .Y(_260_)
);

AOI21X1 _429_ (
    .A(_257_),
    .B(_258_),
    .C(_260_),
    .Y(_261_)
);

OAI21X1 _430_ (
    .A(_250_),
    .B(_251_),
    .C(_261_),
    .Y(_262_)
);

NAND2X1 _431_ (
    .A(_262_),
    .B(_253_),
    .Y(_263_)
);

OAI21X1 _432_ (
    .A(acc_reg[16]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_264_)
);

AOI21X1 _433_ (
    .A(_263_),
    .B(RdyCtl_6_bF$buf2),
    .C(_264_),
    .Y(_23_)
);

AOI21X1 _434_ (
    .A(_249_),
    .B(_252_),
    .C(_250_),
    .Y(_265_)
);

AND2X2 _435_ (
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_266_)
);

NOR2X1 _436_ (
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_267_)
);

NOR2X1 _437_ (
    .A(_267_),
    .B(_266_),
    .Y(_268_)
);

OR2X2 _438_ (
    .A(_265_),
    .B(_268_),
    .Y(_269_)
);

AOI21X1 _439_ (
    .A(_265_),
    .B(_268_),
    .C(_73__bF$buf4),
    .Y(_270_)
);

OAI21X1 _440_ (
    .A(acc_reg[17]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf1),
    .Y(_271_)
);

AOI21X1 _441_ (
    .A(_269_),
    .B(_270_),
    .C(_271_),
    .Y(_24_)
);

NAND2X1 _442_ (
    .A(_252_),
    .B(_268_),
    .Y(_272_)
);

AOI21X1 _443_ (
    .A(_268_),
    .B(_250_),
    .C(_266_),
    .Y(_273_)
);

OAI21X1 _444_ (
    .A(_272_),
    .B(_261_),
    .C(_273_),
    .Y(_274_)
);

INVX1 _445_ (
    .A(FCW[18]),
    .Y(_275_)
);

NOR2X1 _446_ (
    .A(_68_),
    .B(_275_),
    .Y(_276_)
);

NOR2X1 _447_ (
    .A(acc_reg[18]),
    .B(FCW[18]),
    .Y(_277_)
);

NOR2X1 _448_ (
    .A(_277_),
    .B(_276_),
    .Y(_278_)
);

NAND2X1 _449_ (
    .A(_278_),
    .B(_274_),
    .Y(_279_)
);

INVX1 _450_ (
    .A(_272_),
    .Y(_280_)
);

INVX1 _451_ (
    .A(_273_),
    .Y(_281_)
);

AOI21X1 _452_ (
    .A(_249_),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

OAI21X1 _453_ (
    .A(_276_),
    .B(_277_),
    .C(_282_),
    .Y(_283_)
);

NAND2X1 _454_ (
    .A(_279_),
    .B(_283_),
    .Y(_284_)
);

OAI21X1 _455_ (
    .A(acc_reg[18]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_285_)
);

AOI21X1 _456_ (
    .A(_284_),
    .B(RdyCtl_6_bF$buf4),
    .C(_285_),
    .Y(_25_)
);

INVX1 _457_ (
    .A(_0_),
    .Y(_286_)
);

NAND2X1 _458_ (
    .A(acc_reg[19]),
    .B(En_bF$buf4),
    .Y(_287_)
);

INVX1 _459_ (
    .A(_276_),
    .Y(_288_)
);

OAI21X1 _460_ (
    .A(_277_),
    .B(_282_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _461_ (
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_290_)
);

OR2X2 _462_ (
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_291_)
);

NAND2X1 _463_ (
    .A(_290_),
    .B(_291_),
    .Y(_292_)
);

NAND2X1 _464_ (
    .A(_292_),
    .B(_289_),
    .Y(_293_)
);

AOI21X1 _465_ (
    .A(_274_),
    .B(_278_),
    .C(_276_),
    .Y(_294_)
);

INVX1 _466_ (
    .A(_292_),
    .Y(_295_)
);

AOI21X1 _467_ (
    .A(_294_),
    .B(_295_),
    .C(_73__bF$buf3),
    .Y(_296_)
);

AOI22X1 _468_ (
    .A(_286_),
    .B(_287_),
    .C(_296_),
    .D(_293_),
    .Y(_26_)
);

NOR2X1 _469_ (
    .A(Atmp[0]),
    .B(RdyCtl_6_bF$buf3),
    .Y(_297_)
);

OAI21X1 _470_ (
    .A(acc_reg[8]),
    .B(_73__bF$buf2),
    .C(En_bF$buf3),
    .Y(_298_)
);

NOR2X1 _471_ (
    .A(_297_),
    .B(_298_),
    .Y(_27_)
);

NOR2X1 _472_ (
    .A(Atmp[1]),
    .B(RdyCtl_6_bF$buf2),
    .Y(_299_)
);

OAI21X1 _473_ (
    .A(acc_reg[9]),
    .B(_73__bF$buf1),
    .C(En_bF$buf2),
    .Y(_300_)
);

NOR2X1 _474_ (
    .A(_299_),
    .B(_300_),
    .Y(_28_)
);

OAI21X1 _475_ (
    .A(acc_reg[10]),
    .B(_73__bF$buf0),
    .C(En_bF$buf1),
    .Y(_301_)
);

AOI21X1 _476_ (
    .A(_51_),
    .B(_73__bF$buf4),
    .C(_301_),
    .Y(_29_)
);

OAI21X1 _477_ (
    .A(acc_reg[11]),
    .B(_73__bF$buf3),
    .C(En_bF$buf0),
    .Y(_302_)
);

AOI21X1 _478_ (
    .A(_62_),
    .B(_73__bF$buf2),
    .C(_302_),
    .Y(_30_)
);

OAI21X1 _479_ (
    .A(acc_reg[12]),
    .B(_73__bF$buf1),
    .C(En_bF$buf4),
    .Y(_303_)
);

AOI21X1 _480_ (
    .A(_39_),
    .B(_73__bF$buf0),
    .C(_303_),
    .Y(_31_)
);

OAI21X1 _481_ (
    .A(acc_reg[13]),
    .B(_73__bF$buf4),
    .C(En_bF$buf3),
    .Y(_304_)
);

AOI21X1 _482_ (
    .A(_55_),
    .B(_73__bF$buf3),
    .C(_304_),
    .Y(_32_)
);

OAI21X1 _483_ (
    .A(acc_reg[14]),
    .B(_73__bF$buf2),
    .C(En_bF$buf2),
    .Y(_305_)
);

AOI21X1 _484_ (
    .A(_41_),
    .B(_73__bF$buf1),
    .C(_305_),
    .Y(_33_)
);

OAI21X1 _485_ (
    .A(acc_reg[15]),
    .B(_73__bF$buf0),
    .C(En_bF$buf1),
    .Y(_306_)
);

AOI21X1 _486_ (
    .A(_58_),
    .B(_73__bF$buf4),
    .C(_306_),
    .Y(_34_)
);

OAI21X1 _487_ (
    .A(acc_reg[16]),
    .B(_73__bF$buf3),
    .C(En_bF$buf0),
    .Y(_307_)
);

AOI21X1 _488_ (
    .A(_43_),
    .B(_73__bF$buf2),
    .C(_307_),
    .Y(_35_)
);

OAI21X1 _489_ (
    .A(acc_reg[17]),
    .B(_73__bF$buf1),
    .C(En_bF$buf4),
    .Y(_308_)
);

AOI21X1 _490_ (
    .A(_56_),
    .B(_73__bF$buf0),
    .C(_308_),
    .Y(_36_)
);

NOR2X1 _491_ (
    .A(Atmp[11]),
    .B(RdyCtl_6_bF$buf1),
    .Y(_309_)
);

OAI21X1 _492_ (
    .A(acc_reg[18]),
    .B(_73__bF$buf4),
    .C(En_bF$buf3),
    .Y(_310_)
);

NOR2X1 _493_ (
    .A(_309_),
    .B(_310_),
    .Y(_37_)
);

INVX1 _494_ (
    .A(Atmp[4]),
    .Y(_39_)
);

INVX1 _495_ (
    .A(RdyCtl[2]),
    .Y(_40_)
);

INVX1 _496_ (
    .A(Atmp[6]),
    .Y(_41_)
);

INVX1 _497_ (
    .A(RdyCtl[3]),
    .Y(_42_)
);

INVX1 _498_ (
    .A(Atmp[8]),
    .Y(_43_)
);

INVX1 _499_ (
    .A(RdyCtl[4]),
    .Y(_44_)
);

NAND2X1 _500_ (
    .A(Atmp[11]),
    .B(_44_),
    .Y(_45_)
);

OAI21X1 _501_ (
    .A(_43_),
    .B(_44_),
    .C(_45_),
    .Y(_46_)
);

NAND2X1 _502_ (
    .A(_42_),
    .B(_46_),
    .Y(_47_)
);

OAI21X1 _503_ (
    .A(_41_),
    .B(_42_),
    .C(_47_),
    .Y(_48_)
);

NAND2X1 _504_ (
    .A(_40_),
    .B(_48_),
    .Y(_49_)
);

OAI21X1 _505_ (
    .A(_39_),
    .B(_40_),
    .C(_49_),
    .Y(_50_)
);

INVX1 _506_ (
    .A(Atmp[2]),
    .Y(_51_)
);

NAND2X1 _507_ (
    .A(RdyCtl[1]),
    .B(_51_),
    .Y(_52_)
);

OAI21X1 _508_ (
    .A(RdyCtl[1]),
    .B(_50_),
    .C(_52_),
    .Y(_53_)
);

NAND2X1 _509_ (
    .A(Atmp[0]),
    .B(RdyCtl[0]),
    .Y(_54_)
);

OAI21X1 _510_ (
    .A(RdyCtl[0]),
    .B(_53_),
    .C(_54_),
    .Y(_311_[0])
);

INVX1 _511_ (
    .A(Atmp[5]),
    .Y(_55_)
);

INVX1 _512_ (
    .A(Atmp[9]),
    .Y(_56_)
);

OAI21X1 _513_ (
    .A(_44_),
    .B(_56_),
    .C(_45_),
    .Y(_57_)
);

INVX1 _514_ (
    .A(Atmp[7]),
    .Y(_58_)
);

AOI21X1 _515_ (
    .A(_58_),
    .B(RdyCtl[3]),
    .C(RdyCtl[2]),
    .Y(_59_)
);

OAI21X1 _516_ (
    .A(RdyCtl[3]),
    .B(_57_),
    .C(_59_),
    .Y(_60_)
);

OAI21X1 _517_ (
    .A(_40_),
    .B(_55_),
    .C(_60_),
    .Y(_61_)
);

INVX1 _518_ (
    .A(Atmp[3]),
    .Y(_62_)
);

NAND2X1 _519_ (
    .A(RdyCtl[1]),
    .B(_62_),
    .Y(_63_)
);

OAI21X1 _520_ (
    .A(RdyCtl[1]),
    .B(_61_),
    .C(_63_),
    .Y(_64_)
);

NAND2X1 _521_ (
    .A(RdyCtl[0]),
    .B(Atmp[1]),
    .Y(_65_)
);

OAI21X1 _522_ (
    .A(RdyCtl[0]),
    .B(_64_),
    .C(_65_),
    .Y(_311_[1])
);

INVX1 _523_ (
    .A(RdyCtl[5]),
    .Y(_66_)
);

NAND2X1 _524_ (
    .A(acc_reg[18]),
    .B(acc_reg[19]),
    .Y(_67_)
);

INVX1 _525_ (
    .A(acc_reg[18]),
    .Y(_68_)
);

INVX1 _526_ (
    .A(acc_reg[19]),
    .Y(_69_)
);

NAND2X1 _527_ (
    .A(_68_),
    .B(_69_),
    .Y(_70_)
);

NAND2X1 _528_ (
    .A(_67_),
    .B(_70_),
    .Y(_71_)
);

NAND2X1 _529_ (
    .A(_312_),
    .B(_66_),
    .Y(_72_)
);

OAI21X1 _530_ (
    .A(_66_),
    .B(_71_),
    .C(_72_),
    .Y(_38_)
);

INVX8 _531_ (
    .A(RdyCtl_6_bF$buf0),
    .Y(_73_)
);

INVX2 _532_ (
    .A(En_bF$buf2),
    .Y(_74_)
);

NOR2X1 _533_ (
    .A(_73__bF$buf3),
    .B(_74_),
    .Y(_0_)
);

AND2X2 _534_ (
    .A(RdyCtl[0]),
    .B(En_bF$buf1),
    .Y(_1_)
);

AND2X2 _535_ (
    .A(RdyCtl[1]),
    .B(En_bF$buf0),
    .Y(_2_)
);

NOR2X1 _536_ (
    .A(_40_),
    .B(_74_),
    .Y(_3_)
);

NOR2X1 _537_ (
    .A(_42_),
    .B(_74_),
    .Y(_4_)
);

NAND2X1 _538_ (
    .A(En_bF$buf4),
    .B(_44_),
    .Y(_5_)
);

NOR2X1 _539_ (
    .A(_66_),
    .B(_74_),
    .Y(_6_)
);

INVX1 _540_ (
    .A(acc_reg[0]),
    .Y(_75_)
);

NAND2X1 _541_ (
    .A(FCW[0]),
    .B(RdyCtl_6_bF$buf4),
    .Y(_76_)
);

OAI21X1 _542_ (
    .A(_75_),
    .B(_76_),
    .C(En_bF$buf3),
    .Y(_77_)
);

AOI21X1 _543_ (
    .A(_75_),
    .B(_76_),
    .C(_77_),
    .Y(_7_)
);

NAND2X1 _544_ (
    .A(acc_reg[0]),
    .B(FCW[0]),
    .Y(_78_)
);

NAND2X1 _545_ (
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_79_)
);

INVX1 _546_ (
    .A(_79_),
    .Y(_80_)
);

NOR2X1 _547_ (
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_81_)
);

OAI21X1 _548_ (
    .A(_81_),
    .B(_80_),
    .C(_78_),
    .Y(_82_)
);

OR2X2 _549_ (
    .A(_80_),
    .B(_81_),
    .Y(_83_)
);

NOR2X1 _550_ (
    .A(_78_),
    .B(_83_),
    .Y(_84_)
);

INVX1 _551_ (
    .A(_84_),
    .Y(_85_)
);

NAND2X1 _552_ (
    .A(_82_),
    .B(_85_),
    .Y(_86_)
);

OAI21X1 _553_ (
    .A(acc_reg[1]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_87_)
);

AOI21X1 _554_ (
    .A(_86_),
    .B(RdyCtl_6_bF$buf2),
    .C(_87_),
    .Y(_8_)
);

OAI21X1 _555_ (
    .A(_78_),
    .B(_81_),
    .C(_79_),
    .Y(_88_)
);

AND2X2 _556_ (
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_89_)
);

NOR2X1 _557_ (
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_90_)
);

NOR2X1 _558_ (
    .A(_90_),
    .B(_89_),
    .Y(_91_)
);

AND2X2 _559_ (
    .A(_91_),
    .B(_88_),
    .Y(_92_)
);

NOR2X1 _560_ (
    .A(_73__bF$buf2),
    .B(_92_),
    .Y(_93_)
);

OAI21X1 _561_ (
    .A(_88_),
    .B(_91_),
    .C(_93_),
    .Y(_94_)
);

NAND2X1 _562_ (
    .A(acc_reg[2]),
    .B(_73__bF$buf1),
    .Y(_95_)
);

AOI21X1 _563_ (
    .A(_94_),
    .B(_95_),
    .C(_74_),
    .Y(_9_)
);

OAI21X1 _564_ (
    .A(acc_reg[3]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf1),
    .Y(_96_)
);

AND2X2 _565_ (
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_97_)
);

NOR2X1 _566_ (
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_98_)
);

NOR2X1 _567_ (
    .A(_98_),
    .B(_97_),
    .Y(_99_)
);

OAI21X1 _568_ (
    .A(_89_),
    .B(_92_),
    .C(_99_),
    .Y(_100_)
);

NOR2X1 _569_ (
    .A(_89_),
    .B(_92_),
    .Y(_101_)
);

OAI21X1 _570_ (
    .A(_97_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

NAND2X1 _571_ (
    .A(_100_),
    .B(_102_),
    .Y(_103_)
);

AOI21X1 _572_ (
    .A(_103_),
    .B(RdyCtl_6_bF$buf0),
    .C(_96_),
    .Y(_10_)
);

NAND3X1 _573_ (
    .A(_88_),
    .B(_91_),
    .C(_99_),
    .Y(_104_)
);

INVX1 _574_ (
    .A(_98_),
    .Y(_105_)
);

AOI21X1 _575_ (
    .A(_105_),
    .B(_89_),
    .C(_97_),
    .Y(_106_)
);

AND2X2 _576_ (
    .A(_104_),
    .B(_106_),
    .Y(_107_)
);

AND2X2 _577_ (
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_108_)
);

NOR2X1 _578_ (
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_109_)
);

OAI21X1 _579_ (
    .A(_108_),
    .B(_109_),
    .C(_107_),
    .Y(_110_)
);

NAND2X1 _580_ (
    .A(_106_),
    .B(_104_),
    .Y(_111_)
);

NOR2X1 _581_ (
    .A(_109_),
    .B(_108_),
    .Y(_112_)
);

NAND2X1 _582_ (
    .A(_112_),
    .B(_111_),
    .Y(_113_)
);

NAND2X1 _583_ (
    .A(_113_),
    .B(_110_),
    .Y(_114_)
);

OAI21X1 _584_ (
    .A(acc_reg[4]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf0),
    .Y(_115_)
);

AOI21X1 _585_ (
    .A(_114_),
    .B(RdyCtl_6_bF$buf3),
    .C(_115_),
    .Y(_11_)
);

AOI21X1 _586_ (
    .A(_111_),
    .B(_112_),
    .C(_108_),
    .Y(_116_)
);

AND2X2 _587_ (
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_117_)
);

NOR2X1 _588_ (
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_118_)
);

NOR2X1 _589_ (
    .A(_118_),
    .B(_117_),
    .Y(_119_)
);

NAND2X1 _590_ (
    .A(_119_),
    .B(_116_),
    .Y(_120_)
);

NOR2X1 _591_ (
    .A(_119_),
    .B(_116_),
    .Y(_121_)
);

NOR2X1 _592_ (
    .A(_73__bF$buf0),
    .B(_121_),
    .Y(_122_)
);

OAI21X1 _593_ (
    .A(acc_reg[5]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf4),
    .Y(_123_)
);

AOI21X1 _594_ (
    .A(_122_),
    .B(_120_),
    .C(_123_),
    .Y(_12_)
);

INVX1 _595_ (
    .A(_108_),
    .Y(_124_)
);

INVX1 _596_ (
    .A(_117_),
    .Y(_125_)
);

OAI21X1 _597_ (
    .A(_118_),
    .B(_124_),
    .C(_125_),
    .Y(_126_)
);

AND2X2 _598_ (
    .A(_112_),
    .B(_119_),
    .Y(_127_)
);

AOI21X1 _599_ (
    .A(_111_),
    .B(_127_),
    .C(_126_),
    .Y(_128_)
);

NAND2X1 _600_ (
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_129_)
);

OR2X2 _601_ (
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_130_)
);

NAND2X1 _602_ (
    .A(_129_),
    .B(_130_),
    .Y(_131_)
);

OR2X2 _603_ (
    .A(_128_),
    .B(_131_),
    .Y(_132_)
);

INVX1 _604_ (
    .A(_129_),
    .Y(_133_)
);

INVX1 _605_ (
    .A(_130_),
    .Y(_134_)
);

OAI21X1 _606_ (
    .A(_133_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

NAND2X1 _607_ (
    .A(_135_),
    .B(_132_),
    .Y(_136_)
);

OAI21X1 _608_ (
    .A(acc_reg[6]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf3),
    .Y(_137_)
);

AOI21X1 _609_ (
    .A(_136_),
    .B(RdyCtl_6_bF$buf0),
    .C(_137_),
    .Y(_13_)
);

OAI21X1 _610_ (
    .A(_134_),
    .B(_128_),
    .C(_129_),
    .Y(_138_)
);

NAND2X1 _611_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_139_)
);

OR2X2 _612_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_140_)
);

NAND2X1 _613_ (
    .A(_139_),
    .B(_140_),
    .Y(_141_)
);

OR2X2 _614_ (
    .A(_138_),
    .B(_141_),
    .Y(_142_)
);

AOI21X1 _615_ (
    .A(_138_),
    .B(_141_),
    .C(_73__bF$buf4),
    .Y(_143_)
);

OAI21X1 _616_ (
    .A(acc_reg[7]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf2),
    .Y(_144_)
);

AOI21X1 _617_ (
    .A(_142_),
    .B(_143_),
    .C(_144_),
    .Y(_14_)
);

NAND2X1 _618_ (
    .A(_112_),
    .B(_119_),
    .Y(_145_)
);

AND2X2 _619_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_146_)
);

NOR2X1 _620_ (
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_147_)
);

NOR2X1 _621_ (
    .A(_147_),
    .B(_146_),
    .Y(_148_)
);

NAND3X1 _622_ (
    .A(_129_),
    .B(_130_),
    .C(_148_),
    .Y(_149_)
);

NOR2X1 _623_ (
    .A(_145_),
    .B(_149_),
    .Y(_150_)
);

INVX1 _624_ (
    .A(_118_),
    .Y(_151_)
);

AOI21X1 _625_ (
    .A(_151_),
    .B(_108_),
    .C(_117_),
    .Y(_152_)
);

DFFPOSX1 _626_ (
    .CLK(clk_bF$buf5),
    .D(_0_),
    .Q(RdyCtl[0])
);

DFFPOSX1 _627_ (
    .CLK(clk_bF$buf4),
    .D(_1_),
    .Q(RdyCtl[1])
);

DFFPOSX1 _628_ (
    .CLK(clk_bF$buf3),
    .D(_2_),
    .Q(RdyCtl[2])
);

DFFPOSX1 _629_ (
    .CLK(clk_bF$buf2),
    .D(_3_),
    .Q(RdyCtl[3])
);

DFFPOSX1 _630_ (
    .CLK(clk_bF$buf1),
    .D(_4_),
    .Q(RdyCtl[4])
);

DFFPOSX1 _631_ (
    .CLK(clk_bF$buf0),
    .D(_5_),
    .Q(RdyCtl[5])
);

DFFPOSX1 _632_ (
    .CLK(clk_bF$buf5),
    .D(_6_),
    .Q(RdyCtl[6])
);

DFFPOSX1 _633_ (
    .CLK(clk_bF$buf4),
    .D(_7_),
    .Q(acc_reg[0])
);

DFFPOSX1 _634_ (
    .CLK(clk_bF$buf3),
    .D(_8_),
    .Q(acc_reg[1])
);

DFFPOSX1 _635_ (
    .CLK(clk_bF$buf2),
    .D(_9_),
    .Q(acc_reg[2])
);

DFFPOSX1 _636_ (
    .CLK(clk_bF$buf1),
    .D(_10_),
    .Q(acc_reg[3])
);

DFFPOSX1 _637_ (
    .CLK(clk_bF$buf0),
    .D(_11_),
    .Q(acc_reg[4])
);

DFFPOSX1 _638_ (
    .CLK(clk_bF$buf5),
    .D(_12_),
    .Q(acc_reg[5])
);

DFFPOSX1 _639_ (
    .CLK(clk_bF$buf4),
    .D(_13_),
    .Q(acc_reg[6])
);

DFFPOSX1 _640_ (
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(acc_reg[7])
);

DFFPOSX1 _641_ (
    .CLK(clk_bF$buf2),
    .D(_15_),
    .Q(acc_reg[8])
);

DFFPOSX1 _642_ (
    .CLK(clk_bF$buf1),
    .D(_16_),
    .Q(acc_reg[9])
);

DFFPOSX1 _643_ (
    .CLK(clk_bF$buf0),
    .D(_17_),
    .Q(acc_reg[10])
);

DFFPOSX1 _644_ (
    .CLK(clk_bF$buf5),
    .D(_18_),
    .Q(acc_reg[11])
);

DFFPOSX1 _645_ (
    .CLK(clk_bF$buf4),
    .D(_19_),
    .Q(acc_reg[12])
);

DFFPOSX1 _646_ (
    .CLK(clk_bF$buf3),
    .D(_20_),
    .Q(acc_reg[13])
);

DFFPOSX1 _647_ (
    .CLK(clk_bF$buf2),
    .D(_21_),
    .Q(acc_reg[14])
);

DFFPOSX1 _648_ (
    .CLK(clk_bF$buf1),
    .D(_22_),
    .Q(acc_reg[15])
);

DFFPOSX1 _649_ (
    .CLK(clk_bF$buf0),
    .D(_23_),
    .Q(acc_reg[16])
);

DFFPOSX1 _650_ (
    .CLK(clk_bF$buf5),
    .D(_24_),
    .Q(acc_reg[17])
);

DFFPOSX1 _651_ (
    .CLK(clk_bF$buf4),
    .D(_25_),
    .Q(acc_reg[18])
);

DFFPOSX1 _652_ (
    .CLK(clk_bF$buf3),
    .D(_26_),
    .Q(acc_reg[19])
);

DFFPOSX1 _653_ (
    .CLK(clk_bF$buf2),
    .D(_27_),
    .Q(Atmp[0])
);

DFFPOSX1 _654_ (
    .CLK(clk_bF$buf1),
    .D(_28_),
    .Q(Atmp[1])
);

DFFPOSX1 _655_ (
    .CLK(clk_bF$buf0),
    .D(_29_),
    .Q(Atmp[2])
);

DFFPOSX1 _656_ (
    .CLK(clk_bF$buf5),
    .D(_30_),
    .Q(Atmp[3])
);

DFFPOSX1 _657_ (
    .CLK(clk_bF$buf4),
    .D(_31_),
    .Q(Atmp[4])
);

DFFPOSX1 _658_ (
    .CLK(clk_bF$buf3),
    .D(_32_),
    .Q(Atmp[5])
);

DFFPOSX1 _659_ (
    .CLK(clk_bF$buf2),
    .D(_33_),
    .Q(Atmp[6])
);

DFFPOSX1 _660_ (
    .CLK(clk_bF$buf1),
    .D(_34_),
    .Q(Atmp[7])
);

DFFPOSX1 _661_ (
    .CLK(clk_bF$buf0),
    .D(_35_),
    .Q(Atmp[8])
);

DFFPOSX1 _662_ (
    .CLK(clk_bF$buf5),
    .D(_36_),
    .Q(Atmp[9])
);

DFFPOSX1 _663_ (
    .CLK(clk_bF$buf4),
    .D(_37_),
    .Q(Atmp[11])
);

DFFPOSX1 _664_ (
    .CLK(clk_bF$buf3),
    .D(_38_),
    .Q(_312_)
);

BUFX2 _665_ (
    .A(_311_[0]),
    .Y(Aout[0])
);

BUFX2 _666_ (
    .A(_311_[1]),
    .Y(Aout[1])
);

BUFX2 _667_ (
    .A(_312_),
    .Y(ISout)
);

BUFX2 _668_ (
    .A(RdyCtl_6_bF$buf3),
    .Y(Vld)
);

endmodule
