magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -140 -1950 2540 5180
<< metal2 >>
rect 100 5032 164 5060
use DOUBLE_GUARD$2  DOUBLE_GUARD$2_0
timestamp 1569533753
transform 1 0 0 0 1 1660
box -20 -20 2419 500
use GUARD$2  GUARD$2_0
timestamp 1569533753
transform 1 0 0 0 1 4220
box -20 -20 2419 792
use GUARD1$1  GUARD1$1_0
timestamp 1569533753
transform 1 0 1193 0 1 4220
box -484 36 1167 756
use INV2$2  INV2$2_0
timestamp 1569533753
transform 1 0 114 0 1 4314
box -2 -42 426 646
use METAL_RING$2  METAL_RING$2_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 5012
use NDRV$2  NDRV$2_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 1560
use PAD_80$2  PAD_80$2_0
timestamp 1569533753
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_POB8$1  PAD_METAL_POB8$1_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 5060
use PDRV$2  PDRV$2_0
timestamp 1569533753
transform 1 0 0 0 1 2260
box -20 -20 2420 1580
use SINGLE_GUARD$2  SINGLE_GUARD$2_0
timestamp 1569533753
transform 1 0 0 0 1 3920
box 0 0 2400 200
<< labels >>
flabel m2p s 135 5060 135 5060 0 FreeSans 400 0 0 0 A
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 PAD
flabel m3p s 0 3018 0 3018 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4339 0 4339 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4788 0 4788 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 752 0 752 0 FreeSans 1000 0 0 0 VSS
<< end >>
