/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module phase_accumulator(
    inout vdd,
    inout gnd,
    output [1:0] Aout,
    input En,
    input [19:0] FCW,
    output ISout,
    output Vld,
    input clk
);

wire _168_ ;
wire _60_ ;
wire _19_ ;
wire _57_ ;
wire _130_ ;
wire _95_ ;
wire _224_ ;
wire _262_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _92_ ;
wire _221_ ;
wire _124_ ;
wire _89_ ;
wire _162_ ;
wire _73__bF$buf0 ;
wire _73__bF$buf1 ;
wire _73__bF$buf2 ;
wire _73__bF$buf3 ;
wire _73__bF$buf4 ;
wire _218_ ;
wire _256_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _197_ ;
wire _7_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire ISout ;
wire _86_ ;
wire _215_ ;
wire _253_ ;
wire [11:0] Atmp ;
wire _309_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _156_ ;
wire _194_ ;
wire _288_ ;
wire _4_ ;
wire _45_ ;
wire _83_ ;
wire [19:0] acc_reg ;
wire _212_ ;
wire _250_ ;
wire _306_ ;
wire En_bF$buf0 ;
wire En_bF$buf1 ;
wire En_bF$buf2 ;
wire En_bF$buf3 ;
wire En_bF$buf4 ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _191_ ;
wire _247_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _188_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _112_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _244_ ;
wire _109_ ;
wire _282_ ;
wire _147_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _241_ ;
wire _106_ ;
wire _144_ ;
wire _182_ ;
wire _238_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _103_ ;
wire _68_ ;
wire _141_ ;
wire _235_ ;
wire _273_ ;
wire _138_ ;
wire _30_ ;
wire En ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _232_ ;
wire _270_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _267_ ;
wire _24_ ;
wire _62_ ;
wire _59_ ;
wire _132_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _264_ ;
wire _129_ ;
wire _21_ ;
wire _167_ ;
wire _299_ ;
wire _18_ ;
wire _56_ ;
wire _94_ ;
wire _223_ ;
wire _261_ ;
wire _126_ ;
wire _164_ ;
wire _258_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _123_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _255_ ;
wire _293_ ;
wire _12_ ;
wire _158_ ;
wire _50_ ;
wire _196_ ;
wire _6_ ;
wire [1:0] _311_ ;
wire _47_ ;
wire _120_ ;
wire _85_ ;
wire _214_ ;
wire _252_ ;
wire _308_ ;
wire _117_ ;
wire _290_ ;
wire _155_ ;
wire [1:0] Aout ;
wire _193_ ;
wire _249_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _82_ ;
wire _211_ ;
wire _305_ ;
wire _114_ ;
wire [19:0] FCW ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _190_ ;
wire _246_ ;
wire _284_ ;
wire _0_ ;
wire _149_ ;
wire _41_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _111_ ;
wire _76_ ;
wire _205_ ;
wire _243_ ;
wire _108_ ;
wire RdyCtl_6_bF$buf0 ;
wire RdyCtl_6_bF$buf1 ;
wire RdyCtl_6_bF$buf2 ;
wire RdyCtl_6_bF$buf3 ;
wire RdyCtl_6_bF$buf4 ;
wire _281_ ;
wire _146_ ;
wire _184_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _181_ ;
wire _237_ ;
wire _275_ ;
wire _32_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _102_ ;
wire _67_ ;
wire _140_ ;
wire _234_ ;
wire _272_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _231_ ;
wire _134_ ;
wire _99_ ;
wire _172_ ;
wire Vld ;
wire _228_ ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _58_ ;
wire _131_ ;
wire [6:0] RdyCtl ;
wire _96_ ;
wire _225_ ;
wire _263_ ;
wire _128_ ;
wire _20_ ;
wire _166_ ;
wire _298_ ;
wire _17_ ;
wire _55_ ;
wire _93_ ;
wire _222_ ;
wire _260_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _257_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _198_ ;
wire _90_ ;
wire _8_ ;
wire _49_ ;
wire _122_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _254_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _157_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _310_ ;
wire _46_ ;
wire _84_ ;
wire _213_ ;
wire _251_ ;
wire _307_ ;
wire _116_ ;
wire _154_ ;
wire _192_ ;
wire _248_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _245_ ;
wire _283_ ;
wire _148_ ;
wire _40_ ;
wire _186_ ;
wire _301_ ;
wire _37_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _242_ ;
wire _107_ ;
wire _280_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _104_ ;
wire _69_ ;
wire _142_ ;
wire _180_ ;
wire _236_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _177_ ;
wire _28_ ;
wire _101_ ;
wire _66_ ;
wire _233_ ;
wire _271_ ;
wire _136_ ;
wire _174_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _230_ ;
wire _133_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _265_ ;
wire _22_ ;

FILL FILL_2__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_118_)
);

FILL FILL_1__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .Y(_230_)
);

FILL FILL_5__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[9]),
    .Y(_56_)
);

FILL FILL_4__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_156_),
    .Y(_161_)
);

FILL FILL76050x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_83_),
    .Y(_84_)
);

FILL FILL_5__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

FILL FILL_4__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_245_),
    .Y(_247_)
);

FILL FILL_4__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _644_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[11])
);

FILL FILL_4__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_277_),
    .C(_282_),
    .Y(_283_)
);

FILL FILL_4__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[0]),
    .B(RdyCtl[0]),
    .Y(_54_)
);

FILL FILL_4__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_158_)
);

FILL FILL_1__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[11]),
    .B(RdyCtl_6_bF$buf2),
    .Y(_309_)
);

FILL FILL_5__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_81_)
);

FILL FILL_1__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_191_),
    .C(_73__bF$buf2),
    .Y(_193_)
);

FILL FILL_1__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(RdyCtl_6_bF$buf4),
    .C(_115_),
    .Y(_11_)
);

FILL FILL_2__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(RdyCtl_6_bF$buf1),
    .C(_227_),
    .Y(_21_)
);

FILL FILL_5__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_73__bF$buf3),
    .C(_307_),
    .Y(_35_)
);

FILL FILL_3__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_131_),
    .Y(_132_)
);

FILL FILL_4__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_217_),
    .Y(_244_)
);

FILL FILL_4__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _641_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[8])
);

FILL FILL_5__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .Y(_280_)
);

FILL FILL_5__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[2]),
    .Y(_51_)
);

FILL FILL_4__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_149_),
    .C(_154_),
    .Y(_155_)
);

FILL FILL_7__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[0]),
    .B(FCW[0]),
    .Y(_78_)
);

FILL FILL_4__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_188_),
    .Y(_190_)
);

FILL FILL_5__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_240_),
    .Y(_241_)
);

FILL FILL_1__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_111_),
    .Y(_113_)
);

FILL FILL_2__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _638_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[5])
);

FILL FILL_1__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_222_),
    .C(_220_),
    .Y(_225_)
);

FILL FILL_5__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[18]),
    .B(FCW[18]),
    .Y(_277_)
);

FILL FILL_4__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[15]),
    .B(_73__bF$buf0),
    .C(En_bF$buf3),
    .Y(_306_)
);

FILL FILL_5__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_109_),
    .C(_107_),
    .Y(_110_)
);

FILL FILL_1__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_222_)
);

FILL FILL_1__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_129_)
);

FILL FILL_8__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_42_),
    .C(_47_),
    .Y(_48_)
);

FILL FILL_4__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[0]),
    .B(RdyCtl_6_bF$buf1),
    .Y(_76_)
);

FILL FILL_5__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_182_),
    .Y(_187_)
);

FILL FILL75450x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_237_),
    .C(_238_),
    .Y(_22_)
);

FILL FILL_1__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _635_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[2])
);

FILL FILL_4__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_261_),
    .C(_273_),
    .Y(_274_)
);

FILL FILL_4__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_73__bF$buf4),
    .C(_304_),
    .Y(_32_)
);

FILL FILL_5__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(En_bF$buf3),
    .B(_44_),
    .Y(_5_)
);

FILL FILL_1__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[10]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_185_)
);

FILL FILL_1__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_106_),
    .Y(_107_)
);

FILL FILL_1__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_218_),
    .C(_211_),
    .Y(_219_)
);

FILL FILL_2__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[12]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_303_)
);

FILL FILL_2__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[11]),
    .B(_44_),
    .Y(_45_)
);

FILL FILL_7__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_235_),
    .Y(_236_)
);

FILL FILL_4__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _632_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[6])
);

FILL FILL_4__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_270_),
    .C(_271_),
    .Y(_24_)
);

FILL FILL_5__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[1]),
    .B(En_bF$buf4),
    .Y(_2_)
);

FILL FILL_4__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_178_),
    .Y(_182_)
);

FILL FILL_8__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_91_),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_5__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _629_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[3])
);

FILL FILL_1__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_215_),
    .C(_216_),
    .Y(_20_)
);

FILL FILL_2__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_268_),
    .Y(_269_)
);

FILL FILL_4__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .Y(ISout)
);

FILL FILL_1__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .B(_73__bF$buf1),
    .C(_301_),
    .Y(_29_)
);

FILL FILL_5__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_213_),
    .Y(_214_)
);

FILL FILL_1__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_232_),
    .C(_224_),
    .Y(_233_)
);

FILL FILL_7__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(En_bF$buf1),
    .Y(_74_)
);

FILL FILL_4__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_179_)
);

FILL FILL_1__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_5__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _626_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[0])
);

FILL FILL_1__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_266_)
);

FILL FILL_4__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _664_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .CLK(clk_bF$buf2),
    .Q(_312_)
);

FILL FILL73050x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[9]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_300_)
);

FILL FILL_5__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_66_),
    .Y(_72_)
);

FILL FILL_1__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .Y(_176_)
);

FILL FILL_1__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_97_),
    .Y(_99_)
);

FILL FILL_1__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_211_)
);

FILL FILL_1__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .B(_149_),
    .Y(_150_)
);

FILL FILL_4__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[16]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_264_)
);

FILL FILL_4__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _661_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .CLK(clk_bF$buf3),
    .Q(Atmp[8])
);

FILL FILL_5__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[8]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_298_)
);

FILL FILL_5__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[19]),
    .Y(_69_)
);

FILL FILL_4__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_170_),
    .C(_173_),
    .Y(_16_)
);

FILL FILL_8__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[3]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_96_)
);

FILL FILL75750x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_195_),
    .C(_74_),
    .Y(_19_)
);

FILL FILL_2__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_258_),
    .C(_260_),
    .Y(_261_)
);

FILL FILL_4__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _658_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[5])
);

FILL FILL_1__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_295_),
    .C(_73__bF$buf2),
    .Y(_296_)
);

FILL FILL_4__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_127_),
    .C(_126_),
    .Y(_128_)
);

FILL FILL_1__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_147_)
);

FILL FILL_1__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[5]),
    .Y(_66_)
);

FILL FILL_4__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_164_),
    .Y(_171_)
);

FILL FILL_8__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_91_),
    .C(_93_),
    .Y(_94_)
);

FILL FILL_5__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_143_),
    .C(_144_),
    .Y(_14_)
);

FILL FILL_1__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

FILL FILL_5__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_240_),
    .Y(_258_)
);

FILL FILL_4__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _655_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .CLK(clk_bF$buf4),
    .Q(Atmp[2])
);

FILL FILL_4__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_289_),
    .Y(_293_)
);

FILL FILL_4__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_167_),
    .Y(_168_)
);

FILL FILL_1__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_90_),
    .B(_89_),
    .Y(_91_)
);

FILL FILL_1__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_203_)
);

FILL FILL_1__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .Y(_125_)
);

FILL FILL_1__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf1)
);

FILL FILL_1__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[4]),
    .Y(_44_)
);

FILL FILL_2__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[1]),
    .B(_61_),
    .C(_63_),
    .Y(_64_)
);

FILL FILL_7__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_141_),
    .Y(_142_)
);

FILL FILL_4__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_127_),
    .Y(_255_)
);

FILL FILL_4__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _652_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[19])
);

FILL FILL_4__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_290_)
);

FILL FILL_5__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_55_),
    .C(_60_),
    .Y(_61_)
);

FILL FILL_4__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_165_)
);

FILL FILL_1__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_81_),
    .C(_79_),
    .Y(_88_)
);

FILL FILL_4__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_179_),
    .C(_188_),
    .Y(_200_)
);

FILL FILL_2__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[5]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_123_)
);

FILL FILL_2__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _649_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf5),
    .Q(acc_reg[16])
);

FILL FILL_1__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[19]),
    .B(En_bF$buf4),
    .Y(_287_)
);

FILL FILL_4__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[6]),
    .Y(_41_)
);

FILL FILL_2__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_230_),
    .Y(_232_)
);

FILL FILL_2__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_139_)
);

FILL FILL_2__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_250_),
    .Y(_252_)
);

FILL FILL_7__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[7]),
    .Y(_58_)
);

FILL FILL_4__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[8]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_163_)
);

FILL FILL75150x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_85_),
    .Y(_86_)
);

FILL FILL_4__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[6]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_137_)
);

FILL FILL_4__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_190_),
    .C(_196_),
    .Y(_197_)
);

FILL FILL_5__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_241_),
    .C(_248_),
    .Y(_249_)
);

FILL FILL_1__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_116_),
    .Y(_120_)
);

FILL FILL_5__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _646_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[13])
);

FILL FILL_1__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[18]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf4),
    .Y(_285_)
);

FILL FILL76050x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_310_),
    .Y(_37_)
);

FILL FILL_5__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_81_),
    .Y(_83_)
);

FILL FILL_1__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_193_),
    .C(_194_),
    .Y(_18_)
);

FILL FILL_1__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[5]),
    .B(FCW[5]),
    .Y(_117_)
);

FILL FILL74850x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_229_)
);

FILL FILL_5__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[5]),
    .Y(_55_)
);

FILL FILL_7__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_159_),
    .Y(_160_)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_73__bF$buf0)
);

FILL FILL_7__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .Y(_134_)
);

FILL FILL_4__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_221_),
    .C(_230_),
    .Y(_246_)
);

FILL FILL_4__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _643_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[10])
);

FILL FILL_4__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

FILL FILL_4__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[1]),
    .B(_50_),
    .C(_52_),
    .Y(_53_)
);

FILL FILL_4__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[8]),
    .B(FCW[8]),
    .Y(_157_)
);

FILL FILL_1__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_73__bF$buf3),
    .C(_308_),
    .Y(_36_)
);

FILL FILL_5__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .Y(_80_)
);

FILL FILL_1__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_191_),
    .Y(_192_)
);

FILL FILL_5__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[4]),
    .B(RdyCtl_6_bF$buf4),
    .C(En_bF$buf1),
    .Y(_115_)
);

FILL FILL_2__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[14]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf3),
    .Y(_227_)
);

FILL FILL_5__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_274_),
    .Y(_279_)
);

FILL FILL_4__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[16]),
    .B(_73__bF$buf3),
    .C(En_bF$buf1),
    .Y(_307_)
);

FILL FILL_5__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_130_),
    .Y(_131_)
);

FILL FILL_4__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_236_),
    .Y(_243_)
);

FILL FILL_7__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _640_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[7])
);

FILL FILL_5__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_40_),
    .C(_49_),
    .Y(_50_)
);

FILL FILL_4__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .Y(_154_)
);

FILL FILL_7__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_76_),
    .C(_77_),
    .Y(_7_)
);

FILL FILL_4__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_189_)
);

FILL FILL_5__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(_232_),
    .C(_217_),
    .Y(_240_)
);

FILL FILL_1__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_108_),
    .Y(_112_)
);

FILL FILL_5__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _637_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[4])
);

FILL FILL_1__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_223_),
    .Y(_224_)
);

FILL FILL_5__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_275_),
    .Y(_276_)
);

FILL FILL_4__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_73__bF$buf0),
    .C(_305_),
    .Y(_33_)
);

FILL FILL_5__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_186_)
);

FILL FILL_1__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_109_)
);

FILL FILL_1__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_221_)
);

FILL FILL_1__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_46_),
    .Y(_47_)
);

FILL FILL_4__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[0]),
    .Y(_75_)
);

FILL FILL_5__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[15]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf3),
    .Y(_238_)
);

FILL FILL_4__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _634_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[1])
);

FILL FILL_4__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_250_),
    .C(_266_),
    .Y(_273_)
);

FILL FILL_4__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[13]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_304_)
);

FILL FILL_5__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_74_),
    .Y(_4_)
);

FILL FILL75450x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(_183_),
    .Y(_184_)
);

FILL FILL_1__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_89_),
    .C(_97_),
    .Y(_106_)
);

FILL FILL_5__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_218_)
);

FILL FILL_2__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_73__bF$buf3),
    .C(_302_),
    .Y(_30_)
);

FILL FILL_3__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .Y(_235_)
);

FILL FILL_4__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _631_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf1),
    .Q(RdyCtl[5])
);

FILL FILL_2__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[17]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_271_)
);

FILL FILL_5__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[0]),
    .B(En_bF$buf2),
    .Y(_1_)
);

FILL FILL_4__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_179_),
    .Y(_181_)
);

FILL FILL74250x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(RdyCtl_6_bF$buf4),
    .C(_96_),
    .Y(_10_)
);

FILL FILL_5__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _628_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[2])
);

FILL FILL_1__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[13]),
    .B(RdyCtl_6_bF$buf2),
    .C(En_bF$buf4),
    .Y(_216_)
);

FILL FILL_5__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_266_),
    .Y(_268_)
);

FILL FILL_4__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_[1]),
    .Y(Aout[1])
);

FILL FILL_1__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[10]),
    .B(_73__bF$buf2),
    .C(En_bF$buf2),
    .Y(_301_)
);

FILL FILL_5__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_92_),
    .Y(_101_)
);

FILL FILL_1__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_212_),
    .Y(_213_)
);

FILL FILL_1__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl_6_bF$buf0),
    .Y(_73_)
);

FILL FILL_1__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_156_),
    .C(_176_),
    .Y(_178_)
);

FILL FILL_1__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_108_),
    .C(_117_),
    .Y(_152_)
);

FILL FILL_4__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_252_),
    .C(_250_),
    .Y(_265_)
);

FILL FILL_4__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _663_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[11])
);

FILL FILL_4__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[1]),
    .B(RdyCtl_6_bF$buf0),
    .Y(_299_)
);

FILL FILL_5__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .B(_70_),
    .Y(_71_)
);

FILL FILL_4__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_174_),
    .C(_165_),
    .Y(_175_)
);

FILL FILL73950x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_98_)
);

FILL FILL_1__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_209_),
    .C(_203_),
    .Y(_210_)
);

FILL FILL_2__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[0]),
    .B(RdyCtl_6_bF$buf0),
    .Y(_297_)
);

FILL FILL_4__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_130_),
    .C(_148_),
    .Y(_149_)
);

FILL FILL_4__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .B(_253_),
    .Y(_263_)
);

FILL FILL_1__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _660_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .CLK(clk_bF$buf1),
    .Q(Atmp[7])
);

FILL FILL_5__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[18]),
    .Y(_68_)
);

FILL FILL_4__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[9]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_173_)
);

FILL FILL_6__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_95_),
    .C(_74_),
    .Y(_9_)
);

FILL FILL_4__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_146_)
);

FILL FILL_1__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_207_),
    .C(RdyCtl_6_bF$buf2),
    .Y(_208_)
);

FILL FILL_2__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_201_),
    .C(_259_),
    .Y(_260_)
);

FILL FILL_4__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _657_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .CLK(clk_bF$buf2),
    .Q(Atmp[4])
);

FILL FILL_1__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .Y(_295_)
);

FILL FILL_2_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_204_),
    .Y(_205_)
);

FILL FILL_1__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_119_),
    .Y(_127_)
);

FILL FILL_1__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[0]),
    .B(_64_),
    .C(_65_),
    .Y(_311_[1])
);

FILL FILL_4__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_164_),
    .Y(_170_)
);

FILL FILL_1__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73__bF$buf0),
    .B(_92_),
    .Y(_93_)
);

FILL FILL_5__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[7]),
    .B(RdyCtl_6_bF$buf0),
    .C(En_bF$buf0),
    .Y(_144_)
);

FILL FILL_1__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_107_),
    .C(_256_),
    .Y(_257_)
);

FILL FILL_4__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _654_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .CLK(clk_bF$buf4),
    .Q(Atmp[1])
);

FILL FILL_4__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_291_),
    .Y(_292_)
);

FILL FILL_4__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[1]),
    .B(_62_),
    .Y(_63_)
);

FILL FILL_4__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[9]),
    .Y(_167_)
);

FILL FILL_1__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_90_)
);

FILL FILL_1__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_156_),
    .C(_201_),
    .Y(_202_)
);

FILL FILL_1__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_124_)
);

FILL FILL_2__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[8]),
    .Y(_43_)
);

FILL FILL_2__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_140_),
    .Y(_141_)
);

FILL FILL_4__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_131_),
    .Y(_254_)
);

FILL FILL_4__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _651_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[18])
);

FILL FILL_5__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_282_),
    .C(_288_),
    .Y(_289_)
);

FILL FILL_5__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[3]),
    .B(_57_),
    .C(_59_),
    .Y(_60_)
);

FILL FILL_4__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_156_),
    .C(_157_),
    .Y(_164_)
);

FILL FILL_4_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(RdyCtl_6_bF$buf1),
    .C(_87_),
    .Y(_8_)
);

FILL FILL_4__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .Y(_199_)
);

FILL FILL_2__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_251_)
);

FILL FILL_1__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73__bF$buf3),
    .B(_121_),
    .Y(_122_)
);

FILL FILL_2__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _648_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[15])
);

FILL FILL_1__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_286_)
);

FILL FILL_4__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[2]),
    .Y(_40_)
);

FILL FILL_2__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_117_),
    .Y(_119_)
);

FILL FILL_1__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[15]),
    .B(FCW[15]),
    .Y(_231_)
);

FILL FILL_3__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .B(_128_),
    .C(_129_),
    .Y(_138_)
);

FILL FILL_8__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_56_),
    .C(_45_),
    .Y(_57_)
);

FILL FILL_4__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_160_),
    .Y(_162_)
);

FILL FILL_7__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .Y(_85_)
);

FILL FILL_5__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_132_),
    .Y(_136_)
);

FILL FILL_4__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_169_),
    .Y(_196_)
);

FILL FILL_5__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_242_),
    .C(_247_),
    .Y(_248_)
);

FILL FILL_1__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _645_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf2),
    .Q(acc_reg[12])
);

FILL FILL_4__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_283_),
    .Y(_284_)
);

FILL FILL_4__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_158_),
    .Y(_159_)
);

FILL FILL_1__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[18]),
    .B(_73__bF$buf4),
    .C(En_bF$buf4),
    .Y(_310_)
);

FILL FILL_5__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_80_),
    .C(_78_),
    .Y(_82_)
);

FILL FILL_1__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[11]),
    .B(RdyCtl_6_bF$buf3),
    .C(En_bF$buf2),
    .Y(_194_)
);

FILL FILL_1__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_112_),
    .C(_108_),
    .Y(_116_)
);

FILL FILL_1__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[14]),
    .B(FCW[14]),
    .Y(_228_)
);

FILL FILL_5__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[17]),
    .B(_73__bF$buf3),
    .C(En_bF$buf2),
    .Y(_308_)
);

FILL FILL_2__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[0]),
    .B(_53_),
    .C(_54_),
    .Y(_311_[0])
);

FILL FILL_7__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[6]),
    .Y(RdyCtl_6_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(En),
    .Y(En_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_73__bF$buf4)
);

FILL FILL_7__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_73__bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_73__bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_73__bF$buf1)
);

FILL FILL_1__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .Y(_133_)
);

FILL FILL_4__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_239_),
    .C(_232_),
    .Y(_245_)
);

FILL FILL_4__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _642_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf4),
    .Q(acc_reg[9])
);

FILL FILL_4__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .Y(_281_)
);

FILL FILL_5__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[1]),
    .B(_51_),
    .Y(_52_)
);

FILL FILL_4__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_111_),
    .C(_155_),
    .Y(_156_)
);

FILL FILL_1__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[1]),
    .B(FCW[1]),
    .Y(_79_)
);

FILL FILL_4__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73650x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .Y(_191_)
);

FILL FILL_5__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_110_),
    .Y(_114_)
);

FILL FILL_2__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _639_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[6])
);

FILL FILL_1__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_224_),
    .Y(_226_)
);

FILL FILL_5__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_276_),
    .Y(_278_)
);

FILL FILL_4__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_73__bF$buf0),
    .C(_306_),
    .Y(_34_)
);

FILL FILL_5__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_222_),
    .Y(_223_)
);

FILL FILL_1__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__466_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[6]),
    .B(FCW[6]),
    .Y(_130_)
);

FILL FILL_2__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_198_),
    .Y(_242_)
);

FILL FILL_7__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_48_),
    .Y(_49_)
);

FILL FILL_4__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__598_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_147_),
    .C(_139_),
    .Y(_153_)
);

FILL FILL_7__385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_76_),
    .C(En_bF$buf3),
    .Y(_77_)
);

FILL FILL_4__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[11]),
    .B(FCW[11]),
    .Y(_188_)
);

FILL FILL_5__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_221_),
    .Y(_239_)
);

FILL FILL_1__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__479_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .B(_104_),
    .Y(_111_)
);

FILL FILL_5__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _636_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf3),
    .Q(acc_reg[3])
);

FILL FILL_1__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(FCW[18]),
    .Y(_275_)
);

FILL FILL_4__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[14]),
    .B(_73__bF$buf0),
    .C(En_bF$buf3),
    .Y(_305_)
);

FILL FILL74850x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_74_),
    .Y(_6_)
);

FILL FILL_1__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(RdyCtl_6_bF$buf3),
    .C(_185_),
    .Y(_17_)
);

FILL FILL_1__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[4]),
    .B(FCW[4]),
    .Y(_108_)
);

FILL FILL_1__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_217_),
    .C(_219_),
    .Y(_220_)
);

FILL FILL_1__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__366_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_44_),
    .C(_45_),
    .Y(_46_)
);

FILL FILL_7__573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_236_),
    .C(_73__bF$buf4),
    .Y(_237_)
);

FILL FILL_4__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__498_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _633_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[0])
);

FILL FILL_4__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_268_),
    .Y(_272_)
);

FILL FILL_4__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_73__bF$buf2),
    .C(_303_),
    .Y(_31_)
);

FILL FILL_5__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_74_),
    .Y(_3_)
);

FILL FILL_1__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_181_),
    .Y(_183_)
);

FILL FILL_8__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .Y(_105_)
);

FILL FILL_5__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_213_),
    .Y(_217_)
);

FILL FILL75150x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_268_),
    .C(_73__bF$buf2),
    .Y(_270_)
);

FILL FILL_4__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl_6_bF$buf1),
    .Y(Vld)
);

FILL FILL_1__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[11]),
    .B(_73__bF$buf1),
    .C(En_bF$buf0),
    .Y(_302_)
);

FILL FILL75450x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_220_),
    .C(_228_),
    .Y(_234_)
);

FILL FILL_7__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _630_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf3),
    .Q(RdyCtl[4])
);

FILL FILL_2__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73__bF$buf2),
    .B(_74_),
    .Y(_0_)
);

FILL FILL_4__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[10]),
    .B(FCW[10]),
    .Y(_180_)
);

FILL FILL_8__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_102_),
    .Y(_103_)
);

FILL FILL_5__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _627_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .CLK(clk_bF$buf5),
    .Q(RdyCtl[1])
);

FILL FILL_1__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_213_),
    .C(_73__bF$buf4),
    .Y(_215_)
);

FILL FILL_5__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[17]),
    .B(FCW[17]),
    .Y(_267_)
);

FILL FILL_4__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_[0]),
    .Y(Aout[0])
);

FILL FILL_4__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_300_),
    .Y(_28_)
);

FILL FILL_5__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_159_),
    .Y(_177_)
);

FILL FILL_1__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_92_),
    .C(_99_),
    .Y(_100_)
);

FILL FILL_1__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[13]),
    .B(FCW[13]),
    .Y(_212_)
);

FILL FILL_1__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__429_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_71_),
    .C(_72_),
    .Y(_38_)
);

FILL FILL_1__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74850x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__489_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .Y(_151_)
);

FILL FILL_4__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(RdyCtl_6_bF$buf3),
    .C(_264_),
    .Y(_23_)
);

FILL FILL_4__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _662_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .CLK(clk_bF$buf3),
    .Q(Atmp[9])
);

FILL FILL_4__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_298_),
    .Y(_27_)
);

FILL FILL_5__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_69_),
    .Y(_70_)
);

FILL FILL_4__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[9]),
    .B(FCW[9]),
    .Y(_174_)
);

FILL FILL_1__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[3]),
    .B(FCW[3]),
    .Y(_97_)
);

FILL FILL_4__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .Y(_209_)
);

FILL FILL_2__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__507_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _659_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .CLK(clk_bF$buf0),
    .Q(Atmp[6])
);

FILL FILL_1__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_287_),
    .C(_296_),
    .D(_293_),
    .Y(_26_)
);

FILL FILL_4__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75150x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__486_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_146_),
    .Y(_148_)
);

FILL FILL76050x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_251_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[18]),
    .B(acc_reg[19]),
    .Y(_67_)
);

FILL FILL_4__452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__508_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73__bF$buf1),
    .B(_171_),
    .Y(_172_)
);

FILL FILL_8__347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[2]),
    .B(_73__bF$buf0),
    .Y(_95_)
);

FILL FILL_4__490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_119_),
    .Y(_145_)
);

FILL FILL_1__402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__546_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_205_),
    .Y(_207_)
);

FILL FILL_5__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__568_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_246_),
    .Y(_259_)
);

FILL FILL_4__355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__377_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _656_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .CLK(clk_bF$buf5),
    .Q(Atmp[3])
);

FILL FILL_1__440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_278_),
    .C(_276_),
    .Y(_294_)
);

FILL FILL_4__393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_88_),
    .Y(_92_)
);

FILL FILL_1__343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[12]),
    .B(FCW[12]),
    .Y(_204_)
);

FILL FILL_1__572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_124_),
    .C(_125_),
    .Y(_126_)
);

FILL FILL75450x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73950x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[0]),
    .B(Atmp[1]),
    .Y(_65_)
);

FILL FILL_7__593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__505_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_168_),
    .Y(_169_)
);

FILL FILL_1__378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__336_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_141_),
    .C(_73__bF$buf1),
    .Y(_143_)
);

FILL FILL_4__543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__565_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_126_),
    .C(_153_),
    .Y(_256_)
);

FILL FILL_4__352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__408_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _653_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .CLK(clk_bF$buf5),
    .Q(Atmp[0])
);

FILL FILL_4__581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__488_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[19]),
    .B(FCW[19]),
    .Y(_291_)
);

FILL FILL_2_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[3]),
    .Y(_62_)
);

FILL FILL_4__446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73350x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__468_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[9]),
    .Y(_166_)
);

FILL FILL_1__531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[2]),
    .B(FCW[2]),
    .Y(_89_)
);

FILL FILL_1__340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_200_),
    .Y(_201_)
);

FILL FILL_2__603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__349_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_120_),
    .C(_123_),
    .Y(_12_)
);

FILL FILL_2__412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .Y(_288_)
);

FILL FILL_4__387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__528_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RdyCtl[3]),
    .Y(_42_)
);

FILL FILL_2__315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__608_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_7__361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL76050x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__477_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[7]),
    .B(FCW[7]),
    .Y(_140_)
);

FILL FILL_4__540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75750x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74550x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__562_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_249_),
    .Y(_253_)
);

FILL FILL74550x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__549_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _650_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf5),
    .Q(acc_reg[17])
);

FILL FILL_5__612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__512_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(RdyCtl[3]),
    .C(RdyCtl[2]),
    .Y(_59_)
);

FILL FILL_4__443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__465_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(RdyCtl_6_bF$buf3),
    .C(_163_),
    .Y(_15_)
);

FILL FILL_7__396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__550_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[1]),
    .B(RdyCtl_6_bF$buf1),
    .C(En_bF$buf3),
    .Y(_87_)
);

FILL FILL_4__481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL75450x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__606_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(RdyCtl_6_bF$buf4),
    .C(_137_),
    .Y(_13_)
);

FILL FILL_4__537_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_181_),
    .C(_190_),
    .Y(_198_)
);

FILL FILL_2__600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__559_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[16]),
    .B(FCW[16]),
    .Y(_250_)
);

FILL FILL_1__622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_116_),
    .Y(_121_)
);

FILL FILL_5__553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__368_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _647_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf0),
    .Q(acc_reg[14])
);

FILL FILL74850x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__597_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(RdyCtl_6_bF$buf2),
    .C(_285_),
    .Y(_25_)
);

FILL FILL_4__384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__525_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Atmp[4]),
    .Y(_39_)
);

FILL FILL_5__456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__356_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(acc_reg[12]),
    .B(_73__bF$buf4),
    .Y(_195_)
);

FILL FILL_1__563_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule
