magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -120 -120 5180 5180
<< metal1 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5030
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal2 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5031
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal3 >>
rect 0 2260 1560 5060
rect 2260 4220 3820 5060
rect 4220 4552 4552 5060
rect 4680 5012 5012 5060
tri 5012 5012 5060 5060 sw
rect 4680 4817 5060 5012
tri 4680 4680 4817 4817 ne
rect 4817 4680 5060 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5060 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5060 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5060 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5060 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5060 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5060 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5060 1560
use VIA1$3  VIA1$3_0
timestamp 1569533753
transform 1 0 4744 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_1
timestamp 1569533753
transform 1 0 4872 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_2
timestamp 1569533753
transform 1 0 4808 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_3
timestamp 1569533753
transform 1 0 4680 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_4
timestamp 1569533753
transform 1 0 4680 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_5
timestamp 1569533753
transform 1 0 4744 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_6
timestamp 1569533753
transform 1 0 4744 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_7
timestamp 1569533753
transform 1 0 4872 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_8
timestamp 1569533753
transform 1 0 4680 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_9
timestamp 1569533753
transform 1 0 4808 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_10
timestamp 1569533753
transform 1 0 4872 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_11
timestamp 1569533753
transform 1 0 4680 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_12
timestamp 1569533753
transform 1 0 4808 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_13
timestamp 1569533753
transform 1 0 4744 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_14
timestamp 1569533753
transform 1 0 4680 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_15
timestamp 1569533753
transform 1 0 4808 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_16
timestamp 1569533753
transform 1 0 4808 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_17
timestamp 1569533753
transform 1 0 4872 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_18
timestamp 1569533753
transform 1 0 4744 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_19
timestamp 1569533753
transform 1 0 4872 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_20
timestamp 1569533753
transform 1 0 4552 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_21
timestamp 1569533753
transform 1 0 4488 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_22
timestamp 1569533753
transform 1 0 4616 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_23
timestamp 1569533753
transform 1 0 4552 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_24
timestamp 1569533753
transform 1 0 4616 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_25
timestamp 1569533753
transform 1 0 4488 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_26
timestamp 1569533753
transform 1 0 4424 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_27
timestamp 1569533753
transform 1 0 4616 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_28
timestamp 1569533753
transform 1 0 4552 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_29
timestamp 1569533753
transform 1 0 4488 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_30
timestamp 1569533753
transform 1 0 4424 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_31
timestamp 1569533753
transform 1 0 4424 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_32
timestamp 1569533753
transform 1 0 4552 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_33
timestamp 1569533753
transform 1 0 4616 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_34
timestamp 1569533753
transform 1 0 4424 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_35
timestamp 1569533753
transform 1 0 4424 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_36
timestamp 1569533753
transform 1 0 4552 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_37
timestamp 1569533753
transform 1 0 4488 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_38
timestamp 1569533753
transform 1 0 4488 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_39
timestamp 1569533753
transform 1 0 4616 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_40
timestamp 1569533753
transform 1 0 4616 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_41
timestamp 1569533753
transform 1 0 4424 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_42
timestamp 1569533753
transform 1 0 4424 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_43
timestamp 1569533753
transform 1 0 4552 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_44
timestamp 1569533753
transform 1 0 4488 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_45
timestamp 1569533753
transform 1 0 4488 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_46
timestamp 1569533753
transform 1 0 4552 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_47
timestamp 1569533753
transform 1 0 4424 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_48
timestamp 1569533753
transform 1 0 4552 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_49
timestamp 1569533753
transform 1 0 4616 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_50
timestamp 1569533753
transform 1 0 4552 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_51
timestamp 1569533753
transform 1 0 4616 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_52
timestamp 1569533753
transform 1 0 4616 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_53
timestamp 1569533753
transform 1 0 4488 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_54
timestamp 1569533753
transform 1 0 4488 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_55
timestamp 1569533753
transform 1 0 4424 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_56
timestamp 1569533753
transform 1 0 4872 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_57
timestamp 1569533753
transform 1 0 4680 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_58
timestamp 1569533753
transform 1 0 4808 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_59
timestamp 1569533753
transform 1 0 4872 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_60
timestamp 1569533753
transform 1 0 4808 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_61
timestamp 1569533753
transform 1 0 4744 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_62
timestamp 1569533753
transform 1 0 4744 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_63
timestamp 1569533753
transform 1 0 4808 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_64
timestamp 1569533753
transform 1 0 4680 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_65
timestamp 1569533753
transform 1 0 4872 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_66
timestamp 1569533753
transform 1 0 4808 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_67
timestamp 1569533753
transform 1 0 4744 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_68
timestamp 1569533753
transform 1 0 4872 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_69
timestamp 1569533753
transform 1 0 4680 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_70
timestamp 1569533753
transform 1 0 4680 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_71
timestamp 1569533753
transform 1 0 4744 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_72
timestamp 1569533753
transform 1 0 4232 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_73
timestamp 1569533753
transform 1 0 4168 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_74
timestamp 1569533753
transform 1 0 4168 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_75
timestamp 1569533753
transform 1 0 4296 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_76
timestamp 1569533753
transform 1 0 4296 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_77
timestamp 1569533753
transform 1 0 4296 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_78
timestamp 1569533753
transform 1 0 4232 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_79
timestamp 1569533753
transform 1 0 4104 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_80
timestamp 1569533753
transform 1 0 4168 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_81
timestamp 1569533753
transform 1 0 4168 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_82
timestamp 1569533753
transform 1 0 4232 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_83
timestamp 1569533753
transform 1 0 4104 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_84
timestamp 1569533753
transform 1 0 4104 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_85
timestamp 1569533753
transform 1 0 4104 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_86
timestamp 1569533753
transform 1 0 4232 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_87
timestamp 1569533753
transform 1 0 4232 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_88
timestamp 1569533753
transform 1 0 4104 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_89
timestamp 1569533753
transform 1 0 4296 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_90
timestamp 1569533753
transform 1 0 4296 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_91
timestamp 1569533753
transform 1 0 4168 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_92
timestamp 1569533753
transform 1 0 3784 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_93
timestamp 1569533753
transform 1 0 3848 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_94
timestamp 1569533753
transform 1 0 3912 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_95
timestamp 1569533753
transform 1 0 4040 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_96
timestamp 1569533753
transform 1 0 4040 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_97
timestamp 1569533753
transform 1 0 3912 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_98
timestamp 1569533753
transform 1 0 3848 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_99
timestamp 1569533753
transform 1 0 3976 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_100
timestamp 1569533753
transform 1 0 3784 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_101
timestamp 1569533753
transform 1 0 3912 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_102
timestamp 1569533753
transform 1 0 4040 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_103
timestamp 1569533753
transform 1 0 3976 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_104
timestamp 1569533753
transform 1 0 4040 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_105
timestamp 1569533753
transform 1 0 3848 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_106
timestamp 1569533753
transform 1 0 3848 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_107
timestamp 1569533753
transform 1 0 3912 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_108
timestamp 1569533753
transform 1 0 4040 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_109
timestamp 1569533753
transform 1 0 3976 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_110
timestamp 1569533753
transform 1 0 3912 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_111
timestamp 1569533753
transform 1 0 3784 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_112
timestamp 1569533753
transform 1 0 3848 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_113
timestamp 1569533753
transform 1 0 3784 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_114
timestamp 1569533753
transform 1 0 3784 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_115
timestamp 1569533753
transform 1 0 3976 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_116
timestamp 1569533753
transform 1 0 3976 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_117
timestamp 1569533753
transform 1 0 3784 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_118
timestamp 1569533753
transform 1 0 3912 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_119
timestamp 1569533753
transform 1 0 3976 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_120
timestamp 1569533753
transform 1 0 3848 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_121
timestamp 1569533753
transform 1 0 4040 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_122
timestamp 1569533753
transform 1 0 3912 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_123
timestamp 1569533753
transform 1 0 4040 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_124
timestamp 1569533753
transform 1 0 3976 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_125
timestamp 1569533753
transform 1 0 3976 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_126
timestamp 1569533753
transform 1 0 3912 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_127
timestamp 1569533753
transform 1 0 3976 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_128
timestamp 1569533753
transform 1 0 3848 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_129
timestamp 1569533753
transform 1 0 3784 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_130
timestamp 1569533753
transform 1 0 4040 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_131
timestamp 1569533753
transform 1 0 3912 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_132
timestamp 1569533753
transform 1 0 3784 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_133
timestamp 1569533753
transform 1 0 3848 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_134
timestamp 1569533753
transform 1 0 4040 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_135
timestamp 1569533753
transform 1 0 3848 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_136
timestamp 1569533753
transform 1 0 3784 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_137
timestamp 1569533753
transform 1 0 4104 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_138
timestamp 1569533753
transform 1 0 4296 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_139
timestamp 1569533753
transform 1 0 4168 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_140
timestamp 1569533753
transform 1 0 4168 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_141
timestamp 1569533753
transform 1 0 4104 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_142
timestamp 1569533753
transform 1 0 4104 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_143
timestamp 1569533753
transform 1 0 4232 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_144
timestamp 1569533753
transform 1 0 4232 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_145
timestamp 1569533753
transform 1 0 4232 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_146
timestamp 1569533753
transform 1 0 4168 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_147
timestamp 1569533753
transform 1 0 4168 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_148
timestamp 1569533753
transform 1 0 4232 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_149
timestamp 1569533753
transform 1 0 4104 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_150
timestamp 1569533753
transform 1 0 4296 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_151
timestamp 1569533753
transform 1 0 4296 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_152
timestamp 1569533753
transform 1 0 4296 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_153
timestamp 1569533753
transform 1 0 4232 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_154
timestamp 1569533753
transform 1 0 4104 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_155
timestamp 1569533753
transform 1 0 4232 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_156
timestamp 1569533753
transform 1 0 4168 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_157
timestamp 1569533753
transform 1 0 4168 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_158
timestamp 1569533753
transform 1 0 4168 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_159
timestamp 1569533753
transform 1 0 4168 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_160
timestamp 1569533753
transform 1 0 4232 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_161
timestamp 1569533753
transform 1 0 4104 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_162
timestamp 1569533753
transform 1 0 4296 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_163
timestamp 1569533753
transform 1 0 4296 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_164
timestamp 1569533753
transform 1 0 4232 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_165
timestamp 1569533753
transform 1 0 4296 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_166
timestamp 1569533753
transform 1 0 4104 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_167
timestamp 1569533753
transform 1 0 4296 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_168
timestamp 1569533753
transform 1 0 4104 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_169
timestamp 1569533753
transform 1 0 3976 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_170
timestamp 1569533753
transform 1 0 3976 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_171
timestamp 1569533753
transform 1 0 3912 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_172
timestamp 1569533753
transform 1 0 4040 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_173
timestamp 1569533753
transform 1 0 3848 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_174
timestamp 1569533753
transform 1 0 3848 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_175
timestamp 1569533753
transform 1 0 3784 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_176
timestamp 1569533753
transform 1 0 3784 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_177
timestamp 1569533753
transform 1 0 3912 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_178
timestamp 1569533753
transform 1 0 3848 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_179
timestamp 1569533753
transform 1 0 4040 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_180
timestamp 1569533753
transform 1 0 3784 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_181
timestamp 1569533753
transform 1 0 3912 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_182
timestamp 1569533753
transform 1 0 3976 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_183
timestamp 1569533753
transform 1 0 3912 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_184
timestamp 1569533753
transform 1 0 3976 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_185
timestamp 1569533753
transform 1 0 4040 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_186
timestamp 1569533753
transform 1 0 3784 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_187
timestamp 1569533753
transform 1 0 4040 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_188
timestamp 1569533753
transform 1 0 3848 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_189
timestamp 1569533753
transform 1 0 3848 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_190
timestamp 1569533753
transform 1 0 4040 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_191
timestamp 1569533753
transform 1 0 3848 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_192
timestamp 1569533753
transform 1 0 3784 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_193
timestamp 1569533753
transform 1 0 4040 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_194
timestamp 1569533753
transform 1 0 4040 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_195
timestamp 1569533753
transform 1 0 3848 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_196
timestamp 1569533753
transform 1 0 3976 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_197
timestamp 1569533753
transform 1 0 3848 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_198
timestamp 1569533753
transform 1 0 3976 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_199
timestamp 1569533753
transform 1 0 3784 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_200
timestamp 1569533753
transform 1 0 3976 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_201
timestamp 1569533753
transform 1 0 3912 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_202
timestamp 1569533753
transform 1 0 3784 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_203
timestamp 1569533753
transform 1 0 3912 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_204
timestamp 1569533753
transform 1 0 3784 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_205
timestamp 1569533753
transform 1 0 3912 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_206
timestamp 1569533753
transform 1 0 4040 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_207
timestamp 1569533753
transform 1 0 3976 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_208
timestamp 1569533753
transform 1 0 3912 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_209
timestamp 1569533753
transform 1 0 3784 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_210
timestamp 1569533753
transform 1 0 3848 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_211
timestamp 1569533753
transform 1 0 4040 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_212
timestamp 1569533753
transform 1 0 3976 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_213
timestamp 1569533753
transform 1 0 3912 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_214
timestamp 1569533753
transform 1 0 4104 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_215
timestamp 1569533753
transform 1 0 4104 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_216
timestamp 1569533753
transform 1 0 4296 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_217
timestamp 1569533753
transform 1 0 4104 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_218
timestamp 1569533753
transform 1 0 4104 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_219
timestamp 1569533753
transform 1 0 4104 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_220
timestamp 1569533753
transform 1 0 4296 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_221
timestamp 1569533753
transform 1 0 4296 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_222
timestamp 1569533753
transform 1 0 4168 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_223
timestamp 1569533753
transform 1 0 4296 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_224
timestamp 1569533753
transform 1 0 4168 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_225
timestamp 1569533753
transform 1 0 4168 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_226
timestamp 1569533753
transform 1 0 4168 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_227
timestamp 1569533753
transform 1 0 4168 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_228
timestamp 1569533753
transform 1 0 4296 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_229
timestamp 1569533753
transform 1 0 4232 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_230
timestamp 1569533753
transform 1 0 4232 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_231
timestamp 1569533753
transform 1 0 4232 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_232
timestamp 1569533753
transform 1 0 4232 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_233
timestamp 1569533753
transform 1 0 4232 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_234
timestamp 1569533753
transform 1 0 4680 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_235
timestamp 1569533753
transform 1 0 4744 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_236
timestamp 1569533753
transform 1 0 4808 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_237
timestamp 1569533753
transform 1 0 4808 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_238
timestamp 1569533753
transform 1 0 4808 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_239
timestamp 1569533753
transform 1 0 4744 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_240
timestamp 1569533753
transform 1 0 4872 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_241
timestamp 1569533753
transform 1 0 4680 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_242
timestamp 1569533753
transform 1 0 4744 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_243
timestamp 1569533753
transform 1 0 4744 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_244
timestamp 1569533753
transform 1 0 4872 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_245
timestamp 1569533753
transform 1 0 4808 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_246
timestamp 1569533753
transform 1 0 4680 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_247
timestamp 1569533753
transform 1 0 4872 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_248
timestamp 1569533753
transform 1 0 4872 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_249
timestamp 1569533753
transform 1 0 4680 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_250
timestamp 1569533753
transform 1 0 4616 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_251
timestamp 1569533753
transform 1 0 4488 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_252
timestamp 1569533753
transform 1 0 4552 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_253
timestamp 1569533753
transform 1 0 4424 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_254
timestamp 1569533753
transform 1 0 4424 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_255
timestamp 1569533753
transform 1 0 4424 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_256
timestamp 1569533753
transform 1 0 4488 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_257
timestamp 1569533753
transform 1 0 4616 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_258
timestamp 1569533753
transform 1 0 4616 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_259
timestamp 1569533753
transform 1 0 4552 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_260
timestamp 1569533753
transform 1 0 4616 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_261
timestamp 1569533753
transform 1 0 4488 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_262
timestamp 1569533753
transform 1 0 4552 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_263
timestamp 1569533753
transform 1 0 4424 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_264
timestamp 1569533753
transform 1 0 4552 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_265
timestamp 1569533753
transform 1 0 4488 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_266
timestamp 1569533753
transform 1 0 4488 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_267
timestamp 1569533753
transform 1 0 4488 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_268
timestamp 1569533753
transform 1 0 4488 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_269
timestamp 1569533753
transform 1 0 4552 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_270
timestamp 1569533753
transform 1 0 4424 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_271
timestamp 1569533753
transform 1 0 4424 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_272
timestamp 1569533753
transform 1 0 4616 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_273
timestamp 1569533753
transform 1 0 4424 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_274
timestamp 1569533753
transform 1 0 4488 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_275
timestamp 1569533753
transform 1 0 4616 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_276
timestamp 1569533753
transform 1 0 4488 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_277
timestamp 1569533753
transform 1 0 4424 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_278
timestamp 1569533753
transform 1 0 4616 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_279
timestamp 1569533753
transform 1 0 4552 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_280
timestamp 1569533753
transform 1 0 4552 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_281
timestamp 1569533753
transform 1 0 4552 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_282
timestamp 1569533753
transform 1 0 4424 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_283
timestamp 1569533753
transform 1 0 4552 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_284
timestamp 1569533753
transform 1 0 4616 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_285
timestamp 1569533753
transform 1 0 4616 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_286
timestamp 1569533753
transform 1 0 4680 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_287
timestamp 1569533753
transform 1 0 4680 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_288
timestamp 1569533753
transform 1 0 4680 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_289
timestamp 1569533753
transform 1 0 4680 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_290
timestamp 1569533753
transform 1 0 4744 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_291
timestamp 1569533753
transform 1 0 4744 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_292
timestamp 1569533753
transform 1 0 4744 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_293
timestamp 1569533753
transform 1 0 4744 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_294
timestamp 1569533753
transform 1 0 4744 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_295
timestamp 1569533753
transform 1 0 4808 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_296
timestamp 1569533753
transform 1 0 4808 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_297
timestamp 1569533753
transform 1 0 4808 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_298
timestamp 1569533753
transform 1 0 4808 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_299
timestamp 1569533753
transform 1 0 4808 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_300
timestamp 1569533753
transform 1 0 4872 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_301
timestamp 1569533753
transform 1 0 4872 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_302
timestamp 1569533753
transform 1 0 4872 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_303
timestamp 1569533753
transform 1 0 4872 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_304
timestamp 1569533753
transform 1 0 4872 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_305
timestamp 1569533753
transform 1 0 4680 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_306
timestamp 1569533753
transform 1 0 3976 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_307
timestamp 1569533753
transform 1 0 3784 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_308
timestamp 1569533753
transform 1 0 4424 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_309
timestamp 1569533753
transform 1 0 4616 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_310
timestamp 1569533753
transform 1 0 4360 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_311
timestamp 1569533753
transform 1 0 3848 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_312
timestamp 1569533753
transform 1 0 4488 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_313
timestamp 1569533753
transform 1 0 4104 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_314
timestamp 1569533753
transform 1 0 4744 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_315
timestamp 1569533753
transform 1 0 4360 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_316
timestamp 1569533753
transform 1 0 3912 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_317
timestamp 1569533753
transform 1 0 4552 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_318
timestamp 1569533753
transform 1 0 4232 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_319
timestamp 1569533753
transform 1 0 4872 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_320
timestamp 1569533753
transform 1 0 4360 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_321
timestamp 1569533753
transform 1 0 4040 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_322
timestamp 1569533753
transform 1 0 4680 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_323
timestamp 1569533753
transform 1 0 4360 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_324
timestamp 1569533753
transform 1 0 4296 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_325
timestamp 1569533753
transform 1 0 4360 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_326
timestamp 1569533753
transform 1 0 4360 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_327
timestamp 1569533753
transform 1 0 4360 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_328
timestamp 1569533753
transform 1 0 4360 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_329
timestamp 1569533753
transform 1 0 4360 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_330
timestamp 1569533753
transform 1 0 4360 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_331
timestamp 1569533753
transform 1 0 4360 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_332
timestamp 1569533753
transform 1 0 4360 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_333
timestamp 1569533753
transform 1 0 4360 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_334
timestamp 1569533753
transform 1 0 4360 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_335
timestamp 1569533753
transform 1 0 4360 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_336
timestamp 1569533753
transform 1 0 4168 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_337
timestamp 1569533753
transform 1 0 4360 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_338
timestamp 1569533753
transform 1 0 4360 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_339
timestamp 1569533753
transform 1 0 4808 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_340
timestamp 1569533753
transform 1 0 4360 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_341
timestamp 1569533753
transform 1 0 4360 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_342
timestamp 1569533753
transform 1 0 3592 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_343
timestamp 1569533753
transform 1 0 3656 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_344
timestamp 1569533753
transform 1 0 3592 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_345
timestamp 1569533753
transform 1 0 3592 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_346
timestamp 1569533753
transform 1 0 3464 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_347
timestamp 1569533753
transform 1 0 3592 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_348
timestamp 1569533753
transform 1 0 3656 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_349
timestamp 1569533753
transform 1 0 3720 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_350
timestamp 1569533753
transform 1 0 3656 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_351
timestamp 1569533753
transform 1 0 3720 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_352
timestamp 1569533753
transform 1 0 3720 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_353
timestamp 1569533753
transform 1 0 3656 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_354
timestamp 1569533753
transform 1 0 3592 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_355
timestamp 1569533753
transform 1 0 3528 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_356
timestamp 1569533753
transform 1 0 3528 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_357
timestamp 1569533753
transform 1 0 3464 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_358
timestamp 1569533753
transform 1 0 3720 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_359
timestamp 1569533753
transform 1 0 3528 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_360
timestamp 1569533753
transform 1 0 3464 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_361
timestamp 1569533753
transform 1 0 3464 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_362
timestamp 1569533753
transform 1 0 3528 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_363
timestamp 1569533753
transform 1 0 3656 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_364
timestamp 1569533753
transform 1 0 3720 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_365
timestamp 1569533753
transform 1 0 3464 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_366
timestamp 1569533753
transform 1 0 3528 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_367
timestamp 1569533753
transform 1 0 3400 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_368
timestamp 1569533753
transform 1 0 3336 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_369
timestamp 1569533753
transform 1 0 3336 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_370
timestamp 1569533753
transform 1 0 3272 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_371
timestamp 1569533753
transform 1 0 3400 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_372
timestamp 1569533753
transform 1 0 3400 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_373
timestamp 1569533753
transform 1 0 3144 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_374
timestamp 1569533753
transform 1 0 3144 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_375
timestamp 1569533753
transform 1 0 3272 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_376
timestamp 1569533753
transform 1 0 3336 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_377
timestamp 1569533753
transform 1 0 3144 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_378
timestamp 1569533753
transform 1 0 3144 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_379
timestamp 1569533753
transform 1 0 3144 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_380
timestamp 1569533753
transform 1 0 3272 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_381
timestamp 1569533753
transform 1 0 3272 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_382
timestamp 1569533753
transform 1 0 3400 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_383
timestamp 1569533753
transform 1 0 3208 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_384
timestamp 1569533753
transform 1 0 3336 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_385
timestamp 1569533753
transform 1 0 3208 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_386
timestamp 1569533753
transform 1 0 3208 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_387
timestamp 1569533753
transform 1 0 3336 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_388
timestamp 1569533753
transform 1 0 3400 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_389
timestamp 1569533753
transform 1 0 3208 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_390
timestamp 1569533753
transform 1 0 3208 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_391
timestamp 1569533753
transform 1 0 3272 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_392
timestamp 1569533753
transform 1 0 3336 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_393
timestamp 1569533753
transform 1 0 3272 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_394
timestamp 1569533753
transform 1 0 3272 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_395
timestamp 1569533753
transform 1 0 3208 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_396
timestamp 1569533753
transform 1 0 3272 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_397
timestamp 1569533753
transform 1 0 3336 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_398
timestamp 1569533753
transform 1 0 3144 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_399
timestamp 1569533753
transform 1 0 3208 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_400
timestamp 1569533753
transform 1 0 3208 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_401
timestamp 1569533753
transform 1 0 3400 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_402
timestamp 1569533753
transform 1 0 3208 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_403
timestamp 1569533753
transform 1 0 3272 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_404
timestamp 1569533753
transform 1 0 3400 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_405
timestamp 1569533753
transform 1 0 3144 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_406
timestamp 1569533753
transform 1 0 3144 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_407
timestamp 1569533753
transform 1 0 3336 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_408
timestamp 1569533753
transform 1 0 3400 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_409
timestamp 1569533753
transform 1 0 3336 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_410
timestamp 1569533753
transform 1 0 3400 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_411
timestamp 1569533753
transform 1 0 3144 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_412
timestamp 1569533753
transform 1 0 3656 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_413
timestamp 1569533753
transform 1 0 3720 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_414
timestamp 1569533753
transform 1 0 3656 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_415
timestamp 1569533753
transform 1 0 3656 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_416
timestamp 1569533753
transform 1 0 3656 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_417
timestamp 1569533753
transform 1 0 3464 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_418
timestamp 1569533753
transform 1 0 3464 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_419
timestamp 1569533753
transform 1 0 3528 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_420
timestamp 1569533753
transform 1 0 3592 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_421
timestamp 1569533753
transform 1 0 3528 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_422
timestamp 1569533753
transform 1 0 3464 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_423
timestamp 1569533753
transform 1 0 3592 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_424
timestamp 1569533753
transform 1 0 3528 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_425
timestamp 1569533753
transform 1 0 3528 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_426
timestamp 1569533753
transform 1 0 3592 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_427
timestamp 1569533753
transform 1 0 3720 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_428
timestamp 1569533753
transform 1 0 3720 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_429
timestamp 1569533753
transform 1 0 3592 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_430
timestamp 1569533753
transform 1 0 3464 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_431
timestamp 1569533753
transform 1 0 3720 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_432
timestamp 1569533753
transform 1 0 2824 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_433
timestamp 1569533753
transform 1 0 3016 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_434
timestamp 1569533753
transform 1 0 2888 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_435
timestamp 1569533753
transform 1 0 3080 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_436
timestamp 1569533753
transform 1 0 3016 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_437
timestamp 1569533753
transform 1 0 3016 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_438
timestamp 1569533753
transform 1 0 3080 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_439
timestamp 1569533753
transform 1 0 2888 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_440
timestamp 1569533753
transform 1 0 2952 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_441
timestamp 1569533753
transform 1 0 2888 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_442
timestamp 1569533753
transform 1 0 2824 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_443
timestamp 1569533753
transform 1 0 2888 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_444
timestamp 1569533753
transform 1 0 2952 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_445
timestamp 1569533753
transform 1 0 2952 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_446
timestamp 1569533753
transform 1 0 2888 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_447
timestamp 1569533753
transform 1 0 2824 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_448
timestamp 1569533753
transform 1 0 2824 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_449
timestamp 1569533753
transform 1 0 3080 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_450
timestamp 1569533753
transform 1 0 2824 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_451
timestamp 1569533753
transform 1 0 3016 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_452
timestamp 1569533753
transform 1 0 2952 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_453
timestamp 1569533753
transform 1 0 3080 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_454
timestamp 1569533753
transform 1 0 3080 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_455
timestamp 1569533753
transform 1 0 3016 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_456
timestamp 1569533753
transform 1 0 2952 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_457
timestamp 1569533753
transform 1 0 2760 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_458
timestamp 1569533753
transform 1 0 2632 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_459
timestamp 1569533753
transform 1 0 2568 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_460
timestamp 1569533753
transform 1 0 2568 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_461
timestamp 1569533753
transform 1 0 2632 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_462
timestamp 1569533753
transform 1 0 2760 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_463
timestamp 1569533753
transform 1 0 2696 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_464
timestamp 1569533753
transform 1 0 2696 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_465
timestamp 1569533753
transform 1 0 2696 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_466
timestamp 1569533753
transform 1 0 2760 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_467
timestamp 1569533753
transform 1 0 2696 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_468
timestamp 1569533753
transform 1 0 2760 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_469
timestamp 1569533753
transform 1 0 2632 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_470
timestamp 1569533753
transform 1 0 2568 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_471
timestamp 1569533753
transform 1 0 2696 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_472
timestamp 1569533753
transform 1 0 2632 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_473
timestamp 1569533753
transform 1 0 2632 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_474
timestamp 1569533753
transform 1 0 2760 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_475
timestamp 1569533753
transform 1 0 2568 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_476
timestamp 1569533753
transform 1 0 2568 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_477
timestamp 1569533753
transform 1 0 2696 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_478
timestamp 1569533753
transform 1 0 2760 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_479
timestamp 1569533753
transform 1 0 2568 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_480
timestamp 1569533753
transform 1 0 2568 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_481
timestamp 1569533753
transform 1 0 2632 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_482
timestamp 1569533753
transform 1 0 2568 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_483
timestamp 1569533753
transform 1 0 2568 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_484
timestamp 1569533753
transform 1 0 2696 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_485
timestamp 1569533753
transform 1 0 2632 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_486
timestamp 1569533753
transform 1 0 2696 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_487
timestamp 1569533753
transform 1 0 2760 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_488
timestamp 1569533753
transform 1 0 2632 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_489
timestamp 1569533753
transform 1 0 2760 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_490
timestamp 1569533753
transform 1 0 2696 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_491
timestamp 1569533753
transform 1 0 2760 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_492
timestamp 1569533753
transform 1 0 2632 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_493
timestamp 1569533753
transform 1 0 2888 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_494
timestamp 1569533753
transform 1 0 2824 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_495
timestamp 1569533753
transform 1 0 3016 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_496
timestamp 1569533753
transform 1 0 3016 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_497
timestamp 1569533753
transform 1 0 2824 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_498
timestamp 1569533753
transform 1 0 2952 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_499
timestamp 1569533753
transform 1 0 2952 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_500
timestamp 1569533753
transform 1 0 2824 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_501
timestamp 1569533753
transform 1 0 3016 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_502
timestamp 1569533753
transform 1 0 2952 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_503
timestamp 1569533753
transform 1 0 3080 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_504
timestamp 1569533753
transform 1 0 2952 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_505
timestamp 1569533753
transform 1 0 3016 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_506
timestamp 1569533753
transform 1 0 3080 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_507
timestamp 1569533753
transform 1 0 3080 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_508
timestamp 1569533753
transform 1 0 3080 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_509
timestamp 1569533753
transform 1 0 2888 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_510
timestamp 1569533753
transform 1 0 2824 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_511
timestamp 1569533753
transform 1 0 2888 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_512
timestamp 1569533753
transform 1 0 2888 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_513
timestamp 1569533753
transform 1 0 2888 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_514
timestamp 1569533753
transform 1 0 2888 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_515
timestamp 1569533753
transform 1 0 3016 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_516
timestamp 1569533753
transform 1 0 2952 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_517
timestamp 1569533753
transform 1 0 3080 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_518
timestamp 1569533753
transform 1 0 3080 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_519
timestamp 1569533753
transform 1 0 3080 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_520
timestamp 1569533753
transform 1 0 3080 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_521
timestamp 1569533753
transform 1 0 2952 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_522
timestamp 1569533753
transform 1 0 2824 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_523
timestamp 1569533753
transform 1 0 2824 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_524
timestamp 1569533753
transform 1 0 2824 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_525
timestamp 1569533753
transform 1 0 2952 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_526
timestamp 1569533753
transform 1 0 3016 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_527
timestamp 1569533753
transform 1 0 3016 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_528
timestamp 1569533753
transform 1 0 3016 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_529
timestamp 1569533753
transform 1 0 2888 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_530
timestamp 1569533753
transform 1 0 2824 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_531
timestamp 1569533753
transform 1 0 2888 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_532
timestamp 1569533753
transform 1 0 2952 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_533
timestamp 1569533753
transform 1 0 2568 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_534
timestamp 1569533753
transform 1 0 2696 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_535
timestamp 1569533753
transform 1 0 2632 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_536
timestamp 1569533753
transform 1 0 2760 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_537
timestamp 1569533753
transform 1 0 2760 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_538
timestamp 1569533753
transform 1 0 2696 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_539
timestamp 1569533753
transform 1 0 2632 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_540
timestamp 1569533753
transform 1 0 2568 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_541
timestamp 1569533753
transform 1 0 2696 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_542
timestamp 1569533753
transform 1 0 2568 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_543
timestamp 1569533753
transform 1 0 2632 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_544
timestamp 1569533753
transform 1 0 2760 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_545
timestamp 1569533753
transform 1 0 2632 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_546
timestamp 1569533753
transform 1 0 2696 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_547
timestamp 1569533753
transform 1 0 2568 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_548
timestamp 1569533753
transform 1 0 2760 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_549
timestamp 1569533753
transform 1 0 2760 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_550
timestamp 1569533753
transform 1 0 2632 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_551
timestamp 1569533753
transform 1 0 2760 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_552
timestamp 1569533753
transform 1 0 2760 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_553
timestamp 1569533753
transform 1 0 2696 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_554
timestamp 1569533753
transform 1 0 2696 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_555
timestamp 1569533753
transform 1 0 2568 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_556
timestamp 1569533753
transform 1 0 2632 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_557
timestamp 1569533753
transform 1 0 2632 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_558
timestamp 1569533753
transform 1 0 2760 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_559
timestamp 1569533753
transform 1 0 2568 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_560
timestamp 1569533753
transform 1 0 2696 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_561
timestamp 1569533753
transform 1 0 2568 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_562
timestamp 1569533753
transform 1 0 2696 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_563
timestamp 1569533753
transform 1 0 2568 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_564
timestamp 1569533753
transform 1 0 2632 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_565
timestamp 1569533753
transform 1 0 2696 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_566
timestamp 1569533753
transform 1 0 2568 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_567
timestamp 1569533753
transform 1 0 2760 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_568
timestamp 1569533753
transform 1 0 2632 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_569
timestamp 1569533753
transform 1 0 3080 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_570
timestamp 1569533753
transform 1 0 2824 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_571
timestamp 1569533753
transform 1 0 3080 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_572
timestamp 1569533753
transform 1 0 2824 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_573
timestamp 1569533753
transform 1 0 2824 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_574
timestamp 1569533753
transform 1 0 3080 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_575
timestamp 1569533753
transform 1 0 2824 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_576
timestamp 1569533753
transform 1 0 2824 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_577
timestamp 1569533753
transform 1 0 3080 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_578
timestamp 1569533753
transform 1 0 3080 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_579
timestamp 1569533753
transform 1 0 2888 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_580
timestamp 1569533753
transform 1 0 2888 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_581
timestamp 1569533753
transform 1 0 2888 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_582
timestamp 1569533753
transform 1 0 2888 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_583
timestamp 1569533753
transform 1 0 2888 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_584
timestamp 1569533753
transform 1 0 2952 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_585
timestamp 1569533753
transform 1 0 2952 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_586
timestamp 1569533753
transform 1 0 2952 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_587
timestamp 1569533753
transform 1 0 2952 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_588
timestamp 1569533753
transform 1 0 2952 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_589
timestamp 1569533753
transform 1 0 3016 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_590
timestamp 1569533753
transform 1 0 3016 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_591
timestamp 1569533753
transform 1 0 3016 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_592
timestamp 1569533753
transform 1 0 3016 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_593
timestamp 1569533753
transform 1 0 3016 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_594
timestamp 1569533753
transform 1 0 3656 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_595
timestamp 1569533753
transform 1 0 3592 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_596
timestamp 1569533753
transform 1 0 3592 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_597
timestamp 1569533753
transform 1 0 3720 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_598
timestamp 1569533753
transform 1 0 3528 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_599
timestamp 1569533753
transform 1 0 3720 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_600
timestamp 1569533753
transform 1 0 3464 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_601
timestamp 1569533753
transform 1 0 3464 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_602
timestamp 1569533753
transform 1 0 3720 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_603
timestamp 1569533753
transform 1 0 3656 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_604
timestamp 1569533753
transform 1 0 3720 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_605
timestamp 1569533753
transform 1 0 3656 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_606
timestamp 1569533753
transform 1 0 3592 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_607
timestamp 1569533753
transform 1 0 3464 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_608
timestamp 1569533753
transform 1 0 3528 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_609
timestamp 1569533753
transform 1 0 3528 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_610
timestamp 1569533753
transform 1 0 3656 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_611
timestamp 1569533753
transform 1 0 3464 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_612
timestamp 1569533753
transform 1 0 3528 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_613
timestamp 1569533753
transform 1 0 3592 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_614
timestamp 1569533753
transform 1 0 3272 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_615
timestamp 1569533753
transform 1 0 3336 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_616
timestamp 1569533753
transform 1 0 3400 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_617
timestamp 1569533753
transform 1 0 3400 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_618
timestamp 1569533753
transform 1 0 3336 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_619
timestamp 1569533753
transform 1 0 3208 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_620
timestamp 1569533753
transform 1 0 3144 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_621
timestamp 1569533753
transform 1 0 3144 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_622
timestamp 1569533753
transform 1 0 3272 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_623
timestamp 1569533753
transform 1 0 3400 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_624
timestamp 1569533753
transform 1 0 3144 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_625
timestamp 1569533753
transform 1 0 3208 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_626
timestamp 1569533753
transform 1 0 3144 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_627
timestamp 1569533753
transform 1 0 3208 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_628
timestamp 1569533753
transform 1 0 3272 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_629
timestamp 1569533753
transform 1 0 3208 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_630
timestamp 1569533753
transform 1 0 3400 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_631
timestamp 1569533753
transform 1 0 3336 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_632
timestamp 1569533753
transform 1 0 3272 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_633
timestamp 1569533753
transform 1 0 3336 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_634
timestamp 1569533753
transform 1 0 3400 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_635
timestamp 1569533753
transform 1 0 3400 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_636
timestamp 1569533753
transform 1 0 3400 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_637
timestamp 1569533753
transform 1 0 3208 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_638
timestamp 1569533753
transform 1 0 3208 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_639
timestamp 1569533753
transform 1 0 3208 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_640
timestamp 1569533753
transform 1 0 3272 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_641
timestamp 1569533753
transform 1 0 3336 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_642
timestamp 1569533753
transform 1 0 3272 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_643
timestamp 1569533753
transform 1 0 3144 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_644
timestamp 1569533753
transform 1 0 3144 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_645
timestamp 1569533753
transform 1 0 3144 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_646
timestamp 1569533753
transform 1 0 3144 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_647
timestamp 1569533753
transform 1 0 3272 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_648
timestamp 1569533753
transform 1 0 3208 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_649
timestamp 1569533753
transform 1 0 3144 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_650
timestamp 1569533753
transform 1 0 3272 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_651
timestamp 1569533753
transform 1 0 3336 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_652
timestamp 1569533753
transform 1 0 3336 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_653
timestamp 1569533753
transform 1 0 3336 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_654
timestamp 1569533753
transform 1 0 3272 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_655
timestamp 1569533753
transform 1 0 3400 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_656
timestamp 1569533753
transform 1 0 3336 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_657
timestamp 1569533753
transform 1 0 3208 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_658
timestamp 1569533753
transform 1 0 3400 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_659
timestamp 1569533753
transform 1 0 3464 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_660
timestamp 1569533753
transform 1 0 3464 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_661
timestamp 1569533753
transform 1 0 3464 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_662
timestamp 1569533753
transform 1 0 3464 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_663
timestamp 1569533753
transform 1 0 3464 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_664
timestamp 1569533753
transform 1 0 3528 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_665
timestamp 1569533753
transform 1 0 3528 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_666
timestamp 1569533753
transform 1 0 3528 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_667
timestamp 1569533753
transform 1 0 3528 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_668
timestamp 1569533753
transform 1 0 3528 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_669
timestamp 1569533753
transform 1 0 3592 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_670
timestamp 1569533753
transform 1 0 3592 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_671
timestamp 1569533753
transform 1 0 3592 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_672
timestamp 1569533753
transform 1 0 3592 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_673
timestamp 1569533753
transform 1 0 3592 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_674
timestamp 1569533753
transform 1 0 3656 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_675
timestamp 1569533753
transform 1 0 3656 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_676
timestamp 1569533753
transform 1 0 3656 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_677
timestamp 1569533753
transform 1 0 3656 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_678
timestamp 1569533753
transform 1 0 3656 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_679
timestamp 1569533753
transform 1 0 3720 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_680
timestamp 1569533753
transform 1 0 3720 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_681
timestamp 1569533753
transform 1 0 3720 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_682
timestamp 1569533753
transform 1 0 3720 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_683
timestamp 1569533753
transform 1 0 3720 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_684
timestamp 1569533753
transform 1 0 3080 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_685
timestamp 1569533753
transform 1 0 3720 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_686
timestamp 1569533753
transform 1 0 3144 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_687
timestamp 1569533753
transform 1 0 2568 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_688
timestamp 1569533753
transform 1 0 3208 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_689
timestamp 1569533753
transform 1 0 2632 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_690
timestamp 1569533753
transform 1 0 3272 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_691
timestamp 1569533753
transform 1 0 2888 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_692
timestamp 1569533753
transform 1 0 3528 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_693
timestamp 1569533753
transform 1 0 2696 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_694
timestamp 1569533753
transform 1 0 3336 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_695
timestamp 1569533753
transform 1 0 2760 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_696
timestamp 1569533753
transform 1 0 3400 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_697
timestamp 1569533753
transform 1 0 2952 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_698
timestamp 1569533753
transform 1 0 3592 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_699
timestamp 1569533753
transform 1 0 3016 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_700
timestamp 1569533753
transform 1 0 3656 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_701
timestamp 1569533753
transform 1 0 2824 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_702
timestamp 1569533753
transform 1 0 3464 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_703
timestamp 1569533753
transform 1 0 3144 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_704
timestamp 1569533753
transform 1 0 3208 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_705
timestamp 1569533753
transform 1 0 3400 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_706
timestamp 1569533753
transform 1 0 3592 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_707
timestamp 1569533753
transform 1 0 3144 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_708
timestamp 1569533753
transform 1 0 3400 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_709
timestamp 1569533753
transform 1 0 3656 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_710
timestamp 1569533753
transform 1 0 3592 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_711
timestamp 1569533753
transform 1 0 3720 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_712
timestamp 1569533753
transform 1 0 3400 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_713
timestamp 1569533753
transform 1 0 3208 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_714
timestamp 1569533753
transform 1 0 3272 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_715
timestamp 1569533753
transform 1 0 3400 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_716
timestamp 1569533753
transform 1 0 3656 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_717
timestamp 1569533753
transform 1 0 3144 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_718
timestamp 1569533753
transform 1 0 3144 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_719
timestamp 1569533753
transform 1 0 3336 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_720
timestamp 1569533753
transform 1 0 3336 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_721
timestamp 1569533753
transform 1 0 3464 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_722
timestamp 1569533753
transform 1 0 3656 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_723
timestamp 1569533753
transform 1 0 3592 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_724
timestamp 1569533753
transform 1 0 3464 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_725
timestamp 1569533753
transform 1 0 3720 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_726
timestamp 1569533753
transform 1 0 3272 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_727
timestamp 1569533753
transform 1 0 3464 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_728
timestamp 1569533753
transform 1 0 3464 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_729
timestamp 1569533753
transform 1 0 3208 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_730
timestamp 1569533753
transform 1 0 3528 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_731
timestamp 1569533753
transform 1 0 3592 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_732
timestamp 1569533753
transform 1 0 3528 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_733
timestamp 1569533753
transform 1 0 3272 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_734
timestamp 1569533753
transform 1 0 3528 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_735
timestamp 1569533753
transform 1 0 3528 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_736
timestamp 1569533753
transform 1 0 3720 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_737
timestamp 1569533753
transform 1 0 3272 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_738
timestamp 1569533753
transform 1 0 3336 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_739
timestamp 1569533753
transform 1 0 3656 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_740
timestamp 1569533753
transform 1 0 3720 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_741
timestamp 1569533753
transform 1 0 3336 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_742
timestamp 1569533753
transform 1 0 3208 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_743
timestamp 1569533753
transform 1 0 2824 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_744
timestamp 1569533753
transform 1 0 3016 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_745
timestamp 1569533753
transform 1 0 2888 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_746
timestamp 1569533753
transform 1 0 2952 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_747
timestamp 1569533753
transform 1 0 2952 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_748
timestamp 1569533753
transform 1 0 2952 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_749
timestamp 1569533753
transform 1 0 3016 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_750
timestamp 1569533753
transform 1 0 2888 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_751
timestamp 1569533753
transform 1 0 3080 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_752
timestamp 1569533753
transform 1 0 3080 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_753
timestamp 1569533753
transform 1 0 3016 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_754
timestamp 1569533753
transform 1 0 2824 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_755
timestamp 1569533753
transform 1 0 2824 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_756
timestamp 1569533753
transform 1 0 2824 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_757
timestamp 1569533753
transform 1 0 2888 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_758
timestamp 1569533753
transform 1 0 3016 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_759
timestamp 1569533753
transform 1 0 2888 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_760
timestamp 1569533753
transform 1 0 2888 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_761
timestamp 1569533753
transform 1 0 3080 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_762
timestamp 1569533753
transform 1 0 3080 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_763
timestamp 1569533753
transform 1 0 2952 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_764
timestamp 1569533753
transform 1 0 2824 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_765
timestamp 1569533753
transform 1 0 2696 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_766
timestamp 1569533753
transform 1 0 2760 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_767
timestamp 1569533753
transform 1 0 2760 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_768
timestamp 1569533753
transform 1 0 2632 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_769
timestamp 1569533753
transform 1 0 2760 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_770
timestamp 1569533753
transform 1 0 2568 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_771
timestamp 1569533753
transform 1 0 2568 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_772
timestamp 1569533753
transform 1 0 2632 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_773
timestamp 1569533753
transform 1 0 2632 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_774
timestamp 1569533753
transform 1 0 2568 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_775
timestamp 1569533753
transform 1 0 2696 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_776
timestamp 1569533753
transform 1 0 2696 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_777
timestamp 1569533753
transform 1 0 2696 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_778
timestamp 1569533753
transform 1 0 2632 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_779
timestamp 1569533753
transform 1 0 2568 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_780
timestamp 1569533753
transform 1 0 2696 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_781
timestamp 1569533753
transform 1 0 2760 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_782
timestamp 1569533753
transform 1 0 2760 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_783
timestamp 1569533753
transform 1 0 2568 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_784
timestamp 1569533753
transform 1 0 2632 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_785
timestamp 1569533753
transform 1 0 2568 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_786
timestamp 1569533753
transform 1 0 2632 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_787
timestamp 1569533753
transform 1 0 2632 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_788
timestamp 1569533753
transform 1 0 2632 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_789
timestamp 1569533753
transform 1 0 2632 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_790
timestamp 1569533753
transform 1 0 2568 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_791
timestamp 1569533753
transform 1 0 2568 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_792
timestamp 1569533753
transform 1 0 2696 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_793
timestamp 1569533753
transform 1 0 2696 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_794
timestamp 1569533753
transform 1 0 2696 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_795
timestamp 1569533753
transform 1 0 2760 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_796
timestamp 1569533753
transform 1 0 2760 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_797
timestamp 1569533753
transform 1 0 2568 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_798
timestamp 1569533753
transform 1 0 2568 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_799
timestamp 1569533753
transform 1 0 2824 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_800
timestamp 1569533753
transform 1 0 3400 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_801
timestamp 1569533753
transform 1 0 3720 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_802
timestamp 1569533753
transform 1 0 3464 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_803
timestamp 1569533753
transform 1 0 3528 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_804
timestamp 1569533753
transform 1 0 3272 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_805
timestamp 1569533753
transform 1 0 3592 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_806
timestamp 1569533753
transform 1 0 3656 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_807
timestamp 1569533753
transform 1 0 3336 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_808
timestamp 1569533753
transform 1 0 3592 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_809
timestamp 1569533753
transform 1 0 3336 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_810
timestamp 1569533753
transform 1 0 3656 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_811
timestamp 1569533753
transform 1 0 3400 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_812
timestamp 1569533753
transform 1 0 3720 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_813
timestamp 1569533753
transform 1 0 3464 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_814
timestamp 1569533753
transform 1 0 3464 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_815
timestamp 1569533753
transform 1 0 3528 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_816
timestamp 1569533753
transform 1 0 3592 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_817
timestamp 1569533753
transform 1 0 3528 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_818
timestamp 1569533753
transform 1 0 3400 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_819
timestamp 1569533753
transform 1 0 3656 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_820
timestamp 1569533753
transform 1 0 3720 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_821
timestamp 1569533753
transform 1 0 4744 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_822
timestamp 1569533753
transform 1 0 4680 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_823
timestamp 1569533753
transform 1 0 4680 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_824
timestamp 1569533753
transform 1 0 4872 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_825
timestamp 1569533753
transform 1 0 4552 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_826
timestamp 1569533753
transform 1 0 4424 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_827
timestamp 1569533753
transform 1 0 4616 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_828
timestamp 1569533753
transform 1 0 4488 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_829
timestamp 1569533753
transform 1 0 4424 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_830
timestamp 1569533753
transform 1 0 4744 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_831
timestamp 1569533753
transform 1 0 4744 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_832
timestamp 1569533753
transform 1 0 4680 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_833
timestamp 1569533753
transform 1 0 4808 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_834
timestamp 1569533753
transform 1 0 4488 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_835
timestamp 1569533753
transform 1 0 4808 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_836
timestamp 1569533753
transform 1 0 4424 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_837
timestamp 1569533753
transform 1 0 4808 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_838
timestamp 1569533753
transform 1 0 4552 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_839
timestamp 1569533753
transform 1 0 4616 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_840
timestamp 1569533753
transform 1 0 4616 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_841
timestamp 1569533753
transform 1 0 4552 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_842
timestamp 1569533753
transform 1 0 4680 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_843
timestamp 1569533753
transform 1 0 4744 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_844
timestamp 1569533753
transform 1 0 4616 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_845
timestamp 1569533753
transform 1 0 4488 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_846
timestamp 1569533753
transform 1 0 4808 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_847
timestamp 1569533753
transform 1 0 4552 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_848
timestamp 1569533753
transform 1 0 4872 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_849
timestamp 1569533753
transform 1 0 4488 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_850
timestamp 1569533753
transform 1 0 4872 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_851
timestamp 1569533753
transform 1 0 4424 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_852
timestamp 1569533753
transform 1 0 4872 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_853
timestamp 1569533753
transform 1 0 3848 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_854
timestamp 1569533753
transform 1 0 4040 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_855
timestamp 1569533753
transform 1 0 4040 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_856
timestamp 1569533753
transform 1 0 4232 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_857
timestamp 1569533753
transform 1 0 4040 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_858
timestamp 1569533753
transform 1 0 4232 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_859
timestamp 1569533753
transform 1 0 4232 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_860
timestamp 1569533753
transform 1 0 3848 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_861
timestamp 1569533753
transform 1 0 3848 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_862
timestamp 1569533753
transform 1 0 4232 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_863
timestamp 1569533753
transform 1 0 4104 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_864
timestamp 1569533753
transform 1 0 4104 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_865
timestamp 1569533753
transform 1 0 4104 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_866
timestamp 1569533753
transform 1 0 4168 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_867
timestamp 1569533753
transform 1 0 4168 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_868
timestamp 1569533753
transform 1 0 4168 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_869
timestamp 1569533753
transform 1 0 3912 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_870
timestamp 1569533753
transform 1 0 3976 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_871
timestamp 1569533753
transform 1 0 4040 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_872
timestamp 1569533753
transform 1 0 4104 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_873
timestamp 1569533753
transform 1 0 4168 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_874
timestamp 1569533753
transform 1 0 4296 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_875
timestamp 1569533753
transform 1 0 4296 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_876
timestamp 1569533753
transform 1 0 4296 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_877
timestamp 1569533753
transform 1 0 4296 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_878
timestamp 1569533753
transform 1 0 3976 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_879
timestamp 1569533753
transform 1 0 3976 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_880
timestamp 1569533753
transform 1 0 3912 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_881
timestamp 1569533753
transform 1 0 3784 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_882
timestamp 1569533753
transform 1 0 3848 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_883
timestamp 1569533753
transform 1 0 3912 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_884
timestamp 1569533753
transform 1 0 3784 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_885
timestamp 1569533753
transform 1 0 3784 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_886
timestamp 1569533753
transform 1 0 3784 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_887
timestamp 1569533753
transform 1 0 3912 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_888
timestamp 1569533753
transform 1 0 3976 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_889
timestamp 1569533753
transform 1 0 4168 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_890
timestamp 1569533753
transform 1 0 3912 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_891
timestamp 1569533753
transform 1 0 4296 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_892
timestamp 1569533753
transform 1 0 4232 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_893
timestamp 1569533753
transform 1 0 3976 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_894
timestamp 1569533753
transform 1 0 3784 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_895
timestamp 1569533753
transform 1 0 4296 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_896
timestamp 1569533753
transform 1 0 4040 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_897
timestamp 1569533753
transform 1 0 3848 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_898
timestamp 1569533753
transform 1 0 4040 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_899
timestamp 1569533753
transform 1 0 4104 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_900
timestamp 1569533753
transform 1 0 3912 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_901
timestamp 1569533753
transform 1 0 3848 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_902
timestamp 1569533753
transform 1 0 4168 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_903
timestamp 1569533753
transform 1 0 3976 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_904
timestamp 1569533753
transform 1 0 4232 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_905
timestamp 1569533753
transform 1 0 4040 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_906
timestamp 1569533753
transform 1 0 3784 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_907
timestamp 1569533753
transform 1 0 4296 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_908
timestamp 1569533753
transform 1 0 4104 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_909
timestamp 1569533753
transform 1 0 3848 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_910
timestamp 1569533753
transform 1 0 4232 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_911
timestamp 1569533753
transform 1 0 3784 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_912
timestamp 1569533753
transform 1 0 4168 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_913
timestamp 1569533753
transform 1 0 3912 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_914
timestamp 1569533753
transform 1 0 3976 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_915
timestamp 1569533753
transform 1 0 4104 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_916
timestamp 1569533753
transform 1 0 4680 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_917
timestamp 1569533753
transform 1 0 4488 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_918
timestamp 1569533753
transform 1 0 4744 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_919
timestamp 1569533753
transform 1 0 4552 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_920
timestamp 1569533753
transform 1 0 4808 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_921
timestamp 1569533753
transform 1 0 4616 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_922
timestamp 1569533753
transform 1 0 4552 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_923
timestamp 1569533753
transform 1 0 4872 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_924
timestamp 1569533753
transform 1 0 4680 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_925
timestamp 1569533753
transform 1 0 4424 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_926
timestamp 1569533753
transform 1 0 4744 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_927
timestamp 1569533753
transform 1 0 4488 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_928
timestamp 1569533753
transform 1 0 4808 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_929
timestamp 1569533753
transform 1 0 4552 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_930
timestamp 1569533753
transform 1 0 4872 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_931
timestamp 1569533753
transform 1 0 4616 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_932
timestamp 1569533753
transform 1 0 4680 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_933
timestamp 1569533753
transform 1 0 4424 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_934
timestamp 1569533753
transform 1 0 4424 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_935
timestamp 1569533753
transform 1 0 4872 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_936
timestamp 1569533753
transform 1 0 4616 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_937
timestamp 1569533753
transform 1 0 4744 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_938
timestamp 1569533753
transform 1 0 4488 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_939
timestamp 1569533753
transform 1 0 4808 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_940
timestamp 1569533753
transform 1 0 4360 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_941
timestamp 1569533753
transform 1 0 4360 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_942
timestamp 1569533753
transform 1 0 4360 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_943
timestamp 1569533753
transform 1 0 4360 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_944
timestamp 1569533753
transform 1 0 4360 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_945
timestamp 1569533753
transform 1 0 4360 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_946
timestamp 1569533753
transform 1 0 4360 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_947
timestamp 1569533753
transform 1 0 2376 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_948
timestamp 1569533753
transform 1 0 2312 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_949
timestamp 1569533753
transform 1 0 2440 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_950
timestamp 1569533753
transform 1 0 2248 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_951
timestamp 1569533753
transform 1 0 2312 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_952
timestamp 1569533753
transform 1 0 2248 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_953
timestamp 1569533753
transform 1 0 2312 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_954
timestamp 1569533753
transform 1 0 2376 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_955
timestamp 1569533753
transform 1 0 2312 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_956
timestamp 1569533753
transform 1 0 2440 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_957
timestamp 1569533753
transform 1 0 2376 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_958
timestamp 1569533753
transform 1 0 2440 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_959
timestamp 1569533753
transform 1 0 2248 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_960
timestamp 1569533753
transform 1 0 2312 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_961
timestamp 1569533753
transform 1 0 2248 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_962
timestamp 1569533753
transform 1 0 2376 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_963
timestamp 1569533753
transform 1 0 2440 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_964
timestamp 1569533753
transform 1 0 2376 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_965
timestamp 1569533753
transform 1 0 2440 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_966
timestamp 1569533753
transform 1 0 2248 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_967
timestamp 1569533753
transform 1 0 2184 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_968
timestamp 1569533753
transform 1 0 2056 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_969
timestamp 1569533753
transform 1 0 1928 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_970
timestamp 1569533753
transform 1 0 2120 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_971
timestamp 1569533753
transform 1 0 2120 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_972
timestamp 1569533753
transform 1 0 2120 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_973
timestamp 1569533753
transform 1 0 1928 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_974
timestamp 1569533753
transform 1 0 2120 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_975
timestamp 1569533753
transform 1 0 1928 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_976
timestamp 1569533753
transform 1 0 1992 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_977
timestamp 1569533753
transform 1 0 2120 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_978
timestamp 1569533753
transform 1 0 1928 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_979
timestamp 1569533753
transform 1 0 1992 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_980
timestamp 1569533753
transform 1 0 1992 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_981
timestamp 1569533753
transform 1 0 2184 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_982
timestamp 1569533753
transform 1 0 1992 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_983
timestamp 1569533753
transform 1 0 2184 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_984
timestamp 1569533753
transform 1 0 1992 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_985
timestamp 1569533753
transform 1 0 1928 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_986
timestamp 1569533753
transform 1 0 2056 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_987
timestamp 1569533753
transform 1 0 2056 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_988
timestamp 1569533753
transform 1 0 2184 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_989
timestamp 1569533753
transform 1 0 2056 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_990
timestamp 1569533753
transform 1 0 2056 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_991
timestamp 1569533753
transform 1 0 2184 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_992
timestamp 1569533753
transform 1 0 1928 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_993
timestamp 1569533753
transform 1 0 2120 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_994
timestamp 1569533753
transform 1 0 2184 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_995
timestamp 1569533753
transform 1 0 2120 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_996
timestamp 1569533753
transform 1 0 2120 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_997
timestamp 1569533753
transform 1 0 1928 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_998
timestamp 1569533753
transform 1 0 2120 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_999
timestamp 1569533753
transform 1 0 2056 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1000
timestamp 1569533753
transform 1 0 1928 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1001
timestamp 1569533753
transform 1 0 2056 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1002
timestamp 1569533753
transform 1 0 1992 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1003
timestamp 1569533753
transform 1 0 1992 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1004
timestamp 1569533753
transform 1 0 1992 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1005
timestamp 1569533753
transform 1 0 1928 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1006
timestamp 1569533753
transform 1 0 2184 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1007
timestamp 1569533753
transform 1 0 1992 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1008
timestamp 1569533753
transform 1 0 2184 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1009
timestamp 1569533753
transform 1 0 2056 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1010
timestamp 1569533753
transform 1 0 2056 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1011
timestamp 1569533753
transform 1 0 2184 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1012
timestamp 1569533753
transform 1 0 2376 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1013
timestamp 1569533753
transform 1 0 2440 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1014
timestamp 1569533753
transform 1 0 2376 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1015
timestamp 1569533753
transform 1 0 2376 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1016
timestamp 1569533753
transform 1 0 2376 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1017
timestamp 1569533753
transform 1 0 2312 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1018
timestamp 1569533753
transform 1 0 2312 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1019
timestamp 1569533753
transform 1 0 2312 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1020
timestamp 1569533753
transform 1 0 2312 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1021
timestamp 1569533753
transform 1 0 2440 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1022
timestamp 1569533753
transform 1 0 2440 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1023
timestamp 1569533753
transform 1 0 2248 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1024
timestamp 1569533753
transform 1 0 2248 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1025
timestamp 1569533753
transform 1 0 2248 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1026
timestamp 1569533753
transform 1 0 2248 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1027
timestamp 1569533753
transform 1 0 2440 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1028
timestamp 1569533753
transform 1 0 1864 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1029
timestamp 1569533753
transform 1 0 1864 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_1030
timestamp 1569533753
transform 1 0 1736 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1031
timestamp 1569533753
transform 1 0 1736 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_1032
timestamp 1569533753
transform 1 0 1864 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_1033
timestamp 1569533753
transform 1 0 1800 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_1034
timestamp 1569533753
transform 1 0 1672 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_1035
timestamp 1569533753
transform 1 0 1672 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_1036
timestamp 1569533753
transform 1 0 1672 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1037
timestamp 1569533753
transform 1 0 1672 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1038
timestamp 1569533753
transform 1 0 1736 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1039
timestamp 1569533753
transform 1 0 1800 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_1040
timestamp 1569533753
transform 1 0 1800 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_1041
timestamp 1569533753
transform 1 0 1864 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1042
timestamp 1569533753
transform 1 0 1608 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_1043
timestamp 1569533753
transform 1 0 1608 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1044
timestamp 1569533753
transform 1 0 1608 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1045
timestamp 1569533753
transform 1 0 1736 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_1046
timestamp 1569533753
transform 1 0 1864 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_1047
timestamp 1569533753
transform 1 0 1800 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1048
timestamp 1569533753
transform 1 0 1800 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1049
timestamp 1569533753
transform 1 0 1736 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_1050
timestamp 1569533753
transform 1 0 1544 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_1051
timestamp 1569533753
transform 1 0 1544 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1052
timestamp 1569533753
transform 1 0 1480 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_1053
timestamp 1569533753
transform 1 0 1544 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1054
timestamp 1569533753
transform 1 0 1544 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1055
timestamp 1569533753
transform 1 0 1544 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1056
timestamp 1569533753
transform 1 0 1544 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1057
timestamp 1569533753
transform 1 0 1288 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1058
timestamp 1569533753
transform 1 0 1416 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1059
timestamp 1569533753
transform 1 0 1416 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1060
timestamp 1569533753
transform 1 0 1416 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1061
timestamp 1569533753
transform 1 0 1416 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1062
timestamp 1569533753
transform 1 0 1480 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1063
timestamp 1569533753
transform 1 0 1480 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1064
timestamp 1569533753
transform 1 0 1480 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1065
timestamp 1569533753
transform 1 0 1352 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1066
timestamp 1569533753
transform 1 0 1352 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1067
timestamp 1569533753
transform 1 0 1352 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1068
timestamp 1569533753
transform 1 0 1480 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1069
timestamp 1569533753
transform 1 0 1288 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1070
timestamp 1569533753
transform 1 0 1736 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1071
timestamp 1569533753
transform 1 0 1608 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1072
timestamp 1569533753
transform 1 0 1608 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1073
timestamp 1569533753
transform 1 0 1608 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1074
timestamp 1569533753
transform 1 0 1608 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1075
timestamp 1569533753
transform 1 0 1800 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1076
timestamp 1569533753
transform 1 0 1736 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1077
timestamp 1569533753
transform 1 0 1800 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1078
timestamp 1569533753
transform 1 0 1736 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1079
timestamp 1569533753
transform 1 0 1736 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1080
timestamp 1569533753
transform 1 0 1672 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1081
timestamp 1569533753
transform 1 0 1672 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1082
timestamp 1569533753
transform 1 0 1672 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1083
timestamp 1569533753
transform 1 0 1672 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1084
timestamp 1569533753
transform 1 0 1864 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_1085
timestamp 1569533753
transform 1 0 1864 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_1086
timestamp 1569533753
transform 1 0 1864 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1087
timestamp 1569533753
transform 1 0 1800 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_1088
timestamp 1569533753
transform 1 0 1864 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1089
timestamp 1569533753
transform 1 0 1800 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1090
timestamp 1569533753
transform 1 0 1736 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1091
timestamp 1569533753
transform 1 0 1800 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1092
timestamp 1569533753
transform 1 0 1736 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1093
timestamp 1569533753
transform 1 0 1864 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1094
timestamp 1569533753
transform 1 0 1672 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1095
timestamp 1569533753
transform 1 0 1864 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1096
timestamp 1569533753
transform 1 0 1672 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1097
timestamp 1569533753
transform 1 0 1736 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1098
timestamp 1569533753
transform 1 0 1864 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1099
timestamp 1569533753
transform 1 0 1864 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1100
timestamp 1569533753
transform 1 0 1608 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1101
timestamp 1569533753
transform 1 0 1800 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1102
timestamp 1569533753
transform 1 0 1672 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1103
timestamp 1569533753
transform 1 0 1736 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1104
timestamp 1569533753
transform 1 0 1608 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1105
timestamp 1569533753
transform 1 0 1608 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1106
timestamp 1569533753
transform 1 0 1800 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1107
timestamp 1569533753
transform 1 0 1800 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1108
timestamp 1569533753
transform 1 0 1672 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1109
timestamp 1569533753
transform 1 0 1608 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1110
timestamp 1569533753
transform 1 0 1544 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1111
timestamp 1569533753
transform 1 0 1416 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1112
timestamp 1569533753
transform 1 0 1480 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1113
timestamp 1569533753
transform 1 0 1544 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1114
timestamp 1569533753
transform 1 0 1288 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1115
timestamp 1569533753
transform 1 0 1416 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1116
timestamp 1569533753
transform 1 0 1544 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1117
timestamp 1569533753
transform 1 0 1416 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1118
timestamp 1569533753
transform 1 0 1480 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1119
timestamp 1569533753
transform 1 0 1352 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1120
timestamp 1569533753
transform 1 0 1352 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1121
timestamp 1569533753
transform 1 0 1288 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1122
timestamp 1569533753
transform 1 0 1480 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1123
timestamp 1569533753
transform 1 0 1352 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1124
timestamp 1569533753
transform 1 0 1544 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1125
timestamp 1569533753
transform 1 0 1352 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1126
timestamp 1569533753
transform 1 0 1480 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1127
timestamp 1569533753
transform 1 0 1288 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1128
timestamp 1569533753
transform 1 0 1288 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1129
timestamp 1569533753
transform 1 0 1416 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1130
timestamp 1569533753
transform 1 0 1352 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1131
timestamp 1569533753
transform 1 0 1544 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1132
timestamp 1569533753
transform 1 0 1544 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1133
timestamp 1569533753
transform 1 0 1416 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1134
timestamp 1569533753
transform 1 0 1288 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1135
timestamp 1569533753
transform 1 0 1480 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1136
timestamp 1569533753
transform 1 0 1288 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1137
timestamp 1569533753
transform 1 0 1288 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1138
timestamp 1569533753
transform 1 0 1416 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1139
timestamp 1569533753
transform 1 0 1480 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1140
timestamp 1569533753
transform 1 0 1416 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1141
timestamp 1569533753
transform 1 0 1544 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1142
timestamp 1569533753
transform 1 0 1288 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1143
timestamp 1569533753
transform 1 0 1416 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1144
timestamp 1569533753
transform 1 0 1480 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1145
timestamp 1569533753
transform 1 0 1544 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1146
timestamp 1569533753
transform 1 0 1288 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1147
timestamp 1569533753
transform 1 0 1352 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1148
timestamp 1569533753
transform 1 0 1416 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1149
timestamp 1569533753
transform 1 0 1352 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1150
timestamp 1569533753
transform 1 0 1352 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1151
timestamp 1569533753
transform 1 0 1480 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1152
timestamp 1569533753
transform 1 0 1480 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1153
timestamp 1569533753
transform 1 0 1544 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1154
timestamp 1569533753
transform 1 0 1352 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1155
timestamp 1569533753
transform 1 0 1672 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1156
timestamp 1569533753
transform 1 0 1672 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1157
timestamp 1569533753
transform 1 0 1736 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1158
timestamp 1569533753
transform 1 0 1736 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1159
timestamp 1569533753
transform 1 0 1736 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1160
timestamp 1569533753
transform 1 0 1736 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1161
timestamp 1569533753
transform 1 0 1736 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1162
timestamp 1569533753
transform 1 0 1800 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1163
timestamp 1569533753
transform 1 0 1800 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1164
timestamp 1569533753
transform 1 0 1800 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1165
timestamp 1569533753
transform 1 0 1800 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1166
timestamp 1569533753
transform 1 0 1800 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1167
timestamp 1569533753
transform 1 0 1672 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1168
timestamp 1569533753
transform 1 0 1608 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1169
timestamp 1569533753
transform 1 0 1864 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1170
timestamp 1569533753
transform 1 0 1864 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1171
timestamp 1569533753
transform 1 0 1608 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1172
timestamp 1569533753
transform 1 0 1864 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1173
timestamp 1569533753
transform 1 0 1672 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1174
timestamp 1569533753
transform 1 0 1608 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1175
timestamp 1569533753
transform 1 0 1864 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1176
timestamp 1569533753
transform 1 0 1864 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1177
timestamp 1569533753
transform 1 0 1608 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1178
timestamp 1569533753
transform 1 0 1672 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1179
timestamp 1569533753
transform 1 0 1608 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1180
timestamp 1569533753
transform 1 0 2248 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1181
timestamp 1569533753
transform 1 0 2376 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1182
timestamp 1569533753
transform 1 0 2440 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1183
timestamp 1569533753
transform 1 0 2376 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1184
timestamp 1569533753
transform 1 0 2440 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1185
timestamp 1569533753
transform 1 0 2376 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1186
timestamp 1569533753
transform 1 0 2312 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1187
timestamp 1569533753
transform 1 0 2312 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1188
timestamp 1569533753
transform 1 0 2376 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1189
timestamp 1569533753
transform 1 0 2248 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1190
timestamp 1569533753
transform 1 0 2312 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1191
timestamp 1569533753
transform 1 0 2312 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1192
timestamp 1569533753
transform 1 0 2248 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1193
timestamp 1569533753
transform 1 0 2248 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1194
timestamp 1569533753
transform 1 0 2440 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1195
timestamp 1569533753
transform 1 0 2440 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1196
timestamp 1569533753
transform 1 0 1992 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1197
timestamp 1569533753
transform 1 0 1992 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1198
timestamp 1569533753
transform 1 0 2056 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1199
timestamp 1569533753
transform 1 0 2120 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1200
timestamp 1569533753
transform 1 0 2184 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1201
timestamp 1569533753
transform 1 0 2184 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1202
timestamp 1569533753
transform 1 0 1992 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1203
timestamp 1569533753
transform 1 0 1992 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1204
timestamp 1569533753
transform 1 0 1928 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1205
timestamp 1569533753
transform 1 0 1928 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1206
timestamp 1569533753
transform 1 0 2120 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1207
timestamp 1569533753
transform 1 0 2056 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1208
timestamp 1569533753
transform 1 0 2056 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1209
timestamp 1569533753
transform 1 0 2056 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1210
timestamp 1569533753
transform 1 0 1928 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1211
timestamp 1569533753
transform 1 0 1928 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1212
timestamp 1569533753
transform 1 0 2120 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1213
timestamp 1569533753
transform 1 0 2120 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1214
timestamp 1569533753
transform 1 0 2184 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1215
timestamp 1569533753
transform 1 0 2184 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1216
timestamp 1569533753
transform 1 0 1928 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1217
timestamp 1569533753
transform 1 0 2120 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1218
timestamp 1569533753
transform 1 0 1928 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1219
timestamp 1569533753
transform 1 0 2120 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1220
timestamp 1569533753
transform 1 0 2120 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1221
timestamp 1569533753
transform 1 0 2120 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1222
timestamp 1569533753
transform 1 0 2120 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1223
timestamp 1569533753
transform 1 0 2184 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1224
timestamp 1569533753
transform 1 0 2184 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1225
timestamp 1569533753
transform 1 0 2184 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1226
timestamp 1569533753
transform 1 0 1992 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1227
timestamp 1569533753
transform 1 0 1992 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1228
timestamp 1569533753
transform 1 0 1992 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1229
timestamp 1569533753
transform 1 0 1992 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1230
timestamp 1569533753
transform 1 0 1992 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1231
timestamp 1569533753
transform 1 0 2056 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1232
timestamp 1569533753
transform 1 0 2056 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1233
timestamp 1569533753
transform 1 0 2056 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1234
timestamp 1569533753
transform 1 0 2056 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1235
timestamp 1569533753
transform 1 0 2056 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1236
timestamp 1569533753
transform 1 0 2184 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1237
timestamp 1569533753
transform 1 0 2184 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1238
timestamp 1569533753
transform 1 0 1928 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1239
timestamp 1569533753
transform 1 0 1928 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1240
timestamp 1569533753
transform 1 0 1928 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1241
timestamp 1569533753
transform 1 0 2376 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1242
timestamp 1569533753
transform 1 0 2376 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1243
timestamp 1569533753
transform 1 0 2376 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1244
timestamp 1569533753
transform 1 0 2376 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1245
timestamp 1569533753
transform 1 0 2376 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1246
timestamp 1569533753
transform 1 0 2440 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1247
timestamp 1569533753
transform 1 0 2440 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1248
timestamp 1569533753
transform 1 0 2440 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1249
timestamp 1569533753
transform 1 0 2440 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1250
timestamp 1569533753
transform 1 0 2440 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1251
timestamp 1569533753
transform 1 0 2248 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1252
timestamp 1569533753
transform 1 0 2312 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1253
timestamp 1569533753
transform 1 0 2312 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1254
timestamp 1569533753
transform 1 0 2312 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1255
timestamp 1569533753
transform 1 0 2312 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1256
timestamp 1569533753
transform 1 0 2312 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1257
timestamp 1569533753
transform 1 0 2248 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1258
timestamp 1569533753
transform 1 0 2248 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1259
timestamp 1569533753
transform 1 0 2248 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1260
timestamp 1569533753
transform 1 0 2248 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1261
timestamp 1569533753
transform 1 0 1672 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1262
timestamp 1569533753
transform 1 0 2312 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1263
timestamp 1569533753
transform 1 0 1352 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1264
timestamp 1569533753
transform 1 0 1992 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1265
timestamp 1569533753
transform 1 0 1416 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1266
timestamp 1569533753
transform 1 0 2056 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1267
timestamp 1569533753
transform 1 0 1480 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1268
timestamp 1569533753
transform 1 0 2120 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1269
timestamp 1569533753
transform 1 0 1544 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1270
timestamp 1569533753
transform 1 0 2184 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1271
timestamp 1569533753
transform 1 0 1608 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1272
timestamp 1569533753
transform 1 0 2248 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1273
timestamp 1569533753
transform 1 0 1736 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1274
timestamp 1569533753
transform 1 0 2376 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1275
timestamp 1569533753
transform 1 0 1800 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1276
timestamp 1569533753
transform 1 0 2440 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1277
timestamp 1569533753
transform 1 0 1864 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1278
timestamp 1569533753
transform 1 0 1288 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1279
timestamp 1569533753
transform 1 0 1928 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1280
timestamp 1569533753
transform 1 0 1224 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_1281
timestamp 1569533753
transform 1 0 584 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1282
timestamp 1569533753
transform 1 0 968 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1283
timestamp 1569533753
transform 1 0 968 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1284
timestamp 1569533753
transform 1 0 1160 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1285
timestamp 1569533753
transform 1 0 1224 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1286
timestamp 1569533753
transform 1 0 1224 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1287
timestamp 1569533753
transform 1 0 1032 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1288
timestamp 1569533753
transform 1 0 1096 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1289
timestamp 1569533753
transform 1 0 1096 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_1290
timestamp 1569533753
transform 1 0 1032 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1291
timestamp 1569533753
transform 1 0 1032 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1292
timestamp 1569533753
transform 1 0 1096 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1293
timestamp 1569533753
transform 1 0 1096 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1294
timestamp 1569533753
transform 1 0 1224 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1295
timestamp 1569533753
transform 1 0 1160 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_1296
timestamp 1569533753
transform 1 0 1224 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1297
timestamp 1569533753
transform 1 0 1160 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_1298
timestamp 1569533753
transform 1 0 1160 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1299
timestamp 1569533753
transform 1 0 904 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_1300
timestamp 1569533753
transform 1 0 904 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1301
timestamp 1569533753
transform 1 0 904 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1302
timestamp 1569533753
transform 1 0 904 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1303
timestamp 1569533753
transform 1 0 904 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1304
timestamp 1569533753
transform 1 0 904 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1305
timestamp 1569533753
transform 1 0 840 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1306
timestamp 1569533753
transform 1 0 840 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1307
timestamp 1569533753
transform 1 0 840 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1308
timestamp 1569533753
transform 1 0 840 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1309
timestamp 1569533753
transform 1 0 840 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1310
timestamp 1569533753
transform 1 0 712 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1311
timestamp 1569533753
transform 1 0 712 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1312
timestamp 1569533753
transform 1 0 712 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1313
timestamp 1569533753
transform 1 0 776 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1314
timestamp 1569533753
transform 1 0 776 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1315
timestamp 1569533753
transform 1 0 776 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1316
timestamp 1569533753
transform 1 0 776 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1317
timestamp 1569533753
transform 1 0 1032 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1318
timestamp 1569533753
transform 1 0 1032 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1319
timestamp 1569533753
transform 1 0 1032 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1320
timestamp 1569533753
transform 1 0 1096 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1321
timestamp 1569533753
transform 1 0 1096 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1322
timestamp 1569533753
transform 1 0 1096 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1323
timestamp 1569533753
transform 1 0 1096 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1324
timestamp 1569533753
transform 1 0 1096 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1325
timestamp 1569533753
transform 1 0 1160 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1326
timestamp 1569533753
transform 1 0 1160 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1327
timestamp 1569533753
transform 1 0 1160 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1328
timestamp 1569533753
transform 1 0 1160 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1329
timestamp 1569533753
transform 1 0 1160 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1330
timestamp 1569533753
transform 1 0 968 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1331
timestamp 1569533753
transform 1 0 968 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1332
timestamp 1569533753
transform 1 0 968 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1333
timestamp 1569533753
transform 1 0 968 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1334
timestamp 1569533753
transform 1 0 968 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1335
timestamp 1569533753
transform 1 0 1224 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1336
timestamp 1569533753
transform 1 0 1224 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1337
timestamp 1569533753
transform 1 0 1224 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_1338
timestamp 1569533753
transform 1 0 1224 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1339
timestamp 1569533753
transform 1 0 1224 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1340
timestamp 1569533753
transform 1 0 1032 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_1341
timestamp 1569533753
transform 1 0 1032 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_1342
timestamp 1569533753
transform 1 0 648 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_1343
timestamp 1569533753
transform 1 0 648 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_1344
timestamp 1569533753
transform 1 0 1160 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1345
timestamp 1569533753
transform 1 0 1224 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_1346
timestamp 1569533753
transform 1 0 1160 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1347
timestamp 1569533753
transform 1 0 1096 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1348
timestamp 1569533753
transform 1 0 1160 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1349
timestamp 1569533753
transform 1 0 1096 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1350
timestamp 1569533753
transform 1 0 1032 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1351
timestamp 1569533753
transform 1 0 968 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1352
timestamp 1569533753
transform 1 0 1160 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1353
timestamp 1569533753
transform 1 0 1160 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1354
timestamp 1569533753
transform 1 0 1096 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1355
timestamp 1569533753
transform 1 0 968 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1356
timestamp 1569533753
transform 1 0 1096 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1357
timestamp 1569533753
transform 1 0 1096 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1358
timestamp 1569533753
transform 1 0 1032 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1359
timestamp 1569533753
transform 1 0 968 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1360
timestamp 1569533753
transform 1 0 1224 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1361
timestamp 1569533753
transform 1 0 1032 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1362
timestamp 1569533753
transform 1 0 968 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1363
timestamp 1569533753
transform 1 0 1224 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1364
timestamp 1569533753
transform 1 0 968 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1365
timestamp 1569533753
transform 1 0 1224 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1366
timestamp 1569533753
transform 1 0 1032 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1367
timestamp 1569533753
transform 1 0 1224 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1368
timestamp 1569533753
transform 1 0 1224 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1369
timestamp 1569533753
transform 1 0 1160 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1370
timestamp 1569533753
transform 1 0 1032 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1371
timestamp 1569533753
transform 1 0 776 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1372
timestamp 1569533753
transform 1 0 840 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1373
timestamp 1569533753
transform 1 0 904 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1374
timestamp 1569533753
transform 1 0 840 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1375
timestamp 1569533753
transform 1 0 712 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1376
timestamp 1569533753
transform 1 0 904 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1377
timestamp 1569533753
transform 1 0 776 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1378
timestamp 1569533753
transform 1 0 712 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1379
timestamp 1569533753
transform 1 0 904 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1380
timestamp 1569533753
transform 1 0 712 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1381
timestamp 1569533753
transform 1 0 840 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1382
timestamp 1569533753
transform 1 0 904 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1383
timestamp 1569533753
transform 1 0 712 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1384
timestamp 1569533753
transform 1 0 840 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1385
timestamp 1569533753
transform 1 0 904 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1386
timestamp 1569533753
transform 1 0 712 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1387
timestamp 1569533753
transform 1 0 840 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1388
timestamp 1569533753
transform 1 0 776 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1389
timestamp 1569533753
transform 1 0 776 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1390
timestamp 1569533753
transform 1 0 776 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1391
timestamp 1569533753
transform 1 0 776 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1392
timestamp 1569533753
transform 1 0 904 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1393
timestamp 1569533753
transform 1 0 776 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1394
timestamp 1569533753
transform 1 0 840 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1395
timestamp 1569533753
transform 1 0 904 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1396
timestamp 1569533753
transform 1 0 776 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1397
timestamp 1569533753
transform 1 0 840 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1398
timestamp 1569533753
transform 1 0 712 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1399
timestamp 1569533753
transform 1 0 840 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1400
timestamp 1569533753
transform 1 0 776 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1401
timestamp 1569533753
transform 1 0 712 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1402
timestamp 1569533753
transform 1 0 904 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1403
timestamp 1569533753
transform 1 0 840 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1404
timestamp 1569533753
transform 1 0 712 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1405
timestamp 1569533753
transform 1 0 904 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1406
timestamp 1569533753
transform 1 0 712 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1407
timestamp 1569533753
transform 1 0 840 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1408
timestamp 1569533753
transform 1 0 712 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1409
timestamp 1569533753
transform 1 0 776 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1410
timestamp 1569533753
transform 1 0 904 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1411
timestamp 1569533753
transform 1 0 1224 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1412
timestamp 1569533753
transform 1 0 1096 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1413
timestamp 1569533753
transform 1 0 1096 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1414
timestamp 1569533753
transform 1 0 1224 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1415
timestamp 1569533753
transform 1 0 1096 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1416
timestamp 1569533753
transform 1 0 1096 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1417
timestamp 1569533753
transform 1 0 1224 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1418
timestamp 1569533753
transform 1 0 1224 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1419
timestamp 1569533753
transform 1 0 1096 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1420
timestamp 1569533753
transform 1 0 1032 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1421
timestamp 1569533753
transform 1 0 1160 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1422
timestamp 1569533753
transform 1 0 968 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1423
timestamp 1569533753
transform 1 0 1032 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1424
timestamp 1569533753
transform 1 0 1160 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1425
timestamp 1569533753
transform 1 0 968 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1426
timestamp 1569533753
transform 1 0 1160 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1427
timestamp 1569533753
transform 1 0 1032 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1428
timestamp 1569533753
transform 1 0 1160 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1429
timestamp 1569533753
transform 1 0 968 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1430
timestamp 1569533753
transform 1 0 1160 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1431
timestamp 1569533753
transform 1 0 968 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1432
timestamp 1569533753
transform 1 0 1224 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1433
timestamp 1569533753
transform 1 0 968 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1434
timestamp 1569533753
transform 1 0 1032 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1435
timestamp 1569533753
transform 1 0 1032 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1436
timestamp 1569533753
transform 1 0 392 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1437
timestamp 1569533753
transform 1 0 584 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1438
timestamp 1569533753
transform 1 0 520 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1439
timestamp 1569533753
transform 1 0 520 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1440
timestamp 1569533753
transform 1 0 392 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1441
timestamp 1569533753
transform 1 0 456 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1442
timestamp 1569533753
transform 1 0 584 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1443
timestamp 1569533753
transform 1 0 520 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1444
timestamp 1569533753
transform 1 0 456 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1445
timestamp 1569533753
transform 1 0 520 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1446
timestamp 1569533753
transform 1 0 456 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1447
timestamp 1569533753
transform 1 0 584 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1448
timestamp 1569533753
transform 1 0 584 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1449
timestamp 1569533753
transform 1 0 584 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1450
timestamp 1569533753
transform 1 0 392 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1451
timestamp 1569533753
transform 1 0 456 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1452
timestamp 1569533753
transform 1 0 520 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1453
timestamp 1569533753
transform 1 0 328 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1454
timestamp 1569533753
transform 1 0 264 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1455
timestamp 1569533753
transform 1 0 328 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1456
timestamp 1569533753
transform 1 0 328 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1457
timestamp 1569533753
transform 1 0 200 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1458
timestamp 1569533753
transform 1 0 136 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1459
timestamp 1569533753
transform 1 0 264 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1460
timestamp 1569533753
transform 1 0 200 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1461
timestamp 1569533753
transform 1 0 72 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1462
timestamp 1569533753
transform 1 0 72 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1463
timestamp 1569533753
transform 1 0 200 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1464
timestamp 1569533753
transform 1 0 136 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1465
timestamp 1569533753
transform 1 0 328 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1466
timestamp 1569533753
transform 1 0 72 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1467
timestamp 1569533753
transform 1 0 200 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1468
timestamp 1569533753
transform 1 0 328 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1469
timestamp 1569533753
transform 1 0 264 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1470
timestamp 1569533753
transform 1 0 136 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1471
timestamp 1569533753
transform 1 0 264 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1472
timestamp 1569533753
transform 1 0 328 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1473
timestamp 1569533753
transform 1 0 328 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1474
timestamp 1569533753
transform 1 0 264 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1475
timestamp 1569533753
transform 1 0 136 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1476
timestamp 1569533753
transform 1 0 264 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1477
timestamp 1569533753
transform 1 0 200 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1478
timestamp 1569533753
transform 1 0 456 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1479
timestamp 1569533753
transform 1 0 584 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1480
timestamp 1569533753
transform 1 0 456 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1481
timestamp 1569533753
transform 1 0 456 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1482
timestamp 1569533753
transform 1 0 456 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1483
timestamp 1569533753
transform 1 0 584 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1484
timestamp 1569533753
transform 1 0 456 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1485
timestamp 1569533753
transform 1 0 392 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1486
timestamp 1569533753
transform 1 0 392 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1487
timestamp 1569533753
transform 1 0 520 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1488
timestamp 1569533753
transform 1 0 584 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1489
timestamp 1569533753
transform 1 0 520 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1490
timestamp 1569533753
transform 1 0 520 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1491
timestamp 1569533753
transform 1 0 392 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1492
timestamp 1569533753
transform 1 0 520 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1493
timestamp 1569533753
transform 1 0 520 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1494
timestamp 1569533753
transform 1 0 392 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1495
timestamp 1569533753
transform 1 0 584 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1496
timestamp 1569533753
transform 1 0 584 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1497
timestamp 1569533753
transform 1 0 392 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1498
timestamp 1569533753
transform 1 0 392 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1499
timestamp 1569533753
transform 1 0 392 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1500
timestamp 1569533753
transform 1 0 456 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1501
timestamp 1569533753
transform 1 0 520 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1502
timestamp 1569533753
transform 1 0 456 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1503
timestamp 1569533753
transform 1 0 520 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1504
timestamp 1569533753
transform 1 0 456 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1505
timestamp 1569533753
transform 1 0 456 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1506
timestamp 1569533753
transform 1 0 392 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1507
timestamp 1569533753
transform 1 0 584 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1508
timestamp 1569533753
transform 1 0 520 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1509
timestamp 1569533753
transform 1 0 584 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1510
timestamp 1569533753
transform 1 0 520 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1511
timestamp 1569533753
transform 1 0 584 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1512
timestamp 1569533753
transform 1 0 456 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1513
timestamp 1569533753
transform 1 0 392 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1514
timestamp 1569533753
transform 1 0 520 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1515
timestamp 1569533753
transform 1 0 584 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1516
timestamp 1569533753
transform 1 0 392 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1517
timestamp 1569533753
transform 1 0 584 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1518
timestamp 1569533753
transform 1 0 200 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1519
timestamp 1569533753
transform 1 0 200 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1520
timestamp 1569533753
transform 1 0 328 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1521
timestamp 1569533753
transform 1 0 72 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1522
timestamp 1569533753
transform 1 0 136 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1523
timestamp 1569533753
transform 1 0 72 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1524
timestamp 1569533753
transform 1 0 264 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1525
timestamp 1569533753
transform 1 0 200 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1526
timestamp 1569533753
transform 1 0 136 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1527
timestamp 1569533753
transform 1 0 328 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1528
timestamp 1569533753
transform 1 0 328 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1529
timestamp 1569533753
transform 1 0 136 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1530
timestamp 1569533753
transform 1 0 72 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1531
timestamp 1569533753
transform 1 0 136 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1532
timestamp 1569533753
transform 1 0 72 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1533
timestamp 1569533753
transform 1 0 328 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1534
timestamp 1569533753
transform 1 0 264 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1535
timestamp 1569533753
transform 1 0 264 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1536
timestamp 1569533753
transform 1 0 200 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1537
timestamp 1569533753
transform 1 0 72 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1538
timestamp 1569533753
transform 1 0 328 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1539
timestamp 1569533753
transform 1 0 200 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1540
timestamp 1569533753
transform 1 0 264 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1541
timestamp 1569533753
transform 1 0 264 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1542
timestamp 1569533753
transform 1 0 136 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1543
timestamp 1569533753
transform 1 0 136 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1544
timestamp 1569533753
transform 1 0 200 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1545
timestamp 1569533753
transform 1 0 264 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1546
timestamp 1569533753
transform 1 0 72 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1547
timestamp 1569533753
transform 1 0 136 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1548
timestamp 1569533753
transform 1 0 328 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1549
timestamp 1569533753
transform 1 0 264 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1550
timestamp 1569533753
transform 1 0 200 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1551
timestamp 1569533753
transform 1 0 328 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1552
timestamp 1569533753
transform 1 0 72 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1553
timestamp 1569533753
transform 1 0 328 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1554
timestamp 1569533753
transform 1 0 200 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1555
timestamp 1569533753
transform 1 0 136 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1556
timestamp 1569533753
transform 1 0 264 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1557
timestamp 1569533753
transform 1 0 328 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1558
timestamp 1569533753
transform 1 0 264 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1559
timestamp 1569533753
transform 1 0 72 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1560
timestamp 1569533753
transform 1 0 72 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1561
timestamp 1569533753
transform 1 0 136 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1562
timestamp 1569533753
transform 1 0 200 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1563
timestamp 1569533753
transform 1 0 392 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1564
timestamp 1569533753
transform 1 0 456 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1565
timestamp 1569533753
transform 1 0 456 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1566
timestamp 1569533753
transform 1 0 584 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1567
timestamp 1569533753
transform 1 0 456 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1568
timestamp 1569533753
transform 1 0 584 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1569
timestamp 1569533753
transform 1 0 520 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1570
timestamp 1569533753
transform 1 0 456 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1571
timestamp 1569533753
transform 1 0 584 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1572
timestamp 1569533753
transform 1 0 392 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1573
timestamp 1569533753
transform 1 0 584 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1574
timestamp 1569533753
transform 1 0 392 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1575
timestamp 1569533753
transform 1 0 520 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1576
timestamp 1569533753
transform 1 0 392 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1577
timestamp 1569533753
transform 1 0 520 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1578
timestamp 1569533753
transform 1 0 520 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1579
timestamp 1569533753
transform 1 0 968 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1580
timestamp 1569533753
transform 1 0 1096 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1581
timestamp 1569533753
transform 1 0 1096 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1582
timestamp 1569533753
transform 1 0 1096 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1583
timestamp 1569533753
transform 1 0 968 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1584
timestamp 1569533753
transform 1 0 1160 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1585
timestamp 1569533753
transform 1 0 1160 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1586
timestamp 1569533753
transform 1 0 1224 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1587
timestamp 1569533753
transform 1 0 1160 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1588
timestamp 1569533753
transform 1 0 1032 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1589
timestamp 1569533753
transform 1 0 968 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1590
timestamp 1569533753
transform 1 0 1096 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1591
timestamp 1569533753
transform 1 0 1032 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1592
timestamp 1569533753
transform 1 0 1160 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1593
timestamp 1569533753
transform 1 0 1032 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1594
timestamp 1569533753
transform 1 0 968 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1595
timestamp 1569533753
transform 1 0 1224 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1596
timestamp 1569533753
transform 1 0 1096 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1597
timestamp 1569533753
transform 1 0 1032 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1598
timestamp 1569533753
transform 1 0 1224 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1599
timestamp 1569533753
transform 1 0 1160 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1600
timestamp 1569533753
transform 1 0 1224 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1601
timestamp 1569533753
transform 1 0 1224 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1602
timestamp 1569533753
transform 1 0 968 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1603
timestamp 1569533753
transform 1 0 1032 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1604
timestamp 1569533753
transform 1 0 840 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1605
timestamp 1569533753
transform 1 0 776 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1606
timestamp 1569533753
transform 1 0 840 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1607
timestamp 1569533753
transform 1 0 776 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1608
timestamp 1569533753
transform 1 0 712 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1609
timestamp 1569533753
transform 1 0 712 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1610
timestamp 1569533753
transform 1 0 840 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1611
timestamp 1569533753
transform 1 0 712 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1612
timestamp 1569533753
transform 1 0 712 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1613
timestamp 1569533753
transform 1 0 904 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1614
timestamp 1569533753
transform 1 0 776 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1615
timestamp 1569533753
transform 1 0 712 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1616
timestamp 1569533753
transform 1 0 776 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1617
timestamp 1569533753
transform 1 0 904 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1618
timestamp 1569533753
transform 1 0 776 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1619
timestamp 1569533753
transform 1 0 840 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1620
timestamp 1569533753
transform 1 0 904 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1621
timestamp 1569533753
transform 1 0 904 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1622
timestamp 1569533753
transform 1 0 840 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1623
timestamp 1569533753
transform 1 0 904 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1624
timestamp 1569533753
transform 1 0 904 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1625
timestamp 1569533753
transform 1 0 776 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1626
timestamp 1569533753
transform 1 0 840 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1627
timestamp 1569533753
transform 1 0 840 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1628
timestamp 1569533753
transform 1 0 840 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1629
timestamp 1569533753
transform 1 0 776 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1630
timestamp 1569533753
transform 1 0 712 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1631
timestamp 1569533753
transform 1 0 904 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1632
timestamp 1569533753
transform 1 0 840 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1633
timestamp 1569533753
transform 1 0 776 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1634
timestamp 1569533753
transform 1 0 904 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1635
timestamp 1569533753
transform 1 0 712 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1636
timestamp 1569533753
transform 1 0 904 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1637
timestamp 1569533753
transform 1 0 712 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1638
timestamp 1569533753
transform 1 0 712 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1639
timestamp 1569533753
transform 1 0 776 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1640
timestamp 1569533753
transform 1 0 1224 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1641
timestamp 1569533753
transform 1 0 968 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1642
timestamp 1569533753
transform 1 0 1160 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1643
timestamp 1569533753
transform 1 0 1032 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1644
timestamp 1569533753
transform 1 0 1224 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1645
timestamp 1569533753
transform 1 0 968 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1646
timestamp 1569533753
transform 1 0 1096 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1647
timestamp 1569533753
transform 1 0 1032 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1648
timestamp 1569533753
transform 1 0 1096 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1649
timestamp 1569533753
transform 1 0 1032 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1650
timestamp 1569533753
transform 1 0 1032 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1651
timestamp 1569533753
transform 1 0 1096 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1652
timestamp 1569533753
transform 1 0 1096 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1653
timestamp 1569533753
transform 1 0 1160 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1654
timestamp 1569533753
transform 1 0 1160 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1655
timestamp 1569533753
transform 1 0 1160 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1656
timestamp 1569533753
transform 1 0 1224 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1657
timestamp 1569533753
transform 1 0 968 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1658
timestamp 1569533753
transform 1 0 1224 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1659
timestamp 1569533753
transform 1 0 968 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1660
timestamp 1569533753
transform 1 0 648 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1661
timestamp 1569533753
transform 1 0 648 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1662
timestamp 1569533753
transform 1 0 648 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1663
timestamp 1569533753
transform 1 0 648 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1664
timestamp 1569533753
transform 1 0 648 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1665
timestamp 1569533753
transform 1 0 648 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1666
timestamp 1569533753
transform 1 0 648 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1667
timestamp 1569533753
transform 1 0 648 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1668
timestamp 1569533753
transform 1 0 648 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1669
timestamp 1569533753
transform 1 0 648 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1670
timestamp 1569533753
transform 1 0 648 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1671
timestamp 1569533753
transform 1 0 648 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1672
timestamp 1569533753
transform 1 0 648 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1673
timestamp 1569533753
transform 1 0 648 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1674
timestamp 1569533753
transform 1 0 648 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1675
timestamp 1569533753
transform 1 0 648 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1676
timestamp 1569533753
transform 1 0 648 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1677
timestamp 1569533753
transform 1 0 648 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1678
timestamp 1569533753
transform 1 0 648 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1679
timestamp 1569533753
transform 1 0 2248 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1680
timestamp 1569533753
transform 1 0 2376 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1681
timestamp 1569533753
transform 1 0 2376 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1682
timestamp 1569533753
transform 1 0 2312 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1683
timestamp 1569533753
transform 1 0 2248 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1684
timestamp 1569533753
transform 1 0 2440 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1685
timestamp 1569533753
transform 1 0 2248 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1686
timestamp 1569533753
transform 1 0 2312 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1687
timestamp 1569533753
transform 1 0 2248 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1688
timestamp 1569533753
transform 1 0 2440 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1689
timestamp 1569533753
transform 1 0 2312 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1690
timestamp 1569533753
transform 1 0 2376 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1691
timestamp 1569533753
transform 1 0 2440 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1692
timestamp 1569533753
transform 1 0 2312 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1693
timestamp 1569533753
transform 1 0 2376 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1694
timestamp 1569533753
transform 1 0 2440 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1695
timestamp 1569533753
transform 1 0 2376 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1696
timestamp 1569533753
transform 1 0 2248 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1697
timestamp 1569533753
transform 1 0 2312 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1698
timestamp 1569533753
transform 1 0 2440 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1699
timestamp 1569533753
transform 1 0 2056 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1700
timestamp 1569533753
transform 1 0 1928 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1701
timestamp 1569533753
transform 1 0 2056 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1702
timestamp 1569533753
transform 1 0 2056 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1703
timestamp 1569533753
transform 1 0 2056 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1704
timestamp 1569533753
transform 1 0 1928 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1705
timestamp 1569533753
transform 1 0 2120 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1706
timestamp 1569533753
transform 1 0 2120 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1707
timestamp 1569533753
transform 1 0 2184 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1708
timestamp 1569533753
transform 1 0 2120 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1709
timestamp 1569533753
transform 1 0 1992 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1710
timestamp 1569533753
transform 1 0 2120 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1711
timestamp 1569533753
transform 1 0 2120 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1712
timestamp 1569533753
transform 1 0 2184 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1713
timestamp 1569533753
transform 1 0 2184 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1714
timestamp 1569533753
transform 1 0 2056 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1715
timestamp 1569533753
transform 1 0 2184 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1716
timestamp 1569533753
transform 1 0 2184 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1717
timestamp 1569533753
transform 1 0 1928 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1718
timestamp 1569533753
transform 1 0 1992 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1719
timestamp 1569533753
transform 1 0 1992 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1720
timestamp 1569533753
transform 1 0 1928 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1721
timestamp 1569533753
transform 1 0 1928 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1722
timestamp 1569533753
transform 1 0 1992 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1723
timestamp 1569533753
transform 1 0 1992 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1724
timestamp 1569533753
transform 1 0 2056 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1725
timestamp 1569533753
transform 1 0 2184 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1726
timestamp 1569533753
transform 1 0 2056 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1727
timestamp 1569533753
transform 1 0 2056 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1728
timestamp 1569533753
transform 1 0 1928 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1729
timestamp 1569533753
transform 1 0 2056 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1730
timestamp 1569533753
transform 1 0 2056 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1731
timestamp 1569533753
transform 1 0 2184 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1732
timestamp 1569533753
transform 1 0 2184 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1733
timestamp 1569533753
transform 1 0 2184 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1734
timestamp 1569533753
transform 1 0 2184 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1735
timestamp 1569533753
transform 1 0 2120 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1736
timestamp 1569533753
transform 1 0 1992 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1737
timestamp 1569533753
transform 1 0 2120 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1738
timestamp 1569533753
transform 1 0 2120 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1739
timestamp 1569533753
transform 1 0 1928 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1740
timestamp 1569533753
transform 1 0 2120 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1741
timestamp 1569533753
transform 1 0 2120 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1742
timestamp 1569533753
transform 1 0 1928 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1743
timestamp 1569533753
transform 1 0 1928 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1744
timestamp 1569533753
transform 1 0 1928 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1745
timestamp 1569533753
transform 1 0 1992 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1746
timestamp 1569533753
transform 1 0 1992 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1747
timestamp 1569533753
transform 1 0 1992 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1748
timestamp 1569533753
transform 1 0 1992 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1749
timestamp 1569533753
transform 1 0 2376 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1750
timestamp 1569533753
transform 1 0 2440 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1751
timestamp 1569533753
transform 1 0 2440 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1752
timestamp 1569533753
transform 1 0 2376 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1753
timestamp 1569533753
transform 1 0 2440 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1754
timestamp 1569533753
transform 1 0 2440 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1755
timestamp 1569533753
transform 1 0 2440 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1756
timestamp 1569533753
transform 1 0 2312 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1757
timestamp 1569533753
transform 1 0 2248 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1758
timestamp 1569533753
transform 1 0 2248 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1759
timestamp 1569533753
transform 1 0 2312 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1760
timestamp 1569533753
transform 1 0 2248 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1761
timestamp 1569533753
transform 1 0 2248 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1762
timestamp 1569533753
transform 1 0 2312 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1763
timestamp 1569533753
transform 1 0 2248 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1764
timestamp 1569533753
transform 1 0 2312 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1765
timestamp 1569533753
transform 1 0 2312 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1766
timestamp 1569533753
transform 1 0 2376 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1767
timestamp 1569533753
transform 1 0 2376 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1768
timestamp 1569533753
transform 1 0 2376 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1769
timestamp 1569533753
transform 1 0 1672 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1770
timestamp 1569533753
transform 1 0 1672 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1771
timestamp 1569533753
transform 1 0 1608 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1772
timestamp 1569533753
transform 1 0 1608 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1773
timestamp 1569533753
transform 1 0 1800 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1774
timestamp 1569533753
transform 1 0 1800 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1775
timestamp 1569533753
transform 1 0 1672 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1776
timestamp 1569533753
transform 1 0 1672 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1777
timestamp 1569533753
transform 1 0 1672 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1778
timestamp 1569533753
transform 1 0 1736 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1779
timestamp 1569533753
transform 1 0 1864 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1780
timestamp 1569533753
transform 1 0 1736 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1781
timestamp 1569533753
transform 1 0 1736 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1782
timestamp 1569533753
transform 1 0 1800 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1783
timestamp 1569533753
transform 1 0 1800 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1784
timestamp 1569533753
transform 1 0 1800 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1785
timestamp 1569533753
transform 1 0 1736 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1786
timestamp 1569533753
transform 1 0 1736 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1787
timestamp 1569533753
transform 1 0 1864 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1788
timestamp 1569533753
transform 1 0 1864 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1789
timestamp 1569533753
transform 1 0 1864 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1790
timestamp 1569533753
transform 1 0 1864 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1791
timestamp 1569533753
transform 1 0 1608 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1792
timestamp 1569533753
transform 1 0 1608 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1793
timestamp 1569533753
transform 1 0 1608 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1794
timestamp 1569533753
transform 1 0 1544 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1795
timestamp 1569533753
transform 1 0 1544 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1796
timestamp 1569533753
transform 1 0 1288 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1797
timestamp 1569533753
transform 1 0 1288 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1798
timestamp 1569533753
transform 1 0 1288 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1799
timestamp 1569533753
transform 1 0 1288 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1800
timestamp 1569533753
transform 1 0 1288 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1801
timestamp 1569533753
transform 1 0 1480 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1802
timestamp 1569533753
transform 1 0 1416 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1803
timestamp 1569533753
transform 1 0 1416 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1804
timestamp 1569533753
transform 1 0 1480 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1805
timestamp 1569533753
transform 1 0 1352 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1806
timestamp 1569533753
transform 1 0 1352 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1807
timestamp 1569533753
transform 1 0 1352 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1808
timestamp 1569533753
transform 1 0 1416 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1809
timestamp 1569533753
transform 1 0 1416 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1810
timestamp 1569533753
transform 1 0 1416 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1811
timestamp 1569533753
transform 1 0 1480 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1812
timestamp 1569533753
transform 1 0 1480 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1813
timestamp 1569533753
transform 1 0 1480 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1814
timestamp 1569533753
transform 1 0 1544 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_1815
timestamp 1569533753
transform 1 0 1544 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_1816
timestamp 1569533753
transform 1 0 1544 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_1817
timestamp 1569533753
transform 1 0 1352 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_1818
timestamp 1569533753
transform 1 0 1352 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_1819
timestamp 1569533753
transform 1 0 1544 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1820
timestamp 1569533753
transform 1 0 1352 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1821
timestamp 1569533753
transform 1 0 1352 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1822
timestamp 1569533753
transform 1 0 1352 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1823
timestamp 1569533753
transform 1 0 1352 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1824
timestamp 1569533753
transform 1 0 1352 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1825
timestamp 1569533753
transform 1 0 1544 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1826
timestamp 1569533753
transform 1 0 1544 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1827
timestamp 1569533753
transform 1 0 1544 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1828
timestamp 1569533753
transform 1 0 1416 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1829
timestamp 1569533753
transform 1 0 1416 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1830
timestamp 1569533753
transform 1 0 1288 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1831
timestamp 1569533753
transform 1 0 1416 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1832
timestamp 1569533753
transform 1 0 1416 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1833
timestamp 1569533753
transform 1 0 1416 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1834
timestamp 1569533753
transform 1 0 1288 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1835
timestamp 1569533753
transform 1 0 1288 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1836
timestamp 1569533753
transform 1 0 1480 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1837
timestamp 1569533753
transform 1 0 1480 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1838
timestamp 1569533753
transform 1 0 1480 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1839
timestamp 1569533753
transform 1 0 1480 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1840
timestamp 1569533753
transform 1 0 1480 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1841
timestamp 1569533753
transform 1 0 1288 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1842
timestamp 1569533753
transform 1 0 1288 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1843
timestamp 1569533753
transform 1 0 1544 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1844
timestamp 1569533753
transform 1 0 1800 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1845
timestamp 1569533753
transform 1 0 1800 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1846
timestamp 1569533753
transform 1 0 1608 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1847
timestamp 1569533753
transform 1 0 1608 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1848
timestamp 1569533753
transform 1 0 1608 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1849
timestamp 1569533753
transform 1 0 1608 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1850
timestamp 1569533753
transform 1 0 1608 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1851
timestamp 1569533753
transform 1 0 1800 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1852
timestamp 1569533753
transform 1 0 1800 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1853
timestamp 1569533753
transform 1 0 1864 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1854
timestamp 1569533753
transform 1 0 1864 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1855
timestamp 1569533753
transform 1 0 1864 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1856
timestamp 1569533753
transform 1 0 1672 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1857
timestamp 1569533753
transform 1 0 1672 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1858
timestamp 1569533753
transform 1 0 1672 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1859
timestamp 1569533753
transform 1 0 1672 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1860
timestamp 1569533753
transform 1 0 1672 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1861
timestamp 1569533753
transform 1 0 1864 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1862
timestamp 1569533753
transform 1 0 1736 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1863
timestamp 1569533753
transform 1 0 1736 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_1864
timestamp 1569533753
transform 1 0 1736 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_1865
timestamp 1569533753
transform 1 0 1736 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1866
timestamp 1569533753
transform 1 0 1736 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_1867
timestamp 1569533753
transform 1 0 1864 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_1868
timestamp 1569533753
transform 1 0 1800 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_1869
timestamp 1569533753
transform 1 0 1800 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1870
timestamp 1569533753
transform 1 0 1608 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1871
timestamp 1569533753
transform 1 0 1864 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1872
timestamp 1569533753
transform 1 0 1608 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1873
timestamp 1569533753
transform 1 0 1800 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1874
timestamp 1569533753
transform 1 0 1672 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1875
timestamp 1569533753
transform 1 0 1864 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1876
timestamp 1569533753
transform 1 0 1672 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1877
timestamp 1569533753
transform 1 0 1864 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1878
timestamp 1569533753
transform 1 0 1672 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1879
timestamp 1569533753
transform 1 0 1864 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1880
timestamp 1569533753
transform 1 0 1672 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1881
timestamp 1569533753
transform 1 0 1672 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1882
timestamp 1569533753
transform 1 0 1736 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1883
timestamp 1569533753
transform 1 0 1800 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1884
timestamp 1569533753
transform 1 0 1736 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1885
timestamp 1569533753
transform 1 0 1736 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1886
timestamp 1569533753
transform 1 0 1608 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1887
timestamp 1569533753
transform 1 0 1736 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1888
timestamp 1569533753
transform 1 0 1608 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1889
timestamp 1569533753
transform 1 0 1736 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1890
timestamp 1569533753
transform 1 0 1608 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1891
timestamp 1569533753
transform 1 0 1864 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1892
timestamp 1569533753
transform 1 0 1800 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1893
timestamp 1569533753
transform 1 0 1800 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1894
timestamp 1569533753
transform 1 0 1352 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1895
timestamp 1569533753
transform 1 0 1480 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1896
timestamp 1569533753
transform 1 0 1480 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1897
timestamp 1569533753
transform 1 0 1544 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1898
timestamp 1569533753
transform 1 0 1544 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1899
timestamp 1569533753
transform 1 0 1416 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1900
timestamp 1569533753
transform 1 0 1288 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1901
timestamp 1569533753
transform 1 0 1544 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1902
timestamp 1569533753
transform 1 0 1416 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1903
timestamp 1569533753
transform 1 0 1544 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1904
timestamp 1569533753
transform 1 0 1288 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1905
timestamp 1569533753
transform 1 0 1544 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1906
timestamp 1569533753
transform 1 0 1480 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1907
timestamp 1569533753
transform 1 0 1288 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1908
timestamp 1569533753
transform 1 0 1480 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1909
timestamp 1569533753
transform 1 0 1288 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1910
timestamp 1569533753
transform 1 0 1352 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1911
timestamp 1569533753
transform 1 0 1352 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1912
timestamp 1569533753
transform 1 0 1352 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1913
timestamp 1569533753
transform 1 0 1288 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1914
timestamp 1569533753
transform 1 0 1352 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1915
timestamp 1569533753
transform 1 0 1416 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1916
timestamp 1569533753
transform 1 0 1416 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1917
timestamp 1569533753
transform 1 0 1416 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1918
timestamp 1569533753
transform 1 0 1480 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1919
timestamp 1569533753
transform 1 0 1352 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1920
timestamp 1569533753
transform 1 0 1288 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1921
timestamp 1569533753
transform 1 0 1544 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1922
timestamp 1569533753
transform 1 0 1352 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1923
timestamp 1569533753
transform 1 0 1288 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1924
timestamp 1569533753
transform 1 0 1416 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1925
timestamp 1569533753
transform 1 0 1416 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1926
timestamp 1569533753
transform 1 0 1480 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1927
timestamp 1569533753
transform 1 0 1480 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1928
timestamp 1569533753
transform 1 0 1480 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1929
timestamp 1569533753
transform 1 0 1352 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1930
timestamp 1569533753
transform 1 0 1480 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1931
timestamp 1569533753
transform 1 0 1544 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1932
timestamp 1569533753
transform 1 0 1416 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1933
timestamp 1569533753
transform 1 0 1544 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1934
timestamp 1569533753
transform 1 0 1288 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1935
timestamp 1569533753
transform 1 0 1544 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1936
timestamp 1569533753
transform 1 0 1416 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1937
timestamp 1569533753
transform 1 0 1288 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1938
timestamp 1569533753
transform 1 0 1352 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1939
timestamp 1569533753
transform 1 0 1608 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1940
timestamp 1569533753
transform 1 0 1864 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1941
timestamp 1569533753
transform 1 0 1608 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1942
timestamp 1569533753
transform 1 0 1672 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1943
timestamp 1569533753
transform 1 0 1672 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1944
timestamp 1569533753
transform 1 0 1672 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1945
timestamp 1569533753
transform 1 0 1736 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1946
timestamp 1569533753
transform 1 0 1736 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1947
timestamp 1569533753
transform 1 0 1800 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1948
timestamp 1569533753
transform 1 0 1736 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1949
timestamp 1569533753
transform 1 0 1800 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1950
timestamp 1569533753
transform 1 0 1864 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1951
timestamp 1569533753
transform 1 0 1800 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1952
timestamp 1569533753
transform 1 0 1608 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1953
timestamp 1569533753
transform 1 0 1800 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1954
timestamp 1569533753
transform 1 0 1864 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_1955
timestamp 1569533753
transform 1 0 1608 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1956
timestamp 1569533753
transform 1 0 1864 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_1957
timestamp 1569533753
transform 1 0 1672 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1958
timestamp 1569533753
transform 1 0 1736 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_1959
timestamp 1569533753
transform 1 0 2376 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1960
timestamp 1569533753
transform 1 0 2376 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1961
timestamp 1569533753
transform 1 0 2248 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1962
timestamp 1569533753
transform 1 0 2440 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1963
timestamp 1569533753
transform 1 0 2440 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1964
timestamp 1569533753
transform 1 0 2312 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1965
timestamp 1569533753
transform 1 0 2376 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1966
timestamp 1569533753
transform 1 0 2248 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1967
timestamp 1569533753
transform 1 0 2248 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1968
timestamp 1569533753
transform 1 0 2312 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1969
timestamp 1569533753
transform 1 0 2312 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1970
timestamp 1569533753
transform 1 0 2248 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1971
timestamp 1569533753
transform 1 0 2248 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1972
timestamp 1569533753
transform 1 0 2312 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1973
timestamp 1569533753
transform 1 0 1992 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1974
timestamp 1569533753
transform 1 0 1992 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1975
timestamp 1569533753
transform 1 0 1928 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1976
timestamp 1569533753
transform 1 0 2056 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1977
timestamp 1569533753
transform 1 0 2056 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1978
timestamp 1569533753
transform 1 0 1992 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1979
timestamp 1569533753
transform 1 0 2120 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1980
timestamp 1569533753
transform 1 0 2120 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1981
timestamp 1569533753
transform 1 0 2056 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1982
timestamp 1569533753
transform 1 0 2184 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1983
timestamp 1569533753
transform 1 0 2184 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1984
timestamp 1569533753
transform 1 0 2120 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1985
timestamp 1569533753
transform 1 0 2056 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1986
timestamp 1569533753
transform 1 0 2056 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1987
timestamp 1569533753
transform 1 0 2120 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1988
timestamp 1569533753
transform 1 0 2120 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1989
timestamp 1569533753
transform 1 0 2184 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1990
timestamp 1569533753
transform 1 0 1928 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1991
timestamp 1569533753
transform 1 0 2184 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1992
timestamp 1569533753
transform 1 0 1992 0 1 2184
box -8 -8 8 8
use VIA1$3  VIA1$3_1993
timestamp 1569533753
transform 1 0 2184 0 1 2056
box -8 -8 8 8
use VIA1$3  VIA1$3_1994
timestamp 1569533753
transform 1 0 1928 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_1995
timestamp 1569533753
transform 1 0 1928 0 1 1992
box -8 -8 8 8
use VIA1$3  VIA1$3_1996
timestamp 1569533753
transform 1 0 1928 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1997
timestamp 1569533753
transform 1 0 1992 0 1 2120
box -8 -8 8 8
use VIA1$3  VIA1$3_1998
timestamp 1569533753
transform 1 0 2056 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_1999
timestamp 1569533753
transform 1 0 1928 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_2000
timestamp 1569533753
transform 1 0 1928 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_2001
timestamp 1569533753
transform 1 0 1992 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_2002
timestamp 1569533753
transform 1 0 1992 0 1 2440
box -8 -8 8 8
use VIA1$3  VIA1$3_2003
timestamp 1569533753
transform 1 0 2184 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_2004
timestamp 1569533753
transform 1 0 1928 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_2005
timestamp 1569533753
transform 1 0 2056 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_2006
timestamp 1569533753
transform 1 0 1992 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_2007
timestamp 1569533753
transform 1 0 2120 0 1 2248
box -8 -8 8 8
use VIA1$3  VIA1$3_2008
timestamp 1569533753
transform 1 0 2056 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_2009
timestamp 1569533753
transform 1 0 2120 0 1 2312
box -8 -8 8 8
use VIA1$3  VIA1$3_2010
timestamp 1569533753
transform 1 0 1928 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_2011
timestamp 1569533753
transform 1 0 1992 0 1 2376
box -8 -8 8 8
use VIA1$3  VIA1$3_2012
timestamp 1569533753
transform 1 0 1864 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2013
timestamp 1569533753
transform 1 0 1672 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2014
timestamp 1569533753
transform 1 0 1672 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2015
timestamp 1569533753
transform 1 0 1608 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2016
timestamp 1569533753
transform 1 0 1736 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2017
timestamp 1569533753
transform 1 0 1608 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2018
timestamp 1569533753
transform 1 0 1800 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2019
timestamp 1569533753
transform 1 0 1672 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2020
timestamp 1569533753
transform 1 0 1800 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2021
timestamp 1569533753
transform 1 0 1672 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2022
timestamp 1569533753
transform 1 0 1736 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2023
timestamp 1569533753
transform 1 0 1608 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2024
timestamp 1569533753
transform 1 0 1608 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2025
timestamp 1569533753
transform 1 0 1480 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2026
timestamp 1569533753
transform 1 0 1416 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2027
timestamp 1569533753
transform 1 0 1352 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2028
timestamp 1569533753
transform 1 0 1416 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2029
timestamp 1569533753
transform 1 0 1416 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2030
timestamp 1569533753
transform 1 0 1416 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2031
timestamp 1569533753
transform 1 0 1352 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2032
timestamp 1569533753
transform 1 0 1352 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2033
timestamp 1569533753
transform 1 0 1288 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2034
timestamp 1569533753
transform 1 0 1544 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2035
timestamp 1569533753
transform 1 0 1288 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2036
timestamp 1569533753
transform 1 0 1544 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2037
timestamp 1569533753
transform 1 0 1288 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2038
timestamp 1569533753
transform 1 0 1352 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2039
timestamp 1569533753
transform 1 0 1480 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2040
timestamp 1569533753
transform 1 0 1544 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2041
timestamp 1569533753
transform 1 0 1480 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2042
timestamp 1569533753
transform 1 0 1544 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2043
timestamp 1569533753
transform 1 0 1480 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2044
timestamp 1569533753
transform 1 0 1288 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2045
timestamp 1569533753
transform 1 0 1288 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2046
timestamp 1569533753
transform 1 0 1288 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2047
timestamp 1569533753
transform 1 0 1288 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2048
timestamp 1569533753
transform 1 0 1544 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2049
timestamp 1569533753
transform 1 0 1544 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2050
timestamp 1569533753
transform 1 0 1416 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2051
timestamp 1569533753
transform 1 0 1288 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2052
timestamp 1569533753
transform 1 0 1416 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2053
timestamp 1569533753
transform 1 0 1352 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2054
timestamp 1569533753
transform 1 0 1352 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2055
timestamp 1569533753
transform 1 0 1416 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2056
timestamp 1569533753
transform 1 0 1480 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2057
timestamp 1569533753
transform 1 0 1288 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2058
timestamp 1569533753
transform 1 0 1416 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2059
timestamp 1569533753
transform 1 0 1480 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2060
timestamp 1569533753
transform 1 0 1352 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2061
timestamp 1569533753
transform 1 0 1480 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2062
timestamp 1569533753
transform 1 0 1352 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2063
timestamp 1569533753
transform 1 0 1416 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2064
timestamp 1569533753
transform 1 0 1352 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2065
timestamp 1569533753
transform 1 0 1480 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2066
timestamp 1569533753
transform 1 0 1480 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2067
timestamp 1569533753
transform 1 0 1608 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2068
timestamp 1569533753
transform 1 0 1480 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2069
timestamp 1569533753
transform 1 0 1480 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2070
timestamp 1569533753
transform 1 0 1480 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2071
timestamp 1569533753
transform 1 0 1352 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2072
timestamp 1569533753
transform 1 0 1288 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2073
timestamp 1569533753
transform 1 0 1480 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2074
timestamp 1569533753
transform 1 0 1480 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2075
timestamp 1569533753
transform 1 0 1352 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2076
timestamp 1569533753
transform 1 0 1416 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2077
timestamp 1569533753
transform 1 0 1480 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2078
timestamp 1569533753
transform 1 0 1288 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2079
timestamp 1569533753
transform 1 0 1288 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2080
timestamp 1569533753
transform 1 0 1416 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2081
timestamp 1569533753
transform 1 0 1480 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2082
timestamp 1569533753
transform 1 0 1480 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2083
timestamp 1569533753
transform 1 0 1352 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2084
timestamp 1569533753
transform 1 0 1352 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2085
timestamp 1569533753
transform 1 0 1352 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2086
timestamp 1569533753
transform 1 0 1288 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2087
timestamp 1569533753
transform 1 0 1288 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2088
timestamp 1569533753
transform 1 0 1352 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2089
timestamp 1569533753
transform 1 0 1352 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2090
timestamp 1569533753
transform 1 0 1288 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2091
timestamp 1569533753
transform 1 0 1416 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2092
timestamp 1569533753
transform 1 0 1352 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2093
timestamp 1569533753
transform 1 0 1416 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2094
timestamp 1569533753
transform 1 0 1480 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2095
timestamp 1569533753
transform 1 0 1288 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2096
timestamp 1569533753
transform 1 0 1416 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2097
timestamp 1569533753
transform 1 0 1416 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2098
timestamp 1569533753
transform 1 0 1352 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2099
timestamp 1569533753
transform 1 0 1288 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2100
timestamp 1569533753
transform 1 0 1352 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2101
timestamp 1569533753
transform 1 0 1416 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2102
timestamp 1569533753
transform 1 0 1480 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2103
timestamp 1569533753
transform 1 0 1288 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2104
timestamp 1569533753
transform 1 0 1416 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2105
timestamp 1569533753
transform 1 0 1416 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2106
timestamp 1569533753
transform 1 0 1288 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2107
timestamp 1569533753
transform 1 0 1416 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2108
timestamp 1569533753
transform 1 0 2440 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2109
timestamp 1569533753
transform 1 0 2440 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2110
timestamp 1569533753
transform 1 0 2440 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2111
timestamp 1569533753
transform 1 0 2376 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2112
timestamp 1569533753
transform 1 0 2376 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2113
timestamp 1569533753
transform 1 0 2440 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2114
timestamp 1569533753
transform 1 0 2376 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2115
timestamp 1569533753
transform 1 0 2312 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2116
timestamp 1569533753
transform 1 0 2376 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2117
timestamp 1569533753
transform 1 0 2440 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2118
timestamp 1569533753
transform 1 0 2376 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2119
timestamp 1569533753
transform 1 0 2376 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2120
timestamp 1569533753
transform 1 0 2376 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2121
timestamp 1569533753
transform 1 0 2312 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2122
timestamp 1569533753
transform 1 0 2312 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2123
timestamp 1569533753
transform 1 0 2312 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2124
timestamp 1569533753
transform 1 0 2312 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2125
timestamp 1569533753
transform 1 0 2312 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2126
timestamp 1569533753
transform 1 0 2440 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2127
timestamp 1569533753
transform 1 0 2440 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2128
timestamp 1569533753
transform 1 0 2440 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2129
timestamp 1569533753
transform 1 0 1096 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2130
timestamp 1569533753
transform 1 0 1160 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2131
timestamp 1569533753
transform 1 0 968 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2132
timestamp 1569533753
transform 1 0 1096 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2133
timestamp 1569533753
transform 1 0 1032 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2134
timestamp 1569533753
transform 1 0 968 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2135
timestamp 1569533753
transform 1 0 1160 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2136
timestamp 1569533753
transform 1 0 1224 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2137
timestamp 1569533753
transform 1 0 1032 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2138
timestamp 1569533753
transform 1 0 1160 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2139
timestamp 1569533753
transform 1 0 1224 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2140
timestamp 1569533753
transform 1 0 1160 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2141
timestamp 1569533753
transform 1 0 968 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2142
timestamp 1569533753
transform 1 0 1096 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2143
timestamp 1569533753
transform 1 0 1032 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2144
timestamp 1569533753
transform 1 0 1096 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2145
timestamp 1569533753
transform 1 0 1032 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2146
timestamp 1569533753
transform 1 0 1224 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2147
timestamp 1569533753
transform 1 0 1224 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2148
timestamp 1569533753
transform 1 0 968 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2149
timestamp 1569533753
transform 1 0 904 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2150
timestamp 1569533753
transform 1 0 904 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2151
timestamp 1569533753
transform 1 0 840 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2152
timestamp 1569533753
transform 1 0 776 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2153
timestamp 1569533753
transform 1 0 840 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2154
timestamp 1569533753
transform 1 0 712 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2155
timestamp 1569533753
transform 1 0 904 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2156
timestamp 1569533753
transform 1 0 712 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2157
timestamp 1569533753
transform 1 0 776 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2158
timestamp 1569533753
transform 1 0 712 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2159
timestamp 1569533753
transform 1 0 776 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2160
timestamp 1569533753
transform 1 0 776 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2161
timestamp 1569533753
transform 1 0 840 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2162
timestamp 1569533753
transform 1 0 904 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2163
timestamp 1569533753
transform 1 0 712 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2164
timestamp 1569533753
transform 1 0 840 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2165
timestamp 1569533753
transform 1 0 840 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2166
timestamp 1569533753
transform 1 0 712 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2167
timestamp 1569533753
transform 1 0 904 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2168
timestamp 1569533753
transform 1 0 776 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2169
timestamp 1569533753
transform 1 0 712 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2170
timestamp 1569533753
transform 1 0 904 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2171
timestamp 1569533753
transform 1 0 904 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2172
timestamp 1569533753
transform 1 0 840 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2173
timestamp 1569533753
transform 1 0 904 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2174
timestamp 1569533753
transform 1 0 840 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2175
timestamp 1569533753
transform 1 0 712 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2176
timestamp 1569533753
transform 1 0 712 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2177
timestamp 1569533753
transform 1 0 776 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2178
timestamp 1569533753
transform 1 0 840 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2179
timestamp 1569533753
transform 1 0 776 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2180
timestamp 1569533753
transform 1 0 840 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2181
timestamp 1569533753
transform 1 0 712 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2182
timestamp 1569533753
transform 1 0 776 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2183
timestamp 1569533753
transform 1 0 776 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2184
timestamp 1569533753
transform 1 0 904 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2185
timestamp 1569533753
transform 1 0 1160 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2186
timestamp 1569533753
transform 1 0 1032 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2187
timestamp 1569533753
transform 1 0 1160 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2188
timestamp 1569533753
transform 1 0 1160 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2189
timestamp 1569533753
transform 1 0 1096 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2190
timestamp 1569533753
transform 1 0 968 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2191
timestamp 1569533753
transform 1 0 1032 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2192
timestamp 1569533753
transform 1 0 1096 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2193
timestamp 1569533753
transform 1 0 1160 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2194
timestamp 1569533753
transform 1 0 968 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2195
timestamp 1569533753
transform 1 0 1224 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2196
timestamp 1569533753
transform 1 0 1224 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2197
timestamp 1569533753
transform 1 0 968 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2198
timestamp 1569533753
transform 1 0 1032 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2199
timestamp 1569533753
transform 1 0 1224 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2200
timestamp 1569533753
transform 1 0 968 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2201
timestamp 1569533753
transform 1 0 1032 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2202
timestamp 1569533753
transform 1 0 1096 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2203
timestamp 1569533753
transform 1 0 1160 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2204
timestamp 1569533753
transform 1 0 1032 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2205
timestamp 1569533753
transform 1 0 968 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2206
timestamp 1569533753
transform 1 0 1096 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2207
timestamp 1569533753
transform 1 0 1224 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2208
timestamp 1569533753
transform 1 0 1096 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2209
timestamp 1569533753
transform 1 0 1224 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2210
timestamp 1569533753
transform 1 0 584 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2211
timestamp 1569533753
transform 1 0 520 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2212
timestamp 1569533753
transform 1 0 392 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2213
timestamp 1569533753
transform 1 0 584 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2214
timestamp 1569533753
transform 1 0 520 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2215
timestamp 1569533753
transform 1 0 392 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2216
timestamp 1569533753
transform 1 0 584 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2217
timestamp 1569533753
transform 1 0 456 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2218
timestamp 1569533753
transform 1 0 392 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2219
timestamp 1569533753
transform 1 0 456 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2220
timestamp 1569533753
transform 1 0 520 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2221
timestamp 1569533753
transform 1 0 520 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2222
timestamp 1569533753
transform 1 0 392 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2223
timestamp 1569533753
transform 1 0 456 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2224
timestamp 1569533753
transform 1 0 456 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2225
timestamp 1569533753
transform 1 0 584 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2226
timestamp 1569533753
transform 1 0 72 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2227
timestamp 1569533753
transform 1 0 328 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2228
timestamp 1569533753
transform 1 0 72 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2229
timestamp 1569533753
transform 1 0 264 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2230
timestamp 1569533753
transform 1 0 264 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2231
timestamp 1569533753
transform 1 0 136 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2232
timestamp 1569533753
transform 1 0 328 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2233
timestamp 1569533753
transform 1 0 200 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2234
timestamp 1569533753
transform 1 0 136 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2235
timestamp 1569533753
transform 1 0 264 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2236
timestamp 1569533753
transform 1 0 328 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2237
timestamp 1569533753
transform 1 0 72 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2238
timestamp 1569533753
transform 1 0 200 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2239
timestamp 1569533753
transform 1 0 72 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2240
timestamp 1569533753
transform 1 0 200 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2241
timestamp 1569533753
transform 1 0 136 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2242
timestamp 1569533753
transform 1 0 264 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2243
timestamp 1569533753
transform 1 0 136 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2244
timestamp 1569533753
transform 1 0 328 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2245
timestamp 1569533753
transform 1 0 200 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2246
timestamp 1569533753
transform 1 0 264 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2247
timestamp 1569533753
transform 1 0 264 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2248
timestamp 1569533753
transform 1 0 136 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2249
timestamp 1569533753
transform 1 0 264 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2250
timestamp 1569533753
transform 1 0 264 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2251
timestamp 1569533753
transform 1 0 200 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2252
timestamp 1569533753
transform 1 0 136 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2253
timestamp 1569533753
transform 1 0 328 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2254
timestamp 1569533753
transform 1 0 136 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2255
timestamp 1569533753
transform 1 0 72 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2256
timestamp 1569533753
transform 1 0 200 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2257
timestamp 1569533753
transform 1 0 136 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2258
timestamp 1569533753
transform 1 0 72 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2259
timestamp 1569533753
transform 1 0 328 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2260
timestamp 1569533753
transform 1 0 328 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2261
timestamp 1569533753
transform 1 0 328 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2262
timestamp 1569533753
transform 1 0 72 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2263
timestamp 1569533753
transform 1 0 328 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2264
timestamp 1569533753
transform 1 0 72 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2265
timestamp 1569533753
transform 1 0 200 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2266
timestamp 1569533753
transform 1 0 200 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2267
timestamp 1569533753
transform 1 0 136 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2268
timestamp 1569533753
transform 1 0 264 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2269
timestamp 1569533753
transform 1 0 200 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2270
timestamp 1569533753
transform 1 0 72 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2271
timestamp 1569533753
transform 1 0 520 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2272
timestamp 1569533753
transform 1 0 392 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2273
timestamp 1569533753
transform 1 0 392 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2274
timestamp 1569533753
transform 1 0 392 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2275
timestamp 1569533753
transform 1 0 520 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2276
timestamp 1569533753
transform 1 0 584 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2277
timestamp 1569533753
transform 1 0 584 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2278
timestamp 1569533753
transform 1 0 456 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2279
timestamp 1569533753
transform 1 0 456 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2280
timestamp 1569533753
transform 1 0 520 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2281
timestamp 1569533753
transform 1 0 520 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2282
timestamp 1569533753
transform 1 0 520 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2283
timestamp 1569533753
transform 1 0 456 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2284
timestamp 1569533753
transform 1 0 392 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2285
timestamp 1569533753
transform 1 0 584 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2286
timestamp 1569533753
transform 1 0 584 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2287
timestamp 1569533753
transform 1 0 584 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2288
timestamp 1569533753
transform 1 0 456 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2289
timestamp 1569533753
transform 1 0 456 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2290
timestamp 1569533753
transform 1 0 392 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2291
timestamp 1569533753
transform 1 0 392 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2292
timestamp 1569533753
transform 1 0 584 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2293
timestamp 1569533753
transform 1 0 520 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2294
timestamp 1569533753
transform 1 0 392 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2295
timestamp 1569533753
transform 1 0 584 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2296
timestamp 1569533753
transform 1 0 392 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2297
timestamp 1569533753
transform 1 0 456 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2298
timestamp 1569533753
transform 1 0 456 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2299
timestamp 1569533753
transform 1 0 456 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2300
timestamp 1569533753
transform 1 0 392 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2301
timestamp 1569533753
transform 1 0 584 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2302
timestamp 1569533753
transform 1 0 520 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2303
timestamp 1569533753
transform 1 0 520 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2304
timestamp 1569533753
transform 1 0 456 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2305
timestamp 1569533753
transform 1 0 584 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2306
timestamp 1569533753
transform 1 0 520 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2307
timestamp 1569533753
transform 1 0 584 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2308
timestamp 1569533753
transform 1 0 520 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2309
timestamp 1569533753
transform 1 0 456 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2310
timestamp 1569533753
transform 1 0 392 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2311
timestamp 1569533753
transform 1 0 264 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2312
timestamp 1569533753
transform 1 0 200 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2313
timestamp 1569533753
transform 1 0 72 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2314
timestamp 1569533753
transform 1 0 72 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2315
timestamp 1569533753
transform 1 0 264 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2316
timestamp 1569533753
transform 1 0 264 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2317
timestamp 1569533753
transform 1 0 200 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2318
timestamp 1569533753
transform 1 0 200 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2319
timestamp 1569533753
transform 1 0 72 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2320
timestamp 1569533753
transform 1 0 328 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2321
timestamp 1569533753
transform 1 0 200 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2322
timestamp 1569533753
transform 1 0 136 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2323
timestamp 1569533753
transform 1 0 136 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2324
timestamp 1569533753
transform 1 0 328 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2325
timestamp 1569533753
transform 1 0 72 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2326
timestamp 1569533753
transform 1 0 136 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2327
timestamp 1569533753
transform 1 0 328 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2328
timestamp 1569533753
transform 1 0 72 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2329
timestamp 1569533753
transform 1 0 136 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2330
timestamp 1569533753
transform 1 0 136 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2331
timestamp 1569533753
transform 1 0 328 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2332
timestamp 1569533753
transform 1 0 200 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2333
timestamp 1569533753
transform 1 0 264 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2334
timestamp 1569533753
transform 1 0 264 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2335
timestamp 1569533753
transform 1 0 328 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2336
timestamp 1569533753
transform 1 0 328 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2337
timestamp 1569533753
transform 1 0 328 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2338
timestamp 1569533753
transform 1 0 72 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2339
timestamp 1569533753
transform 1 0 200 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2340
timestamp 1569533753
transform 1 0 72 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2341
timestamp 1569533753
transform 1 0 136 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2342
timestamp 1569533753
transform 1 0 136 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2343
timestamp 1569533753
transform 1 0 72 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2344
timestamp 1569533753
transform 1 0 136 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2345
timestamp 1569533753
transform 1 0 72 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2346
timestamp 1569533753
transform 1 0 136 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2347
timestamp 1569533753
transform 1 0 328 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2348
timestamp 1569533753
transform 1 0 200 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2349
timestamp 1569533753
transform 1 0 136 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2350
timestamp 1569533753
transform 1 0 72 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2351
timestamp 1569533753
transform 1 0 200 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2352
timestamp 1569533753
transform 1 0 328 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2353
timestamp 1569533753
transform 1 0 264 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2354
timestamp 1569533753
transform 1 0 264 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2355
timestamp 1569533753
transform 1 0 264 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2356
timestamp 1569533753
transform 1 0 264 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2357
timestamp 1569533753
transform 1 0 264 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2358
timestamp 1569533753
transform 1 0 200 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2359
timestamp 1569533753
transform 1 0 200 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2360
timestamp 1569533753
transform 1 0 328 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2361
timestamp 1569533753
transform 1 0 392 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2362
timestamp 1569533753
transform 1 0 456 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2363
timestamp 1569533753
transform 1 0 392 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2364
timestamp 1569533753
transform 1 0 456 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2365
timestamp 1569533753
transform 1 0 584 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2366
timestamp 1569533753
transform 1 0 456 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2367
timestamp 1569533753
transform 1 0 456 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2368
timestamp 1569533753
transform 1 0 456 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2369
timestamp 1569533753
transform 1 0 584 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2370
timestamp 1569533753
transform 1 0 584 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2371
timestamp 1569533753
transform 1 0 520 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2372
timestamp 1569533753
transform 1 0 520 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2373
timestamp 1569533753
transform 1 0 520 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2374
timestamp 1569533753
transform 1 0 520 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2375
timestamp 1569533753
transform 1 0 584 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2376
timestamp 1569533753
transform 1 0 392 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2377
timestamp 1569533753
transform 1 0 584 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2378
timestamp 1569533753
transform 1 0 520 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2379
timestamp 1569533753
transform 1 0 392 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2380
timestamp 1569533753
transform 1 0 392 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2381
timestamp 1569533753
transform 1 0 1224 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2382
timestamp 1569533753
transform 1 0 968 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2383
timestamp 1569533753
transform 1 0 1096 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2384
timestamp 1569533753
transform 1 0 968 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2385
timestamp 1569533753
transform 1 0 968 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2386
timestamp 1569533753
transform 1 0 968 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2387
timestamp 1569533753
transform 1 0 1224 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2388
timestamp 1569533753
transform 1 0 1160 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2389
timestamp 1569533753
transform 1 0 1032 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2390
timestamp 1569533753
transform 1 0 1160 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2391
timestamp 1569533753
transform 1 0 1160 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2392
timestamp 1569533753
transform 1 0 1096 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2393
timestamp 1569533753
transform 1 0 1160 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2394
timestamp 1569533753
transform 1 0 1032 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2395
timestamp 1569533753
transform 1 0 1032 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2396
timestamp 1569533753
transform 1 0 1160 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2397
timestamp 1569533753
transform 1 0 1032 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2398
timestamp 1569533753
transform 1 0 1224 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2399
timestamp 1569533753
transform 1 0 968 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2400
timestamp 1569533753
transform 1 0 1096 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2401
timestamp 1569533753
transform 1 0 1096 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2402
timestamp 1569533753
transform 1 0 1224 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2403
timestamp 1569533753
transform 1 0 1032 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2404
timestamp 1569533753
transform 1 0 1224 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2405
timestamp 1569533753
transform 1 0 1096 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2406
timestamp 1569533753
transform 1 0 840 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2407
timestamp 1569533753
transform 1 0 840 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2408
timestamp 1569533753
transform 1 0 840 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2409
timestamp 1569533753
transform 1 0 712 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2410
timestamp 1569533753
transform 1 0 904 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2411
timestamp 1569533753
transform 1 0 904 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2412
timestamp 1569533753
transform 1 0 904 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2413
timestamp 1569533753
transform 1 0 904 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2414
timestamp 1569533753
transform 1 0 712 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2415
timestamp 1569533753
transform 1 0 776 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2416
timestamp 1569533753
transform 1 0 840 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2417
timestamp 1569533753
transform 1 0 776 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2418
timestamp 1569533753
transform 1 0 776 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2419
timestamp 1569533753
transform 1 0 776 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2420
timestamp 1569533753
transform 1 0 776 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2421
timestamp 1569533753
transform 1 0 712 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2422
timestamp 1569533753
transform 1 0 904 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2423
timestamp 1569533753
transform 1 0 712 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2424
timestamp 1569533753
transform 1 0 840 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2425
timestamp 1569533753
transform 1 0 712 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2426
timestamp 1569533753
transform 1 0 712 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2427
timestamp 1569533753
transform 1 0 712 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2428
timestamp 1569533753
transform 1 0 712 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2429
timestamp 1569533753
transform 1 0 712 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2430
timestamp 1569533753
transform 1 0 776 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2431
timestamp 1569533753
transform 1 0 776 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2432
timestamp 1569533753
transform 1 0 712 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2433
timestamp 1569533753
transform 1 0 840 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2434
timestamp 1569533753
transform 1 0 840 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2435
timestamp 1569533753
transform 1 0 776 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2436
timestamp 1569533753
transform 1 0 776 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2437
timestamp 1569533753
transform 1 0 776 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2438
timestamp 1569533753
transform 1 0 904 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2439
timestamp 1569533753
transform 1 0 840 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2440
timestamp 1569533753
transform 1 0 840 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2441
timestamp 1569533753
transform 1 0 904 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2442
timestamp 1569533753
transform 1 0 840 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2443
timestamp 1569533753
transform 1 0 904 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2444
timestamp 1569533753
transform 1 0 904 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2445
timestamp 1569533753
transform 1 0 904 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2446
timestamp 1569533753
transform 1 0 1096 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2447
timestamp 1569533753
transform 1 0 1096 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2448
timestamp 1569533753
transform 1 0 1096 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2449
timestamp 1569533753
transform 1 0 1224 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2450
timestamp 1569533753
transform 1 0 1096 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2451
timestamp 1569533753
transform 1 0 1096 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2452
timestamp 1569533753
transform 1 0 1224 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2453
timestamp 1569533753
transform 1 0 1160 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2454
timestamp 1569533753
transform 1 0 1160 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2455
timestamp 1569533753
transform 1 0 1160 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2456
timestamp 1569533753
transform 1 0 968 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2457
timestamp 1569533753
transform 1 0 968 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2458
timestamp 1569533753
transform 1 0 968 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2459
timestamp 1569533753
transform 1 0 1032 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2460
timestamp 1569533753
transform 1 0 1032 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2461
timestamp 1569533753
transform 1 0 1032 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2462
timestamp 1569533753
transform 1 0 1224 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2463
timestamp 1569533753
transform 1 0 1224 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2464
timestamp 1569533753
transform 1 0 1224 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2465
timestamp 1569533753
transform 1 0 1160 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2466
timestamp 1569533753
transform 1 0 968 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2467
timestamp 1569533753
transform 1 0 968 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2468
timestamp 1569533753
transform 1 0 1160 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2469
timestamp 1569533753
transform 1 0 1032 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2470
timestamp 1569533753
transform 1 0 1032 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2471
timestamp 1569533753
transform 1 0 648 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2472
timestamp 1569533753
transform 1 0 648 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_2473
timestamp 1569533753
transform 1 0 648 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2474
timestamp 1569533753
transform 1 0 648 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2475
timestamp 1569533753
transform 1 0 648 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2476
timestamp 1569533753
transform 1 0 648 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2477
timestamp 1569533753
transform 1 0 648 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_2478
timestamp 1569533753
transform 1 0 648 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_2479
timestamp 1569533753
transform 1 0 648 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2480
timestamp 1569533753
transform 1 0 648 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_2481
timestamp 1569533753
transform 1 0 648 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2482
timestamp 1569533753
transform 1 0 648 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2483
timestamp 1569533753
transform 1 0 648 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_2484
timestamp 1569533753
transform 1 0 648 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_2485
timestamp 1569533753
transform 1 0 648 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_2486
timestamp 1569533753
transform 1 0 648 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_2487
timestamp 1569533753
transform 1 0 648 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2488
timestamp 1569533753
transform 1 0 648 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_2489
timestamp 1569533753
transform 1 0 648 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_2490
timestamp 1569533753
transform 1 0 1096 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2491
timestamp 1569533753
transform 1 0 1032 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2492
timestamp 1569533753
transform 1 0 1096 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2493
timestamp 1569533753
transform 1 0 1032 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2494
timestamp 1569533753
transform 1 0 968 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2495
timestamp 1569533753
transform 1 0 1160 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2496
timestamp 1569533753
transform 1 0 1160 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2497
timestamp 1569533753
transform 1 0 1096 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2498
timestamp 1569533753
transform 1 0 1096 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2499
timestamp 1569533753
transform 1 0 1224 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2500
timestamp 1569533753
transform 1 0 1224 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2501
timestamp 1569533753
transform 1 0 1224 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2502
timestamp 1569533753
transform 1 0 1160 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2503
timestamp 1569533753
transform 1 0 1224 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2504
timestamp 1569533753
transform 1 0 1224 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2505
timestamp 1569533753
transform 1 0 968 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2506
timestamp 1569533753
transform 1 0 968 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2507
timestamp 1569533753
transform 1 0 968 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2508
timestamp 1569533753
transform 1 0 1032 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2509
timestamp 1569533753
transform 1 0 968 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2510
timestamp 1569533753
transform 1 0 1160 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2511
timestamp 1569533753
transform 1 0 1160 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2512
timestamp 1569533753
transform 1 0 1032 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2513
timestamp 1569533753
transform 1 0 1096 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2514
timestamp 1569533753
transform 1 0 1032 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2515
timestamp 1569533753
transform 1 0 712 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2516
timestamp 1569533753
transform 1 0 840 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2517
timestamp 1569533753
transform 1 0 840 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2518
timestamp 1569533753
transform 1 0 776 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2519
timestamp 1569533753
transform 1 0 776 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2520
timestamp 1569533753
transform 1 0 840 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2521
timestamp 1569533753
transform 1 0 712 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2522
timestamp 1569533753
transform 1 0 904 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2523
timestamp 1569533753
transform 1 0 904 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2524
timestamp 1569533753
transform 1 0 712 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2525
timestamp 1569533753
transform 1 0 904 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2526
timestamp 1569533753
transform 1 0 904 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2527
timestamp 1569533753
transform 1 0 776 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2528
timestamp 1569533753
transform 1 0 712 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2529
timestamp 1569533753
transform 1 0 840 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2530
timestamp 1569533753
transform 1 0 904 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2531
timestamp 1569533753
transform 1 0 776 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2532
timestamp 1569533753
transform 1 0 712 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2533
timestamp 1569533753
transform 1 0 776 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2534
timestamp 1569533753
transform 1 0 840 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2535
timestamp 1569533753
transform 1 0 840 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2536
timestamp 1569533753
transform 1 0 840 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2537
timestamp 1569533753
transform 1 0 712 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2538
timestamp 1569533753
transform 1 0 840 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2539
timestamp 1569533753
transform 1 0 840 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2540
timestamp 1569533753
transform 1 0 712 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2541
timestamp 1569533753
transform 1 0 712 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2542
timestamp 1569533753
transform 1 0 776 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2543
timestamp 1569533753
transform 1 0 776 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2544
timestamp 1569533753
transform 1 0 776 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2545
timestamp 1569533753
transform 1 0 904 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2546
timestamp 1569533753
transform 1 0 776 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2547
timestamp 1569533753
transform 1 0 904 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2548
timestamp 1569533753
transform 1 0 904 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2549
timestamp 1569533753
transform 1 0 712 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2550
timestamp 1569533753
transform 1 0 904 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2551
timestamp 1569533753
transform 1 0 1032 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2552
timestamp 1569533753
transform 1 0 1032 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2553
timestamp 1569533753
transform 1 0 1160 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2554
timestamp 1569533753
transform 1 0 1160 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2555
timestamp 1569533753
transform 1 0 1224 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2556
timestamp 1569533753
transform 1 0 1160 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2557
timestamp 1569533753
transform 1 0 1096 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2558
timestamp 1569533753
transform 1 0 1160 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2559
timestamp 1569533753
transform 1 0 1224 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2560
timestamp 1569533753
transform 1 0 1096 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2561
timestamp 1569533753
transform 1 0 1224 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2562
timestamp 1569533753
transform 1 0 1096 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2563
timestamp 1569533753
transform 1 0 1224 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2564
timestamp 1569533753
transform 1 0 1096 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2565
timestamp 1569533753
transform 1 0 968 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2566
timestamp 1569533753
transform 1 0 968 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2567
timestamp 1569533753
transform 1 0 968 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2568
timestamp 1569533753
transform 1 0 968 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2569
timestamp 1569533753
transform 1 0 1032 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2570
timestamp 1569533753
transform 1 0 1032 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2571
timestamp 1569533753
transform 1 0 392 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2572
timestamp 1569533753
transform 1 0 584 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2573
timestamp 1569533753
transform 1 0 584 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2574
timestamp 1569533753
transform 1 0 392 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2575
timestamp 1569533753
transform 1 0 456 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2576
timestamp 1569533753
transform 1 0 584 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2577
timestamp 1569533753
transform 1 0 392 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2578
timestamp 1569533753
transform 1 0 520 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2579
timestamp 1569533753
transform 1 0 520 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2580
timestamp 1569533753
transform 1 0 392 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2581
timestamp 1569533753
transform 1 0 584 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2582
timestamp 1569533753
transform 1 0 520 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2583
timestamp 1569533753
transform 1 0 456 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2584
timestamp 1569533753
transform 1 0 392 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2585
timestamp 1569533753
transform 1 0 584 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2586
timestamp 1569533753
transform 1 0 520 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2587
timestamp 1569533753
transform 1 0 456 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2588
timestamp 1569533753
transform 1 0 520 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2589
timestamp 1569533753
transform 1 0 456 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2590
timestamp 1569533753
transform 1 0 456 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2591
timestamp 1569533753
transform 1 0 200 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2592
timestamp 1569533753
transform 1 0 72 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2593
timestamp 1569533753
transform 1 0 200 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2594
timestamp 1569533753
transform 1 0 72 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2595
timestamp 1569533753
transform 1 0 72 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2596
timestamp 1569533753
transform 1 0 136 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2597
timestamp 1569533753
transform 1 0 264 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2598
timestamp 1569533753
transform 1 0 136 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2599
timestamp 1569533753
transform 1 0 72 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2600
timestamp 1569533753
transform 1 0 328 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2601
timestamp 1569533753
transform 1 0 264 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2602
timestamp 1569533753
transform 1 0 136 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2603
timestamp 1569533753
transform 1 0 72 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2604
timestamp 1569533753
transform 1 0 136 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2605
timestamp 1569533753
transform 1 0 264 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2606
timestamp 1569533753
transform 1 0 264 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2607
timestamp 1569533753
transform 1 0 136 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2608
timestamp 1569533753
transform 1 0 264 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2609
timestamp 1569533753
transform 1 0 200 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2610
timestamp 1569533753
transform 1 0 328 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2611
timestamp 1569533753
transform 1 0 328 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2612
timestamp 1569533753
transform 1 0 200 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2613
timestamp 1569533753
transform 1 0 200 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2614
timestamp 1569533753
transform 1 0 328 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2615
timestamp 1569533753
transform 1 0 328 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2616
timestamp 1569533753
transform 1 0 136 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2617
timestamp 1569533753
transform 1 0 136 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2618
timestamp 1569533753
transform 1 0 136 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2619
timestamp 1569533753
transform 1 0 136 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2620
timestamp 1569533753
transform 1 0 72 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2621
timestamp 1569533753
transform 1 0 72 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2622
timestamp 1569533753
transform 1 0 200 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2623
timestamp 1569533753
transform 1 0 200 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2624
timestamp 1569533753
transform 1 0 200 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2625
timestamp 1569533753
transform 1 0 200 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2626
timestamp 1569533753
transform 1 0 72 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2627
timestamp 1569533753
transform 1 0 264 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2628
timestamp 1569533753
transform 1 0 264 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2629
timestamp 1569533753
transform 1 0 264 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2630
timestamp 1569533753
transform 1 0 264 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2631
timestamp 1569533753
transform 1 0 328 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2632
timestamp 1569533753
transform 1 0 328 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2633
timestamp 1569533753
transform 1 0 328 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2634
timestamp 1569533753
transform 1 0 328 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2635
timestamp 1569533753
transform 1 0 72 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2636
timestamp 1569533753
transform 1 0 520 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2637
timestamp 1569533753
transform 1 0 520 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2638
timestamp 1569533753
transform 1 0 456 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2639
timestamp 1569533753
transform 1 0 456 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2640
timestamp 1569533753
transform 1 0 392 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2641
timestamp 1569533753
transform 1 0 392 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2642
timestamp 1569533753
transform 1 0 392 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2643
timestamp 1569533753
transform 1 0 392 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2644
timestamp 1569533753
transform 1 0 456 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2645
timestamp 1569533753
transform 1 0 456 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2646
timestamp 1569533753
transform 1 0 584 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2647
timestamp 1569533753
transform 1 0 584 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2648
timestamp 1569533753
transform 1 0 584 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2649
timestamp 1569533753
transform 1 0 520 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2650
timestamp 1569533753
transform 1 0 520 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2651
timestamp 1569533753
transform 1 0 584 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2652
timestamp 1569533753
transform 1 0 584 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2653
timestamp 1569533753
transform 1 0 392 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2654
timestamp 1569533753
transform 1 0 520 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2655
timestamp 1569533753
transform 1 0 520 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2656
timestamp 1569533753
transform 1 0 584 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2657
timestamp 1569533753
transform 1 0 520 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2658
timestamp 1569533753
transform 1 0 456 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2659
timestamp 1569533753
transform 1 0 456 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2660
timestamp 1569533753
transform 1 0 584 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2661
timestamp 1569533753
transform 1 0 520 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2662
timestamp 1569533753
transform 1 0 392 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2663
timestamp 1569533753
transform 1 0 584 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2664
timestamp 1569533753
transform 1 0 392 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2665
timestamp 1569533753
transform 1 0 456 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2666
timestamp 1569533753
transform 1 0 456 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2667
timestamp 1569533753
transform 1 0 392 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2668
timestamp 1569533753
transform 1 0 136 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2669
timestamp 1569533753
transform 1 0 328 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2670
timestamp 1569533753
transform 1 0 264 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2671
timestamp 1569533753
transform 1 0 264 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2672
timestamp 1569533753
transform 1 0 72 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2673
timestamp 1569533753
transform 1 0 200 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2674
timestamp 1569533753
transform 1 0 328 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2675
timestamp 1569533753
transform 1 0 136 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2676
timestamp 1569533753
transform 1 0 328 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2677
timestamp 1569533753
transform 1 0 72 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2678
timestamp 1569533753
transform 1 0 264 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2679
timestamp 1569533753
transform 1 0 328 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2680
timestamp 1569533753
transform 1 0 136 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2681
timestamp 1569533753
transform 1 0 264 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2682
timestamp 1569533753
transform 1 0 136 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2683
timestamp 1569533753
transform 1 0 72 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2684
timestamp 1569533753
transform 1 0 200 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2685
timestamp 1569533753
transform 1 0 200 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2686
timestamp 1569533753
transform 1 0 200 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2687
timestamp 1569533753
transform 1 0 72 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2688
timestamp 1569533753
transform 1 0 264 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2689
timestamp 1569533753
transform 1 0 264 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2690
timestamp 1569533753
transform 1 0 200 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2691
timestamp 1569533753
transform 1 0 136 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2692
timestamp 1569533753
transform 1 0 136 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2693
timestamp 1569533753
transform 1 0 136 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2694
timestamp 1569533753
transform 1 0 136 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2695
timestamp 1569533753
transform 1 0 72 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2696
timestamp 1569533753
transform 1 0 328 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2697
timestamp 1569533753
transform 1 0 328 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2698
timestamp 1569533753
transform 1 0 328 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2699
timestamp 1569533753
transform 1 0 328 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2700
timestamp 1569533753
transform 1 0 72 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2701
timestamp 1569533753
transform 1 0 72 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2702
timestamp 1569533753
transform 1 0 264 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2703
timestamp 1569533753
transform 1 0 200 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2704
timestamp 1569533753
transform 1 0 200 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2705
timestamp 1569533753
transform 1 0 200 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2706
timestamp 1569533753
transform 1 0 264 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2707
timestamp 1569533753
transform 1 0 72 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2708
timestamp 1569533753
transform 1 0 392 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2709
timestamp 1569533753
transform 1 0 392 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2710
timestamp 1569533753
transform 1 0 392 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2711
timestamp 1569533753
transform 1 0 392 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2712
timestamp 1569533753
transform 1 0 456 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2713
timestamp 1569533753
transform 1 0 456 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2714
timestamp 1569533753
transform 1 0 456 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2715
timestamp 1569533753
transform 1 0 456 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2716
timestamp 1569533753
transform 1 0 520 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2717
timestamp 1569533753
transform 1 0 520 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2718
timestamp 1569533753
transform 1 0 520 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2719
timestamp 1569533753
transform 1 0 520 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2720
timestamp 1569533753
transform 1 0 584 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2721
timestamp 1569533753
transform 1 0 584 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2722
timestamp 1569533753
transform 1 0 584 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2723
timestamp 1569533753
transform 1 0 584 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2724
timestamp 1569533753
transform 1 0 1096 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2725
timestamp 1569533753
transform 1 0 1160 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2726
timestamp 1569533753
transform 1 0 968 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2727
timestamp 1569533753
transform 1 0 1096 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2728
timestamp 1569533753
transform 1 0 1224 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2729
timestamp 1569533753
transform 1 0 968 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2730
timestamp 1569533753
transform 1 0 1096 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2731
timestamp 1569533753
transform 1 0 1224 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2732
timestamp 1569533753
transform 1 0 1096 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2733
timestamp 1569533753
transform 1 0 1224 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2734
timestamp 1569533753
transform 1 0 968 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2735
timestamp 1569533753
transform 1 0 968 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2736
timestamp 1569533753
transform 1 0 1160 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2737
timestamp 1569533753
transform 1 0 1160 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2738
timestamp 1569533753
transform 1 0 1032 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2739
timestamp 1569533753
transform 1 0 1032 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2740
timestamp 1569533753
transform 1 0 1032 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2741
timestamp 1569533753
transform 1 0 1032 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2742
timestamp 1569533753
transform 1 0 1224 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2743
timestamp 1569533753
transform 1 0 1160 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2744
timestamp 1569533753
transform 1 0 712 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2745
timestamp 1569533753
transform 1 0 840 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2746
timestamp 1569533753
transform 1 0 776 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2747
timestamp 1569533753
transform 1 0 776 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2748
timestamp 1569533753
transform 1 0 904 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2749
timestamp 1569533753
transform 1 0 776 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2750
timestamp 1569533753
transform 1 0 904 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2751
timestamp 1569533753
transform 1 0 840 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2752
timestamp 1569533753
transform 1 0 840 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2753
timestamp 1569533753
transform 1 0 840 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2754
timestamp 1569533753
transform 1 0 904 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2755
timestamp 1569533753
transform 1 0 776 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2756
timestamp 1569533753
transform 1 0 904 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2757
timestamp 1569533753
transform 1 0 712 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2758
timestamp 1569533753
transform 1 0 712 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2759
timestamp 1569533753
transform 1 0 712 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2760
timestamp 1569533753
transform 1 0 904 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2761
timestamp 1569533753
transform 1 0 904 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2762
timestamp 1569533753
transform 1 0 904 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2763
timestamp 1569533753
transform 1 0 776 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2764
timestamp 1569533753
transform 1 0 840 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2765
timestamp 1569533753
transform 1 0 776 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2766
timestamp 1569533753
transform 1 0 776 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2767
timestamp 1569533753
transform 1 0 776 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2768
timestamp 1569533753
transform 1 0 840 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2769
timestamp 1569533753
transform 1 0 712 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2770
timestamp 1569533753
transform 1 0 712 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2771
timestamp 1569533753
transform 1 0 840 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2772
timestamp 1569533753
transform 1 0 712 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2773
timestamp 1569533753
transform 1 0 712 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2774
timestamp 1569533753
transform 1 0 904 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2775
timestamp 1569533753
transform 1 0 840 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2776
timestamp 1569533753
transform 1 0 968 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2777
timestamp 1569533753
transform 1 0 968 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2778
timestamp 1569533753
transform 1 0 968 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2779
timestamp 1569533753
transform 1 0 968 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2780
timestamp 1569533753
transform 1 0 1032 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2781
timestamp 1569533753
transform 1 0 1032 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2782
timestamp 1569533753
transform 1 0 1032 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2783
timestamp 1569533753
transform 1 0 1032 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2784
timestamp 1569533753
transform 1 0 1096 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2785
timestamp 1569533753
transform 1 0 1096 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2786
timestamp 1569533753
transform 1 0 1096 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2787
timestamp 1569533753
transform 1 0 1096 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2788
timestamp 1569533753
transform 1 0 1160 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2789
timestamp 1569533753
transform 1 0 1160 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2790
timestamp 1569533753
transform 1 0 1160 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2791
timestamp 1569533753
transform 1 0 1160 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2792
timestamp 1569533753
transform 1 0 1224 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2793
timestamp 1569533753
transform 1 0 1224 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2794
timestamp 1569533753
transform 1 0 1224 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2795
timestamp 1569533753
transform 1 0 1224 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2796
timestamp 1569533753
transform 1 0 456 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2797
timestamp 1569533753
transform 1 0 1096 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2798
timestamp 1569533753
transform 1 0 136 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2799
timestamp 1569533753
transform 1 0 776 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2800
timestamp 1569533753
transform 1 0 520 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2801
timestamp 1569533753
transform 1 0 1160 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2802
timestamp 1569533753
transform 1 0 200 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2803
timestamp 1569533753
transform 1 0 840 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2804
timestamp 1569533753
transform 1 0 264 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2805
timestamp 1569533753
transform 1 0 904 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2806
timestamp 1569533753
transform 1 0 328 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2807
timestamp 1569533753
transform 1 0 968 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2808
timestamp 1569533753
transform 1 0 392 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2809
timestamp 1569533753
transform 1 0 1032 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2810
timestamp 1569533753
transform 1 0 648 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2811
timestamp 1569533753
transform 1 0 584 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2812
timestamp 1569533753
transform 1 0 1224 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2813
timestamp 1569533753
transform 1 0 648 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2814
timestamp 1569533753
transform 1 0 648 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2815
timestamp 1569533753
transform 1 0 648 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2816
timestamp 1569533753
transform 1 0 648 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2817
timestamp 1569533753
transform 1 0 648 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2818
timestamp 1569533753
transform 1 0 648 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2819
timestamp 1569533753
transform 1 0 648 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2820
timestamp 1569533753
transform 1 0 648 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2821
timestamp 1569533753
transform 1 0 648 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2822
timestamp 1569533753
transform 1 0 648 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2823
timestamp 1569533753
transform 1 0 648 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2824
timestamp 1569533753
transform 1 0 648 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2825
timestamp 1569533753
transform 1 0 72 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2826
timestamp 1569533753
transform 1 0 712 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2827
timestamp 1569533753
transform 1 0 648 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2828
timestamp 1569533753
transform 1 0 648 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2829
timestamp 1569533753
transform 1 0 648 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2830
timestamp 1569533753
transform 1 0 648 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2831
timestamp 1569533753
transform 1 0 648 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2832
timestamp 1569533753
transform 1 0 2376 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2833
timestamp 1569533753
transform 1 0 2440 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2834
timestamp 1569533753
transform 1 0 2376 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2835
timestamp 1569533753
transform 1 0 2376 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2836
timestamp 1569533753
transform 1 0 2376 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2837
timestamp 1569533753
transform 1 0 2376 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2838
timestamp 1569533753
transform 1 0 2376 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2839
timestamp 1569533753
transform 1 0 2376 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2840
timestamp 1569533753
transform 1 0 2440 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2841
timestamp 1569533753
transform 1 0 2440 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2842
timestamp 1569533753
transform 1 0 2312 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2843
timestamp 1569533753
transform 1 0 2312 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2844
timestamp 1569533753
transform 1 0 2312 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2845
timestamp 1569533753
transform 1 0 2312 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2846
timestamp 1569533753
transform 1 0 2312 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2847
timestamp 1569533753
transform 1 0 2440 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2848
timestamp 1569533753
transform 1 0 2440 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2849
timestamp 1569533753
transform 1 0 2440 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2850
timestamp 1569533753
transform 1 0 2440 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2851
timestamp 1569533753
transform 1 0 2440 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2852
timestamp 1569533753
transform 1 0 2312 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2853
timestamp 1569533753
transform 1 0 2312 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2854
timestamp 1569533753
transform 1 0 2312 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2855
timestamp 1569533753
transform 1 0 2312 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2856
timestamp 1569533753
transform 1 0 2440 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2857
timestamp 1569533753
transform 1 0 2376 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2858
timestamp 1569533753
transform 1 0 2376 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2859
timestamp 1569533753
transform 1 0 1352 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2860
timestamp 1569533753
transform 1 0 1352 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2861
timestamp 1569533753
transform 1 0 1352 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2862
timestamp 1569533753
transform 1 0 1352 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2863
timestamp 1569533753
transform 1 0 1288 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2864
timestamp 1569533753
transform 1 0 1352 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2865
timestamp 1569533753
transform 1 0 1352 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2866
timestamp 1569533753
transform 1 0 1416 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2867
timestamp 1569533753
transform 1 0 1352 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2868
timestamp 1569533753
transform 1 0 1416 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2869
timestamp 1569533753
transform 1 0 1416 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2870
timestamp 1569533753
transform 1 0 1416 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2871
timestamp 1569533753
transform 1 0 1416 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2872
timestamp 1569533753
transform 1 0 1480 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2873
timestamp 1569533753
transform 1 0 1480 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2874
timestamp 1569533753
transform 1 0 1288 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2875
timestamp 1569533753
transform 1 0 1480 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2876
timestamp 1569533753
transform 1 0 1480 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2877
timestamp 1569533753
transform 1 0 1352 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2878
timestamp 1569533753
transform 1 0 1288 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2879
timestamp 1569533753
transform 1 0 1416 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2880
timestamp 1569533753
transform 1 0 1416 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2881
timestamp 1569533753
transform 1 0 1416 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2882
timestamp 1569533753
transform 1 0 1416 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2883
timestamp 1569533753
transform 1 0 1288 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2884
timestamp 1569533753
transform 1 0 1480 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_2885
timestamp 1569533753
transform 1 0 1480 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_2886
timestamp 1569533753
transform 1 0 1480 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_2887
timestamp 1569533753
transform 1 0 1480 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_2888
timestamp 1569533753
transform 1 0 1352 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2889
timestamp 1569533753
transform 1 0 1288 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2890
timestamp 1569533753
transform 1 0 1480 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_2891
timestamp 1569533753
transform 1 0 1288 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_2892
timestamp 1569533753
transform 1 0 1288 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_2893
timestamp 1569533753
transform 1 0 1288 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_2894
timestamp 1569533753
transform 1 0 1288 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_2895
timestamp 1569533753
transform 1 0 1352 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2896
timestamp 1569533753
transform 1 0 1480 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2897
timestamp 1569533753
transform 1 0 1480 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2898
timestamp 1569533753
transform 1 0 1416 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2899
timestamp 1569533753
transform 1 0 1416 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2900
timestamp 1569533753
transform 1 0 1480 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2901
timestamp 1569533753
transform 1 0 1480 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2902
timestamp 1569533753
transform 1 0 1352 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2903
timestamp 1569533753
transform 1 0 1352 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2904
timestamp 1569533753
transform 1 0 1352 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2905
timestamp 1569533753
transform 1 0 1352 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2906
timestamp 1569533753
transform 1 0 1352 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2907
timestamp 1569533753
transform 1 0 1480 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2908
timestamp 1569533753
transform 1 0 1352 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2909
timestamp 1569533753
transform 1 0 1480 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2910
timestamp 1569533753
transform 1 0 1352 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2911
timestamp 1569533753
transform 1 0 1416 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2912
timestamp 1569533753
transform 1 0 1416 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2913
timestamp 1569533753
transform 1 0 1480 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2914
timestamp 1569533753
transform 1 0 1416 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2915
timestamp 1569533753
transform 1 0 1416 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2916
timestamp 1569533753
transform 1 0 1416 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2917
timestamp 1569533753
transform 1 0 1288 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2918
timestamp 1569533753
transform 1 0 1288 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2919
timestamp 1569533753
transform 1 0 1416 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2920
timestamp 1569533753
transform 1 0 1288 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2921
timestamp 1569533753
transform 1 0 1288 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2922
timestamp 1569533753
transform 1 0 1288 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2923
timestamp 1569533753
transform 1 0 1288 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2924
timestamp 1569533753
transform 1 0 1288 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2925
timestamp 1569533753
transform 1 0 1288 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2926
timestamp 1569533753
transform 1 0 1480 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2927
timestamp 1569533753
transform 1 0 2376 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2928
timestamp 1569533753
transform 1 0 2312 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2929
timestamp 1569533753
transform 1 0 2312 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2930
timestamp 1569533753
transform 1 0 2312 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2931
timestamp 1569533753
transform 1 0 2312 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2932
timestamp 1569533753
transform 1 0 2312 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2933
timestamp 1569533753
transform 1 0 2312 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2934
timestamp 1569533753
transform 1 0 2376 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2935
timestamp 1569533753
transform 1 0 2376 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2936
timestamp 1569533753
transform 1 0 2376 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2937
timestamp 1569533753
transform 1 0 2376 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2938
timestamp 1569533753
transform 1 0 2376 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2939
timestamp 1569533753
transform 1 0 2440 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_2940
timestamp 1569533753
transform 1 0 2440 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_2941
timestamp 1569533753
transform 1 0 2440 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_2942
timestamp 1569533753
transform 1 0 2440 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_2943
timestamp 1569533753
transform 1 0 2440 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_2944
timestamp 1569533753
transform 1 0 2312 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2945
timestamp 1569533753
transform 1 0 2440 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_2946
timestamp 1569533753
transform 1 0 2376 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2947
timestamp 1569533753
transform 1 0 2312 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2948
timestamp 1569533753
transform 1 0 2440 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_2949
timestamp 1569533753
transform 1 0 2376 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2950
timestamp 1569533753
transform 1 0 2440 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_2951
timestamp 1569533753
transform 1 0 1416 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2952
timestamp 1569533753
transform 1 0 1480 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2953
timestamp 1569533753
transform 1 0 2312 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2954
timestamp 1569533753
transform 1 0 2376 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2955
timestamp 1569533753
transform 1 0 2440 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2956
timestamp 1569533753
transform 1 0 1288 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2957
timestamp 1569533753
transform 1 0 1352 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_2958
timestamp 1569533753
transform 1 0 4680 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2959
timestamp 1569533753
transform 1 0 4744 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2960
timestamp 1569533753
transform 1 0 4872 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2961
timestamp 1569533753
transform 1 0 4872 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2962
timestamp 1569533753
transform 1 0 4744 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2963
timestamp 1569533753
transform 1 0 4680 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2964
timestamp 1569533753
transform 1 0 4680 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2965
timestamp 1569533753
transform 1 0 4744 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2966
timestamp 1569533753
transform 1 0 4680 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2967
timestamp 1569533753
transform 1 0 4808 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2968
timestamp 1569533753
transform 1 0 4744 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2969
timestamp 1569533753
transform 1 0 4872 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2970
timestamp 1569533753
transform 1 0 4808 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2971
timestamp 1569533753
transform 1 0 4808 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2972
timestamp 1569533753
transform 1 0 4808 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2973
timestamp 1569533753
transform 1 0 4872 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2974
timestamp 1569533753
transform 1 0 4616 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2975
timestamp 1569533753
transform 1 0 4488 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2976
timestamp 1569533753
transform 1 0 4424 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2977
timestamp 1569533753
transform 1 0 4424 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2978
timestamp 1569533753
transform 1 0 4488 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2979
timestamp 1569533753
transform 1 0 4616 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2980
timestamp 1569533753
transform 1 0 4488 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2981
timestamp 1569533753
transform 1 0 4616 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2982
timestamp 1569533753
transform 1 0 4616 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2983
timestamp 1569533753
transform 1 0 4552 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2984
timestamp 1569533753
transform 1 0 4552 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_2985
timestamp 1569533753
transform 1 0 4552 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2986
timestamp 1569533753
transform 1 0 4424 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2987
timestamp 1569533753
transform 1 0 4552 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_2988
timestamp 1569533753
transform 1 0 4424 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_2989
timestamp 1569533753
transform 1 0 4488 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_2990
timestamp 1569533753
transform 1 0 4616 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_2991
timestamp 1569533753
transform 1 0 4552 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2992
timestamp 1569533753
transform 1 0 4424 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2993
timestamp 1569533753
transform 1 0 4616 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_2994
timestamp 1569533753
transform 1 0 4488 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_2995
timestamp 1569533753
transform 1 0 4616 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2996
timestamp 1569533753
transform 1 0 4616 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2997
timestamp 1569533753
transform 1 0 4488 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_2998
timestamp 1569533753
transform 1 0 4488 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_2999
timestamp 1569533753
transform 1 0 4488 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3000
timestamp 1569533753
transform 1 0 4552 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3001
timestamp 1569533753
transform 1 0 4424 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3002
timestamp 1569533753
transform 1 0 4424 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3003
timestamp 1569533753
transform 1 0 4488 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3004
timestamp 1569533753
transform 1 0 4424 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3005
timestamp 1569533753
transform 1 0 4552 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3006
timestamp 1569533753
transform 1 0 4424 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3007
timestamp 1569533753
transform 1 0 4552 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3008
timestamp 1569533753
transform 1 0 4552 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3009
timestamp 1569533753
transform 1 0 4616 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3010
timestamp 1569533753
transform 1 0 4872 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3011
timestamp 1569533753
transform 1 0 4744 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3012
timestamp 1569533753
transform 1 0 4872 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3013
timestamp 1569533753
transform 1 0 4744 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3014
timestamp 1569533753
transform 1 0 4872 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3015
timestamp 1569533753
transform 1 0 4808 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3016
timestamp 1569533753
transform 1 0 4744 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3017
timestamp 1569533753
transform 1 0 4680 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3018
timestamp 1569533753
transform 1 0 4808 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3019
timestamp 1569533753
transform 1 0 4680 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3020
timestamp 1569533753
transform 1 0 4808 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3021
timestamp 1569533753
transform 1 0 4808 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3022
timestamp 1569533753
transform 1 0 4680 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3023
timestamp 1569533753
transform 1 0 4872 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3024
timestamp 1569533753
transform 1 0 4872 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3025
timestamp 1569533753
transform 1 0 4680 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3026
timestamp 1569533753
transform 1 0 4680 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3027
timestamp 1569533753
transform 1 0 4744 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3028
timestamp 1569533753
transform 1 0 4808 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3029
timestamp 1569533753
transform 1 0 4744 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3030
timestamp 1569533753
transform 1 0 4104 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3031
timestamp 1569533753
transform 1 0 4232 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3032
timestamp 1569533753
transform 1 0 4104 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3033
timestamp 1569533753
transform 1 0 4232 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3034
timestamp 1569533753
transform 1 0 4168 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3035
timestamp 1569533753
transform 1 0 4296 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3036
timestamp 1569533753
transform 1 0 4296 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3037
timestamp 1569533753
transform 1 0 4168 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3038
timestamp 1569533753
transform 1 0 4296 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3039
timestamp 1569533753
transform 1 0 4104 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3040
timestamp 1569533753
transform 1 0 4232 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3041
timestamp 1569533753
transform 1 0 4168 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3042
timestamp 1569533753
transform 1 0 4168 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3043
timestamp 1569533753
transform 1 0 4232 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3044
timestamp 1569533753
transform 1 0 4104 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3045
timestamp 1569533753
transform 1 0 4296 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3046
timestamp 1569533753
transform 1 0 3848 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3047
timestamp 1569533753
transform 1 0 3976 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3048
timestamp 1569533753
transform 1 0 3912 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3049
timestamp 1569533753
transform 1 0 3976 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3050
timestamp 1569533753
transform 1 0 3784 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3051
timestamp 1569533753
transform 1 0 3848 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3052
timestamp 1569533753
transform 1 0 3976 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3053
timestamp 1569533753
transform 1 0 3784 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3054
timestamp 1569533753
transform 1 0 4040 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3055
timestamp 1569533753
transform 1 0 3976 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3056
timestamp 1569533753
transform 1 0 3912 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3057
timestamp 1569533753
transform 1 0 3912 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3058
timestamp 1569533753
transform 1 0 3848 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3059
timestamp 1569533753
transform 1 0 3848 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3060
timestamp 1569533753
transform 1 0 3784 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3061
timestamp 1569533753
transform 1 0 4040 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3062
timestamp 1569533753
transform 1 0 4040 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3063
timestamp 1569533753
transform 1 0 3912 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3064
timestamp 1569533753
transform 1 0 4040 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3065
timestamp 1569533753
transform 1 0 3784 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3066
timestamp 1569533753
transform 1 0 3912 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3067
timestamp 1569533753
transform 1 0 3784 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3068
timestamp 1569533753
transform 1 0 3848 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3069
timestamp 1569533753
transform 1 0 4040 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3070
timestamp 1569533753
transform 1 0 3848 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3071
timestamp 1569533753
transform 1 0 3976 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3072
timestamp 1569533753
transform 1 0 3976 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3073
timestamp 1569533753
transform 1 0 3848 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3074
timestamp 1569533753
transform 1 0 3976 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3075
timestamp 1569533753
transform 1 0 3912 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3076
timestamp 1569533753
transform 1 0 3784 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3077
timestamp 1569533753
transform 1 0 3976 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3078
timestamp 1569533753
transform 1 0 4040 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3079
timestamp 1569533753
transform 1 0 3784 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3080
timestamp 1569533753
transform 1 0 3912 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3081
timestamp 1569533753
transform 1 0 4040 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3082
timestamp 1569533753
transform 1 0 3784 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3083
timestamp 1569533753
transform 1 0 3848 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3084
timestamp 1569533753
transform 1 0 4040 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3085
timestamp 1569533753
transform 1 0 4040 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3086
timestamp 1569533753
transform 1 0 3912 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3087
timestamp 1569533753
transform 1 0 3848 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3088
timestamp 1569533753
transform 1 0 3784 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3089
timestamp 1569533753
transform 1 0 3976 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3090
timestamp 1569533753
transform 1 0 3912 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3091
timestamp 1569533753
transform 1 0 4104 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3092
timestamp 1569533753
transform 1 0 4104 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3093
timestamp 1569533753
transform 1 0 4232 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3094
timestamp 1569533753
transform 1 0 4104 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3095
timestamp 1569533753
transform 1 0 4232 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3096
timestamp 1569533753
transform 1 0 4168 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3097
timestamp 1569533753
transform 1 0 4296 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3098
timestamp 1569533753
transform 1 0 4168 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3099
timestamp 1569533753
transform 1 0 4232 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3100
timestamp 1569533753
transform 1 0 4296 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3101
timestamp 1569533753
transform 1 0 4168 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3102
timestamp 1569533753
transform 1 0 4104 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3103
timestamp 1569533753
transform 1 0 4104 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3104
timestamp 1569533753
transform 1 0 4168 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3105
timestamp 1569533753
transform 1 0 4168 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3106
timestamp 1569533753
transform 1 0 4232 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3107
timestamp 1569533753
transform 1 0 4232 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3108
timestamp 1569533753
transform 1 0 4296 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3109
timestamp 1569533753
transform 1 0 4296 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3110
timestamp 1569533753
transform 1 0 4296 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3111
timestamp 1569533753
transform 1 0 4168 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3112
timestamp 1569533753
transform 1 0 4232 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3113
timestamp 1569533753
transform 1 0 4104 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3114
timestamp 1569533753
transform 1 0 4104 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3115
timestamp 1569533753
transform 1 0 4232 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3116
timestamp 1569533753
transform 1 0 4168 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3117
timestamp 1569533753
transform 1 0 4232 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3118
timestamp 1569533753
transform 1 0 4104 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3119
timestamp 1569533753
transform 1 0 4104 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3120
timestamp 1569533753
transform 1 0 4168 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3121
timestamp 1569533753
transform 1 0 4104 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3122
timestamp 1569533753
transform 1 0 4296 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3123
timestamp 1569533753
transform 1 0 4232 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3124
timestamp 1569533753
transform 1 0 4168 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3125
timestamp 1569533753
transform 1 0 4232 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3126
timestamp 1569533753
transform 1 0 4296 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3127
timestamp 1569533753
transform 1 0 4296 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3128
timestamp 1569533753
transform 1 0 4296 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3129
timestamp 1569533753
transform 1 0 4296 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3130
timestamp 1569533753
transform 1 0 4168 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3131
timestamp 1569533753
transform 1 0 3848 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3132
timestamp 1569533753
transform 1 0 4040 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3133
timestamp 1569533753
transform 1 0 3912 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3134
timestamp 1569533753
transform 1 0 3848 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3135
timestamp 1569533753
transform 1 0 3784 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3136
timestamp 1569533753
transform 1 0 3784 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3137
timestamp 1569533753
transform 1 0 3848 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3138
timestamp 1569533753
transform 1 0 3784 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3139
timestamp 1569533753
transform 1 0 3912 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3140
timestamp 1569533753
transform 1 0 3976 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3141
timestamp 1569533753
transform 1 0 3912 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3142
timestamp 1569533753
transform 1 0 3848 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3143
timestamp 1569533753
transform 1 0 3976 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3144
timestamp 1569533753
transform 1 0 3976 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3145
timestamp 1569533753
transform 1 0 3784 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3146
timestamp 1569533753
transform 1 0 3976 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3147
timestamp 1569533753
transform 1 0 3976 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3148
timestamp 1569533753
transform 1 0 3784 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3149
timestamp 1569533753
transform 1 0 4040 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3150
timestamp 1569533753
transform 1 0 3912 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3151
timestamp 1569533753
transform 1 0 4040 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3152
timestamp 1569533753
transform 1 0 3848 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3153
timestamp 1569533753
transform 1 0 4040 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3154
timestamp 1569533753
transform 1 0 3912 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3155
timestamp 1569533753
transform 1 0 4040 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3156
timestamp 1569533753
transform 1 0 4040 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3157
timestamp 1569533753
transform 1 0 3784 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3158
timestamp 1569533753
transform 1 0 3784 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3159
timestamp 1569533753
transform 1 0 3784 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3160
timestamp 1569533753
transform 1 0 3784 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3161
timestamp 1569533753
transform 1 0 4040 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3162
timestamp 1569533753
transform 1 0 3912 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3163
timestamp 1569533753
transform 1 0 3912 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3164
timestamp 1569533753
transform 1 0 3976 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3165
timestamp 1569533753
transform 1 0 3976 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3166
timestamp 1569533753
transform 1 0 3976 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3167
timestamp 1569533753
transform 1 0 3848 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3168
timestamp 1569533753
transform 1 0 3976 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3169
timestamp 1569533753
transform 1 0 3976 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3170
timestamp 1569533753
transform 1 0 3848 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3171
timestamp 1569533753
transform 1 0 3848 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3172
timestamp 1569533753
transform 1 0 3848 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3173
timestamp 1569533753
transform 1 0 4040 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3174
timestamp 1569533753
transform 1 0 3912 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3175
timestamp 1569533753
transform 1 0 4040 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3176
timestamp 1569533753
transform 1 0 3912 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3177
timestamp 1569533753
transform 1 0 3912 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3178
timestamp 1569533753
transform 1 0 3848 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3179
timestamp 1569533753
transform 1 0 4040 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3180
timestamp 1569533753
transform 1 0 3784 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3181
timestamp 1569533753
transform 1 0 4232 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3182
timestamp 1569533753
transform 1 0 4232 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3183
timestamp 1569533753
transform 1 0 4232 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3184
timestamp 1569533753
transform 1 0 4104 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3185
timestamp 1569533753
transform 1 0 4296 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3186
timestamp 1569533753
transform 1 0 4296 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3187
timestamp 1569533753
transform 1 0 4296 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3188
timestamp 1569533753
transform 1 0 4104 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3189
timestamp 1569533753
transform 1 0 4168 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3190
timestamp 1569533753
transform 1 0 4104 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3191
timestamp 1569533753
transform 1 0 4104 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3192
timestamp 1569533753
transform 1 0 4296 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3193
timestamp 1569533753
transform 1 0 4296 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3194
timestamp 1569533753
transform 1 0 4168 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3195
timestamp 1569533753
transform 1 0 4168 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3196
timestamp 1569533753
transform 1 0 4232 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3197
timestamp 1569533753
transform 1 0 4232 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3198
timestamp 1569533753
transform 1 0 4168 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3199
timestamp 1569533753
transform 1 0 4168 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3200
timestamp 1569533753
transform 1 0 4104 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3201
timestamp 1569533753
transform 1 0 4744 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3202
timestamp 1569533753
transform 1 0 4744 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3203
timestamp 1569533753
transform 1 0 4744 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3204
timestamp 1569533753
transform 1 0 4744 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3205
timestamp 1569533753
transform 1 0 4744 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3206
timestamp 1569533753
transform 1 0 4808 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3207
timestamp 1569533753
transform 1 0 4808 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3208
timestamp 1569533753
transform 1 0 4808 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3209
timestamp 1569533753
transform 1 0 4872 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3210
timestamp 1569533753
transform 1 0 4680 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3211
timestamp 1569533753
transform 1 0 4808 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3212
timestamp 1569533753
transform 1 0 4808 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3213
timestamp 1569533753
transform 1 0 4872 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3214
timestamp 1569533753
transform 1 0 4680 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3215
timestamp 1569533753
transform 1 0 4680 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3216
timestamp 1569533753
transform 1 0 4872 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3217
timestamp 1569533753
transform 1 0 4680 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3218
timestamp 1569533753
transform 1 0 4680 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3219
timestamp 1569533753
transform 1 0 4872 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3220
timestamp 1569533753
transform 1 0 4872 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3221
timestamp 1569533753
transform 1 0 4552 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3222
timestamp 1569533753
transform 1 0 4488 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3223
timestamp 1569533753
transform 1 0 4488 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3224
timestamp 1569533753
transform 1 0 4488 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3225
timestamp 1569533753
transform 1 0 4616 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3226
timestamp 1569533753
transform 1 0 4552 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3227
timestamp 1569533753
transform 1 0 4424 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3228
timestamp 1569533753
transform 1 0 4616 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3229
timestamp 1569533753
transform 1 0 4616 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3230
timestamp 1569533753
transform 1 0 4616 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3231
timestamp 1569533753
transform 1 0 4616 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3232
timestamp 1569533753
transform 1 0 4552 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3233
timestamp 1569533753
transform 1 0 4552 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3234
timestamp 1569533753
transform 1 0 4552 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3235
timestamp 1569533753
transform 1 0 4424 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3236
timestamp 1569533753
transform 1 0 4424 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3237
timestamp 1569533753
transform 1 0 4424 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3238
timestamp 1569533753
transform 1 0 4424 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3239
timestamp 1569533753
transform 1 0 4488 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3240
timestamp 1569533753
transform 1 0 4488 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3241
timestamp 1569533753
transform 1 0 4552 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3242
timestamp 1569533753
transform 1 0 4616 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3243
timestamp 1569533753
transform 1 0 4616 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3244
timestamp 1569533753
transform 1 0 4424 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3245
timestamp 1569533753
transform 1 0 4424 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3246
timestamp 1569533753
transform 1 0 4424 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3247
timestamp 1569533753
transform 1 0 4424 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3248
timestamp 1569533753
transform 1 0 4424 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3249
timestamp 1569533753
transform 1 0 4488 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3250
timestamp 1569533753
transform 1 0 4616 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3251
timestamp 1569533753
transform 1 0 4616 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3252
timestamp 1569533753
transform 1 0 4616 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3253
timestamp 1569533753
transform 1 0 4488 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3254
timestamp 1569533753
transform 1 0 4488 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3255
timestamp 1569533753
transform 1 0 4488 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3256
timestamp 1569533753
transform 1 0 4488 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3257
timestamp 1569533753
transform 1 0 4552 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3258
timestamp 1569533753
transform 1 0 4552 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3259
timestamp 1569533753
transform 1 0 4552 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3260
timestamp 1569533753
transform 1 0 4552 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3261
timestamp 1569533753
transform 1 0 4680 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3262
timestamp 1569533753
transform 1 0 4680 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3263
timestamp 1569533753
transform 1 0 4744 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3264
timestamp 1569533753
transform 1 0 4744 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3265
timestamp 1569533753
transform 1 0 4808 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3266
timestamp 1569533753
transform 1 0 4808 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3267
timestamp 1569533753
transform 1 0 4872 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3268
timestamp 1569533753
transform 1 0 4872 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3269
timestamp 1569533753
transform 1 0 4680 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3270
timestamp 1569533753
transform 1 0 4680 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3271
timestamp 1569533753
transform 1 0 4680 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3272
timestamp 1569533753
transform 1 0 4744 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3273
timestamp 1569533753
transform 1 0 4744 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3274
timestamp 1569533753
transform 1 0 4744 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3275
timestamp 1569533753
transform 1 0 4808 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3276
timestamp 1569533753
transform 1 0 4808 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3277
timestamp 1569533753
transform 1 0 4808 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3278
timestamp 1569533753
transform 1 0 4872 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3279
timestamp 1569533753
transform 1 0 4872 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3280
timestamp 1569533753
transform 1 0 4872 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3281
timestamp 1569533753
transform 1 0 4360 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3282
timestamp 1569533753
transform 1 0 4360 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3283
timestamp 1569533753
transform 1 0 4360 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3284
timestamp 1569533753
transform 1 0 4360 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3285
timestamp 1569533753
transform 1 0 4360 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3286
timestamp 1569533753
transform 1 0 4360 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3287
timestamp 1569533753
transform 1 0 4360 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3288
timestamp 1569533753
transform 1 0 4360 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3289
timestamp 1569533753
transform 1 0 4360 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3290
timestamp 1569533753
transform 1 0 4360 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3291
timestamp 1569533753
transform 1 0 4360 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3292
timestamp 1569533753
transform 1 0 4360 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3293
timestamp 1569533753
transform 1 0 4360 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3294
timestamp 1569533753
transform 1 0 4360 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3295
timestamp 1569533753
transform 1 0 4360 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3296
timestamp 1569533753
transform 1 0 4360 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3297
timestamp 1569533753
transform 1 0 4360 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3298
timestamp 1569533753
transform 1 0 4360 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3299
timestamp 1569533753
transform 1 0 4360 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3300
timestamp 1569533753
transform 1 0 3464 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3301
timestamp 1569533753
transform 1 0 3720 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3302
timestamp 1569533753
transform 1 0 3592 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3303
timestamp 1569533753
transform 1 0 3720 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3304
timestamp 1569533753
transform 1 0 3464 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3305
timestamp 1569533753
transform 1 0 3592 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3306
timestamp 1569533753
transform 1 0 3464 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3307
timestamp 1569533753
transform 1 0 3656 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3308
timestamp 1569533753
transform 1 0 3528 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3309
timestamp 1569533753
transform 1 0 3656 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3310
timestamp 1569533753
transform 1 0 3720 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3311
timestamp 1569533753
transform 1 0 3528 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3312
timestamp 1569533753
transform 1 0 3592 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3313
timestamp 1569533753
transform 1 0 3528 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3314
timestamp 1569533753
transform 1 0 3528 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3315
timestamp 1569533753
transform 1 0 3656 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3316
timestamp 1569533753
transform 1 0 3656 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3317
timestamp 1569533753
transform 1 0 3592 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3318
timestamp 1569533753
transform 1 0 3464 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3319
timestamp 1569533753
transform 1 0 3720 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3320
timestamp 1569533753
transform 1 0 3336 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3321
timestamp 1569533753
transform 1 0 3336 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3322
timestamp 1569533753
transform 1 0 3208 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3323
timestamp 1569533753
transform 1 0 3336 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3324
timestamp 1569533753
transform 1 0 3400 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3325
timestamp 1569533753
transform 1 0 3144 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3326
timestamp 1569533753
transform 1 0 3400 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3327
timestamp 1569533753
transform 1 0 3208 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3328
timestamp 1569533753
transform 1 0 3272 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3329
timestamp 1569533753
transform 1 0 3400 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3330
timestamp 1569533753
transform 1 0 3144 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3331
timestamp 1569533753
transform 1 0 3144 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3332
timestamp 1569533753
transform 1 0 3208 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3333
timestamp 1569533753
transform 1 0 3144 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3334
timestamp 1569533753
transform 1 0 3400 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3335
timestamp 1569533753
transform 1 0 3272 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3336
timestamp 1569533753
transform 1 0 3208 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3337
timestamp 1569533753
transform 1 0 3272 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3338
timestamp 1569533753
transform 1 0 3336 0 1 2568
box -8 -8 8 8
use VIA1$3  VIA1$3_3339
timestamp 1569533753
transform 1 0 3272 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3340
timestamp 1569533753
transform 1 0 3336 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3341
timestamp 1569533753
transform 1 0 3208 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3342
timestamp 1569533753
transform 1 0 3272 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3343
timestamp 1569533753
transform 1 0 3208 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3344
timestamp 1569533753
transform 1 0 3144 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3345
timestamp 1569533753
transform 1 0 3400 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3346
timestamp 1569533753
transform 1 0 3400 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3347
timestamp 1569533753
transform 1 0 3272 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3348
timestamp 1569533753
transform 1 0 3336 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3349
timestamp 1569533753
transform 1 0 3272 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3350
timestamp 1569533753
transform 1 0 3208 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3351
timestamp 1569533753
transform 1 0 3336 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3352
timestamp 1569533753
transform 1 0 3272 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3353
timestamp 1569533753
transform 1 0 3336 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3354
timestamp 1569533753
transform 1 0 3208 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3355
timestamp 1569533753
transform 1 0 3400 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3356
timestamp 1569533753
transform 1 0 3400 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3357
timestamp 1569533753
transform 1 0 3144 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3358
timestamp 1569533753
transform 1 0 3144 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3359
timestamp 1569533753
transform 1 0 3400 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3360
timestamp 1569533753
transform 1 0 3144 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3361
timestamp 1569533753
transform 1 0 3336 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3362
timestamp 1569533753
transform 1 0 3144 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3363
timestamp 1569533753
transform 1 0 3272 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3364
timestamp 1569533753
transform 1 0 3208 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3365
timestamp 1569533753
transform 1 0 3592 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3366
timestamp 1569533753
transform 1 0 3720 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3367
timestamp 1569533753
transform 1 0 3464 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3368
timestamp 1569533753
transform 1 0 3720 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3369
timestamp 1569533753
transform 1 0 3464 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3370
timestamp 1569533753
transform 1 0 3656 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3371
timestamp 1569533753
transform 1 0 3528 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3372
timestamp 1569533753
transform 1 0 3528 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3373
timestamp 1569533753
transform 1 0 3592 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3374
timestamp 1569533753
transform 1 0 3592 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3375
timestamp 1569533753
transform 1 0 3528 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3376
timestamp 1569533753
transform 1 0 3656 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3377
timestamp 1569533753
transform 1 0 3656 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3378
timestamp 1569533753
transform 1 0 3656 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3379
timestamp 1569533753
transform 1 0 3528 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3380
timestamp 1569533753
transform 1 0 3528 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3381
timestamp 1569533753
transform 1 0 3464 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3382
timestamp 1569533753
transform 1 0 3720 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3383
timestamp 1569533753
transform 1 0 3592 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3384
timestamp 1569533753
transform 1 0 3464 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3385
timestamp 1569533753
transform 1 0 3720 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3386
timestamp 1569533753
transform 1 0 3464 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3387
timestamp 1569533753
transform 1 0 3720 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3388
timestamp 1569533753
transform 1 0 3656 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3389
timestamp 1569533753
transform 1 0 3592 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3390
timestamp 1569533753
transform 1 0 3080 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3391
timestamp 1569533753
transform 1 0 3080 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3392
timestamp 1569533753
transform 1 0 2952 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3393
timestamp 1569533753
transform 1 0 2696 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3394
timestamp 1569533753
transform 1 0 2952 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3395
timestamp 1569533753
transform 1 0 3016 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3396
timestamp 1569533753
transform 1 0 2888 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3397
timestamp 1569533753
transform 1 0 3016 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3398
timestamp 1569533753
transform 1 0 2760 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3399
timestamp 1569533753
transform 1 0 3016 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3400
timestamp 1569533753
transform 1 0 2952 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3401
timestamp 1569533753
transform 1 0 3080 0 1 2696
box -8 -8 8 8
use VIA1$3  VIA1$3_3402
timestamp 1569533753
transform 1 0 2824 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3403
timestamp 1569533753
transform 1 0 3080 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3404
timestamp 1569533753
transform 1 0 2824 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3405
timestamp 1569533753
transform 1 0 3080 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3406
timestamp 1569533753
transform 1 0 2952 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3407
timestamp 1569533753
transform 1 0 2952 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3408
timestamp 1569533753
transform 1 0 2888 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3409
timestamp 1569533753
transform 1 0 2888 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3410
timestamp 1569533753
transform 1 0 2632 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3411
timestamp 1569533753
transform 1 0 2952 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3412
timestamp 1569533753
transform 1 0 2696 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3413
timestamp 1569533753
transform 1 0 2888 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3414
timestamp 1569533753
transform 1 0 3016 0 1 2760
box -8 -8 8 8
use VIA1$3  VIA1$3_3415
timestamp 1569533753
transform 1 0 3016 0 1 2824
box -8 -8 8 8
use VIA1$3  VIA1$3_3416
timestamp 1569533753
transform 1 0 3016 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3417
timestamp 1569533753
transform 1 0 2760 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3418
timestamp 1569533753
transform 1 0 3016 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3419
timestamp 1569533753
transform 1 0 2760 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3420
timestamp 1569533753
transform 1 0 2888 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3421
timestamp 1569533753
transform 1 0 3080 0 1 2888
box -8 -8 8 8
use VIA1$3  VIA1$3_3422
timestamp 1569533753
transform 1 0 2824 0 1 2952
box -8 -8 8 8
use VIA1$3  VIA1$3_3423
timestamp 1569533753
transform 1 0 3080 0 1 3016
box -8 -8 8 8
use VIA1$3  VIA1$3_3424
timestamp 1569533753
transform 1 0 2824 0 1 3080
box -8 -8 8 8
use VIA1$3  VIA1$3_3425
timestamp 1569533753
transform 1 0 3080 0 1 2632
box -8 -8 8 8
use VIA1$3  VIA1$3_3426
timestamp 1569533753
transform 1 0 2888 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3427
timestamp 1569533753
transform 1 0 3016 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3428
timestamp 1569533753
transform 1 0 3080 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3429
timestamp 1569533753
transform 1 0 2888 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3430
timestamp 1569533753
transform 1 0 2824 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3431
timestamp 1569533753
transform 1 0 2888 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3432
timestamp 1569533753
transform 1 0 2888 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3433
timestamp 1569533753
transform 1 0 2888 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3434
timestamp 1569533753
transform 1 0 3016 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3435
timestamp 1569533753
transform 1 0 3080 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3436
timestamp 1569533753
transform 1 0 3080 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3437
timestamp 1569533753
transform 1 0 2952 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3438
timestamp 1569533753
transform 1 0 2952 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3439
timestamp 1569533753
transform 1 0 2952 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3440
timestamp 1569533753
transform 1 0 2952 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3441
timestamp 1569533753
transform 1 0 3016 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3442
timestamp 1569533753
transform 1 0 3016 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3443
timestamp 1569533753
transform 1 0 3080 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3444
timestamp 1569533753
transform 1 0 2824 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3445
timestamp 1569533753
transform 1 0 2824 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3446
timestamp 1569533753
transform 1 0 3016 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3447
timestamp 1569533753
transform 1 0 2824 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3448
timestamp 1569533753
transform 1 0 2824 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3449
timestamp 1569533753
transform 1 0 2952 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3450
timestamp 1569533753
transform 1 0 3080 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3451
timestamp 1569533753
transform 1 0 2696 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3452
timestamp 1569533753
transform 1 0 2568 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3453
timestamp 1569533753
transform 1 0 2760 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3454
timestamp 1569533753
transform 1 0 2632 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3455
timestamp 1569533753
transform 1 0 2696 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3456
timestamp 1569533753
transform 1 0 2696 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3457
timestamp 1569533753
transform 1 0 2696 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3458
timestamp 1569533753
transform 1 0 2696 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3459
timestamp 1569533753
transform 1 0 2632 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3460
timestamp 1569533753
transform 1 0 2632 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3461
timestamp 1569533753
transform 1 0 2568 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3462
timestamp 1569533753
transform 1 0 2760 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3463
timestamp 1569533753
transform 1 0 2760 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3464
timestamp 1569533753
transform 1 0 2760 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3465
timestamp 1569533753
transform 1 0 2632 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3466
timestamp 1569533753
transform 1 0 2760 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3467
timestamp 1569533753
transform 1 0 2568 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3468
timestamp 1569533753
transform 1 0 2568 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3469
timestamp 1569533753
transform 1 0 2568 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3470
timestamp 1569533753
transform 1 0 2632 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3471
timestamp 1569533753
transform 1 0 2568 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3472
timestamp 1569533753
transform 1 0 2632 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3473
timestamp 1569533753
transform 1 0 2632 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3474
timestamp 1569533753
transform 1 0 2632 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3475
timestamp 1569533753
transform 1 0 2760 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3476
timestamp 1569533753
transform 1 0 2760 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3477
timestamp 1569533753
transform 1 0 2696 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3478
timestamp 1569533753
transform 1 0 2696 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3479
timestamp 1569533753
transform 1 0 2760 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3480
timestamp 1569533753
transform 1 0 2760 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3481
timestamp 1569533753
transform 1 0 2760 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3482
timestamp 1569533753
transform 1 0 2632 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3483
timestamp 1569533753
transform 1 0 2568 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3484
timestamp 1569533753
transform 1 0 2632 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3485
timestamp 1569533753
transform 1 0 2568 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3486
timestamp 1569533753
transform 1 0 2568 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3487
timestamp 1569533753
transform 1 0 2568 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3488
timestamp 1569533753
transform 1 0 2696 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3489
timestamp 1569533753
transform 1 0 2696 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3490
timestamp 1569533753
transform 1 0 2696 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3491
timestamp 1569533753
transform 1 0 3080 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3492
timestamp 1569533753
transform 1 0 3016 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3493
timestamp 1569533753
transform 1 0 3080 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3494
timestamp 1569533753
transform 1 0 3016 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3495
timestamp 1569533753
transform 1 0 2824 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3496
timestamp 1569533753
transform 1 0 2824 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3497
timestamp 1569533753
transform 1 0 2888 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3498
timestamp 1569533753
transform 1 0 2888 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3499
timestamp 1569533753
transform 1 0 3080 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3500
timestamp 1569533753
transform 1 0 2952 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3501
timestamp 1569533753
transform 1 0 2952 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3502
timestamp 1569533753
transform 1 0 3080 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3503
timestamp 1569533753
transform 1 0 3016 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3504
timestamp 1569533753
transform 1 0 3080 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3505
timestamp 1569533753
transform 1 0 2824 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3506
timestamp 1569533753
transform 1 0 2824 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3507
timestamp 1569533753
transform 1 0 2824 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3508
timestamp 1569533753
transform 1 0 2888 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3509
timestamp 1569533753
transform 1 0 2888 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3510
timestamp 1569533753
transform 1 0 2888 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3511
timestamp 1569533753
transform 1 0 3016 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3512
timestamp 1569533753
transform 1 0 2952 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3513
timestamp 1569533753
transform 1 0 2952 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3514
timestamp 1569533753
transform 1 0 2952 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3515
timestamp 1569533753
transform 1 0 3016 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3516
timestamp 1569533753
transform 1 0 3656 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3517
timestamp 1569533753
transform 1 0 3720 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3518
timestamp 1569533753
transform 1 0 3720 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3519
timestamp 1569533753
transform 1 0 3720 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3520
timestamp 1569533753
transform 1 0 3720 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3521
timestamp 1569533753
transform 1 0 3720 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3522
timestamp 1569533753
transform 1 0 3464 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3523
timestamp 1569533753
transform 1 0 3464 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3524
timestamp 1569533753
transform 1 0 3464 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3525
timestamp 1569533753
transform 1 0 3464 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3526
timestamp 1569533753
transform 1 0 3464 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3527
timestamp 1569533753
transform 1 0 3528 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3528
timestamp 1569533753
transform 1 0 3528 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3529
timestamp 1569533753
transform 1 0 3528 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3530
timestamp 1569533753
transform 1 0 3528 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3531
timestamp 1569533753
transform 1 0 3528 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3532
timestamp 1569533753
transform 1 0 3592 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3533
timestamp 1569533753
transform 1 0 3592 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3534
timestamp 1569533753
transform 1 0 3592 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3535
timestamp 1569533753
transform 1 0 3592 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3536
timestamp 1569533753
transform 1 0 3592 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3537
timestamp 1569533753
transform 1 0 3656 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3538
timestamp 1569533753
transform 1 0 3656 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3539
timestamp 1569533753
transform 1 0 3656 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3540
timestamp 1569533753
transform 1 0 3656 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3541
timestamp 1569533753
transform 1 0 3208 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3542
timestamp 1569533753
transform 1 0 3272 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3543
timestamp 1569533753
transform 1 0 3336 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3544
timestamp 1569533753
transform 1 0 3400 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3545
timestamp 1569533753
transform 1 0 3336 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3546
timestamp 1569533753
transform 1 0 3336 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3547
timestamp 1569533753
transform 1 0 3336 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3548
timestamp 1569533753
transform 1 0 3336 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3549
timestamp 1569533753
transform 1 0 3144 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3550
timestamp 1569533753
transform 1 0 3400 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3551
timestamp 1569533753
transform 1 0 3400 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3552
timestamp 1569533753
transform 1 0 3400 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3553
timestamp 1569533753
transform 1 0 3400 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3554
timestamp 1569533753
transform 1 0 3208 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3555
timestamp 1569533753
transform 1 0 3208 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3556
timestamp 1569533753
transform 1 0 3208 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3557
timestamp 1569533753
transform 1 0 3208 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3558
timestamp 1569533753
transform 1 0 3144 0 1 3144
box -8 -8 8 8
use VIA1$3  VIA1$3_3559
timestamp 1569533753
transform 1 0 3272 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3560
timestamp 1569533753
transform 1 0 3272 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3561
timestamp 1569533753
transform 1 0 3272 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3562
timestamp 1569533753
transform 1 0 3272 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_3563
timestamp 1569533753
transform 1 0 3144 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_3564
timestamp 1569533753
transform 1 0 3144 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_3565
timestamp 1569533753
transform 1 0 3144 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_3566
timestamp 1569533753
transform 1 0 3336 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3567
timestamp 1569533753
transform 1 0 3336 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3568
timestamp 1569533753
transform 1 0 3400 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3569
timestamp 1569533753
transform 1 0 3400 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3570
timestamp 1569533753
transform 1 0 3272 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3571
timestamp 1569533753
transform 1 0 3272 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3572
timestamp 1569533753
transform 1 0 3336 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3573
timestamp 1569533753
transform 1 0 3336 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3574
timestamp 1569533753
transform 1 0 3336 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3575
timestamp 1569533753
transform 1 0 3272 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3576
timestamp 1569533753
transform 1 0 3272 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3577
timestamp 1569533753
transform 1 0 3400 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3578
timestamp 1569533753
transform 1 0 3400 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3579
timestamp 1569533753
transform 1 0 3400 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3580
timestamp 1569533753
transform 1 0 3272 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3581
timestamp 1569533753
transform 1 0 3144 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3582
timestamp 1569533753
transform 1 0 3144 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3583
timestamp 1569533753
transform 1 0 3144 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3584
timestamp 1569533753
transform 1 0 3208 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3585
timestamp 1569533753
transform 1 0 3208 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3586
timestamp 1569533753
transform 1 0 3208 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3587
timestamp 1569533753
transform 1 0 3144 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3588
timestamp 1569533753
transform 1 0 3144 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3589
timestamp 1569533753
transform 1 0 3208 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3590
timestamp 1569533753
transform 1 0 3208 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3591
timestamp 1569533753
transform 1 0 3464 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3592
timestamp 1569533753
transform 1 0 3464 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3593
timestamp 1569533753
transform 1 0 3528 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3594
timestamp 1569533753
transform 1 0 3528 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3595
timestamp 1569533753
transform 1 0 3592 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3596
timestamp 1569533753
transform 1 0 3592 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3597
timestamp 1569533753
transform 1 0 3720 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3598
timestamp 1569533753
transform 1 0 3464 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3599
timestamp 1569533753
transform 1 0 3464 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3600
timestamp 1569533753
transform 1 0 3464 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3601
timestamp 1569533753
transform 1 0 3528 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3602
timestamp 1569533753
transform 1 0 3528 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3603
timestamp 1569533753
transform 1 0 3528 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3604
timestamp 1569533753
transform 1 0 3592 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3605
timestamp 1569533753
transform 1 0 3592 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3606
timestamp 1569533753
transform 1 0 3592 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3607
timestamp 1569533753
transform 1 0 3720 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3608
timestamp 1569533753
transform 1 0 3720 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3609
timestamp 1569533753
transform 1 0 3656 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3610
timestamp 1569533753
transform 1 0 3656 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3611
timestamp 1569533753
transform 1 0 3720 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_3612
timestamp 1569533753
transform 1 0 3720 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_3613
timestamp 1569533753
transform 1 0 3656 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_3614
timestamp 1569533753
transform 1 0 3656 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_3615
timestamp 1569533753
transform 1 0 3656 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_3616
timestamp 1569533753
transform 1 0 3592 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3617
timestamp 1569533753
transform 1 0 3720 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3618
timestamp 1569533753
transform 1 0 3720 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3619
timestamp 1569533753
transform 1 0 3720 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3620
timestamp 1569533753
transform 1 0 3592 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3621
timestamp 1569533753
transform 1 0 3592 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3622
timestamp 1569533753
transform 1 0 3656 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3623
timestamp 1569533753
transform 1 0 3720 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3624
timestamp 1569533753
transform 1 0 3656 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3625
timestamp 1569533753
transform 1 0 3592 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3626
timestamp 1569533753
transform 1 0 3528 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3627
timestamp 1569533753
transform 1 0 3464 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3628
timestamp 1569533753
transform 1 0 3464 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3629
timestamp 1569533753
transform 1 0 3464 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3630
timestamp 1569533753
transform 1 0 3656 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3631
timestamp 1569533753
transform 1 0 3464 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3632
timestamp 1569533753
transform 1 0 3656 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3633
timestamp 1569533753
transform 1 0 3464 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3634
timestamp 1569533753
transform 1 0 3528 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3635
timestamp 1569533753
transform 1 0 3720 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3636
timestamp 1569533753
transform 1 0 3528 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3637
timestamp 1569533753
transform 1 0 3528 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3638
timestamp 1569533753
transform 1 0 3528 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3639
timestamp 1569533753
transform 1 0 3656 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3640
timestamp 1569533753
transform 1 0 3592 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3641
timestamp 1569533753
transform 1 0 3336 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3642
timestamp 1569533753
transform 1 0 3336 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3643
timestamp 1569533753
transform 1 0 3336 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3644
timestamp 1569533753
transform 1 0 3272 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3645
timestamp 1569533753
transform 1 0 3336 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3646
timestamp 1569533753
transform 1 0 3272 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3647
timestamp 1569533753
transform 1 0 3400 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3648
timestamp 1569533753
transform 1 0 3144 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3649
timestamp 1569533753
transform 1 0 3400 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3650
timestamp 1569533753
transform 1 0 3400 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3651
timestamp 1569533753
transform 1 0 3272 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3652
timestamp 1569533753
transform 1 0 3144 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3653
timestamp 1569533753
transform 1 0 3400 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3654
timestamp 1569533753
transform 1 0 3400 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3655
timestamp 1569533753
transform 1 0 3144 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3656
timestamp 1569533753
transform 1 0 3144 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3657
timestamp 1569533753
transform 1 0 3272 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3658
timestamp 1569533753
transform 1 0 3208 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3659
timestamp 1569533753
transform 1 0 3208 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3660
timestamp 1569533753
transform 1 0 3336 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3661
timestamp 1569533753
transform 1 0 3208 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3662
timestamp 1569533753
transform 1 0 3208 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3663
timestamp 1569533753
transform 1 0 3208 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3664
timestamp 1569533753
transform 1 0 3272 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3665
timestamp 1569533753
transform 1 0 3144 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3666
timestamp 1569533753
transform 1 0 3272 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3667
timestamp 1569533753
transform 1 0 3272 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3668
timestamp 1569533753
transform 1 0 3272 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3669
timestamp 1569533753
transform 1 0 3272 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3670
timestamp 1569533753
transform 1 0 3144 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3671
timestamp 1569533753
transform 1 0 3336 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3672
timestamp 1569533753
transform 1 0 3336 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3673
timestamp 1569533753
transform 1 0 3336 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3674
timestamp 1569533753
transform 1 0 3336 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3675
timestamp 1569533753
transform 1 0 3208 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3676
timestamp 1569533753
transform 1 0 3144 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3677
timestamp 1569533753
transform 1 0 3400 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3678
timestamp 1569533753
transform 1 0 3400 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3679
timestamp 1569533753
transform 1 0 3400 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3680
timestamp 1569533753
transform 1 0 3400 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3681
timestamp 1569533753
transform 1 0 3208 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3682
timestamp 1569533753
transform 1 0 3208 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3683
timestamp 1569533753
transform 1 0 3144 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3684
timestamp 1569533753
transform 1 0 3144 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3685
timestamp 1569533753
transform 1 0 3208 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3686
timestamp 1569533753
transform 1 0 3592 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3687
timestamp 1569533753
transform 1 0 3656 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3688
timestamp 1569533753
transform 1 0 3656 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3689
timestamp 1569533753
transform 1 0 3656 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3690
timestamp 1569533753
transform 1 0 3464 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3691
timestamp 1569533753
transform 1 0 3656 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3692
timestamp 1569533753
transform 1 0 3464 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3693
timestamp 1569533753
transform 1 0 3464 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3694
timestamp 1569533753
transform 1 0 3464 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3695
timestamp 1569533753
transform 1 0 3720 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3696
timestamp 1569533753
transform 1 0 3528 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3697
timestamp 1569533753
transform 1 0 3720 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3698
timestamp 1569533753
transform 1 0 3528 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3699
timestamp 1569533753
transform 1 0 3528 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3700
timestamp 1569533753
transform 1 0 3720 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3701
timestamp 1569533753
transform 1 0 3528 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3702
timestamp 1569533753
transform 1 0 3720 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3703
timestamp 1569533753
transform 1 0 3592 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3704
timestamp 1569533753
transform 1 0 3592 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3705
timestamp 1569533753
transform 1 0 3592 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3706
timestamp 1569533753
transform 1 0 2824 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3707
timestamp 1569533753
transform 1 0 3080 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3708
timestamp 1569533753
transform 1 0 2824 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3709
timestamp 1569533753
transform 1 0 2824 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3710
timestamp 1569533753
transform 1 0 2824 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3711
timestamp 1569533753
transform 1 0 2824 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3712
timestamp 1569533753
transform 1 0 2888 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3713
timestamp 1569533753
transform 1 0 2888 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3714
timestamp 1569533753
transform 1 0 2888 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3715
timestamp 1569533753
transform 1 0 2888 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3716
timestamp 1569533753
transform 1 0 2952 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3717
timestamp 1569533753
transform 1 0 2952 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3718
timestamp 1569533753
transform 1 0 2952 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3719
timestamp 1569533753
transform 1 0 2952 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3720
timestamp 1569533753
transform 1 0 2888 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3721
timestamp 1569533753
transform 1 0 3016 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3722
timestamp 1569533753
transform 1 0 3016 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3723
timestamp 1569533753
transform 1 0 3016 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3724
timestamp 1569533753
transform 1 0 3016 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3725
timestamp 1569533753
transform 1 0 3016 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3726
timestamp 1569533753
transform 1 0 3080 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3727
timestamp 1569533753
transform 1 0 3080 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3728
timestamp 1569533753
transform 1 0 2952 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3729
timestamp 1569533753
transform 1 0 3080 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3730
timestamp 1569533753
transform 1 0 3080 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3731
timestamp 1569533753
transform 1 0 2696 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3732
timestamp 1569533753
transform 1 0 2696 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3733
timestamp 1569533753
transform 1 0 2696 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3734
timestamp 1569533753
transform 1 0 2696 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3735
timestamp 1569533753
transform 1 0 2760 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3736
timestamp 1569533753
transform 1 0 2760 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3737
timestamp 1569533753
transform 1 0 2760 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3738
timestamp 1569533753
transform 1 0 2760 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3739
timestamp 1569533753
transform 1 0 2696 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3740
timestamp 1569533753
transform 1 0 2568 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3741
timestamp 1569533753
transform 1 0 2568 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3742
timestamp 1569533753
transform 1 0 2760 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3743
timestamp 1569533753
transform 1 0 2568 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3744
timestamp 1569533753
transform 1 0 2568 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3745
timestamp 1569533753
transform 1 0 2632 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3746
timestamp 1569533753
transform 1 0 2568 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3747
timestamp 1569533753
transform 1 0 2632 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3748
timestamp 1569533753
transform 1 0 2632 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3749
timestamp 1569533753
transform 1 0 2632 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3750
timestamp 1569533753
transform 1 0 2632 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3751
timestamp 1569533753
transform 1 0 2696 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3752
timestamp 1569533753
transform 1 0 2696 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3753
timestamp 1569533753
transform 1 0 2696 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3754
timestamp 1569533753
transform 1 0 2696 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3755
timestamp 1569533753
transform 1 0 2760 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3756
timestamp 1569533753
transform 1 0 2760 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3757
timestamp 1569533753
transform 1 0 2760 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3758
timestamp 1569533753
transform 1 0 2760 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3759
timestamp 1569533753
transform 1 0 2632 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3760
timestamp 1569533753
transform 1 0 2632 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3761
timestamp 1569533753
transform 1 0 2632 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3762
timestamp 1569533753
transform 1 0 2632 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3763
timestamp 1569533753
transform 1 0 2568 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3764
timestamp 1569533753
transform 1 0 2568 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3765
timestamp 1569533753
transform 1 0 2568 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3766
timestamp 1569533753
transform 1 0 2568 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3767
timestamp 1569533753
transform 1 0 2824 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3768
timestamp 1569533753
transform 1 0 2824 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3769
timestamp 1569533753
transform 1 0 2824 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3770
timestamp 1569533753
transform 1 0 2824 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3771
timestamp 1569533753
transform 1 0 2888 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3772
timestamp 1569533753
transform 1 0 2888 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3773
timestamp 1569533753
transform 1 0 2888 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3774
timestamp 1569533753
transform 1 0 2888 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3775
timestamp 1569533753
transform 1 0 2952 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3776
timestamp 1569533753
transform 1 0 2952 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3777
timestamp 1569533753
transform 1 0 2952 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3778
timestamp 1569533753
transform 1 0 2952 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3779
timestamp 1569533753
transform 1 0 3016 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3780
timestamp 1569533753
transform 1 0 3016 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3781
timestamp 1569533753
transform 1 0 3016 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3782
timestamp 1569533753
transform 1 0 3016 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3783
timestamp 1569533753
transform 1 0 3080 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3784
timestamp 1569533753
transform 1 0 3080 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3785
timestamp 1569533753
transform 1 0 3080 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_3786
timestamp 1569533753
transform 1 0 3080 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3787
timestamp 1569533753
transform 1 0 3016 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3788
timestamp 1569533753
transform 1 0 2888 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3789
timestamp 1569533753
transform 1 0 3080 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3790
timestamp 1569533753
transform 1 0 2952 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3791
timestamp 1569533753
transform 1 0 2824 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3792
timestamp 1569533753
transform 1 0 2824 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3793
timestamp 1569533753
transform 1 0 3080 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3794
timestamp 1569533753
transform 1 0 3080 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3795
timestamp 1569533753
transform 1 0 3016 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3796
timestamp 1569533753
transform 1 0 2888 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3797
timestamp 1569533753
transform 1 0 2824 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3798
timestamp 1569533753
transform 1 0 2888 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3799
timestamp 1569533753
transform 1 0 3016 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3800
timestamp 1569533753
transform 1 0 2952 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3801
timestamp 1569533753
transform 1 0 2952 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3802
timestamp 1569533753
transform 1 0 2888 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3803
timestamp 1569533753
transform 1 0 2824 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3804
timestamp 1569533753
transform 1 0 2952 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3805
timestamp 1569533753
transform 1 0 3016 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3806
timestamp 1569533753
transform 1 0 3080 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3807
timestamp 1569533753
transform 1 0 2760 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3808
timestamp 1569533753
transform 1 0 2696 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3809
timestamp 1569533753
transform 1 0 2632 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3810
timestamp 1569533753
transform 1 0 2568 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3811
timestamp 1569533753
transform 1 0 2632 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3812
timestamp 1569533753
transform 1 0 2760 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3813
timestamp 1569533753
transform 1 0 2632 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3814
timestamp 1569533753
transform 1 0 2696 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3815
timestamp 1569533753
transform 1 0 2760 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3816
timestamp 1569533753
transform 1 0 2568 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3817
timestamp 1569533753
transform 1 0 2568 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3818
timestamp 1569533753
transform 1 0 2696 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3819
timestamp 1569533753
transform 1 0 2696 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3820
timestamp 1569533753
transform 1 0 2760 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3821
timestamp 1569533753
transform 1 0 2568 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3822
timestamp 1569533753
transform 1 0 2632 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3823
timestamp 1569533753
transform 1 0 2696 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3824
timestamp 1569533753
transform 1 0 2632 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3825
timestamp 1569533753
transform 1 0 2760 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3826
timestamp 1569533753
transform 1 0 2760 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3827
timestamp 1569533753
transform 1 0 2760 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3828
timestamp 1569533753
transform 1 0 2696 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3829
timestamp 1569533753
transform 1 0 2696 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3830
timestamp 1569533753
transform 1 0 2760 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3831
timestamp 1569533753
transform 1 0 2696 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3832
timestamp 1569533753
transform 1 0 2568 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3833
timestamp 1569533753
transform 1 0 2568 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3834
timestamp 1569533753
transform 1 0 2568 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3835
timestamp 1569533753
transform 1 0 2632 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3836
timestamp 1569533753
transform 1 0 2568 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3837
timestamp 1569533753
transform 1 0 2632 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3838
timestamp 1569533753
transform 1 0 2632 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3839
timestamp 1569533753
transform 1 0 2824 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3840
timestamp 1569533753
transform 1 0 2952 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3841
timestamp 1569533753
transform 1 0 2952 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3842
timestamp 1569533753
transform 1 0 2824 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3843
timestamp 1569533753
transform 1 0 2952 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3844
timestamp 1569533753
transform 1 0 2952 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3845
timestamp 1569533753
transform 1 0 2824 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3846
timestamp 1569533753
transform 1 0 3016 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3847
timestamp 1569533753
transform 1 0 3016 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3848
timestamp 1569533753
transform 1 0 2824 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3849
timestamp 1569533753
transform 1 0 3016 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3850
timestamp 1569533753
transform 1 0 3016 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3851
timestamp 1569533753
transform 1 0 3080 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3852
timestamp 1569533753
transform 1 0 3080 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3853
timestamp 1569533753
transform 1 0 3080 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3854
timestamp 1569533753
transform 1 0 3080 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3855
timestamp 1569533753
transform 1 0 2888 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3856
timestamp 1569533753
transform 1 0 2888 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3857
timestamp 1569533753
transform 1 0 2888 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3858
timestamp 1569533753
transform 1 0 2888 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3859
timestamp 1569533753
transform 1 0 3464 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3860
timestamp 1569533753
transform 1 0 3656 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3861
timestamp 1569533753
transform 1 0 3464 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3862
timestamp 1569533753
transform 1 0 3464 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3863
timestamp 1569533753
transform 1 0 3528 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3864
timestamp 1569533753
transform 1 0 3592 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3865
timestamp 1569533753
transform 1 0 3720 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3866
timestamp 1569533753
transform 1 0 3592 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3867
timestamp 1569533753
transform 1 0 3592 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3868
timestamp 1569533753
transform 1 0 3720 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3869
timestamp 1569533753
transform 1 0 3528 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3870
timestamp 1569533753
transform 1 0 3464 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3871
timestamp 1569533753
transform 1 0 3592 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3872
timestamp 1569533753
transform 1 0 3528 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3873
timestamp 1569533753
transform 1 0 3656 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3874
timestamp 1569533753
transform 1 0 3656 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3875
timestamp 1569533753
transform 1 0 3720 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3876
timestamp 1569533753
transform 1 0 3656 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3877
timestamp 1569533753
transform 1 0 3528 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3878
timestamp 1569533753
transform 1 0 3720 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3879
timestamp 1569533753
transform 1 0 3336 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3880
timestamp 1569533753
transform 1 0 3208 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3881
timestamp 1569533753
transform 1 0 3400 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3882
timestamp 1569533753
transform 1 0 3336 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3883
timestamp 1569533753
transform 1 0 3208 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3884
timestamp 1569533753
transform 1 0 3336 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3885
timestamp 1569533753
transform 1 0 3208 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3886
timestamp 1569533753
transform 1 0 3272 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3887
timestamp 1569533753
transform 1 0 3400 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3888
timestamp 1569533753
transform 1 0 3144 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3889
timestamp 1569533753
transform 1 0 3272 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3890
timestamp 1569533753
transform 1 0 3272 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3891
timestamp 1569533753
transform 1 0 3272 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3892
timestamp 1569533753
transform 1 0 3144 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3893
timestamp 1569533753
transform 1 0 3400 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3894
timestamp 1569533753
transform 1 0 3400 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3895
timestamp 1569533753
transform 1 0 3144 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_3896
timestamp 1569533753
transform 1 0 3336 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3897
timestamp 1569533753
transform 1 0 3208 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_3898
timestamp 1569533753
transform 1 0 3144 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3899
timestamp 1569533753
transform 1 0 3272 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3900
timestamp 1569533753
transform 1 0 3272 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3901
timestamp 1569533753
transform 1 0 3272 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3902
timestamp 1569533753
transform 1 0 3336 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3903
timestamp 1569533753
transform 1 0 3336 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3904
timestamp 1569533753
transform 1 0 3336 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3905
timestamp 1569533753
transform 1 0 3336 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3906
timestamp 1569533753
transform 1 0 3400 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3907
timestamp 1569533753
transform 1 0 3400 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3908
timestamp 1569533753
transform 1 0 3400 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3909
timestamp 1569533753
transform 1 0 3144 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3910
timestamp 1569533753
transform 1 0 3144 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3911
timestamp 1569533753
transform 1 0 3400 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3912
timestamp 1569533753
transform 1 0 3144 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3913
timestamp 1569533753
transform 1 0 3144 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3914
timestamp 1569533753
transform 1 0 3208 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3915
timestamp 1569533753
transform 1 0 3208 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3916
timestamp 1569533753
transform 1 0 3208 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3917
timestamp 1569533753
transform 1 0 3208 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3918
timestamp 1569533753
transform 1 0 3272 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3919
timestamp 1569533753
transform 1 0 3464 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3920
timestamp 1569533753
transform 1 0 3592 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3921
timestamp 1569533753
transform 1 0 3592 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3922
timestamp 1569533753
transform 1 0 3592 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3923
timestamp 1569533753
transform 1 0 3592 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3924
timestamp 1569533753
transform 1 0 3656 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3925
timestamp 1569533753
transform 1 0 3656 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3926
timestamp 1569533753
transform 1 0 3656 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3927
timestamp 1569533753
transform 1 0 3656 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3928
timestamp 1569533753
transform 1 0 3720 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3929
timestamp 1569533753
transform 1 0 3720 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3930
timestamp 1569533753
transform 1 0 3720 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3931
timestamp 1569533753
transform 1 0 3464 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3932
timestamp 1569533753
transform 1 0 3720 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3933
timestamp 1569533753
transform 1 0 3464 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3934
timestamp 1569533753
transform 1 0 3528 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3935
timestamp 1569533753
transform 1 0 3528 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3936
timestamp 1569533753
transform 1 0 3528 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3937
timestamp 1569533753
transform 1 0 3528 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3938
timestamp 1569533753
transform 1 0 3464 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3939
timestamp 1569533753
transform 1 0 2696 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3940
timestamp 1569533753
transform 1 0 3336 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3941
timestamp 1569533753
transform 1 0 2760 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3942
timestamp 1569533753
transform 1 0 3400 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3943
timestamp 1569533753
transform 1 0 2824 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3944
timestamp 1569533753
transform 1 0 3464 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3945
timestamp 1569533753
transform 1 0 2888 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3946
timestamp 1569533753
transform 1 0 3528 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3947
timestamp 1569533753
transform 1 0 2952 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3948
timestamp 1569533753
transform 1 0 3592 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3949
timestamp 1569533753
transform 1 0 3016 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3950
timestamp 1569533753
transform 1 0 3656 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3951
timestamp 1569533753
transform 1 0 3080 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3952
timestamp 1569533753
transform 1 0 3720 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3953
timestamp 1569533753
transform 1 0 3144 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3954
timestamp 1569533753
transform 1 0 2568 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3955
timestamp 1569533753
transform 1 0 3208 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3956
timestamp 1569533753
transform 1 0 2632 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3957
timestamp 1569533753
transform 1 0 3272 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_3958
timestamp 1569533753
transform 1 0 4616 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3959
timestamp 1569533753
transform 1 0 4680 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3960
timestamp 1569533753
transform 1 0 4744 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3961
timestamp 1569533753
transform 1 0 4808 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3962
timestamp 1569533753
transform 1 0 4872 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3963
timestamp 1569533753
transform 1 0 4488 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3964
timestamp 1569533753
transform 1 0 4552 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_3965
timestamp 1569533753
transform 1 0 3976 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3966
timestamp 1569533753
transform 1 0 3976 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3967
timestamp 1569533753
transform 1 0 3976 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3968
timestamp 1569533753
transform 1 0 3976 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3969
timestamp 1569533753
transform 1 0 4040 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3970
timestamp 1569533753
transform 1 0 4040 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3971
timestamp 1569533753
transform 1 0 4040 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3972
timestamp 1569533753
transform 1 0 4104 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3973
timestamp 1569533753
transform 1 0 4104 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3974
timestamp 1569533753
transform 1 0 4168 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3975
timestamp 1569533753
transform 1 0 3848 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3976
timestamp 1569533753
transform 1 0 3848 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3977
timestamp 1569533753
transform 1 0 3912 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3978
timestamp 1569533753
transform 1 0 3912 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3979
timestamp 1569533753
transform 1 0 3912 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3980
timestamp 1569533753
transform 1 0 3912 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3981
timestamp 1569533753
transform 1 0 3784 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3982
timestamp 1569533753
transform 1 0 3784 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3983
timestamp 1569533753
transform 1 0 3784 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_3984
timestamp 1569533753
transform 1 0 3848 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3985
timestamp 1569533753
transform 1 0 3848 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_3986
timestamp 1569533753
transform 1 0 3912 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_3987
timestamp 1569533753
transform 1 0 3784 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3988
timestamp 1569533753
transform 1 0 3784 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3989
timestamp 1569533753
transform 1 0 3784 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_3990
timestamp 1569533753
transform 1 0 3784 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_3991
timestamp 1569533753
transform 1 0 3848 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_3992
timestamp 1569533753
transform 1 0 3848 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_3993
timestamp 1569533753
transform 1 0 4296 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_3994
timestamp 1569533753
transform 1 0 4296 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_3995
timestamp 1569533753
transform 1 0 4296 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_3996
timestamp 1569533753
transform 1 0 4296 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_3997
timestamp 1569533753
transform 1 0 4296 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_3998
timestamp 1569533753
transform 1 0 4296 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_3999
timestamp 1569533753
transform 1 0 4296 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4000
timestamp 1569533753
transform 1 0 4616 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4001
timestamp 1569533753
transform 1 0 4680 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4002
timestamp 1569533753
transform 1 0 4744 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4003
timestamp 1569533753
transform 1 0 4808 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4004
timestamp 1569533753
transform 1 0 4872 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4005
timestamp 1569533753
transform 1 0 4936 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4006
timestamp 1569533753
transform 1 0 4936 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4007
timestamp 1569533753
transform 1 0 4936 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4008
timestamp 1569533753
transform 1 0 4936 0 1 4936
box -8 -8 8 8
use VIA1$3  VIA1$3_4009
timestamp 1569533753
transform 1 0 4424 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4010
timestamp 1569533753
transform 1 0 4488 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4011
timestamp 1569533753
transform 1 0 4424 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_4012
timestamp 1569533753
transform 1 0 4424 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_4013
timestamp 1569533753
transform 1 0 4424 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4014
timestamp 1569533753
transform 1 0 4424 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4015
timestamp 1569533753
transform 1 0 4424 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4016
timestamp 1569533753
transform 1 0 4488 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4017
timestamp 1569533753
transform 1 0 4616 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4018
timestamp 1569533753
transform 1 0 4552 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4019
timestamp 1569533753
transform 1 0 4488 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_4020
timestamp 1569533753
transform 1 0 4424 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4021
timestamp 1569533753
transform 1 0 4488 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4022
timestamp 1569533753
transform 1 0 4552 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4023
timestamp 1569533753
transform 1 0 4744 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4024
timestamp 1569533753
transform 1 0 4744 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4025
timestamp 1569533753
transform 1 0 4744 0 1 4936
box -8 -8 8 8
use VIA1$3  VIA1$3_4026
timestamp 1569533753
transform 1 0 4808 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4027
timestamp 1569533753
transform 1 0 4808 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4028
timestamp 1569533753
transform 1 0 4808 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4029
timestamp 1569533753
transform 1 0 4808 0 1 4936
box -8 -8 8 8
use VIA1$3  VIA1$3_4030
timestamp 1569533753
transform 1 0 4424 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4031
timestamp 1569533753
transform 1 0 4552 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4032
timestamp 1569533753
transform 1 0 4872 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4033
timestamp 1569533753
transform 1 0 4872 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4034
timestamp 1569533753
transform 1 0 4872 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4035
timestamp 1569533753
transform 1 0 4872 0 1 4936
box -8 -8 8 8
use VIA1$3  VIA1$3_4036
timestamp 1569533753
transform 1 0 4616 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4037
timestamp 1569533753
transform 1 0 4680 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4038
timestamp 1569533753
transform 1 0 4744 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4039
timestamp 1569533753
transform 1 0 4808 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4040
timestamp 1569533753
transform 1 0 4872 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4041
timestamp 1569533753
transform 1 0 4360 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4042
timestamp 1569533753
transform 1 0 4360 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_4043
timestamp 1569533753
transform 1 0 4360 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_4044
timestamp 1569533753
transform 1 0 4360 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4045
timestamp 1569533753
transform 1 0 4360 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4046
timestamp 1569533753
transform 1 0 4360 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4047
timestamp 1569533753
transform 1 0 4360 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4048
timestamp 1569533753
transform 1 0 4360 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4049
timestamp 1569533753
transform 1 0 4424 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4050
timestamp 1569533753
transform 1 0 4488 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4051
timestamp 1569533753
transform 1 0 4552 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4052
timestamp 1569533753
transform 1 0 2504 0 1 4616
box -8 -8 8 8
use VIA1$3  VIA1$3_4053
timestamp 1569533753
transform 1 0 2504 0 1 4680
box -8 -8 8 8
use VIA1$3  VIA1$3_4054
timestamp 1569533753
transform 1 0 2504 0 1 4744
box -8 -8 8 8
use VIA1$3  VIA1$3_4055
timestamp 1569533753
transform 1 0 2504 0 1 4808
box -8 -8 8 8
use VIA1$3  VIA1$3_4056
timestamp 1569533753
transform 1 0 2504 0 1 4872
box -8 -8 8 8
use VIA1$3  VIA1$3_4057
timestamp 1569533753
transform 1 0 2504 0 1 136
box -8 -8 8 8
use VIA1$3  VIA1$3_4058
timestamp 1569533753
transform 1 0 2504 0 1 200
box -8 -8 8 8
use VIA1$3  VIA1$3_4059
timestamp 1569533753
transform 1 0 2504 0 1 264
box -8 -8 8 8
use VIA1$3  VIA1$3_4060
timestamp 1569533753
transform 1 0 2504 0 1 328
box -8 -8 8 8
use VIA1$3  VIA1$3_4061
timestamp 1569533753
transform 1 0 2504 0 1 392
box -8 -8 8 8
use VIA1$3  VIA1$3_4062
timestamp 1569533753
transform 1 0 2504 0 1 456
box -8 -8 8 8
use VIA1$3  VIA1$3_4063
timestamp 1569533753
transform 1 0 2504 0 1 520
box -8 -8 8 8
use VIA1$3  VIA1$3_4064
timestamp 1569533753
transform 1 0 2504 0 1 584
box -8 -8 8 8
use VIA1$3  VIA1$3_4065
timestamp 1569533753
transform 1 0 2504 0 1 648
box -8 -8 8 8
use VIA1$3  VIA1$3_4066
timestamp 1569533753
transform 1 0 2504 0 1 712
box -8 -8 8 8
use VIA1$3  VIA1$3_4067
timestamp 1569533753
transform 1 0 2504 0 1 776
box -8 -8 8 8
use VIA1$3  VIA1$3_4068
timestamp 1569533753
transform 1 0 2504 0 1 840
box -8 -8 8 8
use VIA1$3  VIA1$3_4069
timestamp 1569533753
transform 1 0 2504 0 1 904
box -8 -8 8 8
use VIA1$3  VIA1$3_4070
timestamp 1569533753
transform 1 0 2504 0 1 968
box -8 -8 8 8
use VIA1$3  VIA1$3_4071
timestamp 1569533753
transform 1 0 2504 0 1 1032
box -8 -8 8 8
use VIA1$3  VIA1$3_4072
timestamp 1569533753
transform 1 0 2504 0 1 1096
box -8 -8 8 8
use VIA1$3  VIA1$3_4073
timestamp 1569533753
transform 1 0 2504 0 1 1160
box -8 -8 8 8
use VIA1$3  VIA1$3_4074
timestamp 1569533753
transform 1 0 2504 0 1 1224
box -8 -8 8 8
use VIA1$3  VIA1$3_4075
timestamp 1569533753
transform 1 0 2504 0 1 1288
box -8 -8 8 8
use VIA1$3  VIA1$3_4076
timestamp 1569533753
transform 1 0 2504 0 1 1352
box -8 -8 8 8
use VIA1$3  VIA1$3_4077
timestamp 1569533753
transform 1 0 2504 0 1 1416
box -8 -8 8 8
use VIA1$3  VIA1$3_4078
timestamp 1569533753
transform 1 0 2504 0 1 1480
box -8 -8 8 8
use VIA1$3  VIA1$3_4079
timestamp 1569533753
transform 1 0 2504 0 1 1544
box -8 -8 8 8
use VIA1$3  VIA1$3_4080
timestamp 1569533753
transform 1 0 2504 0 1 1608
box -8 -8 8 8
use VIA1$3  VIA1$3_4081
timestamp 1569533753
transform 1 0 2504 0 1 1672
box -8 -8 8 8
use VIA1$3  VIA1$3_4082
timestamp 1569533753
transform 1 0 2504 0 1 1736
box -8 -8 8 8
use VIA1$3  VIA1$3_4083
timestamp 1569533753
transform 1 0 2504 0 1 1800
box -8 -8 8 8
use VIA1$3  VIA1$3_4084
timestamp 1569533753
transform 1 0 2504 0 1 1864
box -8 -8 8 8
use VIA1$3  VIA1$3_4085
timestamp 1569533753
transform 1 0 2504 0 1 1928
box -8 -8 8 8
use VIA1$3  VIA1$3_4086
timestamp 1569533753
transform 1 0 392 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4087
timestamp 1569533753
transform 1 0 1160 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4088
timestamp 1569533753
transform 1 0 1928 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4089
timestamp 1569533753
transform 1 0 3464 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4090
timestamp 1569533753
transform 1 0 4232 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4091
timestamp 1569533753
transform 1 0 456 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4092
timestamp 1569533753
transform 1 0 1224 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4093
timestamp 1569533753
transform 1 0 3528 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4094
timestamp 1569533753
transform 1 0 4296 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4095
timestamp 1569533753
transform 1 0 520 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4096
timestamp 1569533753
transform 1 0 1288 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4097
timestamp 1569533753
transform 1 0 3592 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4098
timestamp 1569533753
transform 1 0 4360 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4099
timestamp 1569533753
transform 1 0 584 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4100
timestamp 1569533753
transform 1 0 1352 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4101
timestamp 1569533753
transform 1 0 3656 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4102
timestamp 1569533753
transform 1 0 4424 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4103
timestamp 1569533753
transform 1 0 648 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4104
timestamp 1569533753
transform 1 0 1416 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4105
timestamp 1569533753
transform 1 0 3720 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4106
timestamp 1569533753
transform 1 0 4488 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4107
timestamp 1569533753
transform 1 0 712 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4108
timestamp 1569533753
transform 1 0 1480 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4109
timestamp 1569533753
transform 1 0 3784 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4110
timestamp 1569533753
transform 1 0 4552 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4111
timestamp 1569533753
transform 1 0 2504 0 1 3208
box -8 -8 8 8
use VIA1$3  VIA1$3_4112
timestamp 1569533753
transform 1 0 2504 0 1 3272
box -8 -8 8 8
use VIA1$3  VIA1$3_4113
timestamp 1569533753
transform 1 0 2504 0 1 3336
box -8 -8 8 8
use VIA1$3  VIA1$3_4114
timestamp 1569533753
transform 1 0 2504 0 1 3400
box -8 -8 8 8
use VIA1$3  VIA1$3_4115
timestamp 1569533753
transform 1 0 2504 0 1 3464
box -8 -8 8 8
use VIA1$3  VIA1$3_4116
timestamp 1569533753
transform 1 0 2504 0 1 3528
box -8 -8 8 8
use VIA1$3  VIA1$3_4117
timestamp 1569533753
transform 1 0 2504 0 1 3592
box -8 -8 8 8
use VIA1$3  VIA1$3_4118
timestamp 1569533753
transform 1 0 2504 0 1 3656
box -8 -8 8 8
use VIA1$3  VIA1$3_4119
timestamp 1569533753
transform 1 0 2504 0 1 3720
box -8 -8 8 8
use VIA1$3  VIA1$3_4120
timestamp 1569533753
transform 1 0 2504 0 1 3784
box -8 -8 8 8
use VIA1$3  VIA1$3_4121
timestamp 1569533753
transform 1 0 2504 0 1 3848
box -8 -8 8 8
use VIA1$3  VIA1$3_4122
timestamp 1569533753
transform 1 0 2504 0 1 3912
box -8 -8 8 8
use VIA1$3  VIA1$3_4123
timestamp 1569533753
transform 1 0 2504 0 1 3976
box -8 -8 8 8
use VIA1$3  VIA1$3_4124
timestamp 1569533753
transform 1 0 2504 0 1 4040
box -8 -8 8 8
use VIA1$3  VIA1$3_4125
timestamp 1569533753
transform 1 0 2504 0 1 4104
box -8 -8 8 8
use VIA1$3  VIA1$3_4126
timestamp 1569533753
transform 1 0 2504 0 1 4168
box -8 -8 8 8
use VIA1$3  VIA1$3_4127
timestamp 1569533753
transform 1 0 2504 0 1 4232
box -8 -8 8 8
use VIA1$3  VIA1$3_4128
timestamp 1569533753
transform 1 0 2504 0 1 4296
box -8 -8 8 8
use VIA1$3  VIA1$3_4129
timestamp 1569533753
transform 1 0 2504 0 1 4360
box -8 -8 8 8
use VIA1$3  VIA1$3_4130
timestamp 1569533753
transform 1 0 2504 0 1 4424
box -8 -8 8 8
use VIA1$3  VIA1$3_4131
timestamp 1569533753
transform 1 0 2504 0 1 4488
box -8 -8 8 8
use VIA1$3  VIA1$3_4132
timestamp 1569533753
transform 1 0 2504 0 1 4552
box -8 -8 8 8
use VIA1$3  VIA1$3_4133
timestamp 1569533753
transform 1 0 2504 0 1 72
box -8 -8 8 8
use VIA1$3  VIA1$3_4134
timestamp 1569533753
transform 1 0 776 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4135
timestamp 1569533753
transform 1 0 1544 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4136
timestamp 1569533753
transform 1 0 3848 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4137
timestamp 1569533753
transform 1 0 4616 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4138
timestamp 1569533753
transform 1 0 72 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4139
timestamp 1569533753
transform 1 0 840 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4140
timestamp 1569533753
transform 1 0 1608 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4141
timestamp 1569533753
transform 1 0 3912 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4142
timestamp 1569533753
transform 1 0 4680 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4143
timestamp 1569533753
transform 1 0 136 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4144
timestamp 1569533753
transform 1 0 904 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4145
timestamp 1569533753
transform 1 0 1672 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4146
timestamp 1569533753
transform 1 0 3208 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4147
timestamp 1569533753
transform 1 0 3976 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4148
timestamp 1569533753
transform 1 0 4744 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4149
timestamp 1569533753
transform 1 0 200 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4150
timestamp 1569533753
transform 1 0 968 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4151
timestamp 1569533753
transform 1 0 1736 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4152
timestamp 1569533753
transform 1 0 3272 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4153
timestamp 1569533753
transform 1 0 4040 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4154
timestamp 1569533753
transform 1 0 4808 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4155
timestamp 1569533753
transform 1 0 264 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4156
timestamp 1569533753
transform 1 0 1032 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4157
timestamp 1569533753
transform 1 0 1800 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4158
timestamp 1569533753
transform 1 0 3336 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4159
timestamp 1569533753
transform 1 0 4104 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4160
timestamp 1569533753
transform 1 0 4872 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4161
timestamp 1569533753
transform 1 0 328 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4162
timestamp 1569533753
transform 1 0 1096 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4163
timestamp 1569533753
transform 1 0 1864 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4164
timestamp 1569533753
transform 1 0 3400 0 1 2504
box -8 -8 8 8
use VIA1$3  VIA1$3_4165
timestamp 1569533753
transform 1 0 4168 0 1 2504
box -8 -8 8 8
use VIA2$3  VIA2$3_0
timestamp 1569533753
transform 1 0 4840 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1
timestamp 1569533753
transform 1 0 4776 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_2
timestamp 1569533753
transform 1 0 4712 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_3
timestamp 1569533753
transform 1 0 4712 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_4
timestamp 1569533753
transform 1 0 4712 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_5
timestamp 1569533753
transform 1 0 4776 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_6
timestamp 1569533753
transform 1 0 4904 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_7
timestamp 1569533753
transform 1 0 4776 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_8
timestamp 1569533753
transform 1 0 4904 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_9
timestamp 1569533753
transform 1 0 4712 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_10
timestamp 1569533753
transform 1 0 4904 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_11
timestamp 1569533753
transform 1 0 4840 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_12
timestamp 1569533753
transform 1 0 4712 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_13
timestamp 1569533753
transform 1 0 4776 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_14
timestamp 1569533753
transform 1 0 4904 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_15
timestamp 1569533753
transform 1 0 4840 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_16
timestamp 1569533753
transform 1 0 4904 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_17
timestamp 1569533753
transform 1 0 4776 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_18
timestamp 1569533753
transform 1 0 4840 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_19
timestamp 1569533753
transform 1 0 4840 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_20
timestamp 1569533753
transform 1 0 4584 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_21
timestamp 1569533753
transform 1 0 4520 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_22
timestamp 1569533753
transform 1 0 4584 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_23
timestamp 1569533753
transform 1 0 4456 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_24
timestamp 1569533753
transform 1 0 4648 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_25
timestamp 1569533753
transform 1 0 4648 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_26
timestamp 1569533753
transform 1 0 4456 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_27
timestamp 1569533753
transform 1 0 4456 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_28
timestamp 1569533753
transform 1 0 4584 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_29
timestamp 1569533753
transform 1 0 4392 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_30
timestamp 1569533753
transform 1 0 4520 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_31
timestamp 1569533753
transform 1 0 4648 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_32
timestamp 1569533753
transform 1 0 4584 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_33
timestamp 1569533753
transform 1 0 4520 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_34
timestamp 1569533753
transform 1 0 4520 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_35
timestamp 1569533753
transform 1 0 4584 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_36
timestamp 1569533753
transform 1 0 4392 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_37
timestamp 1569533753
transform 1 0 4456 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_38
timestamp 1569533753
transform 1 0 4392 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_39
timestamp 1569533753
transform 1 0 4392 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_40
timestamp 1569533753
transform 1 0 4648 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_41
timestamp 1569533753
transform 1 0 4520 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_42
timestamp 1569533753
transform 1 0 4648 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_43
timestamp 1569533753
transform 1 0 4456 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_44
timestamp 1569533753
transform 1 0 4392 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_45
timestamp 1569533753
transform 1 0 4584 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_46
timestamp 1569533753
transform 1 0 4456 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_47
timestamp 1569533753
transform 1 0 4520 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_48
timestamp 1569533753
transform 1 0 4456 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_49
timestamp 1569533753
transform 1 0 4584 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_50
timestamp 1569533753
transform 1 0 4392 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_51
timestamp 1569533753
transform 1 0 4584 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_52
timestamp 1569533753
transform 1 0 4648 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_53
timestamp 1569533753
transform 1 0 4520 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_54
timestamp 1569533753
transform 1 0 4456 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_55
timestamp 1569533753
transform 1 0 4520 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_56
timestamp 1569533753
transform 1 0 4456 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_57
timestamp 1569533753
transform 1 0 4648 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_58
timestamp 1569533753
transform 1 0 4648 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_59
timestamp 1569533753
transform 1 0 4520 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_60
timestamp 1569533753
transform 1 0 4584 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_61
timestamp 1569533753
transform 1 0 4648 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_62
timestamp 1569533753
transform 1 0 4392 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_63
timestamp 1569533753
transform 1 0 4520 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_64
timestamp 1569533753
transform 1 0 4392 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_65
timestamp 1569533753
transform 1 0 4648 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_66
timestamp 1569533753
transform 1 0 4392 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_67
timestamp 1569533753
transform 1 0 4456 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_68
timestamp 1569533753
transform 1 0 4392 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_69
timestamp 1569533753
transform 1 0 4584 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_70
timestamp 1569533753
transform 1 0 4776 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_71
timestamp 1569533753
transform 1 0 4712 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_72
timestamp 1569533753
transform 1 0 4840 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_73
timestamp 1569533753
transform 1 0 4904 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_74
timestamp 1569533753
transform 1 0 4904 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_75
timestamp 1569533753
transform 1 0 4904 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_76
timestamp 1569533753
transform 1 0 4840 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_77
timestamp 1569533753
transform 1 0 4776 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_78
timestamp 1569533753
transform 1 0 4904 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_79
timestamp 1569533753
transform 1 0 4776 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_80
timestamp 1569533753
transform 1 0 4840 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_81
timestamp 1569533753
transform 1 0 4712 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_82
timestamp 1569533753
transform 1 0 4712 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_83
timestamp 1569533753
transform 1 0 4840 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_84
timestamp 1569533753
transform 1 0 4904 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_85
timestamp 1569533753
transform 1 0 4776 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_86
timestamp 1569533753
transform 1 0 4712 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_87
timestamp 1569533753
transform 1 0 4840 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_88
timestamp 1569533753
transform 1 0 4712 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_89
timestamp 1569533753
transform 1 0 4776 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_90
timestamp 1569533753
transform 1 0 4136 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_91
timestamp 1569533753
transform 1 0 4264 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_92
timestamp 1569533753
transform 1 0 4200 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_93
timestamp 1569533753
transform 1 0 4200 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_94
timestamp 1569533753
transform 1 0 4200 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_95
timestamp 1569533753
transform 1 0 4072 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_96
timestamp 1569533753
transform 1 0 4072 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_97
timestamp 1569533753
transform 1 0 4136 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_98
timestamp 1569533753
transform 1 0 4200 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_99
timestamp 1569533753
transform 1 0 4072 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_100
timestamp 1569533753
transform 1 0 4072 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_101
timestamp 1569533753
transform 1 0 4328 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_102
timestamp 1569533753
transform 1 0 4136 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_103
timestamp 1569533753
transform 1 0 4328 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_104
timestamp 1569533753
transform 1 0 4264 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_105
timestamp 1569533753
transform 1 0 4200 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_106
timestamp 1569533753
transform 1 0 4136 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_107
timestamp 1569533753
transform 1 0 4328 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_108
timestamp 1569533753
transform 1 0 4328 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_109
timestamp 1569533753
transform 1 0 4264 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_110
timestamp 1569533753
transform 1 0 4264 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_111
timestamp 1569533753
transform 1 0 4264 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_112
timestamp 1569533753
transform 1 0 4072 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_113
timestamp 1569533753
transform 1 0 4136 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_114
timestamp 1569533753
transform 1 0 4328 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_115
timestamp 1569533753
transform 1 0 3816 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_116
timestamp 1569533753
transform 1 0 3880 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_117
timestamp 1569533753
transform 1 0 4008 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_118
timestamp 1569533753
transform 1 0 3816 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_119
timestamp 1569533753
transform 1 0 3944 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_120
timestamp 1569533753
transform 1 0 3752 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_121
timestamp 1569533753
transform 1 0 3944 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_122
timestamp 1569533753
transform 1 0 3880 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_123
timestamp 1569533753
transform 1 0 4008 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_124
timestamp 1569533753
transform 1 0 3944 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_125
timestamp 1569533753
transform 1 0 3944 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_126
timestamp 1569533753
transform 1 0 3880 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_127
timestamp 1569533753
transform 1 0 3752 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_128
timestamp 1569533753
transform 1 0 4008 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_129
timestamp 1569533753
transform 1 0 3752 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_130
timestamp 1569533753
transform 1 0 4008 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_131
timestamp 1569533753
transform 1 0 3944 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_132
timestamp 1569533753
transform 1 0 3880 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_133
timestamp 1569533753
transform 1 0 3816 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_134
timestamp 1569533753
transform 1 0 4008 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_135
timestamp 1569533753
transform 1 0 3752 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_136
timestamp 1569533753
transform 1 0 3752 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_137
timestamp 1569533753
transform 1 0 3816 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_138
timestamp 1569533753
transform 1 0 3880 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_139
timestamp 1569533753
transform 1 0 3816 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_140
timestamp 1569533753
transform 1 0 3752 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_141
timestamp 1569533753
transform 1 0 3880 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_142
timestamp 1569533753
transform 1 0 3944 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_143
timestamp 1569533753
transform 1 0 3752 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_144
timestamp 1569533753
transform 1 0 3816 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_145
timestamp 1569533753
transform 1 0 3752 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_146
timestamp 1569533753
transform 1 0 3944 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_147
timestamp 1569533753
transform 1 0 4008 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_148
timestamp 1569533753
transform 1 0 4008 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_149
timestamp 1569533753
transform 1 0 3880 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_150
timestamp 1569533753
transform 1 0 4008 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_151
timestamp 1569533753
transform 1 0 3944 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_152
timestamp 1569533753
transform 1 0 3880 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_153
timestamp 1569533753
transform 1 0 4008 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_154
timestamp 1569533753
transform 1 0 3880 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_155
timestamp 1569533753
transform 1 0 3752 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_156
timestamp 1569533753
transform 1 0 3816 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_157
timestamp 1569533753
transform 1 0 4008 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_158
timestamp 1569533753
transform 1 0 3944 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_159
timestamp 1569533753
transform 1 0 3816 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_160
timestamp 1569533753
transform 1 0 3816 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_161
timestamp 1569533753
transform 1 0 3944 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_162
timestamp 1569533753
transform 1 0 3752 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_163
timestamp 1569533753
transform 1 0 3816 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_164
timestamp 1569533753
transform 1 0 3880 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_165
timestamp 1569533753
transform 1 0 4200 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_166
timestamp 1569533753
transform 1 0 4072 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_167
timestamp 1569533753
transform 1 0 4200 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_168
timestamp 1569533753
transform 1 0 4264 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_169
timestamp 1569533753
transform 1 0 4072 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_170
timestamp 1569533753
transform 1 0 4136 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_171
timestamp 1569533753
transform 1 0 4200 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_172
timestamp 1569533753
transform 1 0 4264 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_173
timestamp 1569533753
transform 1 0 4328 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_174
timestamp 1569533753
transform 1 0 4136 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_175
timestamp 1569533753
transform 1 0 4136 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_176
timestamp 1569533753
transform 1 0 4328 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_177
timestamp 1569533753
transform 1 0 4072 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_178
timestamp 1569533753
transform 1 0 4328 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_179
timestamp 1569533753
transform 1 0 4200 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_180
timestamp 1569533753
transform 1 0 4328 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_181
timestamp 1569533753
transform 1 0 4264 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_182
timestamp 1569533753
transform 1 0 4328 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_183
timestamp 1569533753
transform 1 0 4200 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_184
timestamp 1569533753
transform 1 0 4264 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_185
timestamp 1569533753
transform 1 0 4072 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_186
timestamp 1569533753
transform 1 0 4136 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_187
timestamp 1569533753
transform 1 0 4264 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_188
timestamp 1569533753
transform 1 0 4072 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_189
timestamp 1569533753
transform 1 0 4136 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_190
timestamp 1569533753
transform 1 0 4136 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_191
timestamp 1569533753
transform 1 0 4264 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_192
timestamp 1569533753
transform 1 0 4200 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_193
timestamp 1569533753
transform 1 0 4072 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_194
timestamp 1569533753
transform 1 0 4264 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_195
timestamp 1569533753
transform 1 0 4328 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_196
timestamp 1569533753
transform 1 0 4072 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_197
timestamp 1569533753
transform 1 0 4328 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_198
timestamp 1569533753
transform 1 0 4136 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_199
timestamp 1569533753
transform 1 0 4200 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_200
timestamp 1569533753
transform 1 0 4136 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_201
timestamp 1569533753
transform 1 0 4264 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_202
timestamp 1569533753
transform 1 0 4328 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_203
timestamp 1569533753
transform 1 0 4200 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_204
timestamp 1569533753
transform 1 0 4072 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_205
timestamp 1569533753
transform 1 0 4136 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_206
timestamp 1569533753
transform 1 0 4200 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_207
timestamp 1569533753
transform 1 0 4264 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_208
timestamp 1569533753
transform 1 0 4072 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_209
timestamp 1569533753
transform 1 0 4136 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_210
timestamp 1569533753
transform 1 0 4328 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_211
timestamp 1569533753
transform 1 0 4264 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_212
timestamp 1569533753
transform 1 0 4328 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_213
timestamp 1569533753
transform 1 0 4072 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_214
timestamp 1569533753
transform 1 0 4200 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_215
timestamp 1569533753
transform 1 0 3816 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_216
timestamp 1569533753
transform 1 0 4008 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_217
timestamp 1569533753
transform 1 0 4008 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_218
timestamp 1569533753
transform 1 0 3752 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_219
timestamp 1569533753
transform 1 0 3880 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_220
timestamp 1569533753
transform 1 0 3816 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_221
timestamp 1569533753
transform 1 0 3944 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_222
timestamp 1569533753
transform 1 0 3752 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_223
timestamp 1569533753
transform 1 0 3944 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_224
timestamp 1569533753
transform 1 0 3816 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_225
timestamp 1569533753
transform 1 0 3816 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_226
timestamp 1569533753
transform 1 0 3752 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_227
timestamp 1569533753
transform 1 0 3752 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_228
timestamp 1569533753
transform 1 0 3944 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_229
timestamp 1569533753
transform 1 0 4008 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_230
timestamp 1569533753
transform 1 0 3880 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_231
timestamp 1569533753
transform 1 0 4008 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_232
timestamp 1569533753
transform 1 0 4008 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_233
timestamp 1569533753
transform 1 0 3816 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_234
timestamp 1569533753
transform 1 0 3880 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_235
timestamp 1569533753
transform 1 0 3944 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_236
timestamp 1569533753
transform 1 0 3944 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_237
timestamp 1569533753
transform 1 0 3880 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_238
timestamp 1569533753
transform 1 0 3752 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_239
timestamp 1569533753
transform 1 0 3880 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_240
timestamp 1569533753
transform 1 0 3816 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_241
timestamp 1569533753
transform 1 0 4008 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_242
timestamp 1569533753
transform 1 0 3880 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_243
timestamp 1569533753
transform 1 0 3944 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_244
timestamp 1569533753
transform 1 0 3944 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_245
timestamp 1569533753
transform 1 0 3816 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_246
timestamp 1569533753
transform 1 0 3880 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_247
timestamp 1569533753
transform 1 0 4008 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_248
timestamp 1569533753
transform 1 0 3880 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_249
timestamp 1569533753
transform 1 0 3816 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_250
timestamp 1569533753
transform 1 0 3816 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_251
timestamp 1569533753
transform 1 0 4008 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_252
timestamp 1569533753
transform 1 0 3944 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_253
timestamp 1569533753
transform 1 0 3944 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_254
timestamp 1569533753
transform 1 0 3944 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_255
timestamp 1569533753
transform 1 0 3752 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_256
timestamp 1569533753
transform 1 0 3816 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_257
timestamp 1569533753
transform 1 0 3752 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_258
timestamp 1569533753
transform 1 0 4008 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_259
timestamp 1569533753
transform 1 0 3752 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_260
timestamp 1569533753
transform 1 0 3752 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_261
timestamp 1569533753
transform 1 0 3752 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_262
timestamp 1569533753
transform 1 0 4008 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_263
timestamp 1569533753
transform 1 0 3880 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_264
timestamp 1569533753
transform 1 0 3880 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_265
timestamp 1569533753
transform 1 0 4328 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_266
timestamp 1569533753
transform 1 0 4200 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_267
timestamp 1569533753
transform 1 0 4264 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_268
timestamp 1569533753
transform 1 0 4200 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_269
timestamp 1569533753
transform 1 0 4328 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_270
timestamp 1569533753
transform 1 0 4072 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_271
timestamp 1569533753
transform 1 0 4136 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_272
timestamp 1569533753
transform 1 0 4328 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_273
timestamp 1569533753
transform 1 0 4072 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_274
timestamp 1569533753
transform 1 0 4264 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_275
timestamp 1569533753
transform 1 0 4136 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_276
timestamp 1569533753
transform 1 0 4072 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_277
timestamp 1569533753
transform 1 0 4264 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_278
timestamp 1569533753
transform 1 0 4200 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_279
timestamp 1569533753
transform 1 0 4136 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_280
timestamp 1569533753
transform 1 0 4136 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_281
timestamp 1569533753
transform 1 0 4328 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_282
timestamp 1569533753
transform 1 0 4136 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_283
timestamp 1569533753
transform 1 0 4200 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_284
timestamp 1569533753
transform 1 0 4072 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_285
timestamp 1569533753
transform 1 0 4328 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_286
timestamp 1569533753
transform 1 0 4264 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_287
timestamp 1569533753
transform 1 0 4200 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_288
timestamp 1569533753
transform 1 0 4264 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_289
timestamp 1569533753
transform 1 0 4072 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_290
timestamp 1569533753
transform 1 0 4712 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_291
timestamp 1569533753
transform 1 0 4712 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_292
timestamp 1569533753
transform 1 0 4904 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_293
timestamp 1569533753
transform 1 0 4776 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_294
timestamp 1569533753
transform 1 0 4776 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_295
timestamp 1569533753
transform 1 0 4904 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_296
timestamp 1569533753
transform 1 0 4840 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_297
timestamp 1569533753
transform 1 0 4904 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_298
timestamp 1569533753
transform 1 0 4840 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_299
timestamp 1569533753
transform 1 0 4904 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_300
timestamp 1569533753
transform 1 0 4840 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_301
timestamp 1569533753
transform 1 0 4776 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_302
timestamp 1569533753
transform 1 0 4840 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_303
timestamp 1569533753
transform 1 0 4776 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_304
timestamp 1569533753
transform 1 0 4904 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_305
timestamp 1569533753
transform 1 0 4712 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_306
timestamp 1569533753
transform 1 0 4712 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_307
timestamp 1569533753
transform 1 0 4776 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_308
timestamp 1569533753
transform 1 0 4712 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_309
timestamp 1569533753
transform 1 0 4840 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_310
timestamp 1569533753
transform 1 0 4520 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_311
timestamp 1569533753
transform 1 0 4520 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_312
timestamp 1569533753
transform 1 0 4520 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_313
timestamp 1569533753
transform 1 0 4520 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_314
timestamp 1569533753
transform 1 0 4392 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_315
timestamp 1569533753
transform 1 0 4392 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_316
timestamp 1569533753
transform 1 0 4392 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_317
timestamp 1569533753
transform 1 0 4392 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_318
timestamp 1569533753
transform 1 0 4392 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_319
timestamp 1569533753
transform 1 0 4584 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_320
timestamp 1569533753
transform 1 0 4584 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_321
timestamp 1569533753
transform 1 0 4648 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_322
timestamp 1569533753
transform 1 0 4648 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_323
timestamp 1569533753
transform 1 0 4648 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_324
timestamp 1569533753
transform 1 0 4584 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_325
timestamp 1569533753
transform 1 0 4456 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_326
timestamp 1569533753
transform 1 0 4456 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_327
timestamp 1569533753
transform 1 0 4456 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_328
timestamp 1569533753
transform 1 0 4648 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_329
timestamp 1569533753
transform 1 0 4584 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_330
timestamp 1569533753
transform 1 0 4456 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_331
timestamp 1569533753
transform 1 0 4456 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_332
timestamp 1569533753
transform 1 0 4648 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_333
timestamp 1569533753
transform 1 0 4584 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_334
timestamp 1569533753
transform 1 0 4520 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_335
timestamp 1569533753
transform 1 0 4648 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_336
timestamp 1569533753
transform 1 0 4456 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_337
timestamp 1569533753
transform 1 0 4520 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_338
timestamp 1569533753
transform 1 0 4584 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_339
timestamp 1569533753
transform 1 0 4456 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_340
timestamp 1569533753
transform 1 0 4520 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_341
timestamp 1569533753
transform 1 0 4392 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_342
timestamp 1569533753
transform 1 0 4520 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_343
timestamp 1569533753
transform 1 0 4648 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_344
timestamp 1569533753
transform 1 0 4456 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_345
timestamp 1569533753
transform 1 0 4520 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_346
timestamp 1569533753
transform 1 0 4584 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_347
timestamp 1569533753
transform 1 0 4392 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_348
timestamp 1569533753
transform 1 0 4648 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_349
timestamp 1569533753
transform 1 0 4520 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_350
timestamp 1569533753
transform 1 0 4392 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_351
timestamp 1569533753
transform 1 0 4392 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_352
timestamp 1569533753
transform 1 0 4584 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_353
timestamp 1569533753
transform 1 0 4456 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_354
timestamp 1569533753
transform 1 0 4648 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_355
timestamp 1569533753
transform 1 0 4584 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_356
timestamp 1569533753
transform 1 0 4392 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_357
timestamp 1569533753
transform 1 0 4456 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_358
timestamp 1569533753
transform 1 0 4584 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_359
timestamp 1569533753
transform 1 0 4648 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_360
timestamp 1569533753
transform 1 0 4712 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_361
timestamp 1569533753
transform 1 0 4840 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_362
timestamp 1569533753
transform 1 0 4904 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_363
timestamp 1569533753
transform 1 0 4776 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_364
timestamp 1569533753
transform 1 0 4776 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_365
timestamp 1569533753
transform 1 0 4712 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_366
timestamp 1569533753
transform 1 0 4904 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_367
timestamp 1569533753
transform 1 0 4840 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_368
timestamp 1569533753
transform 1 0 4776 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_369
timestamp 1569533753
transform 1 0 4712 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_370
timestamp 1569533753
transform 1 0 4904 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_371
timestamp 1569533753
transform 1 0 4840 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_372
timestamp 1569533753
transform 1 0 4840 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_373
timestamp 1569533753
transform 1 0 4712 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_374
timestamp 1569533753
transform 1 0 4840 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_375
timestamp 1569533753
transform 1 0 4712 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_376
timestamp 1569533753
transform 1 0 4904 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_377
timestamp 1569533753
transform 1 0 4776 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_378
timestamp 1569533753
transform 1 0 4776 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_379
timestamp 1569533753
transform 1 0 4904 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_380
timestamp 1569533753
transform 1 0 3688 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_381
timestamp 1569533753
transform 1 0 3560 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_382
timestamp 1569533753
transform 1 0 3624 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_383
timestamp 1569533753
transform 1 0 3496 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_384
timestamp 1569533753
transform 1 0 3560 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_385
timestamp 1569533753
transform 1 0 3560 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_386
timestamp 1569533753
transform 1 0 3496 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_387
timestamp 1569533753
transform 1 0 3624 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_388
timestamp 1569533753
transform 1 0 3688 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_389
timestamp 1569533753
transform 1 0 3688 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_390
timestamp 1569533753
transform 1 0 3688 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_391
timestamp 1569533753
transform 1 0 3496 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_392
timestamp 1569533753
transform 1 0 3496 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_393
timestamp 1569533753
transform 1 0 3688 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_394
timestamp 1569533753
transform 1 0 3560 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_395
timestamp 1569533753
transform 1 0 3624 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_396
timestamp 1569533753
transform 1 0 3624 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_397
timestamp 1569533753
transform 1 0 3496 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_398
timestamp 1569533753
transform 1 0 3624 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_399
timestamp 1569533753
transform 1 0 3560 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_400
timestamp 1569533753
transform 1 0 3368 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_401
timestamp 1569533753
transform 1 0 3240 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_402
timestamp 1569533753
transform 1 0 3176 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_403
timestamp 1569533753
transform 1 0 3368 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_404
timestamp 1569533753
transform 1 0 3304 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_405
timestamp 1569533753
transform 1 0 3240 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_406
timestamp 1569533753
transform 1 0 3304 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_407
timestamp 1569533753
transform 1 0 3368 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_408
timestamp 1569533753
transform 1 0 3176 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_409
timestamp 1569533753
transform 1 0 3240 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_410
timestamp 1569533753
transform 1 0 3176 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_411
timestamp 1569533753
transform 1 0 3304 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_412
timestamp 1569533753
transform 1 0 3176 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_413
timestamp 1569533753
transform 1 0 3368 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_414
timestamp 1569533753
transform 1 0 3304 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_415
timestamp 1569533753
transform 1 0 3304 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_416
timestamp 1569533753
transform 1 0 3176 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_417
timestamp 1569533753
transform 1 0 3240 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_418
timestamp 1569533753
transform 1 0 3368 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_419
timestamp 1569533753
transform 1 0 3240 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_420
timestamp 1569533753
transform 1 0 3240 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_421
timestamp 1569533753
transform 1 0 3240 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_422
timestamp 1569533753
transform 1 0 3176 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_423
timestamp 1569533753
transform 1 0 3176 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_424
timestamp 1569533753
transform 1 0 3368 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_425
timestamp 1569533753
transform 1 0 3176 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_426
timestamp 1569533753
transform 1 0 3240 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_427
timestamp 1569533753
transform 1 0 3176 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_428
timestamp 1569533753
transform 1 0 3176 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_429
timestamp 1569533753
transform 1 0 3368 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_430
timestamp 1569533753
transform 1 0 3240 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_431
timestamp 1569533753
transform 1 0 3368 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_432
timestamp 1569533753
transform 1 0 3368 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_433
timestamp 1569533753
transform 1 0 3368 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_434
timestamp 1569533753
transform 1 0 3304 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_435
timestamp 1569533753
transform 1 0 3304 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_436
timestamp 1569533753
transform 1 0 3304 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_437
timestamp 1569533753
transform 1 0 3240 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_438
timestamp 1569533753
transform 1 0 3304 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_439
timestamp 1569533753
transform 1 0 3304 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_440
timestamp 1569533753
transform 1 0 3560 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_441
timestamp 1569533753
transform 1 0 3624 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_442
timestamp 1569533753
transform 1 0 3496 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_443
timestamp 1569533753
transform 1 0 3560 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_444
timestamp 1569533753
transform 1 0 3688 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_445
timestamp 1569533753
transform 1 0 3688 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_446
timestamp 1569533753
transform 1 0 3624 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_447
timestamp 1569533753
transform 1 0 3560 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_448
timestamp 1569533753
transform 1 0 3688 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_449
timestamp 1569533753
transform 1 0 3560 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_450
timestamp 1569533753
transform 1 0 3624 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_451
timestamp 1569533753
transform 1 0 3688 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_452
timestamp 1569533753
transform 1 0 3688 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_453
timestamp 1569533753
transform 1 0 3496 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_454
timestamp 1569533753
transform 1 0 3560 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_455
timestamp 1569533753
transform 1 0 3624 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_456
timestamp 1569533753
transform 1 0 3496 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_457
timestamp 1569533753
transform 1 0 3496 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_458
timestamp 1569533753
transform 1 0 3624 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_459
timestamp 1569533753
transform 1 0 3496 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_460
timestamp 1569533753
transform 1 0 3432 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_461
timestamp 1569533753
transform 1 0 3432 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_462
timestamp 1569533753
transform 1 0 3432 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_463
timestamp 1569533753
transform 1 0 3432 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_464
timestamp 1569533753
transform 1 0 3432 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_465
timestamp 1569533753
transform 1 0 3432 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_466
timestamp 1569533753
transform 1 0 3432 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_467
timestamp 1569533753
transform 1 0 3432 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_468
timestamp 1569533753
transform 1 0 3432 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_469
timestamp 1569533753
transform 1 0 3432 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_470
timestamp 1569533753
transform 1 0 3048 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_471
timestamp 1569533753
transform 1 0 2920 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_472
timestamp 1569533753
transform 1 0 3048 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_473
timestamp 1569533753
transform 1 0 3048 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_474
timestamp 1569533753
transform 1 0 2920 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_475
timestamp 1569533753
transform 1 0 2984 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_476
timestamp 1569533753
transform 1 0 2984 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_477
timestamp 1569533753
transform 1 0 2920 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_478
timestamp 1569533753
transform 1 0 2984 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_479
timestamp 1569533753
transform 1 0 2920 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_480
timestamp 1569533753
transform 1 0 2856 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_481
timestamp 1569533753
transform 1 0 3048 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_482
timestamp 1569533753
transform 1 0 3112 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_483
timestamp 1569533753
transform 1 0 2856 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_484
timestamp 1569533753
transform 1 0 3048 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_485
timestamp 1569533753
transform 1 0 3112 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_486
timestamp 1569533753
transform 1 0 2920 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_487
timestamp 1569533753
transform 1 0 3112 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_488
timestamp 1569533753
transform 1 0 3112 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_489
timestamp 1569533753
transform 1 0 2856 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_490
timestamp 1569533753
transform 1 0 2984 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_491
timestamp 1569533753
transform 1 0 2856 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_492
timestamp 1569533753
transform 1 0 3112 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_493
timestamp 1569533753
transform 1 0 2984 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_494
timestamp 1569533753
transform 1 0 2856 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_495
timestamp 1569533753
transform 1 0 2792 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_496
timestamp 1569533753
transform 1 0 2664 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_497
timestamp 1569533753
transform 1 0 2728 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_498
timestamp 1569533753
transform 1 0 2792 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_499
timestamp 1569533753
transform 1 0 2728 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_500
timestamp 1569533753
transform 1 0 2664 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_501
timestamp 1569533753
transform 1 0 2536 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_502
timestamp 1569533753
transform 1 0 2536 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_503
timestamp 1569533753
transform 1 0 2664 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_504
timestamp 1569533753
transform 1 0 2664 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_505
timestamp 1569533753
transform 1 0 2536 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_506
timestamp 1569533753
transform 1 0 2792 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_507
timestamp 1569533753
transform 1 0 2728 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_508
timestamp 1569533753
transform 1 0 2600 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_509
timestamp 1569533753
transform 1 0 2664 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_510
timestamp 1569533753
transform 1 0 2792 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_511
timestamp 1569533753
transform 1 0 2728 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_512
timestamp 1569533753
transform 1 0 2600 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_513
timestamp 1569533753
transform 1 0 2600 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_514
timestamp 1569533753
transform 1 0 2536 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_515
timestamp 1569533753
transform 1 0 2600 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_516
timestamp 1569533753
transform 1 0 2600 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_517
timestamp 1569533753
transform 1 0 2728 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_518
timestamp 1569533753
transform 1 0 2536 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_519
timestamp 1569533753
transform 1 0 2792 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_520
timestamp 1569533753
transform 1 0 2728 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_521
timestamp 1569533753
transform 1 0 2792 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_522
timestamp 1569533753
transform 1 0 2728 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_523
timestamp 1569533753
transform 1 0 2792 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_524
timestamp 1569533753
transform 1 0 2728 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_525
timestamp 1569533753
transform 1 0 2792 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_526
timestamp 1569533753
transform 1 0 2664 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_527
timestamp 1569533753
transform 1 0 2664 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_528
timestamp 1569533753
transform 1 0 2792 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_529
timestamp 1569533753
transform 1 0 2792 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_530
timestamp 1569533753
transform 1 0 2664 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_531
timestamp 1569533753
transform 1 0 2536 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_532
timestamp 1569533753
transform 1 0 2664 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_533
timestamp 1569533753
transform 1 0 2664 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_534
timestamp 1569533753
transform 1 0 2536 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_535
timestamp 1569533753
transform 1 0 2536 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_536
timestamp 1569533753
transform 1 0 2536 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_537
timestamp 1569533753
transform 1 0 2600 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_538
timestamp 1569533753
transform 1 0 2728 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_539
timestamp 1569533753
transform 1 0 2600 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_540
timestamp 1569533753
transform 1 0 2728 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_541
timestamp 1569533753
transform 1 0 2600 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_542
timestamp 1569533753
transform 1 0 2600 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_543
timestamp 1569533753
transform 1 0 2600 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_544
timestamp 1569533753
transform 1 0 2536 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_545
timestamp 1569533753
transform 1 0 2856 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_546
timestamp 1569533753
transform 1 0 3048 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_547
timestamp 1569533753
transform 1 0 3048 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_548
timestamp 1569533753
transform 1 0 3048 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_549
timestamp 1569533753
transform 1 0 3048 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_550
timestamp 1569533753
transform 1 0 3048 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_551
timestamp 1569533753
transform 1 0 2856 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_552
timestamp 1569533753
transform 1 0 2984 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_553
timestamp 1569533753
transform 1 0 2856 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_554
timestamp 1569533753
transform 1 0 2856 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_555
timestamp 1569533753
transform 1 0 3112 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_556
timestamp 1569533753
transform 1 0 3112 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_557
timestamp 1569533753
transform 1 0 2920 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_558
timestamp 1569533753
transform 1 0 3112 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_559
timestamp 1569533753
transform 1 0 3112 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_560
timestamp 1569533753
transform 1 0 2984 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_561
timestamp 1569533753
transform 1 0 3112 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_562
timestamp 1569533753
transform 1 0 2920 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_563
timestamp 1569533753
transform 1 0 2984 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_564
timestamp 1569533753
transform 1 0 2856 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_565
timestamp 1569533753
transform 1 0 2920 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_566
timestamp 1569533753
transform 1 0 2984 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_567
timestamp 1569533753
transform 1 0 2920 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_568
timestamp 1569533753
transform 1 0 2920 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_569
timestamp 1569533753
transform 1 0 2984 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_570
timestamp 1569533753
transform 1 0 3048 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_571
timestamp 1569533753
transform 1 0 2920 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_572
timestamp 1569533753
transform 1 0 3112 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_573
timestamp 1569533753
transform 1 0 2984 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_574
timestamp 1569533753
transform 1 0 3048 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_575
timestamp 1569533753
transform 1 0 3112 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_576
timestamp 1569533753
transform 1 0 2856 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_577
timestamp 1569533753
transform 1 0 2920 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_578
timestamp 1569533753
transform 1 0 2856 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_579
timestamp 1569533753
transform 1 0 3112 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_580
timestamp 1569533753
transform 1 0 2984 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_581
timestamp 1569533753
transform 1 0 3048 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_582
timestamp 1569533753
transform 1 0 2984 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_583
timestamp 1569533753
transform 1 0 2920 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_584
timestamp 1569533753
transform 1 0 2856 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_585
timestamp 1569533753
transform 1 0 3112 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_586
timestamp 1569533753
transform 1 0 2856 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_587
timestamp 1569533753
transform 1 0 2920 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_588
timestamp 1569533753
transform 1 0 3048 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_589
timestamp 1569533753
transform 1 0 2920 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_590
timestamp 1569533753
transform 1 0 3112 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_591
timestamp 1569533753
transform 1 0 2984 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_592
timestamp 1569533753
transform 1 0 3048 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_593
timestamp 1569533753
transform 1 0 2856 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_594
timestamp 1569533753
transform 1 0 2984 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_595
timestamp 1569533753
transform 1 0 2728 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_596
timestamp 1569533753
transform 1 0 2664 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_597
timestamp 1569533753
transform 1 0 2536 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_598
timestamp 1569533753
transform 1 0 2728 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_599
timestamp 1569533753
transform 1 0 2728 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_600
timestamp 1569533753
transform 1 0 2600 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_601
timestamp 1569533753
transform 1 0 2792 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_602
timestamp 1569533753
transform 1 0 2600 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_603
timestamp 1569533753
transform 1 0 2792 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_604
timestamp 1569533753
transform 1 0 2600 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_605
timestamp 1569533753
transform 1 0 2664 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_606
timestamp 1569533753
transform 1 0 2600 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_607
timestamp 1569533753
transform 1 0 2728 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_608
timestamp 1569533753
transform 1 0 2792 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_609
timestamp 1569533753
transform 1 0 2728 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_610
timestamp 1569533753
transform 1 0 2600 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_611
timestamp 1569533753
transform 1 0 2664 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_612
timestamp 1569533753
transform 1 0 2792 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_613
timestamp 1569533753
transform 1 0 2536 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_614
timestamp 1569533753
transform 1 0 2664 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_615
timestamp 1569533753
transform 1 0 2536 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_616
timestamp 1569533753
transform 1 0 2664 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_617
timestamp 1569533753
transform 1 0 2536 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_618
timestamp 1569533753
transform 1 0 2792 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_619
timestamp 1569533753
transform 1 0 2536 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_620
timestamp 1569533753
transform 1 0 2792 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_621
timestamp 1569533753
transform 1 0 2664 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_622
timestamp 1569533753
transform 1 0 2536 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_623
timestamp 1569533753
transform 1 0 2664 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_624
timestamp 1569533753
transform 1 0 2792 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_625
timestamp 1569533753
transform 1 0 2536 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_626
timestamp 1569533753
transform 1 0 2600 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_627
timestamp 1569533753
transform 1 0 2792 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_628
timestamp 1569533753
transform 1 0 2792 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_629
timestamp 1569533753
transform 1 0 2536 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_630
timestamp 1569533753
transform 1 0 2728 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_631
timestamp 1569533753
transform 1 0 2600 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_632
timestamp 1569533753
transform 1 0 2600 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_633
timestamp 1569533753
transform 1 0 2664 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_634
timestamp 1569533753
transform 1 0 2536 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_635
timestamp 1569533753
transform 1 0 2728 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_636
timestamp 1569533753
transform 1 0 2664 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_637
timestamp 1569533753
transform 1 0 2728 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_638
timestamp 1569533753
transform 1 0 2792 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_639
timestamp 1569533753
transform 1 0 2664 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_640
timestamp 1569533753
transform 1 0 2728 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_641
timestamp 1569533753
transform 1 0 2600 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_642
timestamp 1569533753
transform 1 0 2600 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_643
timestamp 1569533753
transform 1 0 2536 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_644
timestamp 1569533753
transform 1 0 2728 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_645
timestamp 1569533753
transform 1 0 2920 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_646
timestamp 1569533753
transform 1 0 2856 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_647
timestamp 1569533753
transform 1 0 2920 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_648
timestamp 1569533753
transform 1 0 2920 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_649
timestamp 1569533753
transform 1 0 2856 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_650
timestamp 1569533753
transform 1 0 3112 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_651
timestamp 1569533753
transform 1 0 3112 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_652
timestamp 1569533753
transform 1 0 3048 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_653
timestamp 1569533753
transform 1 0 2856 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_654
timestamp 1569533753
transform 1 0 3112 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_655
timestamp 1569533753
transform 1 0 2856 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_656
timestamp 1569533753
transform 1 0 3112 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_657
timestamp 1569533753
transform 1 0 2984 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_658
timestamp 1569533753
transform 1 0 3048 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_659
timestamp 1569533753
transform 1 0 2856 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_660
timestamp 1569533753
transform 1 0 2984 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_661
timestamp 1569533753
transform 1 0 2984 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_662
timestamp 1569533753
transform 1 0 2984 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_663
timestamp 1569533753
transform 1 0 2920 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_664
timestamp 1569533753
transform 1 0 2984 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_665
timestamp 1569533753
transform 1 0 2920 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_666
timestamp 1569533753
transform 1 0 3048 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_667
timestamp 1569533753
transform 1 0 3112 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_668
timestamp 1569533753
transform 1 0 3048 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_669
timestamp 1569533753
transform 1 0 3048 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_670
timestamp 1569533753
transform 1 0 3496 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_671
timestamp 1569533753
transform 1 0 3624 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_672
timestamp 1569533753
transform 1 0 3560 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_673
timestamp 1569533753
transform 1 0 3496 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_674
timestamp 1569533753
transform 1 0 3624 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_675
timestamp 1569533753
transform 1 0 3560 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_676
timestamp 1569533753
transform 1 0 3496 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_677
timestamp 1569533753
transform 1 0 3560 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_678
timestamp 1569533753
transform 1 0 3688 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_679
timestamp 1569533753
transform 1 0 3496 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_680
timestamp 1569533753
transform 1 0 3688 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_681
timestamp 1569533753
transform 1 0 3624 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_682
timestamp 1569533753
transform 1 0 3688 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_683
timestamp 1569533753
transform 1 0 3496 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_684
timestamp 1569533753
transform 1 0 3560 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_685
timestamp 1569533753
transform 1 0 3688 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_686
timestamp 1569533753
transform 1 0 3560 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_687
timestamp 1569533753
transform 1 0 3688 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_688
timestamp 1569533753
transform 1 0 3624 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_689
timestamp 1569533753
transform 1 0 3624 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_690
timestamp 1569533753
transform 1 0 3240 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_691
timestamp 1569533753
transform 1 0 3240 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_692
timestamp 1569533753
transform 1 0 3368 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_693
timestamp 1569533753
transform 1 0 3304 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_694
timestamp 1569533753
transform 1 0 3304 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_695
timestamp 1569533753
transform 1 0 3304 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_696
timestamp 1569533753
transform 1 0 3304 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_697
timestamp 1569533753
transform 1 0 3304 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_698
timestamp 1569533753
transform 1 0 3368 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_699
timestamp 1569533753
transform 1 0 3368 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_700
timestamp 1569533753
transform 1 0 3368 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_701
timestamp 1569533753
transform 1 0 3176 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_702
timestamp 1569533753
transform 1 0 3176 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_703
timestamp 1569533753
transform 1 0 3176 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_704
timestamp 1569533753
transform 1 0 3176 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_705
timestamp 1569533753
transform 1 0 3176 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_706
timestamp 1569533753
transform 1 0 3368 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_707
timestamp 1569533753
transform 1 0 3240 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_708
timestamp 1569533753
transform 1 0 3240 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_709
timestamp 1569533753
transform 1 0 3240 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_710
timestamp 1569533753
transform 1 0 3368 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_711
timestamp 1569533753
transform 1 0 3176 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_712
timestamp 1569533753
transform 1 0 3368 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_713
timestamp 1569533753
transform 1 0 3176 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_714
timestamp 1569533753
transform 1 0 3368 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_715
timestamp 1569533753
transform 1 0 3368 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_716
timestamp 1569533753
transform 1 0 3240 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_717
timestamp 1569533753
transform 1 0 3304 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_718
timestamp 1569533753
transform 1 0 3176 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_719
timestamp 1569533753
transform 1 0 3240 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_720
timestamp 1569533753
transform 1 0 3368 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_721
timestamp 1569533753
transform 1 0 3240 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_722
timestamp 1569533753
transform 1 0 3304 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_723
timestamp 1569533753
transform 1 0 3176 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_724
timestamp 1569533753
transform 1 0 3304 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_725
timestamp 1569533753
transform 1 0 3240 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_726
timestamp 1569533753
transform 1 0 3304 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_727
timestamp 1569533753
transform 1 0 3240 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_728
timestamp 1569533753
transform 1 0 3304 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_729
timestamp 1569533753
transform 1 0 3176 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_730
timestamp 1569533753
transform 1 0 3624 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_731
timestamp 1569533753
transform 1 0 3624 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_732
timestamp 1569533753
transform 1 0 3496 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_733
timestamp 1569533753
transform 1 0 3624 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_734
timestamp 1569533753
transform 1 0 3560 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_735
timestamp 1569533753
transform 1 0 3688 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_736
timestamp 1569533753
transform 1 0 3560 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_737
timestamp 1569533753
transform 1 0 3560 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_738
timestamp 1569533753
transform 1 0 3688 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_739
timestamp 1569533753
transform 1 0 3624 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_740
timestamp 1569533753
transform 1 0 3688 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_741
timestamp 1569533753
transform 1 0 3624 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_742
timestamp 1569533753
transform 1 0 3496 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_743
timestamp 1569533753
transform 1 0 3560 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_744
timestamp 1569533753
transform 1 0 3496 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_745
timestamp 1569533753
transform 1 0 3496 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_746
timestamp 1569533753
transform 1 0 3688 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_747
timestamp 1569533753
transform 1 0 3496 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_748
timestamp 1569533753
transform 1 0 3560 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_749
timestamp 1569533753
transform 1 0 3688 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_750
timestamp 1569533753
transform 1 0 3432 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_751
timestamp 1569533753
transform 1 0 3432 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_752
timestamp 1569533753
transform 1 0 3432 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_753
timestamp 1569533753
transform 1 0 3432 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_754
timestamp 1569533753
transform 1 0 3432 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_755
timestamp 1569533753
transform 1 0 3432 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_756
timestamp 1569533753
transform 1 0 3432 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_757
timestamp 1569533753
transform 1 0 3432 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_758
timestamp 1569533753
transform 1 0 3432 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_759
timestamp 1569533753
transform 1 0 3432 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_760
timestamp 1569533753
transform 1 0 3688 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_761
timestamp 1569533753
transform 1 0 3368 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_762
timestamp 1569533753
transform 1 0 3624 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_763
timestamp 1569533753
transform 1 0 3496 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_764
timestamp 1569533753
transform 1 0 3432 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_765
timestamp 1569533753
transform 1 0 3304 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_766
timestamp 1569533753
transform 1 0 3176 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_767
timestamp 1569533753
transform 1 0 3688 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_768
timestamp 1569533753
transform 1 0 3432 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_769
timestamp 1569533753
transform 1 0 3432 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_770
timestamp 1569533753
transform 1 0 3624 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_771
timestamp 1569533753
transform 1 0 3176 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_772
timestamp 1569533753
transform 1 0 3240 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_773
timestamp 1569533753
transform 1 0 3240 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_774
timestamp 1569533753
transform 1 0 3176 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_775
timestamp 1569533753
transform 1 0 3560 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_776
timestamp 1569533753
transform 1 0 3496 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_777
timestamp 1569533753
transform 1 0 3432 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_778
timestamp 1569533753
transform 1 0 3560 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_779
timestamp 1569533753
transform 1 0 3624 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_780
timestamp 1569533753
transform 1 0 3624 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_781
timestamp 1569533753
transform 1 0 3240 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_782
timestamp 1569533753
transform 1 0 3176 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_783
timestamp 1569533753
transform 1 0 3688 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_784
timestamp 1569533753
transform 1 0 3304 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_785
timestamp 1569533753
transform 1 0 3240 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_786
timestamp 1569533753
transform 1 0 3304 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_787
timestamp 1569533753
transform 1 0 3688 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_788
timestamp 1569533753
transform 1 0 3496 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_789
timestamp 1569533753
transform 1 0 3304 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_790
timestamp 1569533753
transform 1 0 3368 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_791
timestamp 1569533753
transform 1 0 3496 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_792
timestamp 1569533753
transform 1 0 3368 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_793
timestamp 1569533753
transform 1 0 3560 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_794
timestamp 1569533753
transform 1 0 3560 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_795
timestamp 1569533753
transform 1 0 3368 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_796
timestamp 1569533753
transform 1 0 3112 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_797
timestamp 1569533753
transform 1 0 3048 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_798
timestamp 1569533753
transform 1 0 2920 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_799
timestamp 1569533753
transform 1 0 3112 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_800
timestamp 1569533753
transform 1 0 2984 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_801
timestamp 1569533753
transform 1 0 2984 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_802
timestamp 1569533753
transform 1 0 2920 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_803
timestamp 1569533753
transform 1 0 2856 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_804
timestamp 1569533753
transform 1 0 3048 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_805
timestamp 1569533753
transform 1 0 2920 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_806
timestamp 1569533753
transform 1 0 2984 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_807
timestamp 1569533753
transform 1 0 2920 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_808
timestamp 1569533753
transform 1 0 3112 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_809
timestamp 1569533753
transform 1 0 2856 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_810
timestamp 1569533753
transform 1 0 3112 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_811
timestamp 1569533753
transform 1 0 3048 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_812
timestamp 1569533753
transform 1 0 2984 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_813
timestamp 1569533753
transform 1 0 2856 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_814
timestamp 1569533753
transform 1 0 3048 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_815
timestamp 1569533753
transform 1 0 2856 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_816
timestamp 1569533753
transform 1 0 2664 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_817
timestamp 1569533753
transform 1 0 2600 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_818
timestamp 1569533753
transform 1 0 2792 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_819
timestamp 1569533753
transform 1 0 2664 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_820
timestamp 1569533753
transform 1 0 2728 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_821
timestamp 1569533753
transform 1 0 2536 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_822
timestamp 1569533753
transform 1 0 2728 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_823
timestamp 1569533753
transform 1 0 2728 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_824
timestamp 1569533753
transform 1 0 2664 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_825
timestamp 1569533753
transform 1 0 2600 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_826
timestamp 1569533753
transform 1 0 2792 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_827
timestamp 1569533753
transform 1 0 2536 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_828
timestamp 1569533753
transform 1 0 2728 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_829
timestamp 1569533753
transform 1 0 2792 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_830
timestamp 1569533753
transform 1 0 2792 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_831
timestamp 1569533753
transform 1 0 2600 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_832
timestamp 1569533753
transform 1 0 2536 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_833
timestamp 1569533753
transform 1 0 2664 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_834
timestamp 1569533753
transform 1 0 2600 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_835
timestamp 1569533753
transform 1 0 2536 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_836
timestamp 1569533753
transform 1 0 2664 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_837
timestamp 1569533753
transform 1 0 2600 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_838
timestamp 1569533753
transform 1 0 2536 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_839
timestamp 1569533753
transform 1 0 2728 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_840
timestamp 1569533753
transform 1 0 2536 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_841
timestamp 1569533753
transform 1 0 2600 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_842
timestamp 1569533753
transform 1 0 2600 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_843
timestamp 1569533753
transform 1 0 2600 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_844
timestamp 1569533753
transform 1 0 2792 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_845
timestamp 1569533753
transform 1 0 2664 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_846
timestamp 1569533753
transform 1 0 2664 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_847
timestamp 1569533753
transform 1 0 2536 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_848
timestamp 1569533753
transform 1 0 2536 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_849
timestamp 1569533753
transform 1 0 2728 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_850
timestamp 1569533753
transform 1 0 2664 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_851
timestamp 1569533753
transform 1 0 2536 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_852
timestamp 1569533753
transform 1 0 2600 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_853
timestamp 1569533753
transform 1 0 2728 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_854
timestamp 1569533753
transform 1 0 2792 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_855
timestamp 1569533753
transform 1 0 2856 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_856
timestamp 1569533753
transform 1 0 2536 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_857
timestamp 1569533753
transform 1 0 3688 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_858
timestamp 1569533753
transform 1 0 3624 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_859
timestamp 1569533753
transform 1 0 3688 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_860
timestamp 1569533753
transform 1 0 3688 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_861
timestamp 1569533753
transform 1 0 3240 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_862
timestamp 1569533753
transform 1 0 3432 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_863
timestamp 1569533753
transform 1 0 3432 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_864
timestamp 1569533753
transform 1 0 3432 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_865
timestamp 1569533753
transform 1 0 3496 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_866
timestamp 1569533753
transform 1 0 3496 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_867
timestamp 1569533753
transform 1 0 3496 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_868
timestamp 1569533753
transform 1 0 3304 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_869
timestamp 1569533753
transform 1 0 3304 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_870
timestamp 1569533753
transform 1 0 3560 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_871
timestamp 1569533753
transform 1 0 3560 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_872
timestamp 1569533753
transform 1 0 3560 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_873
timestamp 1569533753
transform 1 0 3368 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_874
timestamp 1569533753
transform 1 0 3368 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_875
timestamp 1569533753
transform 1 0 3624 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_876
timestamp 1569533753
transform 1 0 3368 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_877
timestamp 1569533753
transform 1 0 3624 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_878
timestamp 1569533753
transform 1 0 4648 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_879
timestamp 1569533753
transform 1 0 4712 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_880
timestamp 1569533753
transform 1 0 4392 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_881
timestamp 1569533753
transform 1 0 4904 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_882
timestamp 1569533753
transform 1 0 4712 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_883
timestamp 1569533753
transform 1 0 4584 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_884
timestamp 1569533753
transform 1 0 4456 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_885
timestamp 1569533753
transform 1 0 4584 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_886
timestamp 1569533753
transform 1 0 4712 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_887
timestamp 1569533753
transform 1 0 4456 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_888
timestamp 1569533753
transform 1 0 4840 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_889
timestamp 1569533753
transform 1 0 4776 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_890
timestamp 1569533753
transform 1 0 4648 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_891
timestamp 1569533753
transform 1 0 4840 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_892
timestamp 1569533753
transform 1 0 4776 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_893
timestamp 1569533753
transform 1 0 4456 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_894
timestamp 1569533753
transform 1 0 4584 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_895
timestamp 1569533753
transform 1 0 4520 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_896
timestamp 1569533753
transform 1 0 4840 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_897
timestamp 1569533753
transform 1 0 4776 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_898
timestamp 1569533753
transform 1 0 4776 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_899
timestamp 1569533753
transform 1 0 4520 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_900
timestamp 1569533753
transform 1 0 4392 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_901
timestamp 1569533753
transform 1 0 4904 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_902
timestamp 1569533753
transform 1 0 4520 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_903
timestamp 1569533753
transform 1 0 4520 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_904
timestamp 1569533753
transform 1 0 4648 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_905
timestamp 1569533753
transform 1 0 4648 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_906
timestamp 1569533753
transform 1 0 4712 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_907
timestamp 1569533753
transform 1 0 4584 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_908
timestamp 1569533753
transform 1 0 4456 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_909
timestamp 1569533753
transform 1 0 4392 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_910
timestamp 1569533753
transform 1 0 4904 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_911
timestamp 1569533753
transform 1 0 4392 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_912
timestamp 1569533753
transform 1 0 4904 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_913
timestamp 1569533753
transform 1 0 4840 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_914
timestamp 1569533753
transform 1 0 4072 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_915
timestamp 1569533753
transform 1 0 3944 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_916
timestamp 1569533753
transform 1 0 3880 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_917
timestamp 1569533753
transform 1 0 4136 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_918
timestamp 1569533753
transform 1 0 3880 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_919
timestamp 1569533753
transform 1 0 3944 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_920
timestamp 1569533753
transform 1 0 4200 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_921
timestamp 1569533753
transform 1 0 4200 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_922
timestamp 1569533753
transform 1 0 3880 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_923
timestamp 1569533753
transform 1 0 3944 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_924
timestamp 1569533753
transform 1 0 4200 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_925
timestamp 1569533753
transform 1 0 3944 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_926
timestamp 1569533753
transform 1 0 3752 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_927
timestamp 1569533753
transform 1 0 4136 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_928
timestamp 1569533753
transform 1 0 4200 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_929
timestamp 1569533753
transform 1 0 4264 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_930
timestamp 1569533753
transform 1 0 4008 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_931
timestamp 1569533753
transform 1 0 4008 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_932
timestamp 1569533753
transform 1 0 3752 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_933
timestamp 1569533753
transform 1 0 4264 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_934
timestamp 1569533753
transform 1 0 3880 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_935
timestamp 1569533753
transform 1 0 4008 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_936
timestamp 1569533753
transform 1 0 3816 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_937
timestamp 1569533753
transform 1 0 3752 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_938
timestamp 1569533753
transform 1 0 4264 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_939
timestamp 1569533753
transform 1 0 4328 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_940
timestamp 1569533753
transform 1 0 4264 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_941
timestamp 1569533753
transform 1 0 3752 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_942
timestamp 1569533753
transform 1 0 4072 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_943
timestamp 1569533753
transform 1 0 4136 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_944
timestamp 1569533753
transform 1 0 3816 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_945
timestamp 1569533753
transform 1 0 4328 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_946
timestamp 1569533753
transform 1 0 4072 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_947
timestamp 1569533753
transform 1 0 3816 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_948
timestamp 1569533753
transform 1 0 4328 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_949
timestamp 1569533753
transform 1 0 4072 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_950
timestamp 1569533753
transform 1 0 3816 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_951
timestamp 1569533753
transform 1 0 4328 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_952
timestamp 1569533753
transform 1 0 4008 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_953
timestamp 1569533753
transform 1 0 4136 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_954
timestamp 1569533753
transform 1 0 4072 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_955
timestamp 1569533753
transform 1 0 4072 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_956
timestamp 1569533753
transform 1 0 3752 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_957
timestamp 1569533753
transform 1 0 4072 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_958
timestamp 1569533753
transform 1 0 3880 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_959
timestamp 1569533753
transform 1 0 3816 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_960
timestamp 1569533753
transform 1 0 3880 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_961
timestamp 1569533753
transform 1 0 4136 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_962
timestamp 1569533753
transform 1 0 3880 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_963
timestamp 1569533753
transform 1 0 3752 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_964
timestamp 1569533753
transform 1 0 4136 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_965
timestamp 1569533753
transform 1 0 4136 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_966
timestamp 1569533753
transform 1 0 3944 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_967
timestamp 1569533753
transform 1 0 4328 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_968
timestamp 1569533753
transform 1 0 4200 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_969
timestamp 1569533753
transform 1 0 3944 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_970
timestamp 1569533753
transform 1 0 4200 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_971
timestamp 1569533753
transform 1 0 3944 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_972
timestamp 1569533753
transform 1 0 4328 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_973
timestamp 1569533753
transform 1 0 4200 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_974
timestamp 1569533753
transform 1 0 4328 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_975
timestamp 1569533753
transform 1 0 4264 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_976
timestamp 1569533753
transform 1 0 3816 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_977
timestamp 1569533753
transform 1 0 4264 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_978
timestamp 1569533753
transform 1 0 4264 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_979
timestamp 1569533753
transform 1 0 4008 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_980
timestamp 1569533753
transform 1 0 4008 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_981
timestamp 1569533753
transform 1 0 3816 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_982
timestamp 1569533753
transform 1 0 4008 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_983
timestamp 1569533753
transform 1 0 3752 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_984
timestamp 1569533753
transform 1 0 4520 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_985
timestamp 1569533753
transform 1 0 4520 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_986
timestamp 1569533753
transform 1 0 4520 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_987
timestamp 1569533753
transform 1 0 4584 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_988
timestamp 1569533753
transform 1 0 4584 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_989
timestamp 1569533753
transform 1 0 4584 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_990
timestamp 1569533753
transform 1 0 4456 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_991
timestamp 1569533753
transform 1 0 4648 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_992
timestamp 1569533753
transform 1 0 4648 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_993
timestamp 1569533753
transform 1 0 4648 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_994
timestamp 1569533753
transform 1 0 4712 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_995
timestamp 1569533753
transform 1 0 4712 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_996
timestamp 1569533753
transform 1 0 4712 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_997
timestamp 1569533753
transform 1 0 4776 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_998
timestamp 1569533753
transform 1 0 4776 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_999
timestamp 1569533753
transform 1 0 4776 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1000
timestamp 1569533753
transform 1 0 4840 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1001
timestamp 1569533753
transform 1 0 4840 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1002
timestamp 1569533753
transform 1 0 4840 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1003
timestamp 1569533753
transform 1 0 4904 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1004
timestamp 1569533753
transform 1 0 4904 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1005
timestamp 1569533753
transform 1 0 4904 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1006
timestamp 1569533753
transform 1 0 4392 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1007
timestamp 1569533753
transform 1 0 4392 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1008
timestamp 1569533753
transform 1 0 4392 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1009
timestamp 1569533753
transform 1 0 4456 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1010
timestamp 1569533753
transform 1 0 4456 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1011
timestamp 1569533753
transform 1 0 2472 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1012
timestamp 1569533753
transform 1 0 2472 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1013
timestamp 1569533753
transform 1 0 2344 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1014
timestamp 1569533753
transform 1 0 2216 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1015
timestamp 1569533753
transform 1 0 2408 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1016
timestamp 1569533753
transform 1 0 2344 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1017
timestamp 1569533753
transform 1 0 2216 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1018
timestamp 1569533753
transform 1 0 2344 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1019
timestamp 1569533753
transform 1 0 2472 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1020
timestamp 1569533753
transform 1 0 2280 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1021
timestamp 1569533753
transform 1 0 2408 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1022
timestamp 1569533753
transform 1 0 2216 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1023
timestamp 1569533753
transform 1 0 2344 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1024
timestamp 1569533753
transform 1 0 2344 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1025
timestamp 1569533753
transform 1 0 2408 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1026
timestamp 1569533753
transform 1 0 2280 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1027
timestamp 1569533753
transform 1 0 2280 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1028
timestamp 1569533753
transform 1 0 2408 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1029
timestamp 1569533753
transform 1 0 2408 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1030
timestamp 1569533753
transform 1 0 2280 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1031
timestamp 1569533753
transform 1 0 2472 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1032
timestamp 1569533753
transform 1 0 2216 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1033
timestamp 1569533753
transform 1 0 2216 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1034
timestamp 1569533753
transform 1 0 2472 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1035
timestamp 1569533753
transform 1 0 2280 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1036
timestamp 1569533753
transform 1 0 2088 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1037
timestamp 1569533753
transform 1 0 2088 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1038
timestamp 1569533753
transform 1 0 1960 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1039
timestamp 1569533753
transform 1 0 2088 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1040
timestamp 1569533753
transform 1 0 2088 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1041
timestamp 1569533753
transform 1 0 2152 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1042
timestamp 1569533753
transform 1 0 2152 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1043
timestamp 1569533753
transform 1 0 1960 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1044
timestamp 1569533753
transform 1 0 2152 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1045
timestamp 1569533753
transform 1 0 1960 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1046
timestamp 1569533753
transform 1 0 1960 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1047
timestamp 1569533753
transform 1 0 1960 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1048
timestamp 1569533753
transform 1 0 2024 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1049
timestamp 1569533753
transform 1 0 2024 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1050
timestamp 1569533753
transform 1 0 2024 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1051
timestamp 1569533753
transform 1 0 1896 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1052
timestamp 1569533753
transform 1 0 2152 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1053
timestamp 1569533753
transform 1 0 1896 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1054
timestamp 1569533753
transform 1 0 2024 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1055
timestamp 1569533753
transform 1 0 2024 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1056
timestamp 1569533753
transform 1 0 1896 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1057
timestamp 1569533753
transform 1 0 2152 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1058
timestamp 1569533753
transform 1 0 1896 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1059
timestamp 1569533753
transform 1 0 2088 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1060
timestamp 1569533753
transform 1 0 1896 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1061
timestamp 1569533753
transform 1 0 1896 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1062
timestamp 1569533753
transform 1 0 2152 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1063
timestamp 1569533753
transform 1 0 1960 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1064
timestamp 1569533753
transform 1 0 1960 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1065
timestamp 1569533753
transform 1 0 1960 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1066
timestamp 1569533753
transform 1 0 1960 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1067
timestamp 1569533753
transform 1 0 2152 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1068
timestamp 1569533753
transform 1 0 1960 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1069
timestamp 1569533753
transform 1 0 2152 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1070
timestamp 1569533753
transform 1 0 2024 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1071
timestamp 1569533753
transform 1 0 2024 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1072
timestamp 1569533753
transform 1 0 2024 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1073
timestamp 1569533753
transform 1 0 2024 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1074
timestamp 1569533753
transform 1 0 2024 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1075
timestamp 1569533753
transform 1 0 2152 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1076
timestamp 1569533753
transform 1 0 2152 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1077
timestamp 1569533753
transform 1 0 1896 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1078
timestamp 1569533753
transform 1 0 2088 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1079
timestamp 1569533753
transform 1 0 1896 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1080
timestamp 1569533753
transform 1 0 1896 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1081
timestamp 1569533753
transform 1 0 2088 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1082
timestamp 1569533753
transform 1 0 2088 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1083
timestamp 1569533753
transform 1 0 2088 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1084
timestamp 1569533753
transform 1 0 1896 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1085
timestamp 1569533753
transform 1 0 2088 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1086
timestamp 1569533753
transform 1 0 2344 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1087
timestamp 1569533753
transform 1 0 2344 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1088
timestamp 1569533753
transform 1 0 2344 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1089
timestamp 1569533753
transform 1 0 2472 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1090
timestamp 1569533753
transform 1 0 2472 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1091
timestamp 1569533753
transform 1 0 2472 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1092
timestamp 1569533753
transform 1 0 2472 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1093
timestamp 1569533753
transform 1 0 2472 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1094
timestamp 1569533753
transform 1 0 2344 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1095
timestamp 1569533753
transform 1 0 2216 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1096
timestamp 1569533753
transform 1 0 2216 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1097
timestamp 1569533753
transform 1 0 2216 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1098
timestamp 1569533753
transform 1 0 2216 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1099
timestamp 1569533753
transform 1 0 2344 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1100
timestamp 1569533753
transform 1 0 2216 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1101
timestamp 1569533753
transform 1 0 2408 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1102
timestamp 1569533753
transform 1 0 2408 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1103
timestamp 1569533753
transform 1 0 2408 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1104
timestamp 1569533753
transform 1 0 2408 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1105
timestamp 1569533753
transform 1 0 2408 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1106
timestamp 1569533753
transform 1 0 2280 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1107
timestamp 1569533753
transform 1 0 2280 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1108
timestamp 1569533753
transform 1 0 2280 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1109
timestamp 1569533753
transform 1 0 2280 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1110
timestamp 1569533753
transform 1 0 2280 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1111
timestamp 1569533753
transform 1 0 1832 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1112
timestamp 1569533753
transform 1 0 1768 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1113
timestamp 1569533753
transform 1 0 1768 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1114
timestamp 1569533753
transform 1 0 1768 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1115
timestamp 1569533753
transform 1 0 1768 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1116
timestamp 1569533753
transform 1 0 1640 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1117
timestamp 1569533753
transform 1 0 1832 0 1 40
box -8 -8 8 8
use VIA2$3  VIA2$3_1118
timestamp 1569533753
transform 1 0 1832 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1119
timestamp 1569533753
transform 1 0 1832 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1120
timestamp 1569533753
transform 1 0 1768 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1121
timestamp 1569533753
transform 1 0 1832 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1122
timestamp 1569533753
transform 1 0 1704 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1123
timestamp 1569533753
transform 1 0 1704 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1124
timestamp 1569533753
transform 1 0 1640 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1125
timestamp 1569533753
transform 1 0 1640 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1126
timestamp 1569533753
transform 1 0 1704 0 1 104
box -8 -8 8 8
use VIA2$3  VIA2$3_1127
timestamp 1569533753
transform 1 0 1704 0 1 168
box -8 -8 8 8
use VIA2$3  VIA2$3_1128
timestamp 1569533753
transform 1 0 1512 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1129
timestamp 1569533753
transform 1 0 1320 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1130
timestamp 1569533753
transform 1 0 1320 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1131
timestamp 1569533753
transform 1 0 1320 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1132
timestamp 1569533753
transform 1 0 1512 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1133
timestamp 1569533753
transform 1 0 1512 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1134
timestamp 1569533753
transform 1 0 1448 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1135
timestamp 1569533753
transform 1 0 1448 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1136
timestamp 1569533753
transform 1 0 1384 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1137
timestamp 1569533753
transform 1 0 1384 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1138
timestamp 1569533753
transform 1 0 1384 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1139
timestamp 1569533753
transform 1 0 1384 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1140
timestamp 1569533753
transform 1 0 1512 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1141
timestamp 1569533753
transform 1 0 1512 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1142
timestamp 1569533753
transform 1 0 1448 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1143
timestamp 1569533753
transform 1 0 1512 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1144
timestamp 1569533753
transform 1 0 1448 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1145
timestamp 1569533753
transform 1 0 1448 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1146
timestamp 1569533753
transform 1 0 1640 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1147
timestamp 1569533753
transform 1 0 1640 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1148
timestamp 1569533753
transform 1 0 1704 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1149
timestamp 1569533753
transform 1 0 1704 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1150
timestamp 1569533753
transform 1 0 1832 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1151
timestamp 1569533753
transform 1 0 1832 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1152
timestamp 1569533753
transform 1 0 1832 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1153
timestamp 1569533753
transform 1 0 1832 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1154
timestamp 1569533753
transform 1 0 1832 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1155
timestamp 1569533753
transform 1 0 1768 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1156
timestamp 1569533753
transform 1 0 1768 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1157
timestamp 1569533753
transform 1 0 1768 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1158
timestamp 1569533753
transform 1 0 1704 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1159
timestamp 1569533753
transform 1 0 1640 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1160
timestamp 1569533753
transform 1 0 1640 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1161
timestamp 1569533753
transform 1 0 1640 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1162
timestamp 1569533753
transform 1 0 1704 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1163
timestamp 1569533753
transform 1 0 1704 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1164
timestamp 1569533753
transform 1 0 1768 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1165
timestamp 1569533753
transform 1 0 1768 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1166
timestamp 1569533753
transform 1 0 1576 0 1 296
box -8 -8 8 8
use VIA2$3  VIA2$3_1167
timestamp 1569533753
transform 1 0 1576 0 1 360
box -8 -8 8 8
use VIA2$3  VIA2$3_1168
timestamp 1569533753
transform 1 0 1576 0 1 424
box -8 -8 8 8
use VIA2$3  VIA2$3_1169
timestamp 1569533753
transform 1 0 1576 0 1 488
box -8 -8 8 8
use VIA2$3  VIA2$3_1170
timestamp 1569533753
transform 1 0 1576 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1171
timestamp 1569533753
transform 1 0 1576 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1172
timestamp 1569533753
transform 1 0 1576 0 1 232
box -8 -8 8 8
use VIA2$3  VIA2$3_1173
timestamp 1569533753
transform 1 0 1640 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1174
timestamp 1569533753
transform 1 0 1704 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1175
timestamp 1569533753
transform 1 0 1640 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1176
timestamp 1569533753
transform 1 0 1704 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1177
timestamp 1569533753
transform 1 0 1768 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1178
timestamp 1569533753
transform 1 0 1832 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1179
timestamp 1569533753
transform 1 0 1704 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1180
timestamp 1569533753
transform 1 0 1832 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1181
timestamp 1569533753
transform 1 0 1640 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1182
timestamp 1569533753
transform 1 0 1768 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1183
timestamp 1569533753
transform 1 0 1832 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1184
timestamp 1569533753
transform 1 0 1768 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1185
timestamp 1569533753
transform 1 0 1640 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1186
timestamp 1569533753
transform 1 0 1832 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1187
timestamp 1569533753
transform 1 0 1768 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1188
timestamp 1569533753
transform 1 0 1704 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1189
timestamp 1569533753
transform 1 0 1704 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1190
timestamp 1569533753
transform 1 0 1832 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1191
timestamp 1569533753
transform 1 0 1768 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1192
timestamp 1569533753
transform 1 0 1640 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1193
timestamp 1569533753
transform 1 0 1512 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1194
timestamp 1569533753
transform 1 0 1512 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1195
timestamp 1569533753
transform 1 0 1320 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1196
timestamp 1569533753
transform 1 0 1320 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1197
timestamp 1569533753
transform 1 0 1320 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1198
timestamp 1569533753
transform 1 0 1320 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1199
timestamp 1569533753
transform 1 0 1320 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1200
timestamp 1569533753
transform 1 0 1384 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1201
timestamp 1569533753
transform 1 0 1384 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1202
timestamp 1569533753
transform 1 0 1448 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1203
timestamp 1569533753
transform 1 0 1384 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1204
timestamp 1569533753
transform 1 0 1384 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1205
timestamp 1569533753
transform 1 0 1448 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1206
timestamp 1569533753
transform 1 0 1384 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1207
timestamp 1569533753
transform 1 0 1512 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1208
timestamp 1569533753
transform 1 0 1448 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1209
timestamp 1569533753
transform 1 0 1448 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1210
timestamp 1569533753
transform 1 0 1512 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1211
timestamp 1569533753
transform 1 0 1448 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1212
timestamp 1569533753
transform 1 0 1512 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1213
timestamp 1569533753
transform 1 0 1320 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1214
timestamp 1569533753
transform 1 0 1320 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1215
timestamp 1569533753
transform 1 0 1384 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1216
timestamp 1569533753
transform 1 0 1448 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1217
timestamp 1569533753
transform 1 0 1512 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1218
timestamp 1569533753
transform 1 0 1384 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1219
timestamp 1569533753
transform 1 0 1512 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1220
timestamp 1569533753
transform 1 0 1512 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1221
timestamp 1569533753
transform 1 0 1384 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1222
timestamp 1569533753
transform 1 0 1448 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1223
timestamp 1569533753
transform 1 0 1384 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1224
timestamp 1569533753
transform 1 0 1512 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1225
timestamp 1569533753
transform 1 0 1320 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1226
timestamp 1569533753
transform 1 0 1448 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1227
timestamp 1569533753
transform 1 0 1320 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1228
timestamp 1569533753
transform 1 0 1448 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1229
timestamp 1569533753
transform 1 0 1512 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1230
timestamp 1569533753
transform 1 0 1448 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1231
timestamp 1569533753
transform 1 0 1384 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1232
timestamp 1569533753
transform 1 0 1320 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1233
timestamp 1569533753
transform 1 0 1832 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1234
timestamp 1569533753
transform 1 0 1768 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1235
timestamp 1569533753
transform 1 0 1768 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1236
timestamp 1569533753
transform 1 0 1768 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1237
timestamp 1569533753
transform 1 0 1640 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1238
timestamp 1569533753
transform 1 0 1640 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1239
timestamp 1569533753
transform 1 0 1832 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1240
timestamp 1569533753
transform 1 0 1704 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1241
timestamp 1569533753
transform 1 0 1832 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1242
timestamp 1569533753
transform 1 0 1832 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1243
timestamp 1569533753
transform 1 0 1832 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1244
timestamp 1569533753
transform 1 0 1704 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1245
timestamp 1569533753
transform 1 0 1768 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1246
timestamp 1569533753
transform 1 0 1768 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1247
timestamp 1569533753
transform 1 0 1640 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1248
timestamp 1569533753
transform 1 0 1640 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1249
timestamp 1569533753
transform 1 0 1704 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1250
timestamp 1569533753
transform 1 0 1704 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1251
timestamp 1569533753
transform 1 0 1704 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1252
timestamp 1569533753
transform 1 0 1640 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1253
timestamp 1569533753
transform 1 0 1576 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1254
timestamp 1569533753
transform 1 0 1576 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1255
timestamp 1569533753
transform 1 0 1576 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1256
timestamp 1569533753
transform 1 0 1576 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1257
timestamp 1569533753
transform 1 0 1576 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1258
timestamp 1569533753
transform 1 0 1576 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1259
timestamp 1569533753
transform 1 0 1576 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1260
timestamp 1569533753
transform 1 0 1576 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1261
timestamp 1569533753
transform 1 0 1576 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1262
timestamp 1569533753
transform 1 0 1576 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1263
timestamp 1569533753
transform 1 0 2280 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1264
timestamp 1569533753
transform 1 0 2344 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1265
timestamp 1569533753
transform 1 0 2472 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1266
timestamp 1569533753
transform 1 0 2472 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1267
timestamp 1569533753
transform 1 0 2472 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1268
timestamp 1569533753
transform 1 0 2344 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1269
timestamp 1569533753
transform 1 0 2216 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1270
timestamp 1569533753
transform 1 0 2216 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1271
timestamp 1569533753
transform 1 0 2216 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1272
timestamp 1569533753
transform 1 0 2408 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1273
timestamp 1569533753
transform 1 0 2216 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1274
timestamp 1569533753
transform 1 0 2216 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1275
timestamp 1569533753
transform 1 0 2408 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1276
timestamp 1569533753
transform 1 0 2472 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1277
timestamp 1569533753
transform 1 0 2344 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1278
timestamp 1569533753
transform 1 0 2408 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1279
timestamp 1569533753
transform 1 0 2344 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1280
timestamp 1569533753
transform 1 0 2344 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1281
timestamp 1569533753
transform 1 0 2408 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1282
timestamp 1569533753
transform 1 0 2408 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1283
timestamp 1569533753
transform 1 0 2472 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1284
timestamp 1569533753
transform 1 0 2280 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1285
timestamp 1569533753
transform 1 0 2280 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1286
timestamp 1569533753
transform 1 0 2280 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1287
timestamp 1569533753
transform 1 0 2280 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1288
timestamp 1569533753
transform 1 0 1896 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1289
timestamp 1569533753
transform 1 0 1896 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1290
timestamp 1569533753
transform 1 0 1896 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1291
timestamp 1569533753
transform 1 0 1896 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1292
timestamp 1569533753
transform 1 0 2152 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1293
timestamp 1569533753
transform 1 0 1896 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1294
timestamp 1569533753
transform 1 0 1960 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1295
timestamp 1569533753
transform 1 0 1960 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1296
timestamp 1569533753
transform 1 0 1960 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1297
timestamp 1569533753
transform 1 0 1960 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1298
timestamp 1569533753
transform 1 0 1960 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1299
timestamp 1569533753
transform 1 0 2024 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1300
timestamp 1569533753
transform 1 0 2024 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1301
timestamp 1569533753
transform 1 0 2024 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1302
timestamp 1569533753
transform 1 0 2024 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1303
timestamp 1569533753
transform 1 0 2024 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1304
timestamp 1569533753
transform 1 0 2088 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1305
timestamp 1569533753
transform 1 0 2088 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1306
timestamp 1569533753
transform 1 0 2088 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1307
timestamp 1569533753
transform 1 0 2088 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1308
timestamp 1569533753
transform 1 0 2088 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1309
timestamp 1569533753
transform 1 0 2152 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1310
timestamp 1569533753
transform 1 0 2152 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1311
timestamp 1569533753
transform 1 0 2152 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1312
timestamp 1569533753
transform 1 0 2152 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1313
timestamp 1569533753
transform 1 0 2152 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1314
timestamp 1569533753
transform 1 0 1960 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1315
timestamp 1569533753
transform 1 0 2024 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1316
timestamp 1569533753
transform 1 0 2024 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1317
timestamp 1569533753
transform 1 0 1896 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1318
timestamp 1569533753
transform 1 0 2088 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1319
timestamp 1569533753
transform 1 0 2088 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1320
timestamp 1569533753
transform 1 0 2152 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1321
timestamp 1569533753
transform 1 0 1896 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1322
timestamp 1569533753
transform 1 0 2088 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1323
timestamp 1569533753
transform 1 0 2024 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1324
timestamp 1569533753
transform 1 0 2152 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1325
timestamp 1569533753
transform 1 0 2088 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1326
timestamp 1569533753
transform 1 0 2088 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1327
timestamp 1569533753
transform 1 0 2024 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1328
timestamp 1569533753
transform 1 0 2024 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1329
timestamp 1569533753
transform 1 0 1896 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1330
timestamp 1569533753
transform 1 0 2152 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1331
timestamp 1569533753
transform 1 0 1896 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1332
timestamp 1569533753
transform 1 0 2152 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1333
timestamp 1569533753
transform 1 0 1896 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1334
timestamp 1569533753
transform 1 0 1960 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1335
timestamp 1569533753
transform 1 0 1960 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1336
timestamp 1569533753
transform 1 0 1960 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1337
timestamp 1569533753
transform 1 0 1960 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1338
timestamp 1569533753
transform 1 0 2280 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1339
timestamp 1569533753
transform 1 0 2280 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1340
timestamp 1569533753
transform 1 0 2280 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1341
timestamp 1569533753
transform 1 0 2408 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1342
timestamp 1569533753
transform 1 0 2408 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1343
timestamp 1569533753
transform 1 0 2344 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1344
timestamp 1569533753
transform 1 0 2344 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1345
timestamp 1569533753
transform 1 0 2344 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1346
timestamp 1569533753
transform 1 0 2408 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1347
timestamp 1569533753
transform 1 0 2408 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1348
timestamp 1569533753
transform 1 0 2408 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1349
timestamp 1569533753
transform 1 0 2472 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1350
timestamp 1569533753
transform 1 0 2216 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1351
timestamp 1569533753
transform 1 0 2472 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1352
timestamp 1569533753
transform 1 0 2216 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1353
timestamp 1569533753
transform 1 0 2472 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1354
timestamp 1569533753
transform 1 0 2216 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1355
timestamp 1569533753
transform 1 0 2472 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1356
timestamp 1569533753
transform 1 0 2216 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1357
timestamp 1569533753
transform 1 0 2472 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1358
timestamp 1569533753
transform 1 0 2216 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1359
timestamp 1569533753
transform 1 0 2344 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1360
timestamp 1569533753
transform 1 0 2344 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1361
timestamp 1569533753
transform 1 0 2280 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1362
timestamp 1569533753
transform 1 0 2280 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1363
timestamp 1569533753
transform 1 0 1192 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1364
timestamp 1569533753
transform 1 0 1256 0 1 552
box -8 -8 8 8
use VIA2$3  VIA2$3_1365
timestamp 1569533753
transform 1 0 1256 0 1 616
box -8 -8 8 8
use VIA2$3  VIA2$3_1366
timestamp 1569533753
transform 1 0 616 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1367
timestamp 1569533753
transform 1 0 552 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1368
timestamp 1569533753
transform 1 0 616 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1369
timestamp 1569533753
transform 1 0 1256 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1370
timestamp 1569533753
transform 1 0 1256 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1371
timestamp 1569533753
transform 1 0 1256 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1372
timestamp 1569533753
transform 1 0 1256 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1373
timestamp 1569533753
transform 1 0 1256 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1374
timestamp 1569533753
transform 1 0 1064 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1375
timestamp 1569533753
transform 1 0 1064 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1376
timestamp 1569533753
transform 1 0 1192 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1377
timestamp 1569533753
transform 1 0 1192 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1378
timestamp 1569533753
transform 1 0 1192 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1379
timestamp 1569533753
transform 1 0 1192 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1380
timestamp 1569533753
transform 1 0 1064 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1381
timestamp 1569533753
transform 1 0 1128 0 1 744
box -8 -8 8 8
use VIA2$3  VIA2$3_1382
timestamp 1569533753
transform 1 0 1128 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1383
timestamp 1569533753
transform 1 0 1128 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1384
timestamp 1569533753
transform 1 0 1128 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1385
timestamp 1569533753
transform 1 0 1128 0 1 680
box -8 -8 8 8
use VIA2$3  VIA2$3_1386
timestamp 1569533753
transform 1 0 1064 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1387
timestamp 1569533753
transform 1 0 1000 0 1 808
box -8 -8 8 8
use VIA2$3  VIA2$3_1388
timestamp 1569533753
transform 1 0 1192 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1389
timestamp 1569533753
transform 1 0 1000 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1390
timestamp 1569533753
transform 1 0 1000 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1391
timestamp 1569533753
transform 1 0 936 0 1 872
box -8 -8 8 8
use VIA2$3  VIA2$3_1392
timestamp 1569533753
transform 1 0 936 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1393
timestamp 1569533753
transform 1 0 872 0 1 936
box -8 -8 8 8
use VIA2$3  VIA2$3_1394
timestamp 1569533753
transform 1 0 872 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1395
timestamp 1569533753
transform 1 0 744 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1396
timestamp 1569533753
transform 1 0 744 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1397
timestamp 1569533753
transform 1 0 872 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1398
timestamp 1569533753
transform 1 0 808 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1399
timestamp 1569533753
transform 1 0 872 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1400
timestamp 1569533753
transform 1 0 808 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1401
timestamp 1569533753
transform 1 0 936 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1402
timestamp 1569533753
transform 1 0 808 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1403
timestamp 1569533753
transform 1 0 680 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1404
timestamp 1569533753
transform 1 0 744 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1405
timestamp 1569533753
transform 1 0 936 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1406
timestamp 1569533753
transform 1 0 936 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1407
timestamp 1569533753
transform 1 0 808 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1408
timestamp 1569533753
transform 1 0 680 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1409
timestamp 1569533753
transform 1 0 744 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1410
timestamp 1569533753
transform 1 0 808 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1411
timestamp 1569533753
transform 1 0 936 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1412
timestamp 1569533753
transform 1 0 680 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1413
timestamp 1569533753
transform 1 0 872 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1414
timestamp 1569533753
transform 1 0 936 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1415
timestamp 1569533753
transform 1 0 872 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1416
timestamp 1569533753
transform 1 0 1128 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1417
timestamp 1569533753
transform 1 0 1000 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1418
timestamp 1569533753
transform 1 0 1256 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1419
timestamp 1569533753
transform 1 0 1000 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1420
timestamp 1569533753
transform 1 0 1256 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1421
timestamp 1569533753
transform 1 0 1128 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1422
timestamp 1569533753
transform 1 0 1000 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1423
timestamp 1569533753
transform 1 0 1064 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1424
timestamp 1569533753
transform 1 0 1064 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1425
timestamp 1569533753
transform 1 0 1256 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1426
timestamp 1569533753
transform 1 0 1064 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1427
timestamp 1569533753
transform 1 0 1064 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1428
timestamp 1569533753
transform 1 0 1128 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1429
timestamp 1569533753
transform 1 0 1128 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1430
timestamp 1569533753
transform 1 0 1064 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1431
timestamp 1569533753
transform 1 0 1192 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1432
timestamp 1569533753
transform 1 0 1192 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1433
timestamp 1569533753
transform 1 0 1192 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1434
timestamp 1569533753
transform 1 0 1192 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1435
timestamp 1569533753
transform 1 0 1192 0 1 1000
box -8 -8 8 8
use VIA2$3  VIA2$3_1436
timestamp 1569533753
transform 1 0 1128 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1437
timestamp 1569533753
transform 1 0 1256 0 1 1064
box -8 -8 8 8
use VIA2$3  VIA2$3_1438
timestamp 1569533753
transform 1 0 1000 0 1 1128
box -8 -8 8 8
use VIA2$3  VIA2$3_1439
timestamp 1569533753
transform 1 0 1256 0 1 1192
box -8 -8 8 8
use VIA2$3  VIA2$3_1440
timestamp 1569533753
transform 1 0 1000 0 1 1256
box -8 -8 8 8
use VIA2$3  VIA2$3_1441
timestamp 1569533753
transform 1 0 1000 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1442
timestamp 1569533753
transform 1 0 1256 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1443
timestamp 1569533753
transform 1 0 1128 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1444
timestamp 1569533753
transform 1 0 1064 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1445
timestamp 1569533753
transform 1 0 1000 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1446
timestamp 1569533753
transform 1 0 1256 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1447
timestamp 1569533753
transform 1 0 1000 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1448
timestamp 1569533753
transform 1 0 1192 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1449
timestamp 1569533753
transform 1 0 1064 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1450
timestamp 1569533753
transform 1 0 1064 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1451
timestamp 1569533753
transform 1 0 1192 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1452
timestamp 1569533753
transform 1 0 1192 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1453
timestamp 1569533753
transform 1 0 1128 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1454
timestamp 1569533753
transform 1 0 1064 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1455
timestamp 1569533753
transform 1 0 1256 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1456
timestamp 1569533753
transform 1 0 1256 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1457
timestamp 1569533753
transform 1 0 1192 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1458
timestamp 1569533753
transform 1 0 1000 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1459
timestamp 1569533753
transform 1 0 1128 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1460
timestamp 1569533753
transform 1 0 1128 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1461
timestamp 1569533753
transform 1 0 744 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1462
timestamp 1569533753
transform 1 0 680 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1463
timestamp 1569533753
transform 1 0 936 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1464
timestamp 1569533753
transform 1 0 744 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1465
timestamp 1569533753
transform 1 0 680 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1466
timestamp 1569533753
transform 1 0 936 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1467
timestamp 1569533753
transform 1 0 808 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1468
timestamp 1569533753
transform 1 0 936 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1469
timestamp 1569533753
transform 1 0 872 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1470
timestamp 1569533753
transform 1 0 808 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1471
timestamp 1569533753
transform 1 0 744 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1472
timestamp 1569533753
transform 1 0 872 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1473
timestamp 1569533753
transform 1 0 872 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1474
timestamp 1569533753
transform 1 0 808 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1475
timestamp 1569533753
transform 1 0 936 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1476
timestamp 1569533753
transform 1 0 680 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1477
timestamp 1569533753
transform 1 0 872 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1478
timestamp 1569533753
transform 1 0 808 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1479
timestamp 1569533753
transform 1 0 680 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1480
timestamp 1569533753
transform 1 0 744 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1481
timestamp 1569533753
transform 1 0 808 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1482
timestamp 1569533753
transform 1 0 936 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1483
timestamp 1569533753
transform 1 0 872 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1484
timestamp 1569533753
transform 1 0 808 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1485
timestamp 1569533753
transform 1 0 808 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1486
timestamp 1569533753
transform 1 0 936 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1487
timestamp 1569533753
transform 1 0 936 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1488
timestamp 1569533753
transform 1 0 872 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1489
timestamp 1569533753
transform 1 0 680 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1490
timestamp 1569533753
transform 1 0 744 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1491
timestamp 1569533753
transform 1 0 680 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1492
timestamp 1569533753
transform 1 0 680 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1493
timestamp 1569533753
transform 1 0 872 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1494
timestamp 1569533753
transform 1 0 744 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1495
timestamp 1569533753
transform 1 0 744 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1496
timestamp 1569533753
transform 1 0 808 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1497
timestamp 1569533753
transform 1 0 936 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1498
timestamp 1569533753
transform 1 0 744 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1499
timestamp 1569533753
transform 1 0 680 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1500
timestamp 1569533753
transform 1 0 872 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1501
timestamp 1569533753
transform 1 0 1000 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1502
timestamp 1569533753
transform 1 0 1256 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1503
timestamp 1569533753
transform 1 0 1128 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1504
timestamp 1569533753
transform 1 0 1064 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1505
timestamp 1569533753
transform 1 0 1256 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1506
timestamp 1569533753
transform 1 0 1256 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1507
timestamp 1569533753
transform 1 0 1000 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1508
timestamp 1569533753
transform 1 0 1128 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1509
timestamp 1569533753
transform 1 0 1192 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1510
timestamp 1569533753
transform 1 0 1192 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1511
timestamp 1569533753
transform 1 0 1000 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1512
timestamp 1569533753
transform 1 0 1000 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1513
timestamp 1569533753
transform 1 0 1256 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1514
timestamp 1569533753
transform 1 0 1064 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1515
timestamp 1569533753
transform 1 0 1064 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1516
timestamp 1569533753
transform 1 0 1064 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1517
timestamp 1569533753
transform 1 0 1128 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1518
timestamp 1569533753
transform 1 0 1128 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1519
timestamp 1569533753
transform 1 0 1192 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1520
timestamp 1569533753
transform 1 0 1192 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1521
timestamp 1569533753
transform 1 0 872 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1522
timestamp 1569533753
transform 1 0 1128 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1523
timestamp 1569533753
transform 1 0 936 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1524
timestamp 1569533753
transform 1 0 808 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1525
timestamp 1569533753
transform 1 0 1064 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1526
timestamp 1569533753
transform 1 0 680 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1527
timestamp 1569533753
transform 1 0 1000 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1528
timestamp 1569533753
transform 1 0 1192 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1529
timestamp 1569533753
transform 1 0 1256 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1530
timestamp 1569533753
transform 1 0 744 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1531
timestamp 1569533753
transform 1 0 488 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1532
timestamp 1569533753
transform 1 0 488 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1533
timestamp 1569533753
transform 1 0 424 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1534
timestamp 1569533753
transform 1 0 616 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1535
timestamp 1569533753
transform 1 0 552 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1536
timestamp 1569533753
transform 1 0 616 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1537
timestamp 1569533753
transform 1 0 552 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1538
timestamp 1569533753
transform 1 0 424 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1539
timestamp 1569533753
transform 1 0 616 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1540
timestamp 1569533753
transform 1 0 552 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1541
timestamp 1569533753
transform 1 0 616 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1542
timestamp 1569533753
transform 1 0 360 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1543
timestamp 1569533753
transform 1 0 488 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1544
timestamp 1569533753
transform 1 0 360 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1545
timestamp 1569533753
transform 1 0 488 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1546
timestamp 1569533753
transform 1 0 424 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1547
timestamp 1569533753
transform 1 0 552 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1548
timestamp 1569533753
transform 1 0 296 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1549
timestamp 1569533753
transform 1 0 40 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1550
timestamp 1569533753
transform 1 0 296 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1551
timestamp 1569533753
transform 1 0 40 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1552
timestamp 1569533753
transform 1 0 232 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1553
timestamp 1569533753
transform 1 0 168 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1554
timestamp 1569533753
transform 1 0 232 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1555
timestamp 1569533753
transform 1 0 232 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1556
timestamp 1569533753
transform 1 0 104 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1557
timestamp 1569533753
transform 1 0 296 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1558
timestamp 1569533753
transform 1 0 296 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1559
timestamp 1569533753
transform 1 0 168 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1560
timestamp 1569533753
transform 1 0 296 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1561
timestamp 1569533753
transform 1 0 168 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1562
timestamp 1569533753
transform 1 0 104 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1563
timestamp 1569533753
transform 1 0 168 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1564
timestamp 1569533753
transform 1 0 232 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1565
timestamp 1569533753
transform 1 0 104 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1566
timestamp 1569533753
transform 1 0 360 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1567
timestamp 1569533753
transform 1 0 360 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1568
timestamp 1569533753
transform 1 0 616 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1569
timestamp 1569533753
transform 1 0 552 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1570
timestamp 1569533753
transform 1 0 424 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1571
timestamp 1569533753
transform 1 0 360 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1572
timestamp 1569533753
transform 1 0 616 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1573
timestamp 1569533753
transform 1 0 424 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1574
timestamp 1569533753
transform 1 0 488 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1575
timestamp 1569533753
transform 1 0 552 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1576
timestamp 1569533753
transform 1 0 424 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1577
timestamp 1569533753
transform 1 0 424 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1578
timestamp 1569533753
transform 1 0 488 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1579
timestamp 1569533753
transform 1 0 488 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1580
timestamp 1569533753
transform 1 0 360 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1581
timestamp 1569533753
transform 1 0 552 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1582
timestamp 1569533753
transform 1 0 552 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1583
timestamp 1569533753
transform 1 0 488 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1584
timestamp 1569533753
transform 1 0 616 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1585
timestamp 1569533753
transform 1 0 616 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1586
timestamp 1569533753
transform 1 0 488 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1587
timestamp 1569533753
transform 1 0 552 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1588
timestamp 1569533753
transform 1 0 616 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1589
timestamp 1569533753
transform 1 0 232 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1590
timestamp 1569533753
transform 1 0 296 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1591
timestamp 1569533753
transform 1 0 424 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1592
timestamp 1569533753
transform 1 0 360 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1593
timestamp 1569533753
transform 1 0 552 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1594
timestamp 1569533753
transform 1 0 488 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1595
timestamp 1569533753
transform 1 0 424 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1596
timestamp 1569533753
transform 1 0 552 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1597
timestamp 1569533753
transform 1 0 360 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1598
timestamp 1569533753
transform 1 0 616 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1599
timestamp 1569533753
transform 1 0 488 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1600
timestamp 1569533753
transform 1 0 424 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1601
timestamp 1569533753
transform 1 0 360 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1602
timestamp 1569533753
transform 1 0 488 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1603
timestamp 1569533753
transform 1 0 616 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1604
timestamp 1569533753
transform 1 0 360 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1605
timestamp 1569533753
transform 1 0 616 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1606
timestamp 1569533753
transform 1 0 552 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1607
timestamp 1569533753
transform 1 0 424 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1608
timestamp 1569533753
transform 1 0 488 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1609
timestamp 1569533753
transform 1 0 424 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1610
timestamp 1569533753
transform 1 0 488 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1611
timestamp 1569533753
transform 1 0 552 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1612
timestamp 1569533753
transform 1 0 552 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1613
timestamp 1569533753
transform 1 0 360 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1614
timestamp 1569533753
transform 1 0 360 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1615
timestamp 1569533753
transform 1 0 616 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1616
timestamp 1569533753
transform 1 0 424 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1617
timestamp 1569533753
transform 1 0 616 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1618
timestamp 1569533753
transform 1 0 40 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1619
timestamp 1569533753
transform 1 0 168 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1620
timestamp 1569533753
transform 1 0 296 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1621
timestamp 1569533753
transform 1 0 40 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1622
timestamp 1569533753
transform 1 0 232 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1623
timestamp 1569533753
transform 1 0 296 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1624
timestamp 1569533753
transform 1 0 168 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1625
timestamp 1569533753
transform 1 0 296 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1626
timestamp 1569533753
transform 1 0 104 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1627
timestamp 1569533753
transform 1 0 168 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1628
timestamp 1569533753
transform 1 0 168 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1629
timestamp 1569533753
transform 1 0 40 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1630
timestamp 1569533753
transform 1 0 296 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1631
timestamp 1569533753
transform 1 0 168 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1632
timestamp 1569533753
transform 1 0 104 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1633
timestamp 1569533753
transform 1 0 232 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1634
timestamp 1569533753
transform 1 0 104 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1635
timestamp 1569533753
transform 1 0 232 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1636
timestamp 1569533753
transform 1 0 40 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1637
timestamp 1569533753
transform 1 0 296 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1638
timestamp 1569533753
transform 1 0 232 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1639
timestamp 1569533753
transform 1 0 104 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1640
timestamp 1569533753
transform 1 0 232 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1641
timestamp 1569533753
transform 1 0 40 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1642
timestamp 1569533753
transform 1 0 104 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1643
timestamp 1569533753
transform 1 0 296 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1644
timestamp 1569533753
transform 1 0 40 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1645
timestamp 1569533753
transform 1 0 296 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1646
timestamp 1569533753
transform 1 0 296 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1647
timestamp 1569533753
transform 1 0 40 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1648
timestamp 1569533753
transform 1 0 168 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1649
timestamp 1569533753
transform 1 0 232 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1650
timestamp 1569533753
transform 1 0 40 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1651
timestamp 1569533753
transform 1 0 168 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1652
timestamp 1569533753
transform 1 0 104 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1653
timestamp 1569533753
transform 1 0 40 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1654
timestamp 1569533753
transform 1 0 232 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1655
timestamp 1569533753
transform 1 0 104 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1656
timestamp 1569533753
transform 1 0 168 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1657
timestamp 1569533753
transform 1 0 232 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1658
timestamp 1569533753
transform 1 0 40 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1659
timestamp 1569533753
transform 1 0 104 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1660
timestamp 1569533753
transform 1 0 104 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1661
timestamp 1569533753
transform 1 0 296 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1662
timestamp 1569533753
transform 1 0 104 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1663
timestamp 1569533753
transform 1 0 168 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1664
timestamp 1569533753
transform 1 0 232 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1665
timestamp 1569533753
transform 1 0 168 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1666
timestamp 1569533753
transform 1 0 296 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1667
timestamp 1569533753
transform 1 0 232 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1668
timestamp 1569533753
transform 1 0 424 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1669
timestamp 1569533753
transform 1 0 488 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1670
timestamp 1569533753
transform 1 0 424 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1671
timestamp 1569533753
transform 1 0 424 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1672
timestamp 1569533753
transform 1 0 488 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1673
timestamp 1569533753
transform 1 0 616 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1674
timestamp 1569533753
transform 1 0 424 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1675
timestamp 1569533753
transform 1 0 360 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1676
timestamp 1569533753
transform 1 0 616 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1677
timestamp 1569533753
transform 1 0 552 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1678
timestamp 1569533753
transform 1 0 552 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1679
timestamp 1569533753
transform 1 0 616 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1680
timestamp 1569533753
transform 1 0 552 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1681
timestamp 1569533753
transform 1 0 552 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1682
timestamp 1569533753
transform 1 0 488 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1683
timestamp 1569533753
transform 1 0 360 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1684
timestamp 1569533753
transform 1 0 552 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1685
timestamp 1569533753
transform 1 0 616 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1686
timestamp 1569533753
transform 1 0 488 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1687
timestamp 1569533753
transform 1 0 360 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1688
timestamp 1569533753
transform 1 0 616 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1689
timestamp 1569533753
transform 1 0 360 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1690
timestamp 1569533753
transform 1 0 424 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1691
timestamp 1569533753
transform 1 0 360 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1692
timestamp 1569533753
transform 1 0 488 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1693
timestamp 1569533753
transform 1 0 1192 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1694
timestamp 1569533753
transform 1 0 1192 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1695
timestamp 1569533753
transform 1 0 1256 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1696
timestamp 1569533753
transform 1 0 1128 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1697
timestamp 1569533753
transform 1 0 1064 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1698
timestamp 1569533753
transform 1 0 1128 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1699
timestamp 1569533753
transform 1 0 1192 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1700
timestamp 1569533753
transform 1 0 1128 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1701
timestamp 1569533753
transform 1 0 1192 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1702
timestamp 1569533753
transform 1 0 1128 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1703
timestamp 1569533753
transform 1 0 1256 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1704
timestamp 1569533753
transform 1 0 1064 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1705
timestamp 1569533753
transform 1 0 1000 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1706
timestamp 1569533753
transform 1 0 1256 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1707
timestamp 1569533753
transform 1 0 1000 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1708
timestamp 1569533753
transform 1 0 1256 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1709
timestamp 1569533753
transform 1 0 1000 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1710
timestamp 1569533753
transform 1 0 1256 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1711
timestamp 1569533753
transform 1 0 1128 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1712
timestamp 1569533753
transform 1 0 1000 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1713
timestamp 1569533753
transform 1 0 1064 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1714
timestamp 1569533753
transform 1 0 1064 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1715
timestamp 1569533753
transform 1 0 1192 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1716
timestamp 1569533753
transform 1 0 1064 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1717
timestamp 1569533753
transform 1 0 1000 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1718
timestamp 1569533753
transform 1 0 808 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1719
timestamp 1569533753
transform 1 0 680 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1720
timestamp 1569533753
transform 1 0 872 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1721
timestamp 1569533753
transform 1 0 936 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1722
timestamp 1569533753
transform 1 0 872 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1723
timestamp 1569533753
transform 1 0 936 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1724
timestamp 1569533753
transform 1 0 744 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1725
timestamp 1569533753
transform 1 0 744 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1726
timestamp 1569533753
transform 1 0 744 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1727
timestamp 1569533753
transform 1 0 872 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1728
timestamp 1569533753
transform 1 0 744 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1729
timestamp 1569533753
transform 1 0 744 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1730
timestamp 1569533753
transform 1 0 680 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1731
timestamp 1569533753
transform 1 0 808 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1732
timestamp 1569533753
transform 1 0 808 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1733
timestamp 1569533753
transform 1 0 808 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1734
timestamp 1569533753
transform 1 0 808 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1735
timestamp 1569533753
transform 1 0 872 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1736
timestamp 1569533753
transform 1 0 680 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1737
timestamp 1569533753
transform 1 0 680 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1738
timestamp 1569533753
transform 1 0 936 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1739
timestamp 1569533753
transform 1 0 872 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1740
timestamp 1569533753
transform 1 0 936 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1741
timestamp 1569533753
transform 1 0 680 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1742
timestamp 1569533753
transform 1 0 936 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1743
timestamp 1569533753
transform 1 0 936 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1744
timestamp 1569533753
transform 1 0 936 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1745
timestamp 1569533753
transform 1 0 808 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1746
timestamp 1569533753
transform 1 0 680 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1747
timestamp 1569533753
transform 1 0 680 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1748
timestamp 1569533753
transform 1 0 680 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1749
timestamp 1569533753
transform 1 0 872 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1750
timestamp 1569533753
transform 1 0 680 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1751
timestamp 1569533753
transform 1 0 808 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1752
timestamp 1569533753
transform 1 0 744 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1753
timestamp 1569533753
transform 1 0 872 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1754
timestamp 1569533753
transform 1 0 808 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1755
timestamp 1569533753
transform 1 0 872 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1756
timestamp 1569533753
transform 1 0 872 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1757
timestamp 1569533753
transform 1 0 872 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1758
timestamp 1569533753
transform 1 0 936 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1759
timestamp 1569533753
transform 1 0 744 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1760
timestamp 1569533753
transform 1 0 744 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1761
timestamp 1569533753
transform 1 0 936 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1762
timestamp 1569533753
transform 1 0 744 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1763
timestamp 1569533753
transform 1 0 936 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1764
timestamp 1569533753
transform 1 0 808 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1765
timestamp 1569533753
transform 1 0 680 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1766
timestamp 1569533753
transform 1 0 744 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1767
timestamp 1569533753
transform 1 0 808 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1768
timestamp 1569533753
transform 1 0 1064 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1769
timestamp 1569533753
transform 1 0 1064 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1770
timestamp 1569533753
transform 1 0 1128 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1771
timestamp 1569533753
transform 1 0 1000 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1772
timestamp 1569533753
transform 1 0 1192 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1773
timestamp 1569533753
transform 1 0 1192 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1774
timestamp 1569533753
transform 1 0 1192 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1775
timestamp 1569533753
transform 1 0 1192 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1776
timestamp 1569533753
transform 1 0 1192 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1777
timestamp 1569533753
transform 1 0 1064 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1778
timestamp 1569533753
transform 1 0 1000 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1779
timestamp 1569533753
transform 1 0 1064 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1780
timestamp 1569533753
transform 1 0 1000 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1781
timestamp 1569533753
transform 1 0 1064 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1782
timestamp 1569533753
transform 1 0 1128 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1783
timestamp 1569533753
transform 1 0 1000 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1784
timestamp 1569533753
transform 1 0 1128 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1785
timestamp 1569533753
transform 1 0 1000 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1786
timestamp 1569533753
transform 1 0 1256 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1787
timestamp 1569533753
transform 1 0 1256 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1788
timestamp 1569533753
transform 1 0 1256 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_1789
timestamp 1569533753
transform 1 0 1128 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_1790
timestamp 1569533753
transform 1 0 1256 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_1791
timestamp 1569533753
transform 1 0 1256 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_1792
timestamp 1569533753
transform 1 0 1128 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_1793
timestamp 1569533753
transform 1 0 2280 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1794
timestamp 1569533753
transform 1 0 2280 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1795
timestamp 1569533753
transform 1 0 2472 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1796
timestamp 1569533753
transform 1 0 2344 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1797
timestamp 1569533753
transform 1 0 2216 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1798
timestamp 1569533753
transform 1 0 2472 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1799
timestamp 1569533753
transform 1 0 2344 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1800
timestamp 1569533753
transform 1 0 2216 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1801
timestamp 1569533753
transform 1 0 2408 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1802
timestamp 1569533753
transform 1 0 2408 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1803
timestamp 1569533753
transform 1 0 2408 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1804
timestamp 1569533753
transform 1 0 2344 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1805
timestamp 1569533753
transform 1 0 2344 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1806
timestamp 1569533753
transform 1 0 2408 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1807
timestamp 1569533753
transform 1 0 2216 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1808
timestamp 1569533753
transform 1 0 2280 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1809
timestamp 1569533753
transform 1 0 2472 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1810
timestamp 1569533753
transform 1 0 2216 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1811
timestamp 1569533753
transform 1 0 2472 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1812
timestamp 1569533753
transform 1 0 2280 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1813
timestamp 1569533753
transform 1 0 2024 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1814
timestamp 1569533753
transform 1 0 1896 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1815
timestamp 1569533753
transform 1 0 2024 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1816
timestamp 1569533753
transform 1 0 2088 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1817
timestamp 1569533753
transform 1 0 2088 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1818
timestamp 1569533753
transform 1 0 2024 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1819
timestamp 1569533753
transform 1 0 2088 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1820
timestamp 1569533753
transform 1 0 2152 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1821
timestamp 1569533753
transform 1 0 1896 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1822
timestamp 1569533753
transform 1 0 1896 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1823
timestamp 1569533753
transform 1 0 2152 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1824
timestamp 1569533753
transform 1 0 1896 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1825
timestamp 1569533753
transform 1 0 1960 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1826
timestamp 1569533753
transform 1 0 1960 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1827
timestamp 1569533753
transform 1 0 1960 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1828
timestamp 1569533753
transform 1 0 2152 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1829
timestamp 1569533753
transform 1 0 1960 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1830
timestamp 1569533753
transform 1 0 2088 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1831
timestamp 1569533753
transform 1 0 2024 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1832
timestamp 1569533753
transform 1 0 2152 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1833
timestamp 1569533753
transform 1 0 1896 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1834
timestamp 1569533753
transform 1 0 2024 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1835
timestamp 1569533753
transform 1 0 2088 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1836
timestamp 1569533753
transform 1 0 2024 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1837
timestamp 1569533753
transform 1 0 2152 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1838
timestamp 1569533753
transform 1 0 2152 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1839
timestamp 1569533753
transform 1 0 1896 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1840
timestamp 1569533753
transform 1 0 1960 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1841
timestamp 1569533753
transform 1 0 1960 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1842
timestamp 1569533753
transform 1 0 1960 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1843
timestamp 1569533753
transform 1 0 2024 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1844
timestamp 1569533753
transform 1 0 2024 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1845
timestamp 1569533753
transform 1 0 1896 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1846
timestamp 1569533753
transform 1 0 2088 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1847
timestamp 1569533753
transform 1 0 2088 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1848
timestamp 1569533753
transform 1 0 1960 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1849
timestamp 1569533753
transform 1 0 2152 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1850
timestamp 1569533753
transform 1 0 2152 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1851
timestamp 1569533753
transform 1 0 2088 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1852
timestamp 1569533753
transform 1 0 1896 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1853
timestamp 1569533753
transform 1 0 2344 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1854
timestamp 1569533753
transform 1 0 2280 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1855
timestamp 1569533753
transform 1 0 2344 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1856
timestamp 1569533753
transform 1 0 2408 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1857
timestamp 1569533753
transform 1 0 2408 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1858
timestamp 1569533753
transform 1 0 2472 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1859
timestamp 1569533753
transform 1 0 2472 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1860
timestamp 1569533753
transform 1 0 2344 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1861
timestamp 1569533753
transform 1 0 2344 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1862
timestamp 1569533753
transform 1 0 2408 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1863
timestamp 1569533753
transform 1 0 2408 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1864
timestamp 1569533753
transform 1 0 2280 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1865
timestamp 1569533753
transform 1 0 2472 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1866
timestamp 1569533753
transform 1 0 2472 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1867
timestamp 1569533753
transform 1 0 2216 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1868
timestamp 1569533753
transform 1 0 2280 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1869
timestamp 1569533753
transform 1 0 2280 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1870
timestamp 1569533753
transform 1 0 2216 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1871
timestamp 1569533753
transform 1 0 2216 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1872
timestamp 1569533753
transform 1 0 2216 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1873
timestamp 1569533753
transform 1 0 1896 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1874
timestamp 1569533753
transform 1 0 2344 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1875
timestamp 1569533753
transform 1 0 2408 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1876
timestamp 1569533753
transform 1 0 1960 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1877
timestamp 1569533753
transform 1 0 2472 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1878
timestamp 1569533753
transform 1 0 2024 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1879
timestamp 1569533753
transform 1 0 2088 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1880
timestamp 1569533753
transform 1 0 2152 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1881
timestamp 1569533753
transform 1 0 2216 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1882
timestamp 1569533753
transform 1 0 2280 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1883
timestamp 1569533753
transform 1 0 1768 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1884
timestamp 1569533753
transform 1 0 1768 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1885
timestamp 1569533753
transform 1 0 1832 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1886
timestamp 1569533753
transform 1 0 1704 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1887
timestamp 1569533753
transform 1 0 1768 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1888
timestamp 1569533753
transform 1 0 1832 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1889
timestamp 1569533753
transform 1 0 1640 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1890
timestamp 1569533753
transform 1 0 1640 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1891
timestamp 1569533753
transform 1 0 1640 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1892
timestamp 1569533753
transform 1 0 1704 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1893
timestamp 1569533753
transform 1 0 1704 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1894
timestamp 1569533753
transform 1 0 1704 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1895
timestamp 1569533753
transform 1 0 1832 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1896
timestamp 1569533753
transform 1 0 1640 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1897
timestamp 1569533753
transform 1 0 1832 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1898
timestamp 1569533753
transform 1 0 1768 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1899
timestamp 1569533753
transform 1 0 1512 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1900
timestamp 1569533753
transform 1 0 1512 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1901
timestamp 1569533753
transform 1 0 1320 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1902
timestamp 1569533753
transform 1 0 1320 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1903
timestamp 1569533753
transform 1 0 1384 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1904
timestamp 1569533753
transform 1 0 1384 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1905
timestamp 1569533753
transform 1 0 1448 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1906
timestamp 1569533753
transform 1 0 1448 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1907
timestamp 1569533753
transform 1 0 1512 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1908
timestamp 1569533753
transform 1 0 1320 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1909
timestamp 1569533753
transform 1 0 1320 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1910
timestamp 1569533753
transform 1 0 1512 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1911
timestamp 1569533753
transform 1 0 1448 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1912
timestamp 1569533753
transform 1 0 1384 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1913
timestamp 1569533753
transform 1 0 1448 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1914
timestamp 1569533753
transform 1 0 1384 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1915
timestamp 1569533753
transform 1 0 1384 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1916
timestamp 1569533753
transform 1 0 1448 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1917
timestamp 1569533753
transform 1 0 1448 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1918
timestamp 1569533753
transform 1 0 1512 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1919
timestamp 1569533753
transform 1 0 1320 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1920
timestamp 1569533753
transform 1 0 1448 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1921
timestamp 1569533753
transform 1 0 1448 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1922
timestamp 1569533753
transform 1 0 1384 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1923
timestamp 1569533753
transform 1 0 1512 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1924
timestamp 1569533753
transform 1 0 1512 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1925
timestamp 1569533753
transform 1 0 1384 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1926
timestamp 1569533753
transform 1 0 1320 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1927
timestamp 1569533753
transform 1 0 1320 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1928
timestamp 1569533753
transform 1 0 1384 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1929
timestamp 1569533753
transform 1 0 1320 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1930
timestamp 1569533753
transform 1 0 1512 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1931
timestamp 1569533753
transform 1 0 1704 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1932
timestamp 1569533753
transform 1 0 1768 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1933
timestamp 1569533753
transform 1 0 1832 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1934
timestamp 1569533753
transform 1 0 1704 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1935
timestamp 1569533753
transform 1 0 1704 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1936
timestamp 1569533753
transform 1 0 1768 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1937
timestamp 1569533753
transform 1 0 1768 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1938
timestamp 1569533753
transform 1 0 1832 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1939
timestamp 1569533753
transform 1 0 1832 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1940
timestamp 1569533753
transform 1 0 1640 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1941
timestamp 1569533753
transform 1 0 1640 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1942
timestamp 1569533753
transform 1 0 1832 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1943
timestamp 1569533753
transform 1 0 1640 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1944
timestamp 1569533753
transform 1 0 1640 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1945
timestamp 1569533753
transform 1 0 1704 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1946
timestamp 1569533753
transform 1 0 1768 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1947
timestamp 1569533753
transform 1 0 1576 0 1 1320
box -8 -8 8 8
use VIA2$3  VIA2$3_1948
timestamp 1569533753
transform 1 0 1576 0 1 1448
box -8 -8 8 8
use VIA2$3  VIA2$3_1949
timestamp 1569533753
transform 1 0 1320 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1950
timestamp 1569533753
transform 1 0 1640 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1951
timestamp 1569533753
transform 1 0 1448 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1952
timestamp 1569533753
transform 1 0 1704 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1953
timestamp 1569533753
transform 1 0 1576 0 1 1640
box -8 -8 8 8
use VIA2$3  VIA2$3_1954
timestamp 1569533753
transform 1 0 1576 0 1 1768
box -8 -8 8 8
use VIA2$3  VIA2$3_1955
timestamp 1569533753
transform 1 0 1768 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1956
timestamp 1569533753
transform 1 0 1512 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1957
timestamp 1569533753
transform 1 0 1832 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1958
timestamp 1569533753
transform 1 0 1384 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1959
timestamp 1569533753
transform 1 0 1576 0 1 1576
box -8 -8 8 8
use VIA2$3  VIA2$3_1960
timestamp 1569533753
transform 1 0 1576 0 1 1832
box -8 -8 8 8
use VIA2$3  VIA2$3_1961
timestamp 1569533753
transform 1 0 1576 0 1 1384
box -8 -8 8 8
use VIA2$3  VIA2$3_1962
timestamp 1569533753
transform 1 0 1576 0 1 1512
box -8 -8 8 8
use VIA2$3  VIA2$3_1963
timestamp 1569533753
transform 1 0 1576 0 1 1704
box -8 -8 8 8
use VIA2$3  VIA2$3_1964
timestamp 1569533753
transform 1 0 1704 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1965
timestamp 1569533753
transform 1 0 1768 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1966
timestamp 1569533753
transform 1 0 1704 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1967
timestamp 1569533753
transform 1 0 1832 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1968
timestamp 1569533753
transform 1 0 1768 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1969
timestamp 1569533753
transform 1 0 1768 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1970
timestamp 1569533753
transform 1 0 1768 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1971
timestamp 1569533753
transform 1 0 1640 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1972
timestamp 1569533753
transform 1 0 1640 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1973
timestamp 1569533753
transform 1 0 1704 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1974
timestamp 1569533753
transform 1 0 1768 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1975
timestamp 1569533753
transform 1 0 1832 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1976
timestamp 1569533753
transform 1 0 1640 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1977
timestamp 1569533753
transform 1 0 1832 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1978
timestamp 1569533753
transform 1 0 1832 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1979
timestamp 1569533753
transform 1 0 1832 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1980
timestamp 1569533753
transform 1 0 1640 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1981
timestamp 1569533753
transform 1 0 1640 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1982
timestamp 1569533753
transform 1 0 1704 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1983
timestamp 1569533753
transform 1 0 1704 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1984
timestamp 1569533753
transform 1 0 1384 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1985
timestamp 1569533753
transform 1 0 1512 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1986
timestamp 1569533753
transform 1 0 1448 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1987
timestamp 1569533753
transform 1 0 1512 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1988
timestamp 1569533753
transform 1 0 1512 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1989
timestamp 1569533753
transform 1 0 1512 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1990
timestamp 1569533753
transform 1 0 1320 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_1991
timestamp 1569533753
transform 1 0 1320 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1992
timestamp 1569533753
transform 1 0 1384 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1993
timestamp 1569533753
transform 1 0 1320 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1994
timestamp 1569533753
transform 1 0 1384 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_1995
timestamp 1569533753
transform 1 0 1320 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_1996
timestamp 1569533753
transform 1 0 1512 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1997
timestamp 1569533753
transform 1 0 1448 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_1998
timestamp 1569533753
transform 1 0 1448 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_1999
timestamp 1569533753
transform 1 0 1448 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2000
timestamp 1569533753
transform 1 0 1448 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2001
timestamp 1569533753
transform 1 0 1320 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2002
timestamp 1569533753
transform 1 0 1384 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2003
timestamp 1569533753
transform 1 0 1384 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2004
timestamp 1569533753
transform 1 0 1384 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2005
timestamp 1569533753
transform 1 0 1320 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2006
timestamp 1569533753
transform 1 0 1512 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2007
timestamp 1569533753
transform 1 0 1384 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2008
timestamp 1569533753
transform 1 0 1320 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2009
timestamp 1569533753
transform 1 0 1512 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2010
timestamp 1569533753
transform 1 0 1320 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2011
timestamp 1569533753
transform 1 0 1384 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2012
timestamp 1569533753
transform 1 0 1320 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2013
timestamp 1569533753
transform 1 0 1448 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2014
timestamp 1569533753
transform 1 0 1384 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2015
timestamp 1569533753
transform 1 0 1448 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2016
timestamp 1569533753
transform 1 0 1384 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2017
timestamp 1569533753
transform 1 0 1448 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2018
timestamp 1569533753
transform 1 0 1320 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2019
timestamp 1569533753
transform 1 0 1512 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2020
timestamp 1569533753
transform 1 0 1448 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2021
timestamp 1569533753
transform 1 0 1512 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2022
timestamp 1569533753
transform 1 0 1448 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2023
timestamp 1569533753
transform 1 0 1512 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2024
timestamp 1569533753
transform 1 0 1704 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2025
timestamp 1569533753
transform 1 0 1704 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2026
timestamp 1569533753
transform 1 0 1768 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2027
timestamp 1569533753
transform 1 0 1768 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2028
timestamp 1569533753
transform 1 0 1704 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2029
timestamp 1569533753
transform 1 0 1768 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2030
timestamp 1569533753
transform 1 0 1832 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2031
timestamp 1569533753
transform 1 0 1832 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2032
timestamp 1569533753
transform 1 0 1832 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2033
timestamp 1569533753
transform 1 0 1832 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2034
timestamp 1569533753
transform 1 0 1832 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2035
timestamp 1569533753
transform 1 0 1704 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2036
timestamp 1569533753
transform 1 0 1704 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2037
timestamp 1569533753
transform 1 0 1768 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2038
timestamp 1569533753
transform 1 0 1768 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2039
timestamp 1569533753
transform 1 0 1640 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2040
timestamp 1569533753
transform 1 0 1640 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2041
timestamp 1569533753
transform 1 0 1640 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2042
timestamp 1569533753
transform 1 0 1640 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2043
timestamp 1569533753
transform 1 0 1640 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2044
timestamp 1569533753
transform 1 0 1576 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2045
timestamp 1569533753
transform 1 0 1576 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2046
timestamp 1569533753
transform 1 0 1576 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2047
timestamp 1569533753
transform 1 0 1576 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2048
timestamp 1569533753
transform 1 0 1576 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2049
timestamp 1569533753
transform 1 0 1576 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2050
timestamp 1569533753
transform 1 0 1576 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2051
timestamp 1569533753
transform 1 0 1576 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2052
timestamp 1569533753
transform 1 0 1576 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2053
timestamp 1569533753
transform 1 0 1576 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2054
timestamp 1569533753
transform 1 0 2344 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2055
timestamp 1569533753
transform 1 0 2408 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2056
timestamp 1569533753
transform 1 0 2472 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2057
timestamp 1569533753
transform 1 0 2408 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2058
timestamp 1569533753
transform 1 0 2280 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2059
timestamp 1569533753
transform 1 0 2280 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2060
timestamp 1569533753
transform 1 0 2280 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2061
timestamp 1569533753
transform 1 0 2344 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2062
timestamp 1569533753
transform 1 0 2344 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2063
timestamp 1569533753
transform 1 0 2216 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2064
timestamp 1569533753
transform 1 0 2344 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2065
timestamp 1569533753
transform 1 0 2280 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2066
timestamp 1569533753
transform 1 0 2280 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2067
timestamp 1569533753
transform 1 0 2216 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2068
timestamp 1569533753
transform 1 0 2216 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2069
timestamp 1569533753
transform 1 0 2216 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2070
timestamp 1569533753
transform 1 0 2408 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2071
timestamp 1569533753
transform 1 0 2472 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2072
timestamp 1569533753
transform 1 0 2216 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2073
timestamp 1569533753
transform 1 0 1896 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2074
timestamp 1569533753
transform 1 0 2024 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2075
timestamp 1569533753
transform 1 0 2024 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2076
timestamp 1569533753
transform 1 0 2024 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2077
timestamp 1569533753
transform 1 0 1960 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2078
timestamp 1569533753
transform 1 0 2088 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2079
timestamp 1569533753
transform 1 0 2088 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2080
timestamp 1569533753
transform 1 0 2088 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2081
timestamp 1569533753
transform 1 0 1896 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2082
timestamp 1569533753
transform 1 0 1960 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2083
timestamp 1569533753
transform 1 0 2152 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2084
timestamp 1569533753
transform 1 0 2024 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2085
timestamp 1569533753
transform 1 0 2088 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2086
timestamp 1569533753
transform 1 0 2024 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2087
timestamp 1569533753
transform 1 0 1960 0 1 2152
box -8 -8 8 8
use VIA2$3  VIA2$3_2088
timestamp 1569533753
transform 1 0 2088 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2089
timestamp 1569533753
transform 1 0 2152 0 1 1896
box -8 -8 8 8
use VIA2$3  VIA2$3_2090
timestamp 1569533753
transform 1 0 1896 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2091
timestamp 1569533753
transform 1 0 2152 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2092
timestamp 1569533753
transform 1 0 1896 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2093
timestamp 1569533753
transform 1 0 2152 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2094
timestamp 1569533753
transform 1 0 1896 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2095
timestamp 1569533753
transform 1 0 2152 0 1 2088
box -8 -8 8 8
use VIA2$3  VIA2$3_2096
timestamp 1569533753
transform 1 0 1960 0 1 1960
box -8 -8 8 8
use VIA2$3  VIA2$3_2097
timestamp 1569533753
transform 1 0 1960 0 1 2024
box -8 -8 8 8
use VIA2$3  VIA2$3_2098
timestamp 1569533753
transform 1 0 1896 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2099
timestamp 1569533753
transform 1 0 1896 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2100
timestamp 1569533753
transform 1 0 1896 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2101
timestamp 1569533753
transform 1 0 1896 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2102
timestamp 1569533753
transform 1 0 1896 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2103
timestamp 1569533753
transform 1 0 1960 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2104
timestamp 1569533753
transform 1 0 1960 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2105
timestamp 1569533753
transform 1 0 1960 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2106
timestamp 1569533753
transform 1 0 1960 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2107
timestamp 1569533753
transform 1 0 1960 0 1 2472
box -8 -8 8 8
use VIA2$3  VIA2$3_2108
timestamp 1569533753
transform 1 0 2152 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2109
timestamp 1569533753
transform 1 0 2152 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2110
timestamp 1569533753
transform 1 0 2024 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2111
timestamp 1569533753
transform 1 0 2024 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2112
timestamp 1569533753
transform 1 0 2024 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2113
timestamp 1569533753
transform 1 0 2024 0 1 2408
box -8 -8 8 8
use VIA2$3  VIA2$3_2114
timestamp 1569533753
transform 1 0 2088 0 1 2344
box -8 -8 8 8
use VIA2$3  VIA2$3_2115
timestamp 1569533753
transform 1 0 2088 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2116
timestamp 1569533753
transform 1 0 2088 0 1 2280
box -8 -8 8 8
use VIA2$3  VIA2$3_2117
timestamp 1569533753
transform 1 0 2216 0 1 2216
box -8 -8 8 8
use VIA2$3  VIA2$3_2118
timestamp 1569533753
transform 1 0 1896 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2119
timestamp 1569533753
transform 1 0 1640 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2120
timestamp 1569533753
transform 1 0 1768 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2121
timestamp 1569533753
transform 1 0 1704 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2122
timestamp 1569533753
transform 1 0 1768 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2123
timestamp 1569533753
transform 1 0 1832 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2124
timestamp 1569533753
transform 1 0 1704 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2125
timestamp 1569533753
transform 1 0 1640 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2126
timestamp 1569533753
transform 1 0 1704 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2127
timestamp 1569533753
transform 1 0 1768 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2128
timestamp 1569533753
transform 1 0 1640 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2129
timestamp 1569533753
transform 1 0 1640 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2130
timestamp 1569533753
transform 1 0 1704 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2131
timestamp 1569533753
transform 1 0 1832 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2132
timestamp 1569533753
transform 1 0 1640 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2133
timestamp 1569533753
transform 1 0 1384 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2134
timestamp 1569533753
transform 1 0 1448 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2135
timestamp 1569533753
transform 1 0 1512 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2136
timestamp 1569533753
transform 1 0 1512 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2137
timestamp 1569533753
transform 1 0 1448 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2138
timestamp 1569533753
transform 1 0 1384 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2139
timestamp 1569533753
transform 1 0 1320 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2140
timestamp 1569533753
transform 1 0 1448 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2141
timestamp 1569533753
transform 1 0 1320 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2142
timestamp 1569533753
transform 1 0 1448 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2143
timestamp 1569533753
transform 1 0 1320 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2144
timestamp 1569533753
transform 1 0 1384 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2145
timestamp 1569533753
transform 1 0 1512 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2146
timestamp 1569533753
transform 1 0 1512 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2147
timestamp 1569533753
transform 1 0 1448 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2148
timestamp 1569533753
transform 1 0 1384 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2149
timestamp 1569533753
transform 1 0 1384 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2150
timestamp 1569533753
transform 1 0 1320 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2151
timestamp 1569533753
transform 1 0 1320 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2152
timestamp 1569533753
transform 1 0 1512 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2153
timestamp 1569533753
transform 1 0 1512 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2154
timestamp 1569533753
transform 1 0 1448 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2155
timestamp 1569533753
transform 1 0 1384 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2156
timestamp 1569533753
transform 1 0 1512 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2157
timestamp 1569533753
transform 1 0 1512 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2158
timestamp 1569533753
transform 1 0 1384 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2159
timestamp 1569533753
transform 1 0 1384 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2160
timestamp 1569533753
transform 1 0 1448 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2161
timestamp 1569533753
transform 1 0 1512 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2162
timestamp 1569533753
transform 1 0 1512 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2163
timestamp 1569533753
transform 1 0 1384 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2164
timestamp 1569533753
transform 1 0 1320 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2165
timestamp 1569533753
transform 1 0 1320 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2166
timestamp 1569533753
transform 1 0 1384 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2167
timestamp 1569533753
transform 1 0 1448 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2168
timestamp 1569533753
transform 1 0 1448 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2169
timestamp 1569533753
transform 1 0 1448 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2170
timestamp 1569533753
transform 1 0 1320 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2171
timestamp 1569533753
transform 1 0 1320 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2172
timestamp 1569533753
transform 1 0 1320 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2173
timestamp 1569533753
transform 1 0 1576 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2174
timestamp 1569533753
transform 1 0 1576 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2175
timestamp 1569533753
transform 1 0 1576 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2176
timestamp 1569533753
transform 1 0 1576 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2177
timestamp 1569533753
transform 1 0 1576 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2178
timestamp 1569533753
transform 1 0 1576 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2179
timestamp 1569533753
transform 1 0 1320 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2180
timestamp 1569533753
transform 1 0 1384 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2181
timestamp 1569533753
transform 1 0 1320 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2182
timestamp 1569533753
transform 1 0 1512 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2183
timestamp 1569533753
transform 1 0 1384 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2184
timestamp 1569533753
transform 1 0 1320 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2185
timestamp 1569533753
transform 1 0 1512 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2186
timestamp 1569533753
transform 1 0 1384 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2187
timestamp 1569533753
transform 1 0 1320 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2188
timestamp 1569533753
transform 1 0 1512 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2189
timestamp 1569533753
transform 1 0 1448 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2190
timestamp 1569533753
transform 1 0 1512 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2191
timestamp 1569533753
transform 1 0 1384 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2192
timestamp 1569533753
transform 1 0 1320 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2193
timestamp 1569533753
transform 1 0 1448 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2194
timestamp 1569533753
transform 1 0 1384 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2195
timestamp 1569533753
transform 1 0 1320 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2196
timestamp 1569533753
transform 1 0 1384 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2197
timestamp 1569533753
transform 1 0 1384 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2198
timestamp 1569533753
transform 1 0 1384 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2199
timestamp 1569533753
transform 1 0 1320 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2200
timestamp 1569533753
transform 1 0 1512 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2201
timestamp 1569533753
transform 1 0 1448 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2202
timestamp 1569533753
transform 1 0 1512 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2203
timestamp 1569533753
transform 1 0 1320 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2204
timestamp 1569533753
transform 1 0 1384 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2205
timestamp 1569533753
transform 1 0 1448 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2206
timestamp 1569533753
transform 1 0 1448 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2207
timestamp 1569533753
transform 1 0 1512 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2208
timestamp 1569533753
transform 1 0 1512 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2209
timestamp 1569533753
transform 1 0 1448 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2210
timestamp 1569533753
transform 1 0 1320 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2211
timestamp 1569533753
transform 1 0 1512 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2212
timestamp 1569533753
transform 1 0 1448 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2213
timestamp 1569533753
transform 1 0 1448 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2214
timestamp 1569533753
transform 1 0 1448 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2215
timestamp 1569533753
transform 1 0 2472 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2216
timestamp 1569533753
transform 1 0 2344 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2217
timestamp 1569533753
transform 1 0 2344 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2218
timestamp 1569533753
transform 1 0 2472 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2219
timestamp 1569533753
transform 1 0 2472 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2220
timestamp 1569533753
transform 1 0 2472 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2221
timestamp 1569533753
transform 1 0 2472 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2222
timestamp 1569533753
transform 1 0 2344 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2223
timestamp 1569533753
transform 1 0 2408 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2224
timestamp 1569533753
transform 1 0 2472 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2225
timestamp 1569533753
transform 1 0 2408 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2226
timestamp 1569533753
transform 1 0 2472 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2227
timestamp 1569533753
transform 1 0 2408 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2228
timestamp 1569533753
transform 1 0 2344 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2229
timestamp 1569533753
transform 1 0 2408 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2230
timestamp 1569533753
transform 1 0 2408 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2231
timestamp 1569533753
transform 1 0 2408 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2232
timestamp 1569533753
transform 1 0 2344 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2233
timestamp 1569533753
transform 1 0 2408 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2234
timestamp 1569533753
transform 1 0 2344 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2235
timestamp 1569533753
transform 1 0 2472 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2236
timestamp 1569533753
transform 1 0 1256 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2237
timestamp 1569533753
transform 1 0 1064 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2238
timestamp 1569533753
transform 1 0 1000 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2239
timestamp 1569533753
transform 1 0 1256 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2240
timestamp 1569533753
transform 1 0 1000 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2241
timestamp 1569533753
transform 1 0 1128 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2242
timestamp 1569533753
transform 1 0 1064 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2243
timestamp 1569533753
transform 1 0 1192 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2244
timestamp 1569533753
transform 1 0 1064 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2245
timestamp 1569533753
transform 1 0 1192 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2246
timestamp 1569533753
transform 1 0 1256 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2247
timestamp 1569533753
transform 1 0 1064 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2248
timestamp 1569533753
transform 1 0 1000 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2249
timestamp 1569533753
transform 1 0 1128 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2250
timestamp 1569533753
transform 1 0 1000 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2251
timestamp 1569533753
transform 1 0 1192 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2252
timestamp 1569533753
transform 1 0 1128 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2253
timestamp 1569533753
transform 1 0 1256 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2254
timestamp 1569533753
transform 1 0 1192 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2255
timestamp 1569533753
transform 1 0 1256 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2256
timestamp 1569533753
transform 1 0 1064 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2257
timestamp 1569533753
transform 1 0 1128 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2258
timestamp 1569533753
transform 1 0 1128 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2259
timestamp 1569533753
transform 1 0 1192 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2260
timestamp 1569533753
transform 1 0 1000 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2261
timestamp 1569533753
transform 1 0 680 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2262
timestamp 1569533753
transform 1 0 936 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2263
timestamp 1569533753
transform 1 0 808 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2264
timestamp 1569533753
transform 1 0 680 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2265
timestamp 1569533753
transform 1 0 744 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2266
timestamp 1569533753
transform 1 0 744 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2267
timestamp 1569533753
transform 1 0 744 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2268
timestamp 1569533753
transform 1 0 936 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2269
timestamp 1569533753
transform 1 0 680 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2270
timestamp 1569533753
transform 1 0 808 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2271
timestamp 1569533753
transform 1 0 808 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2272
timestamp 1569533753
transform 1 0 808 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2273
timestamp 1569533753
transform 1 0 872 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2274
timestamp 1569533753
transform 1 0 872 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2275
timestamp 1569533753
transform 1 0 936 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2276
timestamp 1569533753
transform 1 0 872 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2277
timestamp 1569533753
transform 1 0 936 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2278
timestamp 1569533753
transform 1 0 680 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2279
timestamp 1569533753
transform 1 0 808 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2280
timestamp 1569533753
transform 1 0 744 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2281
timestamp 1569533753
transform 1 0 680 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2282
timestamp 1569533753
transform 1 0 872 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2283
timestamp 1569533753
transform 1 0 936 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2284
timestamp 1569533753
transform 1 0 744 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2285
timestamp 1569533753
transform 1 0 872 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2286
timestamp 1569533753
transform 1 0 936 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2287
timestamp 1569533753
transform 1 0 808 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2288
timestamp 1569533753
transform 1 0 872 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2289
timestamp 1569533753
transform 1 0 680 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2290
timestamp 1569533753
transform 1 0 872 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2291
timestamp 1569533753
transform 1 0 680 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2292
timestamp 1569533753
transform 1 0 744 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2293
timestamp 1569533753
transform 1 0 744 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2294
timestamp 1569533753
transform 1 0 808 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2295
timestamp 1569533753
transform 1 0 808 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2296
timestamp 1569533753
transform 1 0 936 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2297
timestamp 1569533753
transform 1 0 872 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2298
timestamp 1569533753
transform 1 0 936 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2299
timestamp 1569533753
transform 1 0 808 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2300
timestamp 1569533753
transform 1 0 744 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2301
timestamp 1569533753
transform 1 0 744 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2302
timestamp 1569533753
transform 1 0 808 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2303
timestamp 1569533753
transform 1 0 936 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2304
timestamp 1569533753
transform 1 0 680 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2305
timestamp 1569533753
transform 1 0 680 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2306
timestamp 1569533753
transform 1 0 936 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2307
timestamp 1569533753
transform 1 0 872 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2308
timestamp 1569533753
transform 1 0 744 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2309
timestamp 1569533753
transform 1 0 872 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2310
timestamp 1569533753
transform 1 0 680 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2311
timestamp 1569533753
transform 1 0 1000 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2312
timestamp 1569533753
transform 1 0 1128 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2313
timestamp 1569533753
transform 1 0 1192 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2314
timestamp 1569533753
transform 1 0 1000 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2315
timestamp 1569533753
transform 1 0 1000 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2316
timestamp 1569533753
transform 1 0 1064 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2317
timestamp 1569533753
transform 1 0 1256 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2318
timestamp 1569533753
transform 1 0 1256 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2319
timestamp 1569533753
transform 1 0 1128 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2320
timestamp 1569533753
transform 1 0 1256 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2321
timestamp 1569533753
transform 1 0 1000 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2322
timestamp 1569533753
transform 1 0 1256 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2323
timestamp 1569533753
transform 1 0 1000 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2324
timestamp 1569533753
transform 1 0 1064 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2325
timestamp 1569533753
transform 1 0 1192 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2326
timestamp 1569533753
transform 1 0 1192 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2327
timestamp 1569533753
transform 1 0 1128 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2328
timestamp 1569533753
transform 1 0 1064 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2329
timestamp 1569533753
transform 1 0 1128 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2330
timestamp 1569533753
transform 1 0 1192 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2331
timestamp 1569533753
transform 1 0 1192 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2332
timestamp 1569533753
transform 1 0 1064 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2333
timestamp 1569533753
transform 1 0 1064 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2334
timestamp 1569533753
transform 1 0 1256 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2335
timestamp 1569533753
transform 1 0 1128 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2336
timestamp 1569533753
transform 1 0 488 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2337
timestamp 1569533753
transform 1 0 616 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2338
timestamp 1569533753
transform 1 0 552 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2339
timestamp 1569533753
transform 1 0 616 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2340
timestamp 1569533753
transform 1 0 616 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2341
timestamp 1569533753
transform 1 0 552 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2342
timestamp 1569533753
transform 1 0 488 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2343
timestamp 1569533753
transform 1 0 616 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2344
timestamp 1569533753
transform 1 0 552 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2345
timestamp 1569533753
transform 1 0 552 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2346
timestamp 1569533753
transform 1 0 488 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2347
timestamp 1569533753
transform 1 0 360 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2348
timestamp 1569533753
transform 1 0 424 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2349
timestamp 1569533753
transform 1 0 360 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2350
timestamp 1569533753
transform 1 0 488 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2351
timestamp 1569533753
transform 1 0 552 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2352
timestamp 1569533753
transform 1 0 424 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2353
timestamp 1569533753
transform 1 0 424 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2354
timestamp 1569533753
transform 1 0 360 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2355
timestamp 1569533753
transform 1 0 488 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2356
timestamp 1569533753
transform 1 0 424 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2357
timestamp 1569533753
transform 1 0 360 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2358
timestamp 1569533753
transform 1 0 616 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2359
timestamp 1569533753
transform 1 0 424 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2360
timestamp 1569533753
transform 1 0 360 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2361
timestamp 1569533753
transform 1 0 232 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2362
timestamp 1569533753
transform 1 0 232 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2363
timestamp 1569533753
transform 1 0 296 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2364
timestamp 1569533753
transform 1 0 296 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2365
timestamp 1569533753
transform 1 0 104 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2366
timestamp 1569533753
transform 1 0 232 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2367
timestamp 1569533753
transform 1 0 168 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2368
timestamp 1569533753
transform 1 0 104 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2369
timestamp 1569533753
transform 1 0 296 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2370
timestamp 1569533753
transform 1 0 104 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2371
timestamp 1569533753
transform 1 0 40 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2372
timestamp 1569533753
transform 1 0 232 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2373
timestamp 1569533753
transform 1 0 40 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2374
timestamp 1569533753
transform 1 0 104 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2375
timestamp 1569533753
transform 1 0 168 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2376
timestamp 1569533753
transform 1 0 168 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2377
timestamp 1569533753
transform 1 0 40 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2378
timestamp 1569533753
transform 1 0 296 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2379
timestamp 1569533753
transform 1 0 168 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2380
timestamp 1569533753
transform 1 0 40 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_2381
timestamp 1569533753
transform 1 0 296 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2382
timestamp 1569533753
transform 1 0 104 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_2383
timestamp 1569533753
transform 1 0 40 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_2384
timestamp 1569533753
transform 1 0 232 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_2385
timestamp 1569533753
transform 1 0 168 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_2386
timestamp 1569533753
transform 1 0 232 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2387
timestamp 1569533753
transform 1 0 168 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2388
timestamp 1569533753
transform 1 0 232 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2389
timestamp 1569533753
transform 1 0 232 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2390
timestamp 1569533753
transform 1 0 232 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2391
timestamp 1569533753
transform 1 0 168 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2392
timestamp 1569533753
transform 1 0 40 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2393
timestamp 1569533753
transform 1 0 40 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2394
timestamp 1569533753
transform 1 0 296 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2395
timestamp 1569533753
transform 1 0 232 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2396
timestamp 1569533753
transform 1 0 296 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2397
timestamp 1569533753
transform 1 0 40 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2398
timestamp 1569533753
transform 1 0 168 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2399
timestamp 1569533753
transform 1 0 104 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2400
timestamp 1569533753
transform 1 0 168 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2401
timestamp 1569533753
transform 1 0 104 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2402
timestamp 1569533753
transform 1 0 104 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2403
timestamp 1569533753
transform 1 0 40 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2404
timestamp 1569533753
transform 1 0 296 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2405
timestamp 1569533753
transform 1 0 296 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2406
timestamp 1569533753
transform 1 0 296 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2407
timestamp 1569533753
transform 1 0 104 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2408
timestamp 1569533753
transform 1 0 40 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2409
timestamp 1569533753
transform 1 0 104 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2410
timestamp 1569533753
transform 1 0 168 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2411
timestamp 1569533753
transform 1 0 616 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2412
timestamp 1569533753
transform 1 0 360 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2413
timestamp 1569533753
transform 1 0 616 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2414
timestamp 1569533753
transform 1 0 616 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2415
timestamp 1569533753
transform 1 0 488 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2416
timestamp 1569533753
transform 1 0 616 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2417
timestamp 1569533753
transform 1 0 360 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2418
timestamp 1569533753
transform 1 0 616 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2419
timestamp 1569533753
transform 1 0 488 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2420
timestamp 1569533753
transform 1 0 360 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2421
timestamp 1569533753
transform 1 0 424 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2422
timestamp 1569533753
transform 1 0 552 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2423
timestamp 1569533753
transform 1 0 488 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2424
timestamp 1569533753
transform 1 0 360 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2425
timestamp 1569533753
transform 1 0 424 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2426
timestamp 1569533753
transform 1 0 488 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2427
timestamp 1569533753
transform 1 0 552 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2428
timestamp 1569533753
transform 1 0 488 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2429
timestamp 1569533753
transform 1 0 424 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2430
timestamp 1569533753
transform 1 0 424 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2431
timestamp 1569533753
transform 1 0 552 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_2432
timestamp 1569533753
transform 1 0 552 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_2433
timestamp 1569533753
transform 1 0 552 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_2434
timestamp 1569533753
transform 1 0 360 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_2435
timestamp 1569533753
transform 1 0 424 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_2436
timestamp 1569533753
transform 1 0 616 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2437
timestamp 1569533753
transform 1 0 552 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2438
timestamp 1569533753
transform 1 0 616 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2439
timestamp 1569533753
transform 1 0 424 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2440
timestamp 1569533753
transform 1 0 360 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2441
timestamp 1569533753
transform 1 0 488 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2442
timestamp 1569533753
transform 1 0 552 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2443
timestamp 1569533753
transform 1 0 360 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2444
timestamp 1569533753
transform 1 0 424 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2445
timestamp 1569533753
transform 1 0 424 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2446
timestamp 1569533753
transform 1 0 488 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2447
timestamp 1569533753
transform 1 0 360 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2448
timestamp 1569533753
transform 1 0 488 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2449
timestamp 1569533753
transform 1 0 552 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2450
timestamp 1569533753
transform 1 0 616 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2451
timestamp 1569533753
transform 1 0 424 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2452
timestamp 1569533753
transform 1 0 616 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2453
timestamp 1569533753
transform 1 0 552 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2454
timestamp 1569533753
transform 1 0 488 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2455
timestamp 1569533753
transform 1 0 360 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2456
timestamp 1569533753
transform 1 0 232 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2457
timestamp 1569533753
transform 1 0 104 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2458
timestamp 1569533753
transform 1 0 168 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2459
timestamp 1569533753
transform 1 0 40 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2460
timestamp 1569533753
transform 1 0 168 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2461
timestamp 1569533753
transform 1 0 296 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2462
timestamp 1569533753
transform 1 0 40 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2463
timestamp 1569533753
transform 1 0 232 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2464
timestamp 1569533753
transform 1 0 40 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2465
timestamp 1569533753
transform 1 0 40 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2466
timestamp 1569533753
transform 1 0 104 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2467
timestamp 1569533753
transform 1 0 296 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2468
timestamp 1569533753
transform 1 0 232 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2469
timestamp 1569533753
transform 1 0 168 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2470
timestamp 1569533753
transform 1 0 296 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2471
timestamp 1569533753
transform 1 0 104 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2472
timestamp 1569533753
transform 1 0 296 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2473
timestamp 1569533753
transform 1 0 168 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2474
timestamp 1569533753
transform 1 0 232 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2475
timestamp 1569533753
transform 1 0 104 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2476
timestamp 1569533753
transform 1 0 296 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2477
timestamp 1569533753
transform 1 0 232 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2478
timestamp 1569533753
transform 1 0 40 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2479
timestamp 1569533753
transform 1 0 104 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2480
timestamp 1569533753
transform 1 0 232 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2481
timestamp 1569533753
transform 1 0 168 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2482
timestamp 1569533753
transform 1 0 104 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2483
timestamp 1569533753
transform 1 0 168 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2484
timestamp 1569533753
transform 1 0 232 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2485
timestamp 1569533753
transform 1 0 296 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2486
timestamp 1569533753
transform 1 0 168 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2487
timestamp 1569533753
transform 1 0 104 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2488
timestamp 1569533753
transform 1 0 296 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2489
timestamp 1569533753
transform 1 0 296 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2490
timestamp 1569533753
transform 1 0 40 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2491
timestamp 1569533753
transform 1 0 40 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2492
timestamp 1569533753
transform 1 0 40 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2493
timestamp 1569533753
transform 1 0 168 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2494
timestamp 1569533753
transform 1 0 232 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2495
timestamp 1569533753
transform 1 0 104 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2496
timestamp 1569533753
transform 1 0 552 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2497
timestamp 1569533753
transform 1 0 360 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2498
timestamp 1569533753
transform 1 0 552 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2499
timestamp 1569533753
transform 1 0 616 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2500
timestamp 1569533753
transform 1 0 424 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2501
timestamp 1569533753
transform 1 0 488 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2502
timestamp 1569533753
transform 1 0 424 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2503
timestamp 1569533753
transform 1 0 616 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2504
timestamp 1569533753
transform 1 0 488 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2505
timestamp 1569533753
transform 1 0 424 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2506
timestamp 1569533753
transform 1 0 616 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2507
timestamp 1569533753
transform 1 0 488 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2508
timestamp 1569533753
transform 1 0 616 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2509
timestamp 1569533753
transform 1 0 552 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2510
timestamp 1569533753
transform 1 0 360 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2511
timestamp 1569533753
transform 1 0 552 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2512
timestamp 1569533753
transform 1 0 360 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2513
timestamp 1569533753
transform 1 0 424 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2514
timestamp 1569533753
transform 1 0 488 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2515
timestamp 1569533753
transform 1 0 360 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2516
timestamp 1569533753
transform 1 0 424 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2517
timestamp 1569533753
transform 1 0 40 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2518
timestamp 1569533753
transform 1 0 296 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2519
timestamp 1569533753
transform 1 0 168 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2520
timestamp 1569533753
transform 1 0 616 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2521
timestamp 1569533753
transform 1 0 488 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2522
timestamp 1569533753
transform 1 0 360 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2523
timestamp 1569533753
transform 1 0 232 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2524
timestamp 1569533753
transform 1 0 104 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2525
timestamp 1569533753
transform 1 0 552 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2526
timestamp 1569533753
transform 1 0 1064 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2527
timestamp 1569533753
transform 1 0 1128 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2528
timestamp 1569533753
transform 1 0 1192 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2529
timestamp 1569533753
transform 1 0 1064 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2530
timestamp 1569533753
transform 1 0 1192 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2531
timestamp 1569533753
transform 1 0 1256 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2532
timestamp 1569533753
transform 1 0 1000 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2533
timestamp 1569533753
transform 1 0 1256 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2534
timestamp 1569533753
transform 1 0 1256 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2535
timestamp 1569533753
transform 1 0 1192 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2536
timestamp 1569533753
transform 1 0 1000 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2537
timestamp 1569533753
transform 1 0 1128 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2538
timestamp 1569533753
transform 1 0 1000 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2539
timestamp 1569533753
transform 1 0 1192 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2540
timestamp 1569533753
transform 1 0 1256 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2541
timestamp 1569533753
transform 1 0 1064 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2542
timestamp 1569533753
transform 1 0 1128 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2543
timestamp 1569533753
transform 1 0 1000 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2544
timestamp 1569533753
transform 1 0 1064 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2545
timestamp 1569533753
transform 1 0 1128 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2546
timestamp 1569533753
transform 1 0 872 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2547
timestamp 1569533753
transform 1 0 680 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2548
timestamp 1569533753
transform 1 0 808 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2549
timestamp 1569533753
transform 1 0 808 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2550
timestamp 1569533753
transform 1 0 936 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2551
timestamp 1569533753
transform 1 0 680 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2552
timestamp 1569533753
transform 1 0 872 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2553
timestamp 1569533753
transform 1 0 744 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2554
timestamp 1569533753
transform 1 0 744 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2555
timestamp 1569533753
transform 1 0 872 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2556
timestamp 1569533753
transform 1 0 872 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2557
timestamp 1569533753
transform 1 0 680 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2558
timestamp 1569533753
transform 1 0 808 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2559
timestamp 1569533753
transform 1 0 744 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_2560
timestamp 1569533753
transform 1 0 936 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_2561
timestamp 1569533753
transform 1 0 936 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2562
timestamp 1569533753
transform 1 0 808 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2563
timestamp 1569533753
transform 1 0 744 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_2564
timestamp 1569533753
transform 1 0 936 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2565
timestamp 1569533753
transform 1 0 680 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_2566
timestamp 1569533753
transform 1 0 680 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2567
timestamp 1569533753
transform 1 0 680 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2568
timestamp 1569533753
transform 1 0 744 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2569
timestamp 1569533753
transform 1 0 808 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2570
timestamp 1569533753
transform 1 0 744 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2571
timestamp 1569533753
transform 1 0 808 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2572
timestamp 1569533753
transform 1 0 936 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2573
timestamp 1569533753
transform 1 0 808 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2574
timestamp 1569533753
transform 1 0 872 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2575
timestamp 1569533753
transform 1 0 936 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2576
timestamp 1569533753
transform 1 0 808 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2577
timestamp 1569533753
transform 1 0 872 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2578
timestamp 1569533753
transform 1 0 936 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2579
timestamp 1569533753
transform 1 0 936 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2580
timestamp 1569533753
transform 1 0 680 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2581
timestamp 1569533753
transform 1 0 680 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2582
timestamp 1569533753
transform 1 0 872 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2583
timestamp 1569533753
transform 1 0 744 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2584
timestamp 1569533753
transform 1 0 872 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2585
timestamp 1569533753
transform 1 0 744 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2586
timestamp 1569533753
transform 1 0 1064 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2587
timestamp 1569533753
transform 1 0 1192 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2588
timestamp 1569533753
transform 1 0 1064 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2589
timestamp 1569533753
transform 1 0 1128 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2590
timestamp 1569533753
transform 1 0 1000 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2591
timestamp 1569533753
transform 1 0 1256 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2592
timestamp 1569533753
transform 1 0 1256 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2593
timestamp 1569533753
transform 1 0 1000 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2594
timestamp 1569533753
transform 1 0 1064 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2595
timestamp 1569533753
transform 1 0 1000 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2596
timestamp 1569533753
transform 1 0 1256 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2597
timestamp 1569533753
transform 1 0 1192 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2598
timestamp 1569533753
transform 1 0 1064 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2599
timestamp 1569533753
transform 1 0 1256 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2600
timestamp 1569533753
transform 1 0 1128 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2601
timestamp 1569533753
transform 1 0 1192 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2602
timestamp 1569533753
transform 1 0 1192 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_2603
timestamp 1569533753
transform 1 0 1128 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_2604
timestamp 1569533753
transform 1 0 1000 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_2605
timestamp 1569533753
transform 1 0 1128 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_2606
timestamp 1569533753
transform 1 0 872 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2607
timestamp 1569533753
transform 1 0 1256 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2608
timestamp 1569533753
transform 1 0 1000 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2609
timestamp 1569533753
transform 1 0 680 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2610
timestamp 1569533753
transform 1 0 1192 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2611
timestamp 1569533753
transform 1 0 744 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2612
timestamp 1569533753
transform 1 0 808 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2613
timestamp 1569533753
transform 1 0 1064 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2614
timestamp 1569533753
transform 1 0 1128 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2615
timestamp 1569533753
transform 1 0 936 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_2616
timestamp 1569533753
transform 1 0 1192 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2617
timestamp 1569533753
transform 1 0 1000 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2618
timestamp 1569533753
transform 1 0 1256 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2619
timestamp 1569533753
transform 1 0 1128 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2620
timestamp 1569533753
transform 1 0 1064 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2621
timestamp 1569533753
transform 1 0 1192 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2622
timestamp 1569533753
transform 1 0 1000 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2623
timestamp 1569533753
transform 1 0 1000 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2624
timestamp 1569533753
transform 1 0 1128 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2625
timestamp 1569533753
transform 1 0 1192 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2626
timestamp 1569533753
transform 1 0 1256 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2627
timestamp 1569533753
transform 1 0 1064 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2628
timestamp 1569533753
transform 1 0 1256 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2629
timestamp 1569533753
transform 1 0 1064 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2630
timestamp 1569533753
transform 1 0 1192 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2631
timestamp 1569533753
transform 1 0 1064 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2632
timestamp 1569533753
transform 1 0 1256 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2633
timestamp 1569533753
transform 1 0 1000 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2634
timestamp 1569533753
transform 1 0 1128 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2635
timestamp 1569533753
transform 1 0 1000 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2636
timestamp 1569533753
transform 1 0 1256 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2637
timestamp 1569533753
transform 1 0 1064 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2638
timestamp 1569533753
transform 1 0 1128 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2639
timestamp 1569533753
transform 1 0 1192 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2640
timestamp 1569533753
transform 1 0 1128 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2641
timestamp 1569533753
transform 1 0 744 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2642
timestamp 1569533753
transform 1 0 936 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2643
timestamp 1569533753
transform 1 0 936 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2644
timestamp 1569533753
transform 1 0 936 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2645
timestamp 1569533753
transform 1 0 872 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2646
timestamp 1569533753
transform 1 0 680 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2647
timestamp 1569533753
transform 1 0 936 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2648
timestamp 1569533753
transform 1 0 872 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2649
timestamp 1569533753
transform 1 0 744 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2650
timestamp 1569533753
transform 1 0 808 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2651
timestamp 1569533753
transform 1 0 744 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2652
timestamp 1569533753
transform 1 0 872 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2653
timestamp 1569533753
transform 1 0 808 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2654
timestamp 1569533753
transform 1 0 744 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2655
timestamp 1569533753
transform 1 0 680 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2656
timestamp 1569533753
transform 1 0 680 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2657
timestamp 1569533753
transform 1 0 808 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2658
timestamp 1569533753
transform 1 0 680 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2659
timestamp 1569533753
transform 1 0 936 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2660
timestamp 1569533753
transform 1 0 872 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2661
timestamp 1569533753
transform 1 0 808 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2662
timestamp 1569533753
transform 1 0 744 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2663
timestamp 1569533753
transform 1 0 808 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2664
timestamp 1569533753
transform 1 0 872 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2665
timestamp 1569533753
transform 1 0 680 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2666
timestamp 1569533753
transform 1 0 744 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2667
timestamp 1569533753
transform 1 0 936 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2668
timestamp 1569533753
transform 1 0 872 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2669
timestamp 1569533753
transform 1 0 936 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2670
timestamp 1569533753
transform 1 0 808 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2671
timestamp 1569533753
transform 1 0 808 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2672
timestamp 1569533753
transform 1 0 872 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2673
timestamp 1569533753
transform 1 0 872 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2674
timestamp 1569533753
transform 1 0 808 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2675
timestamp 1569533753
transform 1 0 936 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2676
timestamp 1569533753
transform 1 0 680 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2677
timestamp 1569533753
transform 1 0 872 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2678
timestamp 1569533753
transform 1 0 680 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2679
timestamp 1569533753
transform 1 0 744 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2680
timestamp 1569533753
transform 1 0 680 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2681
timestamp 1569533753
transform 1 0 872 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2682
timestamp 1569533753
transform 1 0 680 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2683
timestamp 1569533753
transform 1 0 744 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2684
timestamp 1569533753
transform 1 0 808 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2685
timestamp 1569533753
transform 1 0 936 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2686
timestamp 1569533753
transform 1 0 936 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2687
timestamp 1569533753
transform 1 0 744 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2688
timestamp 1569533753
transform 1 0 744 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2689
timestamp 1569533753
transform 1 0 808 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2690
timestamp 1569533753
transform 1 0 680 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2691
timestamp 1569533753
transform 1 0 1128 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2692
timestamp 1569533753
transform 1 0 1000 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2693
timestamp 1569533753
transform 1 0 1256 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2694
timestamp 1569533753
transform 1 0 1256 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2695
timestamp 1569533753
transform 1 0 1256 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2696
timestamp 1569533753
transform 1 0 1256 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2697
timestamp 1569533753
transform 1 0 1192 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2698
timestamp 1569533753
transform 1 0 1128 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2699
timestamp 1569533753
transform 1 0 1000 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2700
timestamp 1569533753
transform 1 0 1192 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2701
timestamp 1569533753
transform 1 0 1000 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2702
timestamp 1569533753
transform 1 0 1064 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2703
timestamp 1569533753
transform 1 0 1192 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2704
timestamp 1569533753
transform 1 0 1000 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2705
timestamp 1569533753
transform 1 0 1000 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2706
timestamp 1569533753
transform 1 0 1192 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2707
timestamp 1569533753
transform 1 0 1064 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2708
timestamp 1569533753
transform 1 0 1064 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2709
timestamp 1569533753
transform 1 0 1064 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2710
timestamp 1569533753
transform 1 0 1128 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2711
timestamp 1569533753
transform 1 0 1256 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2712
timestamp 1569533753
transform 1 0 1128 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2713
timestamp 1569533753
transform 1 0 1128 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2714
timestamp 1569533753
transform 1 0 1192 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2715
timestamp 1569533753
transform 1 0 1064 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2716
timestamp 1569533753
transform 1 0 424 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2717
timestamp 1569533753
transform 1 0 424 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2718
timestamp 1569533753
transform 1 0 488 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2719
timestamp 1569533753
transform 1 0 616 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2720
timestamp 1569533753
transform 1 0 552 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2721
timestamp 1569533753
transform 1 0 360 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2722
timestamp 1569533753
transform 1 0 488 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2723
timestamp 1569533753
transform 1 0 360 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2724
timestamp 1569533753
transform 1 0 424 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2725
timestamp 1569533753
transform 1 0 488 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2726
timestamp 1569533753
transform 1 0 424 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2727
timestamp 1569533753
transform 1 0 616 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2728
timestamp 1569533753
transform 1 0 488 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2729
timestamp 1569533753
transform 1 0 616 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2730
timestamp 1569533753
transform 1 0 552 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2731
timestamp 1569533753
transform 1 0 360 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2732
timestamp 1569533753
transform 1 0 360 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2733
timestamp 1569533753
transform 1 0 616 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2734
timestamp 1569533753
transform 1 0 552 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2735
timestamp 1569533753
transform 1 0 424 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2736
timestamp 1569533753
transform 1 0 552 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2737
timestamp 1569533753
transform 1 0 616 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2738
timestamp 1569533753
transform 1 0 552 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2739
timestamp 1569533753
transform 1 0 360 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2740
timestamp 1569533753
transform 1 0 488 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2741
timestamp 1569533753
transform 1 0 104 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2742
timestamp 1569533753
transform 1 0 104 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2743
timestamp 1569533753
transform 1 0 40 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2744
timestamp 1569533753
transform 1 0 232 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2745
timestamp 1569533753
transform 1 0 232 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2746
timestamp 1569533753
transform 1 0 40 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2747
timestamp 1569533753
transform 1 0 40 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2748
timestamp 1569533753
transform 1 0 40 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2749
timestamp 1569533753
transform 1 0 104 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2750
timestamp 1569533753
transform 1 0 168 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2751
timestamp 1569533753
transform 1 0 232 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2752
timestamp 1569533753
transform 1 0 296 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_2753
timestamp 1569533753
transform 1 0 232 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2754
timestamp 1569533753
transform 1 0 104 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2755
timestamp 1569533753
transform 1 0 40 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2756
timestamp 1569533753
transform 1 0 168 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2757
timestamp 1569533753
transform 1 0 296 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2758
timestamp 1569533753
transform 1 0 168 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2759
timestamp 1569533753
transform 1 0 232 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2760
timestamp 1569533753
transform 1 0 296 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2761
timestamp 1569533753
transform 1 0 168 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_2762
timestamp 1569533753
transform 1 0 168 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2763
timestamp 1569533753
transform 1 0 296 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2764
timestamp 1569533753
transform 1 0 104 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_2765
timestamp 1569533753
transform 1 0 296 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_2766
timestamp 1569533753
transform 1 0 232 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2767
timestamp 1569533753
transform 1 0 168 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2768
timestamp 1569533753
transform 1 0 168 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2769
timestamp 1569533753
transform 1 0 232 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2770
timestamp 1569533753
transform 1 0 104 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2771
timestamp 1569533753
transform 1 0 232 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2772
timestamp 1569533753
transform 1 0 168 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2773
timestamp 1569533753
transform 1 0 296 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2774
timestamp 1569533753
transform 1 0 104 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2775
timestamp 1569533753
transform 1 0 40 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2776
timestamp 1569533753
transform 1 0 296 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2777
timestamp 1569533753
transform 1 0 296 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2778
timestamp 1569533753
transform 1 0 296 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2779
timestamp 1569533753
transform 1 0 104 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2780
timestamp 1569533753
transform 1 0 232 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2781
timestamp 1569533753
transform 1 0 40 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2782
timestamp 1569533753
transform 1 0 40 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2783
timestamp 1569533753
transform 1 0 40 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2784
timestamp 1569533753
transform 1 0 168 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2785
timestamp 1569533753
transform 1 0 232 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2786
timestamp 1569533753
transform 1 0 104 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2787
timestamp 1569533753
transform 1 0 104 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2788
timestamp 1569533753
transform 1 0 296 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2789
timestamp 1569533753
transform 1 0 40 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2790
timestamp 1569533753
transform 1 0 168 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2791
timestamp 1569533753
transform 1 0 616 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2792
timestamp 1569533753
transform 1 0 616 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2793
timestamp 1569533753
transform 1 0 424 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2794
timestamp 1569533753
transform 1 0 488 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2795
timestamp 1569533753
transform 1 0 488 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2796
timestamp 1569533753
transform 1 0 424 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2797
timestamp 1569533753
transform 1 0 424 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2798
timestamp 1569533753
transform 1 0 552 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2799
timestamp 1569533753
transform 1 0 360 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2800
timestamp 1569533753
transform 1 0 424 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2801
timestamp 1569533753
transform 1 0 552 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2802
timestamp 1569533753
transform 1 0 360 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2803
timestamp 1569533753
transform 1 0 552 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2804
timestamp 1569533753
transform 1 0 360 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2805
timestamp 1569533753
transform 1 0 360 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2806
timestamp 1569533753
transform 1 0 552 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2807
timestamp 1569533753
transform 1 0 616 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2808
timestamp 1569533753
transform 1 0 616 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2809
timestamp 1569533753
transform 1 0 616 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_2810
timestamp 1569533753
transform 1 0 360 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2811
timestamp 1569533753
transform 1 0 424 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_2812
timestamp 1569533753
transform 1 0 488 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2813
timestamp 1569533753
transform 1 0 488 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2814
timestamp 1569533753
transform 1 0 552 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_2815
timestamp 1569533753
transform 1 0 488 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2816
timestamp 1569533753
transform 1 0 424 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2817
timestamp 1569533753
transform 1 0 424 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2818
timestamp 1569533753
transform 1 0 360 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2819
timestamp 1569533753
transform 1 0 616 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2820
timestamp 1569533753
transform 1 0 488 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2821
timestamp 1569533753
transform 1 0 488 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2822
timestamp 1569533753
transform 1 0 424 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2823
timestamp 1569533753
transform 1 0 360 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2824
timestamp 1569533753
transform 1 0 488 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2825
timestamp 1569533753
transform 1 0 552 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2826
timestamp 1569533753
transform 1 0 552 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2827
timestamp 1569533753
transform 1 0 360 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2828
timestamp 1569533753
transform 1 0 616 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2829
timestamp 1569533753
transform 1 0 616 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2830
timestamp 1569533753
transform 1 0 488 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2831
timestamp 1569533753
transform 1 0 360 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2832
timestamp 1569533753
transform 1 0 360 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2833
timestamp 1569533753
transform 1 0 424 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2834
timestamp 1569533753
transform 1 0 616 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2835
timestamp 1569533753
transform 1 0 552 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2836
timestamp 1569533753
transform 1 0 488 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2837
timestamp 1569533753
transform 1 0 552 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2838
timestamp 1569533753
transform 1 0 424 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2839
timestamp 1569533753
transform 1 0 616 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2840
timestamp 1569533753
transform 1 0 552 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2841
timestamp 1569533753
transform 1 0 40 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2842
timestamp 1569533753
transform 1 0 232 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2843
timestamp 1569533753
transform 1 0 104 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2844
timestamp 1569533753
transform 1 0 232 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2845
timestamp 1569533753
transform 1 0 232 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2846
timestamp 1569533753
transform 1 0 168 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2847
timestamp 1569533753
transform 1 0 296 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2848
timestamp 1569533753
transform 1 0 296 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2849
timestamp 1569533753
transform 1 0 232 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2850
timestamp 1569533753
transform 1 0 40 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2851
timestamp 1569533753
transform 1 0 296 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2852
timestamp 1569533753
transform 1 0 104 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2853
timestamp 1569533753
transform 1 0 296 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2854
timestamp 1569533753
transform 1 0 296 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2855
timestamp 1569533753
transform 1 0 104 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2856
timestamp 1569533753
transform 1 0 232 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2857
timestamp 1569533753
transform 1 0 104 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2858
timestamp 1569533753
transform 1 0 168 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2859
timestamp 1569533753
transform 1 0 104 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2860
timestamp 1569533753
transform 1 0 168 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2861
timestamp 1569533753
transform 1 0 40 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2862
timestamp 1569533753
transform 1 0 168 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2863
timestamp 1569533753
transform 1 0 40 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2864
timestamp 1569533753
transform 1 0 40 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2865
timestamp 1569533753
transform 1 0 168 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2866
timestamp 1569533753
transform 1 0 40 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2867
timestamp 1569533753
transform 1 0 232 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2868
timestamp 1569533753
transform 1 0 296 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2869
timestamp 1569533753
transform 1 0 232 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2870
timestamp 1569533753
transform 1 0 168 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2871
timestamp 1569533753
transform 1 0 168 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2872
timestamp 1569533753
transform 1 0 104 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2873
timestamp 1569533753
transform 1 0 232 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2874
timestamp 1569533753
transform 1 0 296 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2875
timestamp 1569533753
transform 1 0 296 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2876
timestamp 1569533753
transform 1 0 104 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2877
timestamp 1569533753
transform 1 0 296 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2878
timestamp 1569533753
transform 1 0 104 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2879
timestamp 1569533753
transform 1 0 232 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2880
timestamp 1569533753
transform 1 0 168 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2881
timestamp 1569533753
transform 1 0 168 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2882
timestamp 1569533753
transform 1 0 40 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2883
timestamp 1569533753
transform 1 0 40 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2884
timestamp 1569533753
transform 1 0 40 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2885
timestamp 1569533753
transform 1 0 104 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2886
timestamp 1569533753
transform 1 0 552 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2887
timestamp 1569533753
transform 1 0 424 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2888
timestamp 1569533753
transform 1 0 488 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2889
timestamp 1569533753
transform 1 0 424 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2890
timestamp 1569533753
transform 1 0 552 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2891
timestamp 1569533753
transform 1 0 360 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2892
timestamp 1569533753
transform 1 0 616 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2893
timestamp 1569533753
transform 1 0 616 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2894
timestamp 1569533753
transform 1 0 552 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2895
timestamp 1569533753
transform 1 0 616 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2896
timestamp 1569533753
transform 1 0 616 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2897
timestamp 1569533753
transform 1 0 488 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2898
timestamp 1569533753
transform 1 0 424 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2899
timestamp 1569533753
transform 1 0 488 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2900
timestamp 1569533753
transform 1 0 360 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2901
timestamp 1569533753
transform 1 0 360 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2902
timestamp 1569533753
transform 1 0 552 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2903
timestamp 1569533753
transform 1 0 424 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2904
timestamp 1569533753
transform 1 0 488 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2905
timestamp 1569533753
transform 1 0 360 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2906
timestamp 1569533753
transform 1 0 1128 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2907
timestamp 1569533753
transform 1 0 1000 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2908
timestamp 1569533753
transform 1 0 1256 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2909
timestamp 1569533753
transform 1 0 1064 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2910
timestamp 1569533753
transform 1 0 1192 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2911
timestamp 1569533753
transform 1 0 1192 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2912
timestamp 1569533753
transform 1 0 1192 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2913
timestamp 1569533753
transform 1 0 1256 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2914
timestamp 1569533753
transform 1 0 1256 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2915
timestamp 1569533753
transform 1 0 1256 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2916
timestamp 1569533753
transform 1 0 1256 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2917
timestamp 1569533753
transform 1 0 1064 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2918
timestamp 1569533753
transform 1 0 1064 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2919
timestamp 1569533753
transform 1 0 1192 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2920
timestamp 1569533753
transform 1 0 1000 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2921
timestamp 1569533753
transform 1 0 1064 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2922
timestamp 1569533753
transform 1 0 1128 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2923
timestamp 1569533753
transform 1 0 1000 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2924
timestamp 1569533753
transform 1 0 1000 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2925
timestamp 1569533753
transform 1 0 1128 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2926
timestamp 1569533753
transform 1 0 1128 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2927
timestamp 1569533753
transform 1 0 1128 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2928
timestamp 1569533753
transform 1 0 1064 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2929
timestamp 1569533753
transform 1 0 1000 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2930
timestamp 1569533753
transform 1 0 1192 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2931
timestamp 1569533753
transform 1 0 936 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2932
timestamp 1569533753
transform 1 0 808 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2933
timestamp 1569533753
transform 1 0 936 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2934
timestamp 1569533753
transform 1 0 808 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2935
timestamp 1569533753
transform 1 0 872 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2936
timestamp 1569533753
transform 1 0 936 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2937
timestamp 1569533753
transform 1 0 872 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2938
timestamp 1569533753
transform 1 0 872 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2939
timestamp 1569533753
transform 1 0 680 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2940
timestamp 1569533753
transform 1 0 680 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2941
timestamp 1569533753
transform 1 0 680 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2942
timestamp 1569533753
transform 1 0 872 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2943
timestamp 1569533753
transform 1 0 680 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2944
timestamp 1569533753
transform 1 0 680 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2945
timestamp 1569533753
transform 1 0 936 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2946
timestamp 1569533753
transform 1 0 744 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_2947
timestamp 1569533753
transform 1 0 808 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2948
timestamp 1569533753
transform 1 0 744 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2949
timestamp 1569533753
transform 1 0 808 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2950
timestamp 1569533753
transform 1 0 744 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_2951
timestamp 1569533753
transform 1 0 808 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2952
timestamp 1569533753
transform 1 0 744 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_2953
timestamp 1569533753
transform 1 0 744 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2954
timestamp 1569533753
transform 1 0 872 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_2955
timestamp 1569533753
transform 1 0 936 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_2956
timestamp 1569533753
transform 1 0 808 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2957
timestamp 1569533753
transform 1 0 872 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2958
timestamp 1569533753
transform 1 0 936 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2959
timestamp 1569533753
transform 1 0 808 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2960
timestamp 1569533753
transform 1 0 872 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2961
timestamp 1569533753
transform 1 0 872 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2962
timestamp 1569533753
transform 1 0 680 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2963
timestamp 1569533753
transform 1 0 680 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2964
timestamp 1569533753
transform 1 0 680 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2965
timestamp 1569533753
transform 1 0 680 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2966
timestamp 1569533753
transform 1 0 872 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2967
timestamp 1569533753
transform 1 0 808 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2968
timestamp 1569533753
transform 1 0 936 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2969
timestamp 1569533753
transform 1 0 744 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2970
timestamp 1569533753
transform 1 0 744 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2971
timestamp 1569533753
transform 1 0 744 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2972
timestamp 1569533753
transform 1 0 744 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2973
timestamp 1569533753
transform 1 0 936 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2974
timestamp 1569533753
transform 1 0 808 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2975
timestamp 1569533753
transform 1 0 936 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2976
timestamp 1569533753
transform 1 0 1192 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2977
timestamp 1569533753
transform 1 0 1064 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2978
timestamp 1569533753
transform 1 0 1256 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2979
timestamp 1569533753
transform 1 0 1256 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2980
timestamp 1569533753
transform 1 0 1256 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2981
timestamp 1569533753
transform 1 0 1256 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2982
timestamp 1569533753
transform 1 0 1192 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2983
timestamp 1569533753
transform 1 0 1128 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2984
timestamp 1569533753
transform 1 0 1064 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2985
timestamp 1569533753
transform 1 0 1000 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2986
timestamp 1569533753
transform 1 0 1000 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2987
timestamp 1569533753
transform 1 0 1128 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2988
timestamp 1569533753
transform 1 0 1192 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2989
timestamp 1569533753
transform 1 0 1064 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2990
timestamp 1569533753
transform 1 0 1192 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2991
timestamp 1569533753
transform 1 0 1000 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2992
timestamp 1569533753
transform 1 0 1128 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_2993
timestamp 1569533753
transform 1 0 1064 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_2994
timestamp 1569533753
transform 1 0 1000 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_2995
timestamp 1569533753
transform 1 0 1128 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_2996
timestamp 1569533753
transform 1 0 2344 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_2997
timestamp 1569533753
transform 1 0 2344 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_2998
timestamp 1569533753
transform 1 0 2344 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_2999
timestamp 1569533753
transform 1 0 2408 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3000
timestamp 1569533753
transform 1 0 2408 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3001
timestamp 1569533753
transform 1 0 2408 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3002
timestamp 1569533753
transform 1 0 2344 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3003
timestamp 1569533753
transform 1 0 2408 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3004
timestamp 1569533753
transform 1 0 2408 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3005
timestamp 1569533753
transform 1 0 2408 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3006
timestamp 1569533753
transform 1 0 2408 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3007
timestamp 1569533753
transform 1 0 2344 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3008
timestamp 1569533753
transform 1 0 2408 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3009
timestamp 1569533753
transform 1 0 2472 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3010
timestamp 1569533753
transform 1 0 2472 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3011
timestamp 1569533753
transform 1 0 2472 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3012
timestamp 1569533753
transform 1 0 2344 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3013
timestamp 1569533753
transform 1 0 2472 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3014
timestamp 1569533753
transform 1 0 2472 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3015
timestamp 1569533753
transform 1 0 2472 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3016
timestamp 1569533753
transform 1 0 2344 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3017
timestamp 1569533753
transform 1 0 2472 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3018
timestamp 1569533753
transform 1 0 2472 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3019
timestamp 1569533753
transform 1 0 2472 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3020
timestamp 1569533753
transform 1 0 2408 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3021
timestamp 1569533753
transform 1 0 2472 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3022
timestamp 1569533753
transform 1 0 2344 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3023
timestamp 1569533753
transform 1 0 2344 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3024
timestamp 1569533753
transform 1 0 2408 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3025
timestamp 1569533753
transform 1 0 2344 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3026
timestamp 1569533753
transform 1 0 1384 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3027
timestamp 1569533753
transform 1 0 1384 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3028
timestamp 1569533753
transform 1 0 1384 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3029
timestamp 1569533753
transform 1 0 1384 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3030
timestamp 1569533753
transform 1 0 1320 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3031
timestamp 1569533753
transform 1 0 1320 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3032
timestamp 1569533753
transform 1 0 1448 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3033
timestamp 1569533753
transform 1 0 1384 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3034
timestamp 1569533753
transform 1 0 1384 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3035
timestamp 1569533753
transform 1 0 1448 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3036
timestamp 1569533753
transform 1 0 1448 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3037
timestamp 1569533753
transform 1 0 1448 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3038
timestamp 1569533753
transform 1 0 1448 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3039
timestamp 1569533753
transform 1 0 1384 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3040
timestamp 1569533753
transform 1 0 1448 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3041
timestamp 1569533753
transform 1 0 1384 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3042
timestamp 1569533753
transform 1 0 1384 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3043
timestamp 1569533753
transform 1 0 1448 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3044
timestamp 1569533753
transform 1 0 1448 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3045
timestamp 1569533753
transform 1 0 1448 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3046
timestamp 1569533753
transform 1 0 1448 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3047
timestamp 1569533753
transform 1 0 1512 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3048
timestamp 1569533753
transform 1 0 1512 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3049
timestamp 1569533753
transform 1 0 1512 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3050
timestamp 1569533753
transform 1 0 1512 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3051
timestamp 1569533753
transform 1 0 1512 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3052
timestamp 1569533753
transform 1 0 1512 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3053
timestamp 1569533753
transform 1 0 1512 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3054
timestamp 1569533753
transform 1 0 1512 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3055
timestamp 1569533753
transform 1 0 1320 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3056
timestamp 1569533753
transform 1 0 1320 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3057
timestamp 1569533753
transform 1 0 1320 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3058
timestamp 1569533753
transform 1 0 1320 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3059
timestamp 1569533753
transform 1 0 1320 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3060
timestamp 1569533753
transform 1 0 1320 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3061
timestamp 1569533753
transform 1 0 1320 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3062
timestamp 1569533753
transform 1 0 1512 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3063
timestamp 1569533753
transform 1 0 1320 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3064
timestamp 1569533753
transform 1 0 1384 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3065
timestamp 1569533753
transform 1 0 1512 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3066
timestamp 1569533753
transform 1 0 1512 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3067
timestamp 1569533753
transform 1 0 1448 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3068
timestamp 1569533753
transform 1 0 1512 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3069
timestamp 1569533753
transform 1 0 1448 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3070
timestamp 1569533753
transform 1 0 1448 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3071
timestamp 1569533753
transform 1 0 1512 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3072
timestamp 1569533753
transform 1 0 1320 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3073
timestamp 1569533753
transform 1 0 1320 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3074
timestamp 1569533753
transform 1 0 1320 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3075
timestamp 1569533753
transform 1 0 1320 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3076
timestamp 1569533753
transform 1 0 1320 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3077
timestamp 1569533753
transform 1 0 1512 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3078
timestamp 1569533753
transform 1 0 1320 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3079
timestamp 1569533753
transform 1 0 1320 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3080
timestamp 1569533753
transform 1 0 1320 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3081
timestamp 1569533753
transform 1 0 1320 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3082
timestamp 1569533753
transform 1 0 1384 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3083
timestamp 1569533753
transform 1 0 1384 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3084
timestamp 1569533753
transform 1 0 1512 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3085
timestamp 1569533753
transform 1 0 1384 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3086
timestamp 1569533753
transform 1 0 1448 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3087
timestamp 1569533753
transform 1 0 1384 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3088
timestamp 1569533753
transform 1 0 1384 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3089
timestamp 1569533753
transform 1 0 1384 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3090
timestamp 1569533753
transform 1 0 1384 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3091
timestamp 1569533753
transform 1 0 1384 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3092
timestamp 1569533753
transform 1 0 1384 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3093
timestamp 1569533753
transform 1 0 1448 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3094
timestamp 1569533753
transform 1 0 1448 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3095
timestamp 1569533753
transform 1 0 1448 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3096
timestamp 1569533753
transform 1 0 1448 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3097
timestamp 1569533753
transform 1 0 1512 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3098
timestamp 1569533753
transform 1 0 1512 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3099
timestamp 1569533753
transform 1 0 1512 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3100
timestamp 1569533753
transform 1 0 1512 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3101
timestamp 1569533753
transform 1 0 1448 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3102
timestamp 1569533753
transform 1 0 2344 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3103
timestamp 1569533753
transform 1 0 2344 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3104
timestamp 1569533753
transform 1 0 2344 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3105
timestamp 1569533753
transform 1 0 2344 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3106
timestamp 1569533753
transform 1 0 2408 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3107
timestamp 1569533753
transform 1 0 2472 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3108
timestamp 1569533753
transform 1 0 2344 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_3109
timestamp 1569533753
transform 1 0 2344 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3110
timestamp 1569533753
transform 1 0 2472 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3111
timestamp 1569533753
transform 1 0 2472 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3112
timestamp 1569533753
transform 1 0 2344 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3113
timestamp 1569533753
transform 1 0 2344 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3114
timestamp 1569533753
transform 1 0 2344 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3115
timestamp 1569533753
transform 1 0 2472 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3116
timestamp 1569533753
transform 1 0 2472 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3117
timestamp 1569533753
transform 1 0 2408 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3118
timestamp 1569533753
transform 1 0 2408 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3119
timestamp 1569533753
transform 1 0 2408 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3120
timestamp 1569533753
transform 1 0 2408 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3121
timestamp 1569533753
transform 1 0 2408 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3122
timestamp 1569533753
transform 1 0 2408 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_3123
timestamp 1569533753
transform 1 0 2408 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3124
timestamp 1569533753
transform 1 0 2472 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_3125
timestamp 1569533753
transform 1 0 2408 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3126
timestamp 1569533753
transform 1 0 2472 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_3127
timestamp 1569533753
transform 1 0 2472 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3128
timestamp 1569533753
transform 1 0 2472 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3129
timestamp 1569533753
transform 1 0 4840 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3130
timestamp 1569533753
transform 1 0 4840 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3131
timestamp 1569533753
transform 1 0 4904 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3132
timestamp 1569533753
transform 1 0 4712 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3133
timestamp 1569533753
transform 1 0 4776 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3134
timestamp 1569533753
transform 1 0 4904 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3135
timestamp 1569533753
transform 1 0 4840 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3136
timestamp 1569533753
transform 1 0 4904 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3137
timestamp 1569533753
transform 1 0 4776 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3138
timestamp 1569533753
transform 1 0 4776 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3139
timestamp 1569533753
transform 1 0 4840 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3140
timestamp 1569533753
transform 1 0 4712 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3141
timestamp 1569533753
transform 1 0 4712 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3142
timestamp 1569533753
transform 1 0 4776 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3143
timestamp 1569533753
transform 1 0 4712 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3144
timestamp 1569533753
transform 1 0 4712 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3145
timestamp 1569533753
transform 1 0 4840 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3146
timestamp 1569533753
transform 1 0 4904 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3147
timestamp 1569533753
transform 1 0 4776 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3148
timestamp 1569533753
transform 1 0 4904 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3149
timestamp 1569533753
transform 1 0 4520 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3150
timestamp 1569533753
transform 1 0 4648 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3151
timestamp 1569533753
transform 1 0 4456 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3152
timestamp 1569533753
transform 1 0 4456 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3153
timestamp 1569533753
transform 1 0 4648 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3154
timestamp 1569533753
transform 1 0 4392 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3155
timestamp 1569533753
transform 1 0 4584 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3156
timestamp 1569533753
transform 1 0 4392 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3157
timestamp 1569533753
transform 1 0 4520 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3158
timestamp 1569533753
transform 1 0 4648 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3159
timestamp 1569533753
transform 1 0 4584 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3160
timestamp 1569533753
transform 1 0 4456 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3161
timestamp 1569533753
transform 1 0 4584 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3162
timestamp 1569533753
transform 1 0 4648 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3163
timestamp 1569533753
transform 1 0 4392 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3164
timestamp 1569533753
transform 1 0 4520 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3165
timestamp 1569533753
transform 1 0 4520 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3166
timestamp 1569533753
transform 1 0 4520 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3167
timestamp 1569533753
transform 1 0 4456 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3168
timestamp 1569533753
transform 1 0 4584 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3169
timestamp 1569533753
transform 1 0 4392 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3170
timestamp 1569533753
transform 1 0 4392 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3171
timestamp 1569533753
transform 1 0 4456 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3172
timestamp 1569533753
transform 1 0 4584 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3173
timestamp 1569533753
transform 1 0 4648 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3174
timestamp 1569533753
transform 1 0 4392 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3175
timestamp 1569533753
transform 1 0 4456 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3176
timestamp 1569533753
transform 1 0 4520 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3177
timestamp 1569533753
transform 1 0 4392 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3178
timestamp 1569533753
transform 1 0 4584 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3179
timestamp 1569533753
transform 1 0 4392 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3180
timestamp 1569533753
transform 1 0 4520 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3181
timestamp 1569533753
transform 1 0 4584 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3182
timestamp 1569533753
transform 1 0 4392 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3183
timestamp 1569533753
transform 1 0 4392 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3184
timestamp 1569533753
transform 1 0 4456 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3185
timestamp 1569533753
transform 1 0 4456 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3186
timestamp 1569533753
transform 1 0 4648 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3187
timestamp 1569533753
transform 1 0 4584 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3188
timestamp 1569533753
transform 1 0 4456 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3189
timestamp 1569533753
transform 1 0 4520 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3190
timestamp 1569533753
transform 1 0 4584 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3191
timestamp 1569533753
transform 1 0 4520 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3192
timestamp 1569533753
transform 1 0 4648 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3193
timestamp 1569533753
transform 1 0 4648 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3194
timestamp 1569533753
transform 1 0 4648 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3195
timestamp 1569533753
transform 1 0 4584 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3196
timestamp 1569533753
transform 1 0 4520 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3197
timestamp 1569533753
transform 1 0 4456 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3198
timestamp 1569533753
transform 1 0 4648 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3199
timestamp 1569533753
transform 1 0 4776 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3200
timestamp 1569533753
transform 1 0 4904 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3201
timestamp 1569533753
transform 1 0 4904 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3202
timestamp 1569533753
transform 1 0 4840 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3203
timestamp 1569533753
transform 1 0 4712 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3204
timestamp 1569533753
transform 1 0 4904 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3205
timestamp 1569533753
transform 1 0 4712 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3206
timestamp 1569533753
transform 1 0 4776 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3207
timestamp 1569533753
transform 1 0 4840 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3208
timestamp 1569533753
transform 1 0 4712 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3209
timestamp 1569533753
transform 1 0 4904 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3210
timestamp 1569533753
transform 1 0 4776 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3211
timestamp 1569533753
transform 1 0 4776 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3212
timestamp 1569533753
transform 1 0 4840 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3213
timestamp 1569533753
transform 1 0 4712 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3214
timestamp 1569533753
transform 1 0 4776 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3215
timestamp 1569533753
transform 1 0 4840 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3216
timestamp 1569533753
transform 1 0 4904 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3217
timestamp 1569533753
transform 1 0 4840 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3218
timestamp 1569533753
transform 1 0 4712 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3219
timestamp 1569533753
transform 1 0 4328 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3220
timestamp 1569533753
transform 1 0 4136 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3221
timestamp 1569533753
transform 1 0 4200 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3222
timestamp 1569533753
transform 1 0 4264 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3223
timestamp 1569533753
transform 1 0 4264 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3224
timestamp 1569533753
transform 1 0 4264 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3225
timestamp 1569533753
transform 1 0 4072 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3226
timestamp 1569533753
transform 1 0 4328 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3227
timestamp 1569533753
transform 1 0 4264 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3228
timestamp 1569533753
transform 1 0 4200 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3229
timestamp 1569533753
transform 1 0 4136 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3230
timestamp 1569533753
transform 1 0 4136 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3231
timestamp 1569533753
transform 1 0 4072 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3232
timestamp 1569533753
transform 1 0 4328 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3233
timestamp 1569533753
transform 1 0 4200 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3234
timestamp 1569533753
transform 1 0 4072 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3235
timestamp 1569533753
transform 1 0 4072 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3236
timestamp 1569533753
transform 1 0 4264 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3237
timestamp 1569533753
transform 1 0 4200 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3238
timestamp 1569533753
transform 1 0 4136 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3239
timestamp 1569533753
transform 1 0 4328 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3240
timestamp 1569533753
transform 1 0 4136 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3241
timestamp 1569533753
transform 1 0 4200 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3242
timestamp 1569533753
transform 1 0 4328 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3243
timestamp 1569533753
transform 1 0 4072 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3244
timestamp 1569533753
transform 1 0 3816 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3245
timestamp 1569533753
transform 1 0 3880 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3246
timestamp 1569533753
transform 1 0 3752 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3247
timestamp 1569533753
transform 1 0 4008 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3248
timestamp 1569533753
transform 1 0 3752 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3249
timestamp 1569533753
transform 1 0 3880 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3250
timestamp 1569533753
transform 1 0 3944 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3251
timestamp 1569533753
transform 1 0 3944 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3252
timestamp 1569533753
transform 1 0 3944 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3253
timestamp 1569533753
transform 1 0 4008 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3254
timestamp 1569533753
transform 1 0 3752 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3255
timestamp 1569533753
transform 1 0 3944 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3256
timestamp 1569533753
transform 1 0 3944 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3257
timestamp 1569533753
transform 1 0 3752 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3258
timestamp 1569533753
transform 1 0 4008 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3259
timestamp 1569533753
transform 1 0 3880 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3260
timestamp 1569533753
transform 1 0 3816 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3261
timestamp 1569533753
transform 1 0 4008 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3262
timestamp 1569533753
transform 1 0 3816 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3263
timestamp 1569533753
transform 1 0 3880 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3264
timestamp 1569533753
transform 1 0 4008 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3265
timestamp 1569533753
transform 1 0 3816 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3266
timestamp 1569533753
transform 1 0 3816 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3267
timestamp 1569533753
transform 1 0 3752 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3268
timestamp 1569533753
transform 1 0 3880 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3269
timestamp 1569533753
transform 1 0 3944 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3270
timestamp 1569533753
transform 1 0 3752 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3271
timestamp 1569533753
transform 1 0 4008 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3272
timestamp 1569533753
transform 1 0 3880 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3273
timestamp 1569533753
transform 1 0 3752 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3274
timestamp 1569533753
transform 1 0 3944 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3275
timestamp 1569533753
transform 1 0 3880 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3276
timestamp 1569533753
transform 1 0 3752 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3277
timestamp 1569533753
transform 1 0 3752 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3278
timestamp 1569533753
transform 1 0 3944 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3279
timestamp 1569533753
transform 1 0 3816 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3280
timestamp 1569533753
transform 1 0 3944 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3281
timestamp 1569533753
transform 1 0 4008 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3282
timestamp 1569533753
transform 1 0 3880 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3283
timestamp 1569533753
transform 1 0 3816 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3284
timestamp 1569533753
transform 1 0 3816 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3285
timestamp 1569533753
transform 1 0 3816 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3286
timestamp 1569533753
transform 1 0 3816 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3287
timestamp 1569533753
transform 1 0 4008 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3288
timestamp 1569533753
transform 1 0 3752 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3289
timestamp 1569533753
transform 1 0 4008 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3290
timestamp 1569533753
transform 1 0 4008 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3291
timestamp 1569533753
transform 1 0 3944 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3292
timestamp 1569533753
transform 1 0 3880 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3293
timestamp 1569533753
transform 1 0 3880 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3294
timestamp 1569533753
transform 1 0 4136 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3295
timestamp 1569533753
transform 1 0 4200 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3296
timestamp 1569533753
transform 1 0 4136 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3297
timestamp 1569533753
transform 1 0 4264 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3298
timestamp 1569533753
transform 1 0 4264 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3299
timestamp 1569533753
transform 1 0 4072 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3300
timestamp 1569533753
transform 1 0 4200 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3301
timestamp 1569533753
transform 1 0 4072 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3302
timestamp 1569533753
transform 1 0 4136 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3303
timestamp 1569533753
transform 1 0 4264 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3304
timestamp 1569533753
transform 1 0 4072 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3305
timestamp 1569533753
transform 1 0 4136 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3306
timestamp 1569533753
transform 1 0 4264 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3307
timestamp 1569533753
transform 1 0 4136 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3308
timestamp 1569533753
transform 1 0 4200 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3309
timestamp 1569533753
transform 1 0 4264 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3310
timestamp 1569533753
transform 1 0 4328 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3311
timestamp 1569533753
transform 1 0 4328 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3312
timestamp 1569533753
transform 1 0 4328 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3313
timestamp 1569533753
transform 1 0 4200 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3314
timestamp 1569533753
transform 1 0 4328 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3315
timestamp 1569533753
transform 1 0 4328 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3316
timestamp 1569533753
transform 1 0 4072 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3317
timestamp 1569533753
transform 1 0 4200 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3318
timestamp 1569533753
transform 1 0 4072 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3319
timestamp 1569533753
transform 1 0 4328 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3320
timestamp 1569533753
transform 1 0 4264 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3321
timestamp 1569533753
transform 1 0 4072 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3322
timestamp 1569533753
transform 1 0 4200 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3323
timestamp 1569533753
transform 1 0 4200 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3324
timestamp 1569533753
transform 1 0 4136 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3325
timestamp 1569533753
transform 1 0 4264 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3326
timestamp 1569533753
transform 1 0 4136 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3327
timestamp 1569533753
transform 1 0 4136 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3328
timestamp 1569533753
transform 1 0 4072 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3329
timestamp 1569533753
transform 1 0 4200 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3330
timestamp 1569533753
transform 1 0 4328 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3331
timestamp 1569533753
transform 1 0 4072 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3332
timestamp 1569533753
transform 1 0 4072 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3333
timestamp 1569533753
transform 1 0 4264 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3334
timestamp 1569533753
transform 1 0 4328 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3335
timestamp 1569533753
transform 1 0 4264 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3336
timestamp 1569533753
transform 1 0 4200 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3337
timestamp 1569533753
transform 1 0 4136 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3338
timestamp 1569533753
transform 1 0 4328 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3339
timestamp 1569533753
transform 1 0 3816 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3340
timestamp 1569533753
transform 1 0 3880 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3341
timestamp 1569533753
transform 1 0 3944 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3342
timestamp 1569533753
transform 1 0 3944 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3343
timestamp 1569533753
transform 1 0 3880 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3344
timestamp 1569533753
transform 1 0 3752 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3345
timestamp 1569533753
transform 1 0 3944 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3346
timestamp 1569533753
transform 1 0 3944 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3347
timestamp 1569533753
transform 1 0 4008 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3348
timestamp 1569533753
transform 1 0 3816 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3349
timestamp 1569533753
transform 1 0 3752 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3350
timestamp 1569533753
transform 1 0 4008 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3351
timestamp 1569533753
transform 1 0 4008 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3352
timestamp 1569533753
transform 1 0 3816 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3353
timestamp 1569533753
transform 1 0 3880 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3354
timestamp 1569533753
transform 1 0 3752 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3355
timestamp 1569533753
transform 1 0 3752 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3356
timestamp 1569533753
transform 1 0 4008 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3357
timestamp 1569533753
transform 1 0 3816 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3358
timestamp 1569533753
transform 1 0 3880 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3359
timestamp 1569533753
transform 1 0 3752 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3360
timestamp 1569533753
transform 1 0 4008 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3361
timestamp 1569533753
transform 1 0 3880 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3362
timestamp 1569533753
transform 1 0 4008 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3363
timestamp 1569533753
transform 1 0 3752 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3364
timestamp 1569533753
transform 1 0 3880 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3365
timestamp 1569533753
transform 1 0 3880 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3366
timestamp 1569533753
transform 1 0 3944 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3367
timestamp 1569533753
transform 1 0 3944 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3368
timestamp 1569533753
transform 1 0 4008 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3369
timestamp 1569533753
transform 1 0 3816 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3370
timestamp 1569533753
transform 1 0 4008 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3371
timestamp 1569533753
transform 1 0 3880 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3372
timestamp 1569533753
transform 1 0 3944 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3373
timestamp 1569533753
transform 1 0 3816 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3374
timestamp 1569533753
transform 1 0 3816 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3375
timestamp 1569533753
transform 1 0 3816 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3376
timestamp 1569533753
transform 1 0 3752 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3377
timestamp 1569533753
transform 1 0 3752 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3378
timestamp 1569533753
transform 1 0 3944 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3379
timestamp 1569533753
transform 1 0 4072 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3380
timestamp 1569533753
transform 1 0 4264 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3381
timestamp 1569533753
transform 1 0 4264 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3382
timestamp 1569533753
transform 1 0 4200 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3383
timestamp 1569533753
transform 1 0 4072 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3384
timestamp 1569533753
transform 1 0 4136 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3385
timestamp 1569533753
transform 1 0 4328 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3386
timestamp 1569533753
transform 1 0 4072 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3387
timestamp 1569533753
transform 1 0 4200 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3388
timestamp 1569533753
transform 1 0 4136 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3389
timestamp 1569533753
transform 1 0 4328 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3390
timestamp 1569533753
transform 1 0 4328 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3391
timestamp 1569533753
transform 1 0 4264 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3392
timestamp 1569533753
transform 1 0 4328 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3393
timestamp 1569533753
transform 1 0 4200 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3394
timestamp 1569533753
transform 1 0 4136 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3395
timestamp 1569533753
transform 1 0 4200 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3396
timestamp 1569533753
transform 1 0 4072 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3397
timestamp 1569533753
transform 1 0 4264 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3398
timestamp 1569533753
transform 1 0 4136 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3399
timestamp 1569533753
transform 1 0 4264 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3400
timestamp 1569533753
transform 1 0 4072 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3401
timestamp 1569533753
transform 1 0 4328 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3402
timestamp 1569533753
transform 1 0 3944 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3403
timestamp 1569533753
transform 1 0 4200 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3404
timestamp 1569533753
transform 1 0 4136 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3405
timestamp 1569533753
transform 1 0 3752 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3406
timestamp 1569533753
transform 1 0 4008 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3407
timestamp 1569533753
transform 1 0 3816 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3408
timestamp 1569533753
transform 1 0 3880 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3409
timestamp 1569533753
transform 1 0 4776 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3410
timestamp 1569533753
transform 1 0 4840 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3411
timestamp 1569533753
transform 1 0 4712 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3412
timestamp 1569533753
transform 1 0 4840 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3413
timestamp 1569533753
transform 1 0 4712 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3414
timestamp 1569533753
transform 1 0 4776 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3415
timestamp 1569533753
transform 1 0 4904 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3416
timestamp 1569533753
transform 1 0 4776 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3417
timestamp 1569533753
transform 1 0 4904 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3418
timestamp 1569533753
transform 1 0 4840 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3419
timestamp 1569533753
transform 1 0 4840 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3420
timestamp 1569533753
transform 1 0 4712 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3421
timestamp 1569533753
transform 1 0 4904 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3422
timestamp 1569533753
transform 1 0 4776 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3423
timestamp 1569533753
transform 1 0 4712 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3424
timestamp 1569533753
transform 1 0 4904 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3425
timestamp 1569533753
transform 1 0 4648 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3426
timestamp 1569533753
transform 1 0 4584 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3427
timestamp 1569533753
transform 1 0 4456 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3428
timestamp 1569533753
transform 1 0 4456 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3429
timestamp 1569533753
transform 1 0 4648 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3430
timestamp 1569533753
transform 1 0 4456 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3431
timestamp 1569533753
transform 1 0 4456 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3432
timestamp 1569533753
transform 1 0 4584 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3433
timestamp 1569533753
transform 1 0 4584 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3434
timestamp 1569533753
transform 1 0 4520 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3435
timestamp 1569533753
transform 1 0 4520 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3436
timestamp 1569533753
transform 1 0 4392 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3437
timestamp 1569533753
transform 1 0 4520 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3438
timestamp 1569533753
transform 1 0 4520 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3439
timestamp 1569533753
transform 1 0 4392 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3440
timestamp 1569533753
transform 1 0 4392 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3441
timestamp 1569533753
transform 1 0 4392 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3442
timestamp 1569533753
transform 1 0 4584 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3443
timestamp 1569533753
transform 1 0 4648 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3444
timestamp 1569533753
transform 1 0 4648 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3445
timestamp 1569533753
transform 1 0 4392 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3446
timestamp 1569533753
transform 1 0 4392 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3447
timestamp 1569533753
transform 1 0 4648 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3448
timestamp 1569533753
transform 1 0 4520 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3449
timestamp 1569533753
transform 1 0 4584 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3450
timestamp 1569533753
transform 1 0 4520 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3451
timestamp 1569533753
transform 1 0 4392 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3452
timestamp 1569533753
transform 1 0 4456 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3453
timestamp 1569533753
transform 1 0 4520 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3454
timestamp 1569533753
transform 1 0 4392 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3455
timestamp 1569533753
transform 1 0 4456 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3456
timestamp 1569533753
transform 1 0 4648 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3457
timestamp 1569533753
transform 1 0 4456 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3458
timestamp 1569533753
transform 1 0 4584 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3459
timestamp 1569533753
transform 1 0 4648 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3460
timestamp 1569533753
transform 1 0 4584 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3461
timestamp 1569533753
transform 1 0 4456 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3462
timestamp 1569533753
transform 1 0 4648 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3463
timestamp 1569533753
transform 1 0 4584 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3464
timestamp 1569533753
transform 1 0 4520 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3465
timestamp 1569533753
transform 1 0 4712 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3466
timestamp 1569533753
transform 1 0 4904 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3467
timestamp 1569533753
transform 1 0 4776 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3468
timestamp 1569533753
transform 1 0 4840 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3469
timestamp 1569533753
transform 1 0 4712 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3470
timestamp 1569533753
transform 1 0 4840 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3471
timestamp 1569533753
transform 1 0 4712 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3472
timestamp 1569533753
transform 1 0 4904 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3473
timestamp 1569533753
transform 1 0 4712 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3474
timestamp 1569533753
transform 1 0 4904 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3475
timestamp 1569533753
transform 1 0 4904 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3476
timestamp 1569533753
transform 1 0 4840 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3477
timestamp 1569533753
transform 1 0 4776 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3478
timestamp 1569533753
transform 1 0 4840 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3479
timestamp 1569533753
transform 1 0 4776 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3480
timestamp 1569533753
transform 1 0 4776 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3481
timestamp 1569533753
transform 1 0 4840 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3482
timestamp 1569533753
transform 1 0 4712 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3483
timestamp 1569533753
transform 1 0 4392 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3484
timestamp 1569533753
transform 1 0 4776 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3485
timestamp 1569533753
transform 1 0 4456 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3486
timestamp 1569533753
transform 1 0 4520 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3487
timestamp 1569533753
transform 1 0 4904 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3488
timestamp 1569533753
transform 1 0 4584 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3489
timestamp 1569533753
transform 1 0 4648 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3490
timestamp 1569533753
transform 1 0 3624 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3491
timestamp 1569533753
transform 1 0 3496 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3492
timestamp 1569533753
transform 1 0 3496 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3493
timestamp 1569533753
transform 1 0 3496 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3494
timestamp 1569533753
transform 1 0 3624 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3495
timestamp 1569533753
transform 1 0 3560 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3496
timestamp 1569533753
transform 1 0 3560 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3497
timestamp 1569533753
transform 1 0 3624 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3498
timestamp 1569533753
transform 1 0 3624 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3499
timestamp 1569533753
transform 1 0 3560 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3500
timestamp 1569533753
transform 1 0 3688 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3501
timestamp 1569533753
transform 1 0 3688 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3502
timestamp 1569533753
transform 1 0 3688 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3503
timestamp 1569533753
transform 1 0 3560 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3504
timestamp 1569533753
transform 1 0 3688 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3505
timestamp 1569533753
transform 1 0 3688 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3506
timestamp 1569533753
transform 1 0 3560 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3507
timestamp 1569533753
transform 1 0 3496 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3508
timestamp 1569533753
transform 1 0 3624 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3509
timestamp 1569533753
transform 1 0 3496 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3510
timestamp 1569533753
transform 1 0 3368 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3511
timestamp 1569533753
transform 1 0 3368 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3512
timestamp 1569533753
transform 1 0 3304 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3513
timestamp 1569533753
transform 1 0 3176 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3514
timestamp 1569533753
transform 1 0 3176 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3515
timestamp 1569533753
transform 1 0 3176 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3516
timestamp 1569533753
transform 1 0 3176 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3517
timestamp 1569533753
transform 1 0 3176 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3518
timestamp 1569533753
transform 1 0 3304 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3519
timestamp 1569533753
transform 1 0 3240 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3520
timestamp 1569533753
transform 1 0 3240 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3521
timestamp 1569533753
transform 1 0 3240 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3522
timestamp 1569533753
transform 1 0 3240 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3523
timestamp 1569533753
transform 1 0 3240 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3524
timestamp 1569533753
transform 1 0 3304 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3525
timestamp 1569533753
transform 1 0 3304 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3526
timestamp 1569533753
transform 1 0 3304 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3527
timestamp 1569533753
transform 1 0 3368 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3528
timestamp 1569533753
transform 1 0 3368 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3529
timestamp 1569533753
transform 1 0 3368 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3530
timestamp 1569533753
transform 1 0 3176 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3531
timestamp 1569533753
transform 1 0 3240 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3532
timestamp 1569533753
transform 1 0 3304 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3533
timestamp 1569533753
transform 1 0 3368 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3534
timestamp 1569533753
transform 1 0 3304 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3535
timestamp 1569533753
transform 1 0 3304 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3536
timestamp 1569533753
transform 1 0 3176 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3537
timestamp 1569533753
transform 1 0 3368 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3538
timestamp 1569533753
transform 1 0 3368 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3539
timestamp 1569533753
transform 1 0 3368 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3540
timestamp 1569533753
transform 1 0 3176 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3541
timestamp 1569533753
transform 1 0 3368 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3542
timestamp 1569533753
transform 1 0 3304 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3543
timestamp 1569533753
transform 1 0 3240 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3544
timestamp 1569533753
transform 1 0 3240 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3545
timestamp 1569533753
transform 1 0 3240 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3546
timestamp 1569533753
transform 1 0 3240 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3547
timestamp 1569533753
transform 1 0 3304 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3548
timestamp 1569533753
transform 1 0 3176 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3549
timestamp 1569533753
transform 1 0 3176 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3550
timestamp 1569533753
transform 1 0 3688 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3551
timestamp 1569533753
transform 1 0 3624 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3552
timestamp 1569533753
transform 1 0 3688 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3553
timestamp 1569533753
transform 1 0 3496 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3554
timestamp 1569533753
transform 1 0 3496 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3555
timestamp 1569533753
transform 1 0 3688 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3556
timestamp 1569533753
transform 1 0 3496 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3557
timestamp 1569533753
transform 1 0 3496 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3558
timestamp 1569533753
transform 1 0 3688 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3559
timestamp 1569533753
transform 1 0 3688 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3560
timestamp 1569533753
transform 1 0 3560 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3561
timestamp 1569533753
transform 1 0 3496 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3562
timestamp 1569533753
transform 1 0 3560 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3563
timestamp 1569533753
transform 1 0 3560 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3564
timestamp 1569533753
transform 1 0 3560 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3565
timestamp 1569533753
transform 1 0 3560 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3566
timestamp 1569533753
transform 1 0 3624 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3567
timestamp 1569533753
transform 1 0 3624 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3568
timestamp 1569533753
transform 1 0 3624 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3569
timestamp 1569533753
transform 1 0 3624 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3570
timestamp 1569533753
transform 1 0 3432 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3571
timestamp 1569533753
transform 1 0 3432 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3572
timestamp 1569533753
transform 1 0 3432 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3573
timestamp 1569533753
transform 1 0 3432 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3574
timestamp 1569533753
transform 1 0 3432 0 1 2536
box -8 -8 8 8
use VIA2$3  VIA2$3_3575
timestamp 1569533753
transform 1 0 3432 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3576
timestamp 1569533753
transform 1 0 3432 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3577
timestamp 1569533753
transform 1 0 3432 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3578
timestamp 1569533753
transform 1 0 3432 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3579
timestamp 1569533753
transform 1 0 3432 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3580
timestamp 1569533753
transform 1 0 3048 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3581
timestamp 1569533753
transform 1 0 3048 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3582
timestamp 1569533753
transform 1 0 3112 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3583
timestamp 1569533753
transform 1 0 2600 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3584
timestamp 1569533753
transform 1 0 2856 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3585
timestamp 1569533753
transform 1 0 2856 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3586
timestamp 1569533753
transform 1 0 2856 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3587
timestamp 1569533753
transform 1 0 2856 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3588
timestamp 1569533753
transform 1 0 2792 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3589
timestamp 1569533753
transform 1 0 2792 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3590
timestamp 1569533753
transform 1 0 2792 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3591
timestamp 1569533753
transform 1 0 2792 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3592
timestamp 1569533753
transform 1 0 3112 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3593
timestamp 1569533753
transform 1 0 3112 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3594
timestamp 1569533753
transform 1 0 2920 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3595
timestamp 1569533753
transform 1 0 2920 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3596
timestamp 1569533753
transform 1 0 2920 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3597
timestamp 1569533753
transform 1 0 2920 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3598
timestamp 1569533753
transform 1 0 3112 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3599
timestamp 1569533753
transform 1 0 3048 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3600
timestamp 1569533753
transform 1 0 3048 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3601
timestamp 1569533753
transform 1 0 3048 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3602
timestamp 1569533753
transform 1 0 3048 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3603
timestamp 1569533753
transform 1 0 3112 0 1 2600
box -8 -8 8 8
use VIA2$3  VIA2$3_3604
timestamp 1569533753
transform 1 0 2664 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3605
timestamp 1569533753
transform 1 0 2664 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3606
timestamp 1569533753
transform 1 0 3112 0 1 2664
box -8 -8 8 8
use VIA2$3  VIA2$3_3607
timestamp 1569533753
transform 1 0 3112 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3608
timestamp 1569533753
transform 1 0 3112 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3609
timestamp 1569533753
transform 1 0 3112 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3610
timestamp 1569533753
transform 1 0 2856 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3611
timestamp 1569533753
transform 1 0 2920 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3612
timestamp 1569533753
transform 1 0 2920 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3613
timestamp 1569533753
transform 1 0 2984 0 1 2728
box -8 -8 8 8
use VIA2$3  VIA2$3_3614
timestamp 1569533753
transform 1 0 2984 0 1 2792
box -8 -8 8 8
use VIA2$3  VIA2$3_3615
timestamp 1569533753
transform 1 0 2984 0 1 2856
box -8 -8 8 8
use VIA2$3  VIA2$3_3616
timestamp 1569533753
transform 1 0 2728 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3617
timestamp 1569533753
transform 1 0 2728 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3618
timestamp 1569533753
transform 1 0 2984 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3619
timestamp 1569533753
transform 1 0 2984 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3620
timestamp 1569533753
transform 1 0 2984 0 1 3048
box -8 -8 8 8
use VIA2$3  VIA2$3_3621
timestamp 1569533753
transform 1 0 2984 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3622
timestamp 1569533753
transform 1 0 2728 0 1 3112
box -8 -8 8 8
use VIA2$3  VIA2$3_3623
timestamp 1569533753
transform 1 0 3048 0 1 2920
box -8 -8 8 8
use VIA2$3  VIA2$3_3624
timestamp 1569533753
transform 1 0 3048 0 1 2984
box -8 -8 8 8
use VIA2$3  VIA2$3_3625
timestamp 1569533753
transform 1 0 2984 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3626
timestamp 1569533753
transform 1 0 2984 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3627
timestamp 1569533753
transform 1 0 2920 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3628
timestamp 1569533753
transform 1 0 3112 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3629
timestamp 1569533753
transform 1 0 3048 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3630
timestamp 1569533753
transform 1 0 3112 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3631
timestamp 1569533753
transform 1 0 2920 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3632
timestamp 1569533753
transform 1 0 2920 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3633
timestamp 1569533753
transform 1 0 3048 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3634
timestamp 1569533753
transform 1 0 2856 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3635
timestamp 1569533753
transform 1 0 3112 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3636
timestamp 1569533753
transform 1 0 2920 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3637
timestamp 1569533753
transform 1 0 3048 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3638
timestamp 1569533753
transform 1 0 2856 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3639
timestamp 1569533753
transform 1 0 2856 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3640
timestamp 1569533753
transform 1 0 2856 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3641
timestamp 1569533753
transform 1 0 2984 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3642
timestamp 1569533753
transform 1 0 3048 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3643
timestamp 1569533753
transform 1 0 3112 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3644
timestamp 1569533753
transform 1 0 2984 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3645
timestamp 1569533753
transform 1 0 2600 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3646
timestamp 1569533753
transform 1 0 2600 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3647
timestamp 1569533753
transform 1 0 2792 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3648
timestamp 1569533753
transform 1 0 2600 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3649
timestamp 1569533753
transform 1 0 2536 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3650
timestamp 1569533753
transform 1 0 2536 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3651
timestamp 1569533753
transform 1 0 2728 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3652
timestamp 1569533753
transform 1 0 2792 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3653
timestamp 1569533753
transform 1 0 2728 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3654
timestamp 1569533753
transform 1 0 2600 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3655
timestamp 1569533753
transform 1 0 2536 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3656
timestamp 1569533753
transform 1 0 2728 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3657
timestamp 1569533753
transform 1 0 2664 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3658
timestamp 1569533753
transform 1 0 2792 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3659
timestamp 1569533753
transform 1 0 2664 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3660
timestamp 1569533753
transform 1 0 2536 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3661
timestamp 1569533753
transform 1 0 2728 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3662
timestamp 1569533753
transform 1 0 2664 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3663
timestamp 1569533753
transform 1 0 2792 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3664
timestamp 1569533753
transform 1 0 2664 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3665
timestamp 1569533753
transform 1 0 2600 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3666
timestamp 1569533753
transform 1 0 2536 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3667
timestamp 1569533753
transform 1 0 2728 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3668
timestamp 1569533753
transform 1 0 2728 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3669
timestamp 1569533753
transform 1 0 2792 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3670
timestamp 1569533753
transform 1 0 2536 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3671
timestamp 1569533753
transform 1 0 2728 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3672
timestamp 1569533753
transform 1 0 2792 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3673
timestamp 1569533753
transform 1 0 2728 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3674
timestamp 1569533753
transform 1 0 2792 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3675
timestamp 1569533753
transform 1 0 2792 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3676
timestamp 1569533753
transform 1 0 2600 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3677
timestamp 1569533753
transform 1 0 2664 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3678
timestamp 1569533753
transform 1 0 2664 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3679
timestamp 1569533753
transform 1 0 2664 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3680
timestamp 1569533753
transform 1 0 2536 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3681
timestamp 1569533753
transform 1 0 2600 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3682
timestamp 1569533753
transform 1 0 2664 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3683
timestamp 1569533753
transform 1 0 2536 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3684
timestamp 1569533753
transform 1 0 2600 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3685
timestamp 1569533753
transform 1 0 2856 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3686
timestamp 1569533753
transform 1 0 2984 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3687
timestamp 1569533753
transform 1 0 2984 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3688
timestamp 1569533753
transform 1 0 2984 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3689
timestamp 1569533753
transform 1 0 2856 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3690
timestamp 1569533753
transform 1 0 2856 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3691
timestamp 1569533753
transform 1 0 3048 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3692
timestamp 1569533753
transform 1 0 2984 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3693
timestamp 1569533753
transform 1 0 3048 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3694
timestamp 1569533753
transform 1 0 2920 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3695
timestamp 1569533753
transform 1 0 2920 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3696
timestamp 1569533753
transform 1 0 3112 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3697
timestamp 1569533753
transform 1 0 2920 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3698
timestamp 1569533753
transform 1 0 3048 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3699
timestamp 1569533753
transform 1 0 3048 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3700
timestamp 1569533753
transform 1 0 3112 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3701
timestamp 1569533753
transform 1 0 3112 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3702
timestamp 1569533753
transform 1 0 2920 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3703
timestamp 1569533753
transform 1 0 3112 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3704
timestamp 1569533753
transform 1 0 2856 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3705
timestamp 1569533753
transform 1 0 2984 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3706
timestamp 1569533753
transform 1 0 3048 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3707
timestamp 1569533753
transform 1 0 2728 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3708
timestamp 1569533753
transform 1 0 2600 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3709
timestamp 1569533753
transform 1 0 2792 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3710
timestamp 1569533753
transform 1 0 2664 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3711
timestamp 1569533753
transform 1 0 3112 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3712
timestamp 1569533753
transform 1 0 2856 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3713
timestamp 1569533753
transform 1 0 2920 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3714
timestamp 1569533753
transform 1 0 2536 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3715
timestamp 1569533753
transform 1 0 3688 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3716
timestamp 1569533753
transform 1 0 3496 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3717
timestamp 1569533753
transform 1 0 3496 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3718
timestamp 1569533753
transform 1 0 3496 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3719
timestamp 1569533753
transform 1 0 3496 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3720
timestamp 1569533753
transform 1 0 3688 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3721
timestamp 1569533753
transform 1 0 3560 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3722
timestamp 1569533753
transform 1 0 3560 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3723
timestamp 1569533753
transform 1 0 3560 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3724
timestamp 1569533753
transform 1 0 3560 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3725
timestamp 1569533753
transform 1 0 3688 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3726
timestamp 1569533753
transform 1 0 3624 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3727
timestamp 1569533753
transform 1 0 3624 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3728
timestamp 1569533753
transform 1 0 3688 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3729
timestamp 1569533753
transform 1 0 3624 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3730
timestamp 1569533753
transform 1 0 3624 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3731
timestamp 1569533753
transform 1 0 3304 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3732
timestamp 1569533753
transform 1 0 3176 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3733
timestamp 1569533753
transform 1 0 3176 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3734
timestamp 1569533753
transform 1 0 3304 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3735
timestamp 1569533753
transform 1 0 3304 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3736
timestamp 1569533753
transform 1 0 3304 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3737
timestamp 1569533753
transform 1 0 3176 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3738
timestamp 1569533753
transform 1 0 3176 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3739
timestamp 1569533753
transform 1 0 3240 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3740
timestamp 1569533753
transform 1 0 3240 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3741
timestamp 1569533753
transform 1 0 3240 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3742
timestamp 1569533753
transform 1 0 3240 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3743
timestamp 1569533753
transform 1 0 3368 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3744
timestamp 1569533753
transform 1 0 3368 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3745
timestamp 1569533753
transform 1 0 3368 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3746
timestamp 1569533753
transform 1 0 3368 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3747
timestamp 1569533753
transform 1 0 3176 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3748
timestamp 1569533753
transform 1 0 3176 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3749
timestamp 1569533753
transform 1 0 3368 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3750
timestamp 1569533753
transform 1 0 3240 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3751
timestamp 1569533753
transform 1 0 3240 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3752
timestamp 1569533753
transform 1 0 3240 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3753
timestamp 1569533753
transform 1 0 3240 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3754
timestamp 1569533753
transform 1 0 3368 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3755
timestamp 1569533753
transform 1 0 3368 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3756
timestamp 1569533753
transform 1 0 3176 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3757
timestamp 1569533753
transform 1 0 3176 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3758
timestamp 1569533753
transform 1 0 3304 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3759
timestamp 1569533753
transform 1 0 3304 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3760
timestamp 1569533753
transform 1 0 3304 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3761
timestamp 1569533753
transform 1 0 3304 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3762
timestamp 1569533753
transform 1 0 3368 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3763
timestamp 1569533753
transform 1 0 3688 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3764
timestamp 1569533753
transform 1 0 3688 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3765
timestamp 1569533753
transform 1 0 3688 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3766
timestamp 1569533753
transform 1 0 3688 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3767
timestamp 1569533753
transform 1 0 3496 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3768
timestamp 1569533753
transform 1 0 3496 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3769
timestamp 1569533753
transform 1 0 3560 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3770
timestamp 1569533753
transform 1 0 3560 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3771
timestamp 1569533753
transform 1 0 3624 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3772
timestamp 1569533753
transform 1 0 3624 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3773
timestamp 1569533753
transform 1 0 3496 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3774
timestamp 1569533753
transform 1 0 3496 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3775
timestamp 1569533753
transform 1 0 3624 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3776
timestamp 1569533753
transform 1 0 3624 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3777
timestamp 1569533753
transform 1 0 3560 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3778
timestamp 1569533753
transform 1 0 3560 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3779
timestamp 1569533753
transform 1 0 3240 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3780
timestamp 1569533753
transform 1 0 3304 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3781
timestamp 1569533753
transform 1 0 3432 0 1 3560
box -8 -8 8 8
use VIA2$3  VIA2$3_3782
timestamp 1569533753
transform 1 0 3496 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3783
timestamp 1569533753
transform 1 0 3560 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3784
timestamp 1569533753
transform 1 0 3624 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3785
timestamp 1569533753
transform 1 0 3432 0 1 3624
box -8 -8 8 8
use VIA2$3  VIA2$3_3786
timestamp 1569533753
transform 1 0 3432 0 1 3688
box -8 -8 8 8
use VIA2$3  VIA2$3_3787
timestamp 1569533753
transform 1 0 3368 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3788
timestamp 1569533753
transform 1 0 3432 0 1 3176
box -8 -8 8 8
use VIA2$3  VIA2$3_3789
timestamp 1569533753
transform 1 0 3432 0 1 3240
box -8 -8 8 8
use VIA2$3  VIA2$3_3790
timestamp 1569533753
transform 1 0 3432 0 1 3304
box -8 -8 8 8
use VIA2$3  VIA2$3_3791
timestamp 1569533753
transform 1 0 3432 0 1 3368
box -8 -8 8 8
use VIA2$3  VIA2$3_3792
timestamp 1569533753
transform 1 0 3432 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3793
timestamp 1569533753
transform 1 0 3432 0 1 3496
box -8 -8 8 8
use VIA2$3  VIA2$3_3794
timestamp 1569533753
transform 1 0 3688 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3795
timestamp 1569533753
transform 1 0 3176 0 1 3432
box -8 -8 8 8
use VIA2$3  VIA2$3_3796
timestamp 1569533753
transform 1 0 3688 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3797
timestamp 1569533753
transform 1 0 3624 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3798
timestamp 1569533753
transform 1 0 3560 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3799
timestamp 1569533753
transform 1 0 3496 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3800
timestamp 1569533753
transform 1 0 3688 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3801
timestamp 1569533753
transform 1 0 3624 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3802
timestamp 1569533753
transform 1 0 3688 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3803
timestamp 1569533753
transform 1 0 3624 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3804
timestamp 1569533753
transform 1 0 3496 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3805
timestamp 1569533753
transform 1 0 3560 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3806
timestamp 1569533753
transform 1 0 3496 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3807
timestamp 1569533753
transform 1 0 3560 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3808
timestamp 1569533753
transform 1 0 3624 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3809
timestamp 1569533753
transform 1 0 3560 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3810
timestamp 1569533753
transform 1 0 3688 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3811
timestamp 1569533753
transform 1 0 3560 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3812
timestamp 1569533753
transform 1 0 3688 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3813
timestamp 1569533753
transform 1 0 3624 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3814
timestamp 1569533753
transform 1 0 3496 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3815
timestamp 1569533753
transform 1 0 3496 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3816
timestamp 1569533753
transform 1 0 3368 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3817
timestamp 1569533753
transform 1 0 3368 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3818
timestamp 1569533753
transform 1 0 3240 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3819
timestamp 1569533753
transform 1 0 3176 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3820
timestamp 1569533753
transform 1 0 3240 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3821
timestamp 1569533753
transform 1 0 3240 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3822
timestamp 1569533753
transform 1 0 3304 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3823
timestamp 1569533753
transform 1 0 3176 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3824
timestamp 1569533753
transform 1 0 3368 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3825
timestamp 1569533753
transform 1 0 3304 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3826
timestamp 1569533753
transform 1 0 3304 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3827
timestamp 1569533753
transform 1 0 3304 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3828
timestamp 1569533753
transform 1 0 3240 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3829
timestamp 1569533753
transform 1 0 3176 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3830
timestamp 1569533753
transform 1 0 3176 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3831
timestamp 1569533753
transform 1 0 3368 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3832
timestamp 1569533753
transform 1 0 3304 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3833
timestamp 1569533753
transform 1 0 3368 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3834
timestamp 1569533753
transform 1 0 3176 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3835
timestamp 1569533753
transform 1 0 3240 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3836
timestamp 1569533753
transform 1 0 3304 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3837
timestamp 1569533753
transform 1 0 3240 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3838
timestamp 1569533753
transform 1 0 3176 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3839
timestamp 1569533753
transform 1 0 3240 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3840
timestamp 1569533753
transform 1 0 3176 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3841
timestamp 1569533753
transform 1 0 3176 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3842
timestamp 1569533753
transform 1 0 3368 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3843
timestamp 1569533753
transform 1 0 3304 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3844
timestamp 1569533753
transform 1 0 3240 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3845
timestamp 1569533753
transform 1 0 3240 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3846
timestamp 1569533753
transform 1 0 3368 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3847
timestamp 1569533753
transform 1 0 3176 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3848
timestamp 1569533753
transform 1 0 3304 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3849
timestamp 1569533753
transform 1 0 3368 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3850
timestamp 1569533753
transform 1 0 3304 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3851
timestamp 1569533753
transform 1 0 3304 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3852
timestamp 1569533753
transform 1 0 3240 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3853
timestamp 1569533753
transform 1 0 3368 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3854
timestamp 1569533753
transform 1 0 3176 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3855
timestamp 1569533753
transform 1 0 3368 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3856
timestamp 1569533753
transform 1 0 3624 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3857
timestamp 1569533753
transform 1 0 3624 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3858
timestamp 1569533753
transform 1 0 3688 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3859
timestamp 1569533753
transform 1 0 3496 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3860
timestamp 1569533753
transform 1 0 3624 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3861
timestamp 1569533753
transform 1 0 3688 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3862
timestamp 1569533753
transform 1 0 3560 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3863
timestamp 1569533753
transform 1 0 3688 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3864
timestamp 1569533753
transform 1 0 3688 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3865
timestamp 1569533753
transform 1 0 3496 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3866
timestamp 1569533753
transform 1 0 3688 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3867
timestamp 1569533753
transform 1 0 3624 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3868
timestamp 1569533753
transform 1 0 3496 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3869
timestamp 1569533753
transform 1 0 3496 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3870
timestamp 1569533753
transform 1 0 3560 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3871
timestamp 1569533753
transform 1 0 3560 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3872
timestamp 1569533753
transform 1 0 3496 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3873
timestamp 1569533753
transform 1 0 3560 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3874
timestamp 1569533753
transform 1 0 3560 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3875
timestamp 1569533753
transform 1 0 3624 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3876
timestamp 1569533753
transform 1 0 3432 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3877
timestamp 1569533753
transform 1 0 3432 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3878
timestamp 1569533753
transform 1 0 3432 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3879
timestamp 1569533753
transform 1 0 3432 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3880
timestamp 1569533753
transform 1 0 3432 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3881
timestamp 1569533753
transform 1 0 3432 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3882
timestamp 1569533753
transform 1 0 3432 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3883
timestamp 1569533753
transform 1 0 3432 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3884
timestamp 1569533753
transform 1 0 3432 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3885
timestamp 1569533753
transform 1 0 3432 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3886
timestamp 1569533753
transform 1 0 2984 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3887
timestamp 1569533753
transform 1 0 3112 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3888
timestamp 1569533753
transform 1 0 2984 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3889
timestamp 1569533753
transform 1 0 2920 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3890
timestamp 1569533753
transform 1 0 3112 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3891
timestamp 1569533753
transform 1 0 2920 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3892
timestamp 1569533753
transform 1 0 2856 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3893
timestamp 1569533753
transform 1 0 2984 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3894
timestamp 1569533753
transform 1 0 2984 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3895
timestamp 1569533753
transform 1 0 2984 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3896
timestamp 1569533753
transform 1 0 3112 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3897
timestamp 1569533753
transform 1 0 2856 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3898
timestamp 1569533753
transform 1 0 3048 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3899
timestamp 1569533753
transform 1 0 2856 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3900
timestamp 1569533753
transform 1 0 2920 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3901
timestamp 1569533753
transform 1 0 2920 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3902
timestamp 1569533753
transform 1 0 3048 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3903
timestamp 1569533753
transform 1 0 3112 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3904
timestamp 1569533753
transform 1 0 2856 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3905
timestamp 1569533753
transform 1 0 3048 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3906
timestamp 1569533753
transform 1 0 3048 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3907
timestamp 1569533753
transform 1 0 3112 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3908
timestamp 1569533753
transform 1 0 3048 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3909
timestamp 1569533753
transform 1 0 2920 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3910
timestamp 1569533753
transform 1 0 2856 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3911
timestamp 1569533753
transform 1 0 2664 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3912
timestamp 1569533753
transform 1 0 2536 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3913
timestamp 1569533753
transform 1 0 2728 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3914
timestamp 1569533753
transform 1 0 2536 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3915
timestamp 1569533753
transform 1 0 2728 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3916
timestamp 1569533753
transform 1 0 2536 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3917
timestamp 1569533753
transform 1 0 2728 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3918
timestamp 1569533753
transform 1 0 2600 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3919
timestamp 1569533753
transform 1 0 2600 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3920
timestamp 1569533753
transform 1 0 2664 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3921
timestamp 1569533753
transform 1 0 2600 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3922
timestamp 1569533753
transform 1 0 2664 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3923
timestamp 1569533753
transform 1 0 2728 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3924
timestamp 1569533753
transform 1 0 2728 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3925
timestamp 1569533753
transform 1 0 2600 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3926
timestamp 1569533753
transform 1 0 2664 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3927
timestamp 1569533753
transform 1 0 2792 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3928
timestamp 1569533753
transform 1 0 2600 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3929
timestamp 1569533753
transform 1 0 2792 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3930
timestamp 1569533753
transform 1 0 2536 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3931
timestamp 1569533753
transform 1 0 2792 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_3932
timestamp 1569533753
transform 1 0 2664 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_3933
timestamp 1569533753
transform 1 0 2536 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_3934
timestamp 1569533753
transform 1 0 2792 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_3935
timestamp 1569533753
transform 1 0 2792 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_3936
timestamp 1569533753
transform 1 0 2792 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3937
timestamp 1569533753
transform 1 0 2664 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3938
timestamp 1569533753
transform 1 0 2536 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3939
timestamp 1569533753
transform 1 0 2536 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3940
timestamp 1569533753
transform 1 0 2600 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3941
timestamp 1569533753
transform 1 0 2600 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3942
timestamp 1569533753
transform 1 0 2728 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3943
timestamp 1569533753
transform 1 0 2600 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3944
timestamp 1569533753
transform 1 0 2664 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3945
timestamp 1569533753
transform 1 0 2728 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3946
timestamp 1569533753
transform 1 0 2792 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3947
timestamp 1569533753
transform 1 0 2792 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3948
timestamp 1569533753
transform 1 0 2728 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3949
timestamp 1569533753
transform 1 0 2664 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3950
timestamp 1569533753
transform 1 0 2792 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3951
timestamp 1569533753
transform 1 0 2536 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3952
timestamp 1569533753
transform 1 0 2792 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3953
timestamp 1569533753
transform 1 0 2536 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3954
timestamp 1569533753
transform 1 0 2536 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3955
timestamp 1569533753
transform 1 0 2728 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3956
timestamp 1569533753
transform 1 0 2600 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3957
timestamp 1569533753
transform 1 0 2664 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3958
timestamp 1569533753
transform 1 0 2664 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3959
timestamp 1569533753
transform 1 0 2728 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3960
timestamp 1569533753
transform 1 0 2600 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3961
timestamp 1569533753
transform 1 0 2856 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3962
timestamp 1569533753
transform 1 0 2984 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3963
timestamp 1569533753
transform 1 0 2984 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3964
timestamp 1569533753
transform 1 0 3112 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3965
timestamp 1569533753
transform 1 0 3112 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3966
timestamp 1569533753
transform 1 0 2984 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3967
timestamp 1569533753
transform 1 0 2920 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3968
timestamp 1569533753
transform 1 0 2920 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3969
timestamp 1569533753
transform 1 0 3048 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3970
timestamp 1569533753
transform 1 0 3048 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3971
timestamp 1569533753
transform 1 0 2920 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3972
timestamp 1569533753
transform 1 0 2920 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3973
timestamp 1569533753
transform 1 0 2920 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3974
timestamp 1569533753
transform 1 0 2984 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3975
timestamp 1569533753
transform 1 0 2984 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_3976
timestamp 1569533753
transform 1 0 3048 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3977
timestamp 1569533753
transform 1 0 3048 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3978
timestamp 1569533753
transform 1 0 3048 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3979
timestamp 1569533753
transform 1 0 3112 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3980
timestamp 1569533753
transform 1 0 3112 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3981
timestamp 1569533753
transform 1 0 3112 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3982
timestamp 1569533753
transform 1 0 2856 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_3983
timestamp 1569533753
transform 1 0 2856 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_3984
timestamp 1569533753
transform 1 0 2856 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_3985
timestamp 1569533753
transform 1 0 2856 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_3986
timestamp 1569533753
transform 1 0 2856 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3987
timestamp 1569533753
transform 1 0 3112 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3988
timestamp 1569533753
transform 1 0 2920 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3989
timestamp 1569533753
transform 1 0 3048 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3990
timestamp 1569533753
transform 1 0 2920 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_3991
timestamp 1569533753
transform 1 0 3048 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3992
timestamp 1569533753
transform 1 0 3112 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3993
timestamp 1569533753
transform 1 0 3048 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_3994
timestamp 1569533753
transform 1 0 2856 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_3995
timestamp 1569533753
transform 1 0 2920 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3996
timestamp 1569533753
transform 1 0 2984 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_3997
timestamp 1569533753
transform 1 0 2856 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3998
timestamp 1569533753
transform 1 0 3112 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_3999
timestamp 1569533753
transform 1 0 2984 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4000
timestamp 1569533753
transform 1 0 2920 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4001
timestamp 1569533753
transform 1 0 3048 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4002
timestamp 1569533753
transform 1 0 2920 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4003
timestamp 1569533753
transform 1 0 2984 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4004
timestamp 1569533753
transform 1 0 2856 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4005
timestamp 1569533753
transform 1 0 3048 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4006
timestamp 1569533753
transform 1 0 2984 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4007
timestamp 1569533753
transform 1 0 2856 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4008
timestamp 1569533753
transform 1 0 3112 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4009
timestamp 1569533753
transform 1 0 2984 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4010
timestamp 1569533753
transform 1 0 3112 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4011
timestamp 1569533753
transform 1 0 2536 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4012
timestamp 1569533753
transform 1 0 2600 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4013
timestamp 1569533753
transform 1 0 2664 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4014
timestamp 1569533753
transform 1 0 2664 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4015
timestamp 1569533753
transform 1 0 2536 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4016
timestamp 1569533753
transform 1 0 2728 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4017
timestamp 1569533753
transform 1 0 2664 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4018
timestamp 1569533753
transform 1 0 2536 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4019
timestamp 1569533753
transform 1 0 2728 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4020
timestamp 1569533753
transform 1 0 2664 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4021
timestamp 1569533753
transform 1 0 2536 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4022
timestamp 1569533753
transform 1 0 2664 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4023
timestamp 1569533753
transform 1 0 2536 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4024
timestamp 1569533753
transform 1 0 2792 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4025
timestamp 1569533753
transform 1 0 2600 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4026
timestamp 1569533753
transform 1 0 2728 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4027
timestamp 1569533753
transform 1 0 2728 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4028
timestamp 1569533753
transform 1 0 2600 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4029
timestamp 1569533753
transform 1 0 2792 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4030
timestamp 1569533753
transform 1 0 2792 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4031
timestamp 1569533753
transform 1 0 2728 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4032
timestamp 1569533753
transform 1 0 2600 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4033
timestamp 1569533753
transform 1 0 2792 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4034
timestamp 1569533753
transform 1 0 2600 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4035
timestamp 1569533753
transform 1 0 2792 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4036
timestamp 1569533753
transform 1 0 2536 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4037
timestamp 1569533753
transform 1 0 2792 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4038
timestamp 1569533753
transform 1 0 2664 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4039
timestamp 1569533753
transform 1 0 2664 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4040
timestamp 1569533753
transform 1 0 2728 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4041
timestamp 1569533753
transform 1 0 2664 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4042
timestamp 1569533753
transform 1 0 2728 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4043
timestamp 1569533753
transform 1 0 2600 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4044
timestamp 1569533753
transform 1 0 2536 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4045
timestamp 1569533753
transform 1 0 2600 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4046
timestamp 1569533753
transform 1 0 2664 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4047
timestamp 1569533753
transform 1 0 2792 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4048
timestamp 1569533753
transform 1 0 2536 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4049
timestamp 1569533753
transform 1 0 2728 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4050
timestamp 1569533753
transform 1 0 2536 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4051
timestamp 1569533753
transform 1 0 2728 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4052
timestamp 1569533753
transform 1 0 2792 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4053
timestamp 1569533753
transform 1 0 2600 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4054
timestamp 1569533753
transform 1 0 2600 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4055
timestamp 1569533753
transform 1 0 2792 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4056
timestamp 1569533753
transform 1 0 3112 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4057
timestamp 1569533753
transform 1 0 2920 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4058
timestamp 1569533753
transform 1 0 2920 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4059
timestamp 1569533753
transform 1 0 2984 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4060
timestamp 1569533753
transform 1 0 2984 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4061
timestamp 1569533753
transform 1 0 2984 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4062
timestamp 1569533753
transform 1 0 3048 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4063
timestamp 1569533753
transform 1 0 3112 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4064
timestamp 1569533753
transform 1 0 3112 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4065
timestamp 1569533753
transform 1 0 3048 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4066
timestamp 1569533753
transform 1 0 2856 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4067
timestamp 1569533753
transform 1 0 2920 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4068
timestamp 1569533753
transform 1 0 3048 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4069
timestamp 1569533753
transform 1 0 2984 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4070
timestamp 1569533753
transform 1 0 3112 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4071
timestamp 1569533753
transform 1 0 3048 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4072
timestamp 1569533753
transform 1 0 2856 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4073
timestamp 1569533753
transform 1 0 2856 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4074
timestamp 1569533753
transform 1 0 2856 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4075
timestamp 1569533753
transform 1 0 2920 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4076
timestamp 1569533753
transform 1 0 3496 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4077
timestamp 1569533753
transform 1 0 3496 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4078
timestamp 1569533753
transform 1 0 3496 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4079
timestamp 1569533753
transform 1 0 3688 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4080
timestamp 1569533753
transform 1 0 3688 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4081
timestamp 1569533753
transform 1 0 3688 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4082
timestamp 1569533753
transform 1 0 3560 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4083
timestamp 1569533753
transform 1 0 3560 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4084
timestamp 1569533753
transform 1 0 3560 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4085
timestamp 1569533753
transform 1 0 3560 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4086
timestamp 1569533753
transform 1 0 3560 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4087
timestamp 1569533753
transform 1 0 3688 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4088
timestamp 1569533753
transform 1 0 3688 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4089
timestamp 1569533753
transform 1 0 3624 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4090
timestamp 1569533753
transform 1 0 3624 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4091
timestamp 1569533753
transform 1 0 3624 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4092
timestamp 1569533753
transform 1 0 3624 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4093
timestamp 1569533753
transform 1 0 3496 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4094
timestamp 1569533753
transform 1 0 3624 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4095
timestamp 1569533753
transform 1 0 3496 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4096
timestamp 1569533753
transform 1 0 3304 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4097
timestamp 1569533753
transform 1 0 3240 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4098
timestamp 1569533753
transform 1 0 3176 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4099
timestamp 1569533753
transform 1 0 3304 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4100
timestamp 1569533753
transform 1 0 3176 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4101
timestamp 1569533753
transform 1 0 3240 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4102
timestamp 1569533753
transform 1 0 3176 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4103
timestamp 1569533753
transform 1 0 3176 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4104
timestamp 1569533753
transform 1 0 3176 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4105
timestamp 1569533753
transform 1 0 3240 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4106
timestamp 1569533753
transform 1 0 3368 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4107
timestamp 1569533753
transform 1 0 3368 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4108
timestamp 1569533753
transform 1 0 3368 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4109
timestamp 1569533753
transform 1 0 3304 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4110
timestamp 1569533753
transform 1 0 3240 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4111
timestamp 1569533753
transform 1 0 3304 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4112
timestamp 1569533753
transform 1 0 3240 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4113
timestamp 1569533753
transform 1 0 3368 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4114
timestamp 1569533753
transform 1 0 3368 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4115
timestamp 1569533753
transform 1 0 3304 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4116
timestamp 1569533753
transform 1 0 3368 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4117
timestamp 1569533753
transform 1 0 3240 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4118
timestamp 1569533753
transform 1 0 3240 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4119
timestamp 1569533753
transform 1 0 3368 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4120
timestamp 1569533753
transform 1 0 3240 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4121
timestamp 1569533753
transform 1 0 3176 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4122
timestamp 1569533753
transform 1 0 3304 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4123
timestamp 1569533753
transform 1 0 3304 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4124
timestamp 1569533753
transform 1 0 3176 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4125
timestamp 1569533753
transform 1 0 3304 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4126
timestamp 1569533753
transform 1 0 3176 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4127
timestamp 1569533753
transform 1 0 3176 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4128
timestamp 1569533753
transform 1 0 3240 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4129
timestamp 1569533753
transform 1 0 3304 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4130
timestamp 1569533753
transform 1 0 3368 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4131
timestamp 1569533753
transform 1 0 3368 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4132
timestamp 1569533753
transform 1 0 3624 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4133
timestamp 1569533753
transform 1 0 3624 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4134
timestamp 1569533753
transform 1 0 3496 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4135
timestamp 1569533753
transform 1 0 3560 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4136
timestamp 1569533753
transform 1 0 3624 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4137
timestamp 1569533753
transform 1 0 3624 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4138
timestamp 1569533753
transform 1 0 3496 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4139
timestamp 1569533753
transform 1 0 3496 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4140
timestamp 1569533753
transform 1 0 3496 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4141
timestamp 1569533753
transform 1 0 3560 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4142
timestamp 1569533753
transform 1 0 3560 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4143
timestamp 1569533753
transform 1 0 3560 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4144
timestamp 1569533753
transform 1 0 3688 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4145
timestamp 1569533753
transform 1 0 3688 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4146
timestamp 1569533753
transform 1 0 3688 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4147
timestamp 1569533753
transform 1 0 3688 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4148
timestamp 1569533753
transform 1 0 3432 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4149
timestamp 1569533753
transform 1 0 3432 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4150
timestamp 1569533753
transform 1 0 3432 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4151
timestamp 1569533753
transform 1 0 3432 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4152
timestamp 1569533753
transform 1 0 3432 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4153
timestamp 1569533753
transform 1 0 3432 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4154
timestamp 1569533753
transform 1 0 3432 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4155
timestamp 1569533753
transform 1 0 3432 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4156
timestamp 1569533753
transform 1 0 3432 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4157
timestamp 1569533753
transform 1 0 4712 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4158
timestamp 1569533753
transform 1 0 4520 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4159
timestamp 1569533753
transform 1 0 4520 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4160
timestamp 1569533753
transform 1 0 4712 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4161
timestamp 1569533753
transform 1 0 4904 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4162
timestamp 1569533753
transform 1 0 4584 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4163
timestamp 1569533753
transform 1 0 4840 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4164
timestamp 1569533753
transform 1 0 4840 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4165
timestamp 1569533753
transform 1 0 4648 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4166
timestamp 1569533753
transform 1 0 4456 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4167
timestamp 1569533753
transform 1 0 4456 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4168
timestamp 1569533753
transform 1 0 4648 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4169
timestamp 1569533753
transform 1 0 4584 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4170
timestamp 1569533753
transform 1 0 4584 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4171
timestamp 1569533753
transform 1 0 4904 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4172
timestamp 1569533753
transform 1 0 4776 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4173
timestamp 1569533753
transform 1 0 4904 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4174
timestamp 1569533753
transform 1 0 4648 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4175
timestamp 1569533753
transform 1 0 4712 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4176
timestamp 1569533753
transform 1 0 4520 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4177
timestamp 1569533753
transform 1 0 4392 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4178
timestamp 1569533753
transform 1 0 4840 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4179
timestamp 1569533753
transform 1 0 4776 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4180
timestamp 1569533753
transform 1 0 4776 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4181
timestamp 1569533753
transform 1 0 4328 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4182
timestamp 1569533753
transform 1 0 3752 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4183
timestamp 1569533753
transform 1 0 3752 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4184
timestamp 1569533753
transform 1 0 3752 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4185
timestamp 1569533753
transform 1 0 3752 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_4186
timestamp 1569533753
transform 1 0 3752 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_4187
timestamp 1569533753
transform 1 0 3752 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_4188
timestamp 1569533753
transform 1 0 3752 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_4189
timestamp 1569533753
transform 1 0 3752 0 1 4200
box -8 -8 8 8
use VIA2$3  VIA2$3_4190
timestamp 1569533753
transform 1 0 3816 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4191
timestamp 1569533753
transform 1 0 3816 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4192
timestamp 1569533753
transform 1 0 3816 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4193
timestamp 1569533753
transform 1 0 3816 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_4194
timestamp 1569533753
transform 1 0 3816 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_4195
timestamp 1569533753
transform 1 0 3816 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_4196
timestamp 1569533753
transform 1 0 3816 0 1 4136
box -8 -8 8 8
use VIA2$3  VIA2$3_4197
timestamp 1569533753
transform 1 0 3880 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4198
timestamp 1569533753
transform 1 0 3880 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4199
timestamp 1569533753
transform 1 0 3880 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4200
timestamp 1569533753
transform 1 0 3880 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_4201
timestamp 1569533753
transform 1 0 3880 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_4202
timestamp 1569533753
transform 1 0 3880 0 1 4072
box -8 -8 8 8
use VIA2$3  VIA2$3_4203
timestamp 1569533753
transform 1 0 3944 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4204
timestamp 1569533753
transform 1 0 3944 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4205
timestamp 1569533753
transform 1 0 3944 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4206
timestamp 1569533753
transform 1 0 3944 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_4207
timestamp 1569533753
transform 1 0 3944 0 1 4008
box -8 -8 8 8
use VIA2$3  VIA2$3_4208
timestamp 1569533753
transform 1 0 4008 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4209
timestamp 1569533753
transform 1 0 4008 0 1 3944
box -8 -8 8 8
use VIA2$3  VIA2$3_4210
timestamp 1569533753
transform 1 0 4072 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4211
timestamp 1569533753
transform 1 0 4072 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4212
timestamp 1569533753
transform 1 0 4072 0 1 3880
box -8 -8 8 8
use VIA2$3  VIA2$3_4213
timestamp 1569533753
transform 1 0 4136 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4214
timestamp 1569533753
transform 1 0 4136 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4215
timestamp 1569533753
transform 1 0 3752 0 1 4264
box -8 -8 8 8
use VIA2$3  VIA2$3_4216
timestamp 1569533753
transform 1 0 3752 0 1 4328
box -8 -8 8 8
use VIA2$3  VIA2$3_4217
timestamp 1569533753
transform 1 0 4200 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4218
timestamp 1569533753
transform 1 0 4264 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4219
timestamp 1569533753
transform 1 0 4008 0 1 3752
box -8 -8 8 8
use VIA2$3  VIA2$3_4220
timestamp 1569533753
transform 1 0 4008 0 1 3816
box -8 -8 8 8
use VIA2$3  VIA2$3_4221
timestamp 1569533753
transform 1 0 4264 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4222
timestamp 1569533753
transform 1 0 4328 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4223
timestamp 1569533753
transform 1 0 4264 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4224
timestamp 1569533753
transform 1 0 3752 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4225
timestamp 1569533753
transform 1 0 3752 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4226
timestamp 1569533753
transform 1 0 3752 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4227
timestamp 1569533753
transform 1 0 3752 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4228
timestamp 1569533753
transform 1 0 3752 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4229
timestamp 1569533753
transform 1 0 4264 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4230
timestamp 1569533753
transform 1 0 3752 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4231
timestamp 1569533753
transform 1 0 4328 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4232
timestamp 1569533753
transform 1 0 4328 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4233
timestamp 1569533753
transform 1 0 4328 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4234
timestamp 1569533753
transform 1 0 4328 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4235
timestamp 1569533753
transform 1 0 4328 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4236
timestamp 1569533753
transform 1 0 4328 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4237
timestamp 1569533753
transform 1 0 4328 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4238
timestamp 1569533753
transform 1 0 3752 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4239
timestamp 1569533753
transform 1 0 4264 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4240
timestamp 1569533753
transform 1 0 4264 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4241
timestamp 1569533753
transform 1 0 3752 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4242
timestamp 1569533753
transform 1 0 4264 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4243
timestamp 1569533753
transform 1 0 3752 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4244
timestamp 1569533753
transform 1 0 4264 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4245
timestamp 1569533753
transform 1 0 4456 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4246
timestamp 1569533753
transform 1 0 4520 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4247
timestamp 1569533753
transform 1 0 4520 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4248
timestamp 1569533753
transform 1 0 4520 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4249
timestamp 1569533753
transform 1 0 4520 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4250
timestamp 1569533753
transform 1 0 4584 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4251
timestamp 1569533753
transform 1 0 4584 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4252
timestamp 1569533753
transform 1 0 4584 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4253
timestamp 1569533753
transform 1 0 4392 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4254
timestamp 1569533753
transform 1 0 4456 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4255
timestamp 1569533753
transform 1 0 4648 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4256
timestamp 1569533753
transform 1 0 4776 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4257
timestamp 1569533753
transform 1 0 4776 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4258
timestamp 1569533753
transform 1 0 4648 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4259
timestamp 1569533753
transform 1 0 4776 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4260
timestamp 1569533753
transform 1 0 4776 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4261
timestamp 1569533753
transform 1 0 4776 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4262
timestamp 1569533753
transform 1 0 4840 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4263
timestamp 1569533753
transform 1 0 4840 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4264
timestamp 1569533753
transform 1 0 4840 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4265
timestamp 1569533753
transform 1 0 4840 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4266
timestamp 1569533753
transform 1 0 4840 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4267
timestamp 1569533753
transform 1 0 4840 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4268
timestamp 1569533753
transform 1 0 4904 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4269
timestamp 1569533753
transform 1 0 4904 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4270
timestamp 1569533753
transform 1 0 4904 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4271
timestamp 1569533753
transform 1 0 4904 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4272
timestamp 1569533753
transform 1 0 4712 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4273
timestamp 1569533753
transform 1 0 4904 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4274
timestamp 1569533753
transform 1 0 4904 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4275
timestamp 1569533753
transform 1 0 4712 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4276
timestamp 1569533753
transform 1 0 4712 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4277
timestamp 1569533753
transform 1 0 4712 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4278
timestamp 1569533753
transform 1 0 4968 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4279
timestamp 1569533753
transform 1 0 4968 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4280
timestamp 1569533753
transform 1 0 4968 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4281
timestamp 1569533753
transform 1 0 4968 0 1 4904
box -8 -8 8 8
use VIA2$3  VIA2$3_4282
timestamp 1569533753
transform 1 0 4712 0 1 4968
box -8 -8 8 8
use VIA2$3  VIA2$3_4283
timestamp 1569533753
transform 1 0 4776 0 1 4968
box -8 -8 8 8
use VIA2$3  VIA2$3_4284
timestamp 1569533753
transform 1 0 4840 0 1 4968
box -8 -8 8 8
use VIA2$3  VIA2$3_4285
timestamp 1569533753
transform 1 0 4904 0 1 4968
box -8 -8 8 8
use VIA2$3  VIA2$3_4286
timestamp 1569533753
transform 1 0 4968 0 1 4968
box -8 -8 8 8
use VIA2$3  VIA2$3_4287
timestamp 1569533753
transform 1 0 4392 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4288
timestamp 1569533753
transform 1 0 4392 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4289
timestamp 1569533753
transform 1 0 4392 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4290
timestamp 1569533753
transform 1 0 4392 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4291
timestamp 1569533753
transform 1 0 4392 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4292
timestamp 1569533753
transform 1 0 4392 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4293
timestamp 1569533753
transform 1 0 4392 0 1 4776
box -8 -8 8 8
use VIA2$3  VIA2$3_4294
timestamp 1569533753
transform 1 0 4392 0 1 4840
box -8 -8 8 8
use VIA2$3  VIA2$3_4295
timestamp 1569533753
transform 1 0 4456 0 1 4392
box -8 -8 8 8
use VIA2$3  VIA2$3_4296
timestamp 1569533753
transform 1 0 4456 0 1 4456
box -8 -8 8 8
use VIA2$3  VIA2$3_4297
timestamp 1569533753
transform 1 0 4456 0 1 4520
box -8 -8 8 8
use VIA2$3  VIA2$3_4298
timestamp 1569533753
transform 1 0 4456 0 1 4584
box -8 -8 8 8
use VIA2$3  VIA2$3_4299
timestamp 1569533753
transform 1 0 4456 0 1 4648
box -8 -8 8 8
use VIA2$3  VIA2$3_4300
timestamp 1569533753
transform 1 0 4456 0 1 4712
box -8 -8 8 8
use VIA2$3  VIA2$3_4301
timestamp 1569533753
transform 1 0 4456 0 1 4776
box -8 -8 8 8
<< end >>
