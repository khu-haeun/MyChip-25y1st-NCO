magic
tech scmos
magscale 1 3
timestamp 1569533753
<< checkpaint >>
rect -485 -485 485 550
<< metal2 >>
rect -425 425 425 490
use pad80_CDNS_704676826050$1  pad80_CDNS_704676826050$1_0
timestamp 1569533753
transform 1 0 -425 0 1 -425
box 0 0 850 850
<< end >>
