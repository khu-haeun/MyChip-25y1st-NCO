magic
tech scmos
magscale 1 6
timestamp 1569543463
<< checkpaint >>
rect 132 -122 2268 5180
<< metal1 >>
rect 352 4520 2048 4580
rect 394 2960 2007 3020
rect 394 1400 2007 1460
<< metal2 >>
rect 252 4581 2148 5060
rect 252 100 352 1560
rect 394 140 494 4581
rect 516 180 624 4500
rect 646 140 746 4581
rect 768 180 876 4500
rect 898 140 998 4581
rect 1020 180 1128 4500
rect 1150 140 1250 4581
rect 1272 180 1380 4500
rect 1402 140 1502 4581
rect 1524 180 1632 4500
rect 1654 140 1754 4581
rect 1906 4579 2148 4581
rect 1776 180 1884 4500
rect 1906 140 2007 4579
rect 394 100 2007 140
rect 2048 100 2148 1560
rect 252 0 2148 100
rect 1906 -2 1998 0
use VIA2$1  VIA2$1_0
array 0 50 36 0 7 36
timestamp 1569543463
transform 1 0 290 0 1 4712
box -8 -8 8 8
use VIA2$1  VIA2$1_1
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 820 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_2
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 568 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_3
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 1828 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_4
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 1578 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_5
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 1326 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_6
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 570 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_7
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 822 0 1 4260
box -8 -8 8 8
use VIA2$1  VIA2$1_8
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 1578 0 1 4260
box -8 -8 8 8
use VIA2$1  VIA2$1_9
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 1072 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_10
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 1830 0 1 4260
box -8 -8 8 8
use VIA2$1  VIA2$1_11
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 1074 0 1 4260
box -8 -8 8 8
use VIA2$1  VIA2$1_12
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 1074 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_13
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 1830 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_14
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 1576 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_15
array 0 0 0 0 17 36
timestamp 1569543463
transform 1 0 1324 0 1 2304
box -8 -8 8 8
use VIA2$1  VIA2$1_16
array 0 0 0 0 12 36
timestamp 1569543463
transform 1 0 822 0 1 3324
box -8 -8 8 8
use VIA2$1  VIA2$1_17
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 570 0 1 4260
box -8 -8 8 8
use VIA2$1  VIA2$1_18
array 0 0 0 0 6 36
timestamp 1569543463
transform 1 0 1326 0 1 4260
box -8 -8 8 8
use via2_array_CDNS_704676826052$1  via2_array_CDNS_704676826052$1_0
array 0 0 0 0 42 36
timestamp 1569543463
transform 1 0 2078 0 1 4
box 0 0 40 40
use via2_array_CDNS_704676826052$1  via2_array_CDNS_704676826052$1_1
array 0 6 252 0 31 36
timestamp 1569543463
transform 1 0 424 0 1 184
box 0 0 40 40
use via2_array_CDNS_704676826052$1  via2_array_CDNS_704676826052$1_2
array 0 0 0 0 42 36
timestamp 1569543463
transform 1 0 282 0 1 4
box 0 0 40 40
<< end >>
